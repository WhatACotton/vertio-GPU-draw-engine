`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
VeuanPbjmKcok/GWGxwteSf9S+IxCWqpwRfef2ZTZzFuOm/hoC5XKHSBv1pWKlbtJRmRpU2KulnCnG7O8EzueU7hjWx7K/5+vMbJSFYVOkwlu1VT5hxwzGBTsUYGhFkFKKTwLKZI0H6n+liYc7mxvwvPEjGoosg8B7PqOmSRC9ZkM0VysVTE6+BCXo+kzahNpkYpVR0rOd+i2v0Gw68ygRnCnzwd8PC50iM7aEp/GvDL+1bmnT3zFr7yphb/9RwYAK1cxxZODJ51ALDekVs30xZwa4Mc0iDxl/LxNL+KNK6/mbZwO2OuUiZZSC1C180sJ0KV+AjJiUaw+lzuy8DuuN2vjGu0KcdNIiYrpo+RBHEefe6uyQdGvu0M81Y9bYygAcVDSVu4buNjyu9Bafrw60lztdbcLNoKaxAVD5ids7OkiiG7ec4yL9CdBw3PuY7xZi8i7PfdCONH6k3UTiOmpIO5x4/UpmFzVVPZA9DmJDmaWqSqZRoUA64RWdURBdrKK+zTPGpW+xyBr0ddyVqySgCtnRNhqcMDem9XTM12oq3FbpLT8jDX/wJeAxX0bEjkYKoWVUjaAkqWXAZBfoELaEoxhMtCH96mZsrNuSr6/S+Cic5KPkTvIr/CVTjArINs7x3ZEuiwHVg62V5aZAm6LtgWSwb6AwkjcR/HtxxqMnM/5DZIiLTwiA+NKow5i180mXoQObEjDYNtczqV2X3WLfD1xYGk0qwzjKoVwraJQ44x/Pjs6hY6Nl97D8lnCiFQcX0kFNyErLXd6WMHaB7wxDNKBi5NbsFydX8ckSYWwim1mnMCDqI/h1NWhFwc3gta2hHT2MgpbM0b3V2x6Y3NszPTalxP+bKjc4BJPeLC6SeP5113oR7LK2JBs2gsrHZzyqb0YDRD/0GTR/TORQCUbnIpt51HBCyiLHgBukqVhwTBI/vfuJDciZ0g5f3wCb9N/qjbsylbljsLZplhec0HS8IfDhq8FsTp3ZFsPrdLVdlGinR1uUXeVxictMQUVMSywxisRRPKRuQoqWzV42Q0zlOzrgKFPkmSiJs7Hg3oCLVSaGXXUSVorhb6CwmdPMdcisj3MQm7xak9bftK8YCbT2R6PCm9R7XeqtkxpRfO+hAMJScDX19a6hGKfNF5SIInr6qfQXk0Gaa9EqKAJAo0pmrOiwm6HtBCoQwQbfbJzcLb+bikj+glm9MZC1duxtBbQpom5sYRstVDp3IDPup3ZdKM71OdpXxv4FcpFefUsjf9V7hNFmvUFQD3MA1TaOk7kQNW46miLyPVxL9an1MY6gWQnIb8JbYki4FyW2ZvzxuaigjsF014CJu58QJeIgCZzKsOi4eD8wDK553hfMO7c+HChb352Bil8EDllpHQw3EsdbBpLDVLbcvypKQywFvf5T5Xdr+O/2WveUNmJHONKDZQ4+fI+79i+nU+op2d2vc=
`pragma protect end_data_block
`pragma protect digest_block
b11cc712bbf8f7531dc41f91834133dee33365662cfb4380bf13fcce01ac5d05
`pragma protect end_digest_block
`pragma protect end_protected
