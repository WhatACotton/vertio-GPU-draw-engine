`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
X6QP7a0IuzOzl9QyxiPJLP5tTyNm8fdVGtIqB3o6qEj+1GXw9IH6ACmS2Vc4hGdlsfEtXHzMRpChp53FJ9oWoRXIzW37FbLnMt2OvAUBhd6BFD9gaHaPsG75uEd/BDBt7kua/nytzxPr6W6itGnl5YNMDA2Vl6cuDboYyDceopKKJlfIS3ROexAZ1niXBMVaMsgRJS5N19wKmyqX0miuoO/YWchDNWphthT5T+S79616GXoBC1PDrm0c0SlKqiGVin7xnbfm4tFAVeD76xnvPo1Frz0dyb12vApxck6EqaOqIQuvd/S/MD1oC2fxJP4woktv0kY2hanWy2fUy8uhk2pSIjz3bEiah77wLBhdrgDydqUaJh2wRH5GoHja/a2auK1tGMt6NtoBv6UNxXQbRdh67QN3c6G8+LTPxPb0TuXldoZvbgKuo4adVmb0jpmsKryykj+QagAh/bQbNnA5rtM9f+C/FUbtMDBZftdja8xe9f33fag44PA4tDLVsSuXor4WSIpWqJordQD7se8LpH82F6PGc4EfTDfeVqq5v4aOFmEfxCeQk6kWDq4egi7FpAjRxTOSOu4/6ctvwvfp8ireZLzLeei3hb5HIoNXKcD9209UaUauYTyYPq7GsX0v0hRe9L6LMKqW6tZiwsBj8898btI9Fz1wYv1cANv0dhsQv32E+fggixpIZrf39LxL5zp41JqtleaewsUO+1bbL6fJXBo3JUdTffiHoEa81mhGmbtU7CrMTnQXD6MtiNUfT4wdVex3TOrIJO/mVSnJM84Kf77ffaqI1hOkTFjqmXYdeUTZ4k+Hha0yN99+JdB00mx7T2aYuPxUPnU2x1/t2leyEfXhknavtte6r2nyTC/sYjcJsdcWmN5VDv/RECn94oboZANEwYHF0l6JUESfPHMNRT0o7BQk8iDes3MY2L7mYJCB/18H3Ke4YNpEubulWgfmDr1I+gY+dqwdf9Gw/eElvXNuw+YeWvS44W/ixRiKTTS1fLRJ0HHOw017GVrfyhemHLo6AaBx6dkIpdlYhvUNtDeUgIUe4teojvgMMzcsrdiGb3kK6mJGTaMl35ry933TpW6f0zkWtJTu1k9KK4f6sWdtOdocxJGV/I4ngjDxmD0RgEww4PyFA/UTkD5LDEm3Yat00GLVU6Bxe7hhPzOzYVtW4TWZ/yh9wTXOxaGnD41SdNJXhozwM3iTno2qyD6Kr74sjByNMrwprTG+TSqu3hTs5ogYz7lq76gr34GP7QsM6nLECJ0qymZIOgkU5NJK55LXnyW4AXyYwMiDnE0j96k+L6hcGaZY8M6FgbJWgeF/piJEoH1sTTAVk8TmBk4r9OPlnvmvUhNScAcP596i+8GCGmBzJw7++genNQ2MceJXgZ6sN1z6oZNO3//XV9JJFPCKhfpBOI0Vi+AFaRKm+bsDofotllvVapP923KOvDCxEIr8bCk6zNsKJeSznysDiqIva0A4/WF8+ILN67MiqhUlANA6rm2IFCyqnVEHMIE/34qd8T8MMvfayFMNQiI2rMEytnftD30nd8E/jpck3fmLsSnKbFDgvVWaVO6ILaEwQljApVL9XQekKyRRzZzQI3HBiNgz02Z6O6pbdlTv7S5Fud6CxZh5NCs7EjGAI3yKqvizrhxJfSG27knFObA+fz+bOkU66vaU5l8zNr/fLRwEvVE041ukGmzxErJfE9GaCXincpGcGbJA9MXZ0yVYiuRQj2KFSf1o6RJdr6fBAu9VSeFbZ3lBR2WQZ3n9fMkmsBZipnWl3a2iKVJMIIy39z8JQUWJo/bP1FQYGEbqB5M+rzb2lfh3zNhXxjAwcFQnCQBq7RN2kl4+nhjBRYrWpgBw4WESTS86EGB5HaxY6fcLxCY+H0/uXFq6YBOzZbBdnLZHjEpdTy5l2vp2myAdIBdXvgBcXmX3BkZQC4jAmtyXsEFOxzWYRGdr4GNH8B1grAw4V+MT1grUmN4Wt2+vjqacyvGK06onsAsGRvBKHVxYO7cioa8G4fJaa7U5sGNaNHzy7xVfbUIRAYoKxgfYIfJMRz+xSyhK1lpWujRLiI7whH0PN3pHPmhBLstfVQMGAT3inCokGecuPq7HmEihvYJLxvhbBSvYs5T8GZN9HBUS9T1HxPDr1bvMzNUXdmkBdl7rHWjtSXMDuUaLH+TldWTk/kNXs6c6jpj9uhwovrXLF9cdMiDU6ltlPFCg5gXifdozVDBZjcuk1n2HdLG6oJNCN+oxhACjIkQtPnR3YIRGn1A9k/Q6E01WZjxx9V12xO1ro+DCoLEx3k4tEuYWuyHKCMFtVHcgIank6mxRMr+43na81N5A9+/d4o7l84WyLnvaVawOw4MPzjSBxGOHAO3l3Um+DUW8Buzns/HkzT5Q0NTfhkP8pSwLyY1cdRxCegKJF38nAGvF5YJOcibUEhcZJBg8Be+Do0VhseZgU7Ny4puzyMl0Qzl1RUkFHPft93RbvM9UKGZrU50/FPkbfMg4QZraR3cWghsfeW2y2Ie1S3rCtw/KNGAZ3dtamNeAjy6OGeoSW4QZerW6JzqEOsujSPAeIOl1kHQUXbVFQRUj8nNvMX/DTA8FCzToeluMCJh1wijD8X3OhjOLQG6adE1yHFmCgYhmInlJ5dvY0idkc6Lv1lF1U9fFcyomEBubnfJOYJ21iG6ihpMmHC2YxC9wRhx8KA1aBIj4kOhm9R15F6lumhi5gBjJKEkmTVb4L1Fsmdiaf7QGKEmoNN1GVPOpnY9RX3NksZf/5P6Mui2CTmFB08hybu/pGHlYcRSTJAjC8kYK2v33/z4ZxFL7F263ARzh+f0soiSD9rxUa1fzd2/WfE/NCHTeFkM0NC8ETQvQsiMmcgmHbmCsePzihpKX6KLNy4GgEh4aGRp2P1uQnYWnhmeWodCo04acTbxWPZGhY7MJrApymobL/2GQSFsN2LR/0WfmoxGJcBjJCqmh+0FkVr2dnPREzgytk3XxqQlLUg0GS3uIxKXYu3mKLjy74eRVpOGXDDFJMEBcx6De8EigHd8gcXZje3YDEA+jhEnf4SSZBu6GBKaunPdcng8EmD1ARwwhs7YEmCp7KeBYlicNa/lsoT0x7BLCjrDNHv/uMRwqnDa1SBlNr08gy0NmozjF4GskDbwAIb7zXSV7QOTABaZeZowumGJjtpWJG5zrR8YH1M6dQTVS/KI8D/xd7eZyol1xGpaMa/PP81GvK+9EnvUI0S7XmI/b5mgu2TclEhLVYK3seBEXYBRH8GigflAgH1mPsH9nhd2CSfNk0fvL1KUZTtTuJYL6y/MwrQfJrnbMfygXJN1Jb1soiVjv6viAY+31Yyw9goToklwm2NOWCXfax2wE/gW3rFDvQMWMHJGZd7a6Iyuvjik692SZ3l6CNg9lRmJ1GDpnLLIclAl1rcLMXQO8zxuqiFKO2rytRLUHfo6v49xzsCsuaBeulP9c53keZwX4yldlL4K7cclMPkMwEC4toz6UvnLVsMCgRP49CWwm8xSk+oenSq3nNEkOfgf3zZERqpRR8utwFsVG8Co5O+TawvheJ9Gqk+JJnPoiRCywHUMmgJSYZBICnETHvga5gUfcHxrfP7eB90f4KdAcQYzNl+WiJYDMEiVcYxCjryHflEvbus1RezWtIxSaRNxiSZxRcxYh87Ry3KvDA5Sk0YdqwEER7XyZs0B4v57CIXOxnUCBVYvLY0At3oP6Mx8ofCspp8PoC6K7YM5ua8eb4EMm0z62UpX8oioX47buGZ23vMNAqppKvey7xuwsNpjnOac539NEYjSSt+04Qm76uiYaOqmIVqTAsalVbGjpciIEBevABp6dpHJO4m8zN9QiGVw3qlnjhNf8HuHn+JYLZdNNt/Vn65I3ym+uAb/BsJBsYBEpVKkxDNPtcrSCEfFW1cJckUxK9/m9aNUXBuFt3X8o1Qo+tuR0AyWxAEzglrB6ihEVS6GByynNIPKHbBW4s3EaQOjI9J5azqG4hSu5N3NDe03b87VOX5ZBbCVstnuQu/uYPjzPHlalouR5nsIewd4qpr5uaje1V1YOBiru0vYqrWMxElByBZhL2D8nlmX+woBs1JcBD/M899FleIVLtzqG9T/hNtylZxMpwtK78k5gcxHh/yqsh0sl8ThjDagt2IanzQkrlLRrvEEK0wYwAoyZBHLVRsMRBmxPREY0LES/ioONDcLNvcwcAQ64qCq4w6q1HmzUZ4In4L/tVBoKHSwZOhelJ+b9l7Lj0RcBpK0D6orIAHCy1M9jix8japjppGOdC2+69HH9vodPpJsYmsUgTGogdfsnRYmVyz2Vt41H4sR+wWNh+F0R9i45CYvBfwuau7cspXZJ+Re9174qmXAPV+bUmXKOnp9EiJh56+fL5p8+63pw6sssVjEAfycxwWs5l167/6kBLAvt39D6/ofwbMM0QorC6blSwPpOZKejDN7P5xX1xMYOyprDsMeMo2E43qJjQHlAGfuAByNkI0bzF1+1sYdch02UbNTBGnRE6KfrNI4R4RAATw+v8MVcJiDnW6sLIC1U3PSY0DwPeH/bfBaKgipjvSEtN1wMj78Uy3pryCHUPwXxtUvunavIqOHvLSYfmFotHSILd70JENVyCOKRAF9hqA3dkX3Yhb5fqfEro6n5R9wHKpxQqZkRZhAkb+3Xwvi0GKLP3A2ay+GQwPPc0/OcalreY69zHNPxJY31HGoayso2zHHr0/yxURuXyk7qa0o4CQ5RqY2ozfCC4aZcdqyKgOWoy51n7+XWhtE+9twCwuInjZf2mad43eKKBIywGtUC5MHLiRcxMGa1sQI68ukdAoT4x7HSh11VNCkTwTt4MwyZEMp7KeK5pwCVUcoBtbWuVu/bW0G0X283k9W8iYsDxXPTCxNy5XIbtUUC2Rs6msubyghk2bgidI1Dm3RL+VM/77npCES46hrf8funUKuzEyboliqtOF0H1ORaw7AlpaM6KU4LWqhtKSB2yVfYx8ujv+P1VTOvlKQ2WilXkM+o/XU+9tW23jl2MXQSudsVPuu+c3ZrTRX/M0xBRqSiOXAAQhBOkRDSrKRwRsoRkeNdsMiLWDPhZJi5QJgXuJD3y+jKGV5QMIaD8Mra0t3BwxKzzqvEHjm7gJCrikUyKZJF7Lg4KkyVcXHrb7WPro2laSWJMakJajP/EOCV27M79e/eFBgGvEIJjjABTfFmThYCU8azJdLSMJ5U+/NusSnZYeMzGXM9X8Gs9M7/j7w/fbzCRxldQ9Wx3rUVNAcwMefv+Oi5l4KI4OohONOBKc+a2migVXak4radWPtDKAqZBvaJh20Mka9huL1Of1dneKMvionfar6RViW48mlafhTRPtVtw4tUkeITs8BIwCQNLh2Wc7KSXmLpLzHff0EhzGyazBDIz9LOHvWG7NO0YMLv1bFtdJ9aafpxCAfx4Oy2C1NcLiPaPL9rXwc2tzcIUMXs+9i5dcrn45pi4J32tzBP1ZHDIIxnLontvHhQqz8PKlPe0VkZods8PGVWn7MchfeoYpsI46DTox1FzxXJib5WBnWyTiK/SkSP6a/nMTa2tXK0LjdruowKaQh6XGWUHzazN4pI9sfu16t1eun+f564BYpAfrhzSzukB9/LfbSelaIuAiLR8L2HE5/oy+zwv7KcYAZUvEO6ImqwBgi3LOfaZfxR2UV5qi+0ON+iKGKBZuRmhFwPgpiskQ645ZNQk+64aUkQaqxgBruAXFOb8TQlXTqJ2WHBz4k0yt4nqTrg+fq4EzOonuLFKux4tl8B2wVUzUXgzoJo2yKgMRhl+FpHj17fwTkg9sshSJiNKNqRW43Kh2MS7gThcnT21jfzKfxychWp/BSWsrxJ3eUpzyn9wVgzUxdNsQSwdj9HodBH+T1R1q14dcPi3UGpHSlpQDW+W4XnVv52sg9SjWgnW4AwNqVKBaqoZUM1akidtnHZPMemsmNYcRIOEu6sJ/ogzspr8w4a0TbvCDnwJWt4Z2fEFBHIz+aC+wU/2NE6gBlitiF7eM0PJGG+0NcP4CuJgWWnwDFSRcia83KUfPTnEVWN4VoMl7mhcbXOGtExysogJyOfnDbvkUGDuA+AStkUEcvZFjLowOp6Dqyhdo1jYPmH64kcxfCFB72FxGQLUEP1Ep0xggn4pMaMPkzH/wmAIABwTXu2iDsTJzdKspIzqm7/v68W0NnuW5YmCXwiFYzDWIMBe2DylP435H9zNRsVtEdUGgHA7+vekWCLLRnRbgqpkxtMcmbcVQomrGsjOtjBdBcsjhIkQh3850RGm0xMjVlwOflCanK/Lb1iHol+D5YFEvEEEemVuGehWfoUDyHolkQt0wVBNXRbnbQg/l0vGKZMHIRvIw0FHc9g0LWWogGTEBulTkMpyUjFCBbYi4VV5BsnsAqe61w0by3JpexHlWVZw016SjfR8AQCGo4mtcJnUhWhwH0n+lpSU1COAr4YNZvj1nVOHzmD8HbAP4zKe+9Jkmr+1hYAkV/KA/zzV+6X8UZwb1AE3qYK9PJCRPvLebnNIU3wba4bV8WO/pFSylyxnBGEMW1zyWqbYIBTD6i7x01rUAB7kDwPFOsOQZVjvkDch72BoEcHy7pmvaTonfObwdBsf/M6/7Ko7DM44n/38jPTQsTDhzlRbIpbc1wEpBx2PcgE5VOBEAcSvD70/MtD+5qmcK/kpoWwSR3xqa27G+tqu5MPSeX05kf+VwT3uMFyU/iK665M8JfmR+ky8gFqbN21xFg3KUnyKodwae/pAJrMQkW83EFMvDJhStvMVkfM2kkOX4xhYQHpAz/ZG5LSM1QkcFqmTCgAC9WpKTEIMkmWw6JSoRgt+sNxZCW5vRIabdh+sTeySjU7tUVW/gbz5ACq+BgEyMn3uU/bbVoSzAMns2dgUKUsXE+fruO0uXEOQnwOr/tABjZDsAEOwi65wUo33XAV2YhDDKLRsjMwv/Spp40ZH4tbp2O0nLObrCgPINsNVid124sh9ih34f5dqm5kUsRN3bk4V9cAmGx8oXZfS9esu4L/QLxwqvVjHrVrIXitYscf7KNyLv1N1MlATos2mW61VGPpIDK1+E5gRER0mGAAvCVnCvC/PQ1OhcbDr1mzGKcWcZJ/gCjUaqwKFVAahP4WjmNoaU3QbguQqoHR1MUv3/Uhxl3XMlcnnOQV8Mt1Shx7o/7YG9/fOvIDQcG3eJbYv52i+DWIsyeQn7dE4xDqSKnPmAfv8qwTqenEy5IZfg0GEUb5Y/LAwbXYklN4n5vDX0yEwSnKWpm8O9B3NhsT6OgpFWobNxczu0s6iF7LGChzomJYMl27ukZ0a9WbLyHCVE9jq/XyS3bnFoteDXdvLHKzccnr0YUc1xLww/eKstRipsUWlL8IxVOUN2rFJH5tuuuNM0ix+Lur/J5d/PqYOeYRIg0qe8sj4yKs9Up/DeAg+WKRNZMm/1moi/x7MT32viC1CTR0+nURb8eMmA2Ez3YYJ4+wqM93GlJLQUSN9w+exABBkPREekUja2GvILv/YgtjCnnzEgx5GRs2KYNxD/1XiBGEwoJ2HQNEPJERSkTb4GIuYmE2HY6YXpG3Isnw+Gz9/Iy9SjAfuz1TwbI7cX+h6mOgScAPfadIAEY9pDOHoq/lsWEY5GvXqdBTl82at33QRji5mOT4r0nh4R7dKc3jyscOUEFZ95ITk5kNdfz/+hLE64nNXW1WWepDV7e/sdF/PtkU1u2LTDSrqd88LwkiHPe2Db8lvZTpNaxt23aCKYwgZXm/ctHKgTHiZJuQ9QPXbFLPIUG/Sa7axAIBIJYdTXJBX3jM3M9LKx01Y7BenpGZklGXFss847Wj0fZ3ygDn8KEEoeHfi6mQpmn/0OLvACLx3JMXp/yTxfpfKIO26llyM6nQUO24TfyUcyyn8lmvejRChXSLcUL9/p1urXYmxXoefn1+yDR1wQJtySJxYhffVvOtD13KIr5m6zXMvntIW7DquBL/vxnn6cthUJIK1903LRBw7iYOMSo7FigrljWLfklJ03/ZIuSr+QqZwiUOTnAhuT2P1lA/7MojS85abnhwHGsakAH78vdjZHo1sinOMHzgW6D4EBcxvxFaiY+Bx6h0pXHEXr4sobMUzyS4DRf9ZiV0THOv6fnJ5ZcGQYWoMIui/OcKWyyk99ZsY4ds3yOw0d8gt+3Jx+W+pGayopMrs3r5df0RgdXyNUgdqgmp34FoCoyW/+SL7Y3rRx2ZgBi/cveIol+75whDjyp47K05qSt0Li1GZcXmEAvLJre3wGOv51nfAlEt0/5dWro80F1AWejj4GlKbni0M8FBy6X7Rdtqw4NRG4zM1PWF6GmMNTi863Ne99eBohU6D7HItE5to1Hv5r6BDVngp68/brhWSJvKFQ/eOESvusqXRtv5dKQg/KOBwhD7wt3oydOP3SO+x5D3pOxUfCnXqFC3neGkOi9jNXoA3BlIMjqjOdDvzzGE2bXCeD61LOBTp649q1zlvK1iRMIdqufE8HOTmeN/eLJNkVWx09+8bJJWr8nMShOn+/VZRGgvKgUHpQZr3MTFi6v9o4jl8cwdocY51253wuIo8MMQYpc0LTlP4y87imO9aI2MEsUWI0VIpv2v4fOj6fPg0E+BwgCuCl8fS4bLI6lXuSaUnJw17k5izYSVD9cemR1hAHkbUeg1Lyd9MmsRXlYWmTGgzlMdhD0qYxxQSesDcCf69zqLXxMELqZtY35qY9ppOlS7yleA8XxzZQUXqGYAD3/FMJK0LIEg+7kj5s27A9wURsbhM1D3JhpkLpbseZcvOTKPzUHFoWcohEF3PnPlv26WScuV0YZi7/2J9KRAzA87I6O0+TXa1JJpEyZFSkajm6Lci7BsVgk45ncGiCMprwj/gjLnYnfhV8TXyh52XPw8WyKDkG32dsqtchqbvXBl/dXc1j4+zw/5pWV9E/c7l3J7Cmub1DFu/MmuQbTeO3szzKt14mW69Sf19yWqqXaDh6jKvhi6Eo9aF0WTtroI6QPk876YxKW/47XUoQjs8QqiwD1qAhvBWFQ66gZ6Vtx+Gx0sJJ63nqrjp8LXBosS1z1xoypBtPHzyAOMBVSzXTgQ/O534YmEcNxthX7DqjbG/DwMTpT06SSE63a0C36gl52ZbMjcbOUCE93/n6yx+ana0CCNY1Wif4qBxKC5uBg+clET3mvjZ9vky9Sji2Dtt4tRW5elmfDnL3t5IhN5AZ3jGs7vsBIEvWsMfvsW6GYuyguAzNzPCs269dkLgdyrG3C9EOVLduJWFrBrqD481G04lq6eQV0bNVlv9zw8nnlLtpW4L04xPgwZVnP7d8CkTRkJejMZDphiruZzHoj/EgsNA9MH6r5VYt4QndwZllm/afvLfHi2N2Tnr2MFdYyS2PHWWh++EqNwb2xcyT+jo7t9OEa/t856PPZyfn18zfcaS3UxsWkZUodjj98OGcfrb3BhpO84fJcWiv9yPlotOTTCeNGtz0py8im1e4oBdogXm7xgEIW2QbyoWBvznftxjNYfufB0ErLl3qpUHWfEE6+Ra1cvY5xSyDksGxohRHRnAvU1QeksDLNrriTcrn4TcrvprdRYIFEkNSTvcELdfi9CivyGuQgTuuJqCMjsbHncZ1a7u7eps5wdoS78hBgX5tJg5q7uk2BLEYWTRdc43cVLBtN2iRiPn9zEaLQuMQUq4dc4snev3bD2xrCW+OpIarx2TBaqMS3agbtrW3GEpLpumQYBdyRbKiuJi+9OccGkuLMX/zgrLtvalT85zTCF9Ap1QyTF+zQuajCHf9cs7ucBVvXNon+ngmdSQbbFCx2wyyytEGtF260Fw5LZXoAP6LIhQW5mMv2IEfoU2ZIfiaaFgc3w5i+qFMyog9OmGyYx9GUKDKfznHDC9q8ERXkSqy2OlkoKf3akoSy7/SWq21z1oWt/jvPh4tgPqPCRDK62SBMl3LwDQhqPWB5FerbZ5IB88JimOIQrTVR9qwV1Duh1Am6dLaicAIH/SZf+IZCTCws4F+pEj1sKT0llnNoyaj9reKWNGf0VfXFt2N9oN2MtHynAuNWXDaPTKBB9JqRJWq3bRsa3tux6oyvH8td90U9W6uiALY3eREUh35pPy4v8b7i7O3+4Rm1AE/MdQSNPlecbaAL+x6bHDdbgdC1lH/dj6NiwoIaVyn8qOXBtiV1vJyMpLkaZtlyt7duERDzUwQw/VEv4oVN95pO6drV9/wLyhv5RQCElFdIldO/u4eXG9wW1Jma6Bkia6ao4NfQcP64cjIEIRsuzgm+KLtdDRYYX0A3/BoJjKwwOrId7dYq3nkR7RNKX0lsa51JJnxXyYsEc0vF4yI4anO/U04VnrQoJa7mqAiPPZ0owo/CDPGSOWm6BFqZ3UDnwsJwGDzoW15Tgic7IfcLaKUvuBkvl5LO5c2eQDVxpE1tQzgofmnCvaZOYC82DfjtVtaZ7kuq3UxGOLS3YoqhSF+8sY2HRc8zuqfuFEpEYrqOSNIqpP+cpv6/G14oibSml8cppzK7hH27Q8DQXVXxIxPJKUw16iqKxOj+EEbLCRk/vPud0pJXVSji0kMitQZu5Ke4Qlc+rK4gV429eCdfn6flumBK0z2pJ/Xc10nJWJqDast1LSzOtgFf4rJPfby8riDj2RtmiwyhFut75CWpGHHKe+tCGBxnUuEkt/GyKJaVbH3fU+Slq80FiR9jcIWQ+ZSYSO2T9YM+gMEbKEUHlJA2Tk+Zc/UzyZsBzZVJFNB3SZwx7oTgPSqDVjScO4fKP1S+oIuRWOshUhT1tFi5J82EUWtQJsXb3v10LH3odPwfMwmcVBrz7ptlvi+s3ceBNt1BRdruu4wHl6dgr8UBn9NVRMW3jwKj95gW5SX2Ln0oESaScrGbSIK5SOv489f8+ICKze9FsGQx7/41avYqb3so4DKQzqP44uk5V1VJYLvAzcNDOMrp7V1vFoe2XohDn5TCsS7DPewpEiN4MvaXi82s8JaLxJqel5iTdZgUndAdYGBuU1/Yhv+QuI/RL3lC3syLnDPBen3j3un3fhzAW2lM0v7OaK32SidSAyKGKts97jL54Hq2DEHOUtviiW8B5oVoJMaiKWrTGdGyjCScioxrto6Klaw3s14gwiudXAiApf85uWsj6mo7Ttz8TQ2B/TzCs0YsU7oJE32Z2s08kop+bckq8e+ExhF8JPnDhkPtN9KuBF2grg6px53+9f+WWdmm2NwxiQtrd0jgWM3WRKOCuuZqiGXEmZ6WDbA8xny4jow2ew9KHnse3oEJ2DNYCVZvPGMIQyp6d9zRqXHUJpTgMKNOs9D8Qd34JlqtAK0vqtG1HXXv6Fs9V9oIoQI/96+e8hR7yMOPLs3ycZ665mr79Osdm+aR8J2Xh/ZJP+fshMo7e304roJAn9S12mKVs2aAaiukgIfqzcYkvCJk0D0FLjAH1TyCcPvZhuO576qwlDbV9Am8QE4moSCvECfjVOfWPCOGXMG12XG193Ulqzv6GVc/vFT6vmDGgHD+V/Hz13yfc4qNPf8rJ/We9PcLVmlDyAbvVLUJ6NtOhPLieEXnsoer8FLYwK4zGBHVez8xBDOgXI/UGHPmf8YcbQcLkMurSg857HW60h/aX5WNiqZn6IZ0DT07iPymflMXuWpqsUt0znaPNW6qx0L3eSnD63ywlOLsUjhBTe7u2H+zFmlRi66HYrjr7s8t/3UROPUZloTRfk8M4w7e6syKqUAc5vbVeUYXEjd9GM2dpH9WPN20Itjfrx3CUoTmqoppJGxdd+AdvEDRTymIuXSIGY0o2xgJx8iglGi8VG3PAU5LBj5nzMSUdXVotvY9fePVBfzCkl2uLm1bYLXJP0ZjiB+uizJMpZylQbTDS8eBlAeqES1gyO3O7b4E1SdK+rqcCt6wExkt3ymBaqeML306YZYIqXMKYTLpZbBPk4+e+xI3JhTbSSRZ4QB/DozQ24eXkIwXrXm8Shd/3H8QszCK+aFkNpCAc2agPhBt2s3TlO9oQE79UJjtHqZ/Op61mVpTOE9snaTr23eGRZ0EMugvun2EvGKLsmAXM1kVeMJbSLcuJybkkfrnx9juPgckLHuHG5IkkwD5SVKkw8AYeXmx7pkiijHnStdTl5U1QcSzBYyH5DdXBdGpgpOrdXufVWCTMV5yKOARTePGa4ocH2+R8hC+kmm4kocYTh6/3IsZDGWS/ElH10HgEPIHlpVOsCQrm5/JtWzXSmZ5R4BbtSJoxN1NmscQ/yz59A1Tr3sXggMVPyT/QPXaThOZ4AWXisrJEbf2Hlp5ByLihOBfw4ufHnnO17dTUSnPH3GX0PdyJVI8I+Pg/s2IEMNVhSRG99k8JSA6+K7Z3Jgsk1iZJCUShJ5wOkcwjIw2Cv2ui3jKRymSMXdZd8vz5dTyqje+FODgsDfiN0KnbxveSNMTgiojs0TaUd9/BElI7aFSsU+QgEWBvGYKO0UMBTrLoDKIiFSfjKNLwW+HjFR/Fl/Jr7zRzmTuMrlPMCxb3qgh1Xy8yycj/0MRvn7+df1betWxmr5ibIUHbmyxKOUCW3/+YWdulr24W5/M3vQxbApEU+AZm5EZ7QwOX9Up6GLnmkmG/cpHW9WYXD4woYCXRwLXoLKR+rHxv5WShoq7JX98omKUmI3ne4nr61nOWxt4A/FMuuN1/hq/Z90baUBv3/kuZAIt+3FdAQHI+UkUqM3DV9udzDWp8924PF9I8C0Gov6a7byCWAWPfmAehgaJTHpbW+HNtww4struiNXh8i2qbpZyFNWEXa7V2t7FpYv2u/PhGx0zeZHg/nh+VaSOptB+BE3O7nKFteEtXu5kZqmRYPyLex/r0nnWrp4SQb7LsgNKHpaeLPYbBvxkx2LnOCkIILubUJzyu0L60iwNTxpKShWrTYJqi6RoOjh7cyYRrYN071UveupfrKCveLRr0pYnaTe6oKv6E9ms9kTnCtILO43ifdLhNcleMsnWc7s3bt9D5sjHr7EA2s2alhSZyrbDCnWBcx+onhssHLggFPaVdfLngpO4nUefrqW21ebdobVpSCKn6SH3IYCM45+vDRYXEsacvKBXS7Ui7ntnI9X3U1Fwou9pXKfKaeGERzOPSJUk4+wC7OGc6WAQ1hgoVVw8uSjwdMxQxxaeRUxJg9+TdBQisrUNUmvh64kIpC9LkUKucaVuMz/PCciroZEOQcMq505FvSdnTCOvqLZ+IfHPJGdUyHtCTD+ecbi4FFjHumo2BZ2BN5e7GBtESvZTb8JNxkoqWAiBl/l9QIufQDpGiShXA2SxFOaiC4U7EuokLpdDquTLO1rIAMAInHq3rhJ2DvoHYPk+WC3lVjl3tM/DrogrwqgNOW7jlAM5RpjcO1hSJzVYrZqkh+AWJ83jywu9Yu9XcvZdpW5p+ykGh6OWhZGKWE8V1+d68yRgDgQoTjvwQ+lIiDaGfrPcEuNNUXtOPXV2WNvDd0Pt8TipBUaMXyNfbYBcRX2/5knJCrSUwuYsUlp7kbIOokygOtiS6x/Psy7YQaAF97hdGGWMMTjY9kKp6z+HjVgIDDR6RG8lHkfIMBF3kDzfIgAEmNiwJ8Aq5/4O439lJAkP0BTXc50R9tdkvZ3UB1Z0E7g1RiffdNneYAY0z8n3iEMvWJZOYulldAM0PyjhkHpeeiqPQo8jn/RQBGni9iLwGSAQD2OCss0tM8LFULNps1VLhfbUHffSVXIWUTOcD8IW+BkwsTyCQLW+1cDm3RB4dQmKDQ9ZqZS6MDbEumruv4WpIlguUB0hlP5pFheC/sqXsFoWR/UM8wJy7rZ4x/C8TG3mg1nVq2u8DxeQiKWrSTxV5CWfkR0H/XSQ2/kc5pYMQLttYmyYOdUzGzb/Gmjg0REn3M2DcA0Qx3bO37nOO55sL12puDT/5Tbp5hlr9pc9XI7NTxgpu8OTRFRDx6Al6ANAkBm4kOcHCF9hGni+zY+MdKBePreQJ8N9Q2bO9AuznGQn+bYPe7afRCpnzXU7kRuyNEXU62Za133J6tMc7tn9h/C0VHlChp8T/7tfGGmlvzCRbsSFqdM0C2Pc8y629JcHjVv1Xj1PoiJtv70Vln0HHStsKbmT4YFjyi6dCCbPV5HumYYECtj+AQlsMop3J6Sry/jTOFZS+kJkdBxvGOZWzRMb14sYHt1Mv/xMheOSRxXN94Ge0CMJsps/2EKL5VwRMXsDxFZGMGCJge0WREHUduox1/H5oqCyBIs+EPjNGfc5c0eIocOHNBl2/4XIWOH6FzNqqMBmuWBPJms90fhfRbs8P+1oswqzxGxzyyRrixKYCwUhvOt31KxZfHEZ6yFb3SIrqzf8MSR5BIu9+2S89mGM8xQBSEr9E0rcqD8aKSGeVY2GnT8IILRWEUnIOXQ/pDyyjQO+lkDezCtdrPGSkMLuQVnrBVelMijiphL99hKOUHvy7zxsfC/tlzSSUTTkL/ZShY08e7wlXngYLwRrjbCrzJV0pCdiXx9MMBwfLtATcrkbIWCY8Jw1fyWn68lNHh5J9pyI6d+84Q5aM/cAKJWx7WKq/nSlH0wuOsWWN/fyXJ/59AVXXoosaOtv2VQUngsEU/LnhtEHzUHk7x5pLIKxKMiUi6R2l6sV+qTdVlJXLHupVz8AKsLACCS/HP3XvCZeD2Zd3WXFMT2kfYsamOAd9nV5yMfDjYRWlXusU0k+1Wt7khTInJ36cCfkQvYnzt0JZhKfSzIx/89IVl32CKPY1pRfjRB5FPMxXAmGTmOpwbxJDWmdIEX/ZEjyBZWgUedBTKchxQQD0vHcSBtJa9aqB4W2aOy6Ugye8qTRlx4xTUARoJZsJ999fVaCE/Yp6ly7Zxwb5VtVBlWCBFzZ+WCkCKuzH3j0nVwGn4kCy5ebIAJX0D+GWMzveNVab5LykbJeT3z6vRKyV3EyV6EbS/3yLNVyvdn+Rm5paFE1sDFOGrzZpHA6J6XZqIbMeO9E5Y3UosI9lD05Z3RJ+hmwSO3amYabRmfBOzyDE7l3p7tZ0N6sUSHFzw4mqL4Sq2r9vsQ+IR4BYkHwRTTwzuHlsIZ9Em45VW8/w2lLJlH/mCU34i1SDZpBEAVs0LrD9jxX+ragg0DD7+bQDOBvJ2WbGXZhljIWnj3pvnnaJc6qK7UTIshe6Ut+EE6c6BNW5shkE+brb/7Jm0y6NFa+cK+G4QNeJgPNjtY+gRZqbdbFzXYYOKnawgfrsyE3x7U2i1cb3oOzT7pTeHBs/Zpv1boBq0oUagPT/uyBU9R5DbeQrGRK6YReJcobIvKWNGfUv+QlE8rV7UoraaZbBgdRd
`pragma protect end_data_block
`pragma protect digest_block
7725e3d8779ee43048a759f90376d33b09e3d8444af0cc80b0d7aa38df4657aa
`pragma protect end_digest_block
`pragma protect end_protected
