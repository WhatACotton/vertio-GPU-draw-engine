`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
m3ro1OYcgXxg6W2b75ijYnOLCiLhUPJ5V27NWBayRK8ohhpLeL8RTbAZiVDZ1FqW/k4n9Du0ZWppyjqPV6/P3slxA+YrGyv25KwPYYIDxbQV5ou8lIoyDwmgSLKdNcfyOE26TvfKhYhN30todXj8PjCGSh7wYwXI0/9VxH0cGmbtxsThHbQBDRvVASiVlr4Ou2fHw1wnQEUc8D2BP82FvJ9u4M/gQsU1P7v0AezsylKWYSEv4X1jEjaymhIz/kxZSZUAp6jXFaFg0jiF4MreJ04UlvlKoW4G/QmGVvC7sGAHM+YX71ySbvDkBU2vB8uzB2OZwQZFPGbnK3C+UKBNQqcbkPknRqN0R3Z8IZnaK0DAOZdafbUXS6xfRfWLCETR0oRdYdkhSgy00b/fVtX8jttSqf911EtYd9ck6NQMOdS/9IgUO9JlxFYEH4PhxmqHNLQwufrWyCtgT99wVDooyuja6SJDfL/YmNlNon8SlfJKXgBCG+JLy+Qwdz79TUJB0LY9lBnUKyc5lSBVIlXfY/47qXK2atsre2BiYZw5ACEuJ45Cbf+KFPinv2a56QZvsnaQ/BCGgb3VwdZ9RAP/FFf/3I2Ew3i9dz+U9kohn3aQjUnYtULc+oiuMHxCn6JSSKxT2fCHfp3atAeWsYseoz7NZjKcC+msZVOTwgA0ybGgyVXaTBMDPOrhqNULMrXpC4Ww/seJrTaxTuxQaS1cOoSObO2JR63jPW0m8ppDlTZ19oYKJYw7OGQFinGlUG+GQyFG7iiN/g3JQo2ld7u+RhJx7LHQv75t9+ADS2/5OwXW7+wNQTcEg6j06MQrbOTaVsVhpYopWA1eqeicpHSyiw6fiMjsT31uB9DDVIji3ANgOCf7TlMWbIM50StToVt89O6q5d3UZOTFm/gArMXYLqjxlH2WxbZI67P6R1gQdA0MzICKeQUPt/o1Isbu80bMH4Mdnh/f462p+sbJ0l/Lv4qSkQ0pFp7ZUK9CbYPiMQ/NdVyKTebg1b9nlwK9R7SjN+z3qgnZQfiQ6ueKbW2J0UCoWRsq/xeBKEch/lyYZp8rFGLdyfe4cWRAzMAmSrj/7EuHq3WIS4NSjoWwgS5Rie6zQocyA6FMklmOTH65EHEMOp4PczttZ+m77YacVsCAa+FjA+W7kgVskBPr3qQ5gITqzQlXRKlWdgVVwQZrwfjkzsOtL36jmAlA3oc2GD06+arfZbNAmx5xrzO4R1rntdO9fbExn2OKyVsxCl38PqCwysQ1Vk8NBkkjAdSQiO5SnoFKoIBYVxVYhlSjyuZ9Pe0PgB9Sa4qAYlNDnlrncjNa0WHwmDKNQGjaJooMNLY3B6c6suj7gQPGWJbibrmlyyO8Wg6gbjDxmlwAijq83PwWCMxSmrCbW8NzpPSGLx8CbxXnx/NIVKWHAGv6ajrpUt8MOnZkSq+MQSIsK+Pp5rXacOd7rZBouLIsOv27sfTsyRa/j3vQIm6/+R+ho7ZM2scBEBPbKiJRsw09BKOTa+mO9BXFCCeuekEO6Li/juQw+aFhrg46jwACpJpFZlpvoNRCulO3Ff9c1I3YfG5m3gpWnQa9MrK2hTx6uzDOx33ZxS0i3NyMNFXg1qd2YV7zX+GkWknnCQA7YUSr3HX3u+hg/E3wT2mmAd4hgdhFFoG8FhAkzUX4hZ08KJ9YzetJlh41+QJ/mLte0fHMjdAmNXgs1cfzk5DrfH3/xM6Fxtgu8ayVh7zFJiId8GtKV2WsQpHGvMSUFndT1x4oBryesYeuZsDcqGdEc62lu5QWvzMxXnDgKPARxD7rmaaRWzebAw==
`pragma protect end_data_block
`pragma protect digest_block
fcabaf23c0c25fb65f02aa7ccffcf3eb8ef54a68f87d1e659bf37a0fbc9c7e3a
`pragma protect end_digest_block
`pragma protect end_protected
