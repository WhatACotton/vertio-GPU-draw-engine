`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
LWROaFY/3q+iZ8oNgvsN2q8mjJatgcJOvn0ZZYyXqVynufrWx82KXsrAHeFKnvPUcm+mLuJ1GKUJHZB8J7vCtR9iX7I6a0PSPkRbkcy3XJbtrzIJip5y5yvURTe7cSxOUNlBNScToEST35BIRBTOtVp0hrQ6fvsy02IGK+3et9hP20mso8LhLX4TvOIINkUKWPIEYFWCwaOu9GyBTtiApvslVBtRg4m2us0GJalKV0vO4SqyidgaH9ZEeiCyEjg4D+P5LwkWRoN8flLmYdWzXKpNMsZ2Nev3a9s0BzPPsMh69tRSQNre7Sb/XQPMZw2jb5cQY/QgohnoJZzLaQMPUFKLfN6HpKHckKD4NViIwUq0PXk0yy42Fg2kzpu8rQWEcYhCKEl3JMKwDrNcjOqEDn2qSaAh7tLR+aj1X9bzCc9HqLN4WsJszcoI7L/3iNCkTTn3wgWOdliUrd/HgQTSac7D6bzruDzUk0kR2sm6xOjv4txDf8+LRgFS2lvp55QctCMY1gXFXp+ql2XpyCNFWJ8c5A/LfESwUzluClvQdTzx1vTlQa2oDQtjrZLDivcQApibrUQWv9QtlEAWRbmo7OYQPIKTKpo633p5ojbFU1nMKbAPtpQqjqbwmXoQIY0X7CuRkKiQtjlZ7+8unT7jL/dBm3dp8Kwwy5fi8EOJpyDonzpJKQWFTGSWllN0rSMxxCb3npbeB26EtFmfnWJsZbB8o6TxPtLE4j5QoLa4G1mkP/n7KEjwKORIQJRI6kTPfXxmgHJwQuws/IgLT9+RHYr7BQwWzv53KSPZJYt/NVwafx6A3W8f7G2+BzIxLqOXWI7W2diUbr7kmWrTjog7pK/J1mbCZsI8jPmIx79LS2VdjevRrrrbdaJpGWuYfXq1/gddthpIoCnpaQGEsyxEwVF57a2hH/ivP8wDOc75hciaohxCCW7Sgdmy1t7h8KeH5O287JlP9W4O5m9e1/Tbo3Xvs1Ko7cL1urCRQH74UTHPA8lRGS7L9Jc4kiNJThqJbkHcXFra0ZsXYOg3tV4xz12dlPy39EHXT3sEGzYqjW0TbpXuIO2LLragDH0mxD7YNXWDNq/KwEwg/QV7hOtXBacgrijfj/pdrZjBHZs3B99xIdmQkw+xLNEb3rwN2MJs8bH31h+ryQdUsYs8QCRGLurAIuBFVNT9BRR9yX2guKEUU7v21TdzzALr4zrDHeWZvznJ8Vsyf0L/q29E2M8LPSSkv+5AWbrvt/UwV5tB1pAFQNvxwIAQ1ObOqWDmyzU5BjV6mi83Qq5h+lp7a/SGAMjClfMXDevq9SdxwvyIsXr/+LkNxxae7gLcy2R7ThgJ8YGiAEDkl8qIBsjbjqag4HnSOJ4Lqyw4P233wklyuivZcGnnXVqJH2eAWBQF2BV5qKvONBFpuU4mqkqeK+Rz82gLeboggl53tPeEw9fd5n7ePVAE8Eb0vEElkmtscxDuVFjDRHBi8RDcUzirb35lJUoummiMUki5ZCy1qzic7y//NkwCzbuX4eF+PjZCOoDja4UxRPIVRhSl7OZ0heoLbY3ZBnQG3/2BAnSs4pSGOYz79UtBuSy4gQbF8HQI8bIYzdslb71YXxHUG89SCMOJKFYxn0vEbVLVnOvdDBVehCaTHnG3r+vP7h+yDtGbkUy+fXK28vCSQ8weYK4SB+Pu1C6wNJJLOXoXKhzzInvjuL/bwh0dI1BZklHV3hcCiC7fSiDVVovb0zvaanf1WCy+7tXIK7jwAZF4mGcu/GHOu07JGOA7YQuaxMq5v7ulDeGe1SJv3cN80+u2AdOAfLP38RrLpU8Iu7Nss3hsJtURJf/D6CYSVn1t4WWdpdCq3kfyuW7kRxy56b0zpgEZGfoa7uTC85VQkZ53TbKVB5zAMhntDA+3K3DQuvGYEpcvd0k583rv8WDiDuD8YQnITH+UgFvgyYbHucFolZQn/8/wTshuFwpO6V8ipwlto/MMkM8J/9PPCodEGJMYfFSam0i/m+DCGG1tM4UuVXDDRziL2mg6E1qm07h53OtRBhAmzm0+fYPRL5XJYlSJOPOEeM28yiobIg/7KsJiASvfjQKCBEbKalNaapu+zfJNdoqMR7z4yAbNDxCMND+Evlpy8c/kLMUBAl9kHEkx59mQGizNJGdqlnJO/u9r3pFLWAKaRrKMXinhhPqRShab1ZjjxGaHfIRjzI6E8bu2ZQBKKjOHrWx/gt2dEyQXGBdgH3lk0nAxXQT4/TUMRtqOKlzrpCNzU1yMPWxj9o2o/9TOiud4UeYmH/bAOHyYNlDDXUD5uNWYMHEY9XvaRaPjpSD6DgeuXvJM5ywataiTsUxUg+VBIWs2S29Hv+L025XWWc3K0ro+IKae22vADh2mk4di61DDYPFJUdKMiAgmyI3ubdonOAnY14UvUYfaBL8MmpYcrVS2H8wJfnGSjOJ4/rD+9dNiD0K0c+9DR80kwwgg2FxWxSWupxhWGt20HlGzSUKbV/+X5KXLbV5d2WzxvY/4kvCvw2vXoSYwtSFDyJVyieSXARB8kIY2x0xvGzrwrOXTszf60DYovCprYbv2JAeup+2r9e5R8/EE0G3dmLU7nimzYj2QjVCHrKpwccKeDPavlhvg2Pp3eUZ5AuIHAmWbdHKLX6ORuU0u3jbxVN+kc1QZMqCNfcEILxP4qBzm+Tq1Y67i6dqKD5NHftoRGr5UjZR8Ic8GLE5jRltlQSUIoZsTKtYPeXmIUrsNpqIw8ZahcsDrRdgJmBqO5brjbnXZqgFZRhLfdbuHXJjutx3p8w47sX544C4gi6T3kTt9ZLGQTczKaH/Q+RzULJNcuyemymtUEKp6DMch4kXKdsilCRi4hHKV0ByH9Fgy10Rz2xSfEkqNqqFk81/bIe6IIAm03QGGFgXGLlhN0WrJ9WHKHsH83KyMKuXm0zAdXqenpYAzQ8YBNpKb3jr9vAT2NZNDeVQPz3WYNC9ZrgkOEzNbIIQ+nipzBr7h66CAJ23BPKM3+URSFawokKA873J3raQwQQbvGsCtGoTo1QSr3YDV97ebIYpKr5OH3PL9A9TTmo+fLmHHijz4sAEoBGkiW+dSqWdJEaxJI8ErwGWmCsb+0TLMhFaEkKFTFfPtaWgQT22eqn2bRHlffMi4OKS665ubTHHSe4ylSwCRMv3e5wVnIGJ5BDU7LFor+kizbp4rzYJKUOO7L+9spVlB34ICNn75UYpMzoX4DulHAzTmk6vIg/4MvBx2trS1CjZb/WkBE0oYVAJRReEfnugqjbKUhPw5JUbZ4cQlANVI9ITUlFmwVFYXPog028CmYSyQts0KyieUNkWgHiB2InoYUWA39Yf2FJo+PGIiiujIrxt3EsA7pVtDB5BLF45STTAdRBcVI5kRabE6PSe3glXVAtd9WmZSnwauFfxTD9WP4GTw7z93Pg4h43J8nSht/q3mKwGGGBQ0ve3aHawVvW5uoz7aUuEdLbQUvsmML6v2tmv5Q0cnqyM3sm445GG2KcwTA+FbsWdQkgUxsIcdGEL8shaMBsXvTjlDk6fzeOi8nkXaKgMJSiJPOOz2XQA5LTypGpnGvB17QOCi8MrAL6eQSnfxMuCvF76inhL3Fr1EMOtNWFKNRdAHPM/EZSsu6syOSUitw/8KdaA8ogtAOmDeB82RtpQ+iNUf/kIVZOQ6w9Uw8v11P9q4WOhFilDdWaKazTyq2JDOQbZixPSxx1dX/qNmst7/H9DjlfWU9Q2hHgxDr2dVBQ5lZqh7EFJwIE5aJN7OD6IzFhG0uVMU2py7b205XMxaBfCejhUhjuYaGg4MzjnmG8TEASmQkzJOAYtu8AWW+rSrPf25LVpuKm47REFPkf7Zyj2o4q7afS2Dyuc3p62OKGXg8LGHVTvO+ojaZRQFZSEpwXl4570y2/SmpigOCvU+TMe1VCAhyoaR4r6HI4mk5CQT2AAyLrnHL2S+xuByfKdqbXPMb/IAZWLjqVk1tnCdOO+pEegTDiCKUKf4s/4SXDQHR389m4xaeDGJaCNquMHEm2AWDGvP8NnTkJ+o1yCIRZmHIjP+9sHBllGcAlNMJBFKm2+D5XaLG9netwl5srnCBMwLy9TzNHHCyCYCLIq22JmIBh+hEpSHMbSwb01Ed3rM4KOSTczqYaXjolPLD93snQrJG1Cn9L2qysAP2PyUc0WwAIzLUqhY1nLPu9hWyg2wkxfRbPNoeL1D0WSBWUCeESfyIzQ9SlY2i+W7d1NIygYs8zfarela4+U6NjY/HvVNm/kYmOZnHsfDwKaA5ZcsO0ybgNo2Hfmo+5sEBsRMszwiZ/VPlSGFHTmrtI4TQr347/+GKj3/vW8jP8IcP4YuYL32iTo4C4Qq51MJs1DoOWpDs3Xx0IMuaEaapFKGLNYhMHnttvbaROtcnXYVt+1RA3VbHFA9rBair789gs+aksxeKDQbkeGInkBTP/2p3x5rEbVKeIyPOiLTAiSe3HPuOr6rzT6nWnDfButyr0SLK8s5bwADRo93WjzlInKSAKWXCxTZgAOyrKjAgaqaj7mVdsN5oDJg4xHsACd6xqP2Ki61Dvn7ObhkJFblOzMdO+MMJIo3wKG/DiAbZ5EEW3Lh6Mp2GNgbcxibA6taTNMdVMLQ1W9C4Xnt+GYM3+naZxYGzlC+FqRBjaQlyX+wGbMsxndVfihwrDyYLVDN+VCUB6BZtmIZv5bPRw/LuBIg9zR8HP2gtbixiZ3Oh5Z14XkFzLi8zH+LfX0lWfcl/zJAX+Le/69Ey7GlCGDOacl38ITWHwL2lxMmvvdmjeJ7P3WkKG9Qb5dUOdLY3G5k1TLzCej3L8LsHBOaZZUrPSJm9Edut2ClSx4rdvIyui3PqRjJxCE1Y8JfX0x3SHjE0KJbi/pOtXq9+SuQWXRE59+m3NFZ63t6rltMcuyYazmBD+1yWRYIOmFwPhDvRmNTk14WQDj+a37fhySBS6czlevsOdEBgCIkjoFt4N1j5Weqht3RVn+hrqMxtNNi2K8iLQ35Ebk8wC2dnwm+Yu1mWyQbAbL4x7sm614tOizFieBzXKc2vOy1CV1K6w1IFiryHo8XYyUWkK6hASoF/I9okUaiEV9uUI2ztSUedWWgVsEL3/kpXI7quvhB9HrA4iRBHCpScnnnOTvT3JUghCgz03OlJ/c1dk5i241XZ1elv6xtz9De+KjrswMJDWhvGRiRaTag02ntw9JUhuz4F8XByHtqOu4fwyjmuVBVLmWw0U2oZKDY95SABAX0lpu0cvys0i2x+Dz2/359hNfJUabPm1VxmeDbsPqocfxJGe1D63R+Bm5e2SxBYpw4ap4otfFoI0adEDxbA1AMMhejI09zdw+3a+ypMCyUBMj5ym8Q4VtEG7xWXLpoWnLhdByKqNqg0ByyUnTVVs1mbIQ5fZx9kTWBrEDZDdtdBVsJoI5ivkzYhGjwrEQY74E5xADOvffkEzA1Oouf4yYsswogD+pe6FmDMEqEoMpPyzzX8j2tJrQ+llQEI98XNkWBck1CmQV+XnStebqBQCMkNkdPZg6e7LEW27bC9hRGnFKSMrXyj/uRuvFozeek0vFb0ay7wtnDCEhDC8Dd0OMsccpxibj4gg9LniAs5LMwkp8qzUQ2MU2YHS2PDjmWeFGkLQQ/1mW1bFxkqBCA6Ke/JRJ3f/RAk42R5Pc2yQA9j4SaxMaeeWkGjxUmQ71PX3W1oqIjwZJA7/FJY4EfXNGGvNSwScriF5VTnPVRI8wgUZDN0nsWOtevnhnpoDGRU5+znCB0Ri/2UEfdo0APhYYuVIgPYQFZc3jv6kBOmgTyUP1TRrVByFTVK+QCIJxwItRlVOLLpPXt8lTx5iXAEyXGUwuS1suY2EwEUmOfuxgFDpivVb+w/xiHwDZV1bOaBMk7Jq2gaeYTL78FPJ5cI8/e9w/9FVmQNXhMQhBat0Z7yCItmRJfnMRuLxuC8n8VVgdJ2c/nWasVNGC5M2GKNx0EyD+vMLESMYe6L6ulV/MvHLnLRjmkDah1PPCYe/7EDaaLh021NWCsShVpcI3g6j45zr6+ks9w/i/YuRa9PfcKAC30FItCGW/Be6h/2TikjPGAIo31xCoyrqZhuSZNYgL1exgXIxGc1xzGXOUG0AT0oP9RSdq11bBw9Pbp6Q7WtGhUfWzlvI1RzV+bEa/VTw3HtTt/auw8fdbuGmtqyy1YkL9T87yb6SHG1Jl+wt208NI9znvBxnCorDbT0nM9wCfJvuPXAy20nLZAgPlBtXvrJcWocUXeYu7+d6CxOLecq+Voe4OvfvbofO4wEr93+M6rVTUuVBP434Bddb2BJJloKevLl6HWuHZuNLFvx3iscVvONHloGBtvOQXrtvNYMoUvPLAsZYIlkSaL3Rb4sv1GSAJZ0+tuuf0guUJUUVYNSi/XUztvRQC0ftL32bS2OOd/lKBXVCHcmu7cnllEVvH7/GiM+phidd/Uqu7BzjwJEj8GMUeY0D8OUzz+Tzxv24SpU57XI7y/wB3sdelwAFuAID1VaIVGL5e2Sd30n6Vg0JSojWIH+LKW8cW+kSWljulVUava28bqg5gMeRiUBD0C7SWo18CEizyQ4FtT3IAD9AZuVX8fF9qjYnvXUeqtgLz4SwhePS2osvrRvPunox9o+UAVjlacWNm3QrrF0XagP0rY2q0eJV20EIcCe+Gz5YvMITYp6lcH9/1JUa87H1Sg+0aXGBYMATdlg88VI2hzuf99dJ0Z/bjvEBnMmOALiJZyoQfcTstbJolwp+ylmlFUexPwFgIUkpXG1h5N+ejJRO1Vuwz6vFCQILp5Cjq6kczGfbkLs+BwLVXDSxcPKIPcTMzQS7o9hhP/Xgzjf6Ijo+fBLegPHVm4iCXNCjfkqscGjwVb+cAv/eYLZD7IaRe5Gp5Fqt9kvq4Tw1tvxEYB1//xK9MXOYj1mIi7gOvyrMnoCHHLY+K1YLMC9x4CYPOhNzI5OTYNjlXc7D5p6fs0aQjgechbFzcrZoBUqN1aJnWWCnMeUXg8Kh5maCJBZa1jC+DzC8RrEZP/oVRuzXtOz/8lY0DVrOkBWiZHHHgMoYhg4Kb1OtOHUKul0GsCV0HBN+I/CA+v8LHHv5BEtg5fAd954a25u3Qy7iOBboMW42xzw87Fb/6fuXdlfbWK+QOQuCJw5tfvz4bSkFLxcOcIXVG4TVZQTP6GjbDY5yvlVOsAMez2MSAZmfCUCf2/uvXDgTmwvCxJQAYlWbc1Iz055XXehBtR2m//4yftEM768UqilAc2fbJPPX3cuREZ20qIb0/FTOZoBkVqRpE9QD9eWu2UMHOFtGOULSXB1xkzwzWhgP1ySdg71y6HzlzZ/RVw7tM33OLZ4iKIPD3lA5gRJwU6Vwr37NscbteycZruUWouOsdMrL9MTVr+95IPo7aEiWaaOkwRCi2W2VE3Lu2Qqfv7ihGWtrqUXPJi1BkWnKVdAgwTSQ0PamkmGJfFLqto6xOEncrOCFGL2+VvtNQNdC37uuhumxMX+MEuRCbXGqcQVz+yPuHnzGE4xJRX0tYjg9T83BHS6tsq1uUrtrGPSnySH4xShqwPHRvDQTJJYJzVPtnIZbUSLcyDylXQetOZQY1qK9QVMaTb8/t2zVqPfuNWzZh5R/XeWk8vMs6YgWrIGjkAW8O7HkYAF7Mke3f17mwue6GL9QAIZ/MtcZn6oTvcz+KQKzeUnPyfIVkr29UqxY+dYnKDwMY6E3Q3o/8Gh402sdBrfU89hnkJlITgJscX+T+Rrk1VcBBOKftHc8x8Y7BIpriPO7CgS/ZxFIXbJ+8/B/ud5q9RrNeO27tupE5jon86pfLhfoXd/FrGDKXDD4vaMk90Fk6mGyiixswXFioP406+hhESFTZV4+lgnapJUcsPh9Uhj9LX2AXNzPOFula0uKuLgGNvt11LuWqlT7uKWEd9XgsCnsYQqXMdYkAm09WmoZ9O6QOTsSnMbeA9lYtCsrHzWZJQcqFr5ohemkRE8bJVz9K9+iHZSbyLfUH4o4eTL4zixqz+dWw0oei6JFw6ktmbaPfyxfAkxHiSqKwNVJ8acRCCKhN90fmC0ZqAtWEIGFr9Z27YRnbrWS4a3gFe9M7GXCZv3DiFfoDD5ulB/B6dMk9LRbll0p1GL50qXEgNKTsAMlY1yCqH+8c5i1R4sPkiMjB/UilzCmFzop9xlMrxXYwj8G9Q0NM710vUIPlYGUKAFlYlM0VHvTWpEeV2bcc2ghMhgDW25+rOzY9ymCkrpvr1hdKbjm8/xzPjmS6sZ718UYuFH27BgBeVyBMs05B4R+NtSmhqpdpxTdfYmi/LfShJW67TVklzKawaj1xVfx3Q8NtJ/Qx6tUcx4Dr8w9LiTEThsiBzKgxW4pzrnbPRMr+3WFFVlXDDMbH/6cMYTUIVEUOixxDpAtPFu2WUiyd/ltQZmpnRrDKHkvp2O2VJKUD1XhdetnoZ897BcRJjo3m3PMUwj3fbcv31C6hVE6iA9O8/43QjSVzjpXBkz1Q4q61OqeKPNGJ1lePuIMGFqah2//0RETXH2DTvc4pl4JGL6v/lLu9VBClnBrc175U8RmuMaT7Bpp+v+kAuH/99rC5xJqOlQUD2vsyW6TlWE8Jd/2FfMVZ2NEI68d9drx106UkML2dlh2CcvLaN973xoFwR1yyWakKCDvIv9Ik64ye1iWAjDGZuIzKEjI6tI/zQ8O1s2SAmF40DEf/2rcKN4o8ii3jvRkMpHUiLC8NR6isWsC0tQv8luTyLj/rf8EvrxvDhz32zD6+GRSrg/HILOyAXyjD492I2Ffx5gOknqYZBSpXQLFdqL9St/7ULVhp+r4s5BwYBpkN6D+GDx+3HJddFHYt+jnOwz4hQrvToxQLNyg65lZdKcNyYqC8MXmJSzsB5rAcrvqHPNkVmAMNTCIZVX/YI4gZsUCkUbB4CFRkiitaJAREDggD1X2LK0yqRhbvcVLx+J1eJpxPx2R82C2pMRzZk7FHFAYP6bb0WP/Rt8nENYsLjXpuGs13/H0vAzZNVLsiQdWZLoNRWANxYm1Ve32v08qQkDJF8EYfVLNv4ctBqG4j9dknRyr2DjsW1CK7nZ4mRtTX72WFRwFEL/vXmHEo1qkYs6oEthp8xv7HaSRX9dVSEaVMltS1y0mxbQaUI1DC22DAuxtATtvdI/3mo/KjgUe8UxxNRiXK7Q3jw7U4chwIOuxoOvQ6Eht717spsIgWfNCrpLEq+rnR6yx6i8oc7v8Jg01K/aG6hWXgP5voi5loZxw2FSjpctlEFUqvo2fmgkJWVMkraHqBZOTKyk15gtQKSgMT4SJHy+8cOkkZI4pEq+1cvnLlDrx+WShcU5UdpWioROTu8znjHlE27AqLZllWd9Jdvl/jaSlwO9kOCUBCc89nxswgrJIJxBku/Kth0sYcijWrwEWStp0HDsEZKL5PDwUlUFCFHdbqNbG+9qalLxZw8czznQJ2go0/8AR1ndt3PxrnvHMmIns4OzokId6cY8ktVOxMrizRAXGxQb/vwh6gY/ESgs/YbBsGDVAx/ilUaPLLbYlepkc/KyEhUHVdBckRyXXdPytfa2Cs/SSpjP5ht65DfK66a00kZULvvjzhTWS4DSGPuQT3kOHzp3ZMIqWUkIT71TYCelK2IiewNk+FpdJGGTGaqbtInprAKMF5LVoxPW93Evo6anCfOfQuE5F+owF6RVQ+pHKU/FjguzCCbHwD6gF9m0XBtLgfdCIrRIJhPhbooG7IPwsKskCqcOeDSI6ZceI4aPGsiAFInAEd6VAmEv1HAN4L/P+HSV9NcwBewEhC2UeMdegq00hjf2KYidlT2Jqe6RipITH3/6US9piFpI8t1uDI2IEWztaaLqQ0XBXuU/7+iQqAJ+FD3qd99VC5cetIN0PovYcSiS4KAepp7HuzherHhQjO4xCcfCeIcWmJWBT9wAWp2Z+Em4e5oMldbXCJdWO6KkfmqNDvJBhiHjIymcntO/DBeJ0tRwMBOe5ChVA7PWTzofokApmTSIp2Hjf+tS2JHz66cb3XiLvuiA5xbMNDWSpr0xTk5Yw55G9n7kGD7Y/7UqotRBqDS5FP32rBGDeYAHzzipsss/ljx9+0j85zrw7vMkbJkbNTXy9cUH8xif9Vxp7QEG6f4lxDICdTHWNNeGdYh6oRA0caBvb+O1alW/bbFT+1Bt5wuJESmuccbq90mAL25DpmoWhe13ne5D2JknOoIugMYtvmyczSvpWvEoeLQu8UrEuyfTFu+YwvvdS1/XReM4wfKSdlkisYxoloSCOX4zuZRdHF7BPjrR55QmQ0eupoggsAj2zSteEICJaIZkoBY5S88xTvaIkT00UTjpqmGE7D8HKu+K5zG162RsbbkmfUhvpSC3nMcmBcDs1VyiiqPxCx8biskxYXE5ts99v9vXlw6XKrkokdaUbTIOZz2C5rdvAj9OXik85qXKoQzBARPucQDzMJ07W7uRrGmGtOLzkP8sEtoIxB0JoukG1agVGZ3azJ92iCDW/1XGJNJ2qoi52COQAcsThKZ6tSDSYPBDPhy8J/2/9n+9J0EgBgBDdL/B78aKhC73DKMW2uGO/8BPJSyz6trFBgNPPxZKwlyqei6IyeEceUX3MLk5NREGmDfwKiBfXsBDYlV9R87zjr5NNqLf8fabShvf3IWUcwjVf3Wl5rRr9lmrZLSG8oBg9aMFIaUikLxxukEWtHcu567S965DcuqYrIJC+SMewOqbTb+L2h2POXdrrmfUgOLmbUm4ymSBD+KTFxrQ8AC7PshhmoVXoGsfu0erQ8ghCBo3B75Rp3omJXi9YUofXdbRIpUUAp5Nabxi3WNYYNE4IWyH8WVIqhEX8NGh6XQV28xwRK0VB7U3A1zJovVAcUUfXXLB6r24gVXIjX2/yVwEpwOc/C0BgOhvMyE3oMhvFUwpicfT1W5VaMniImSB2mgAVXhNeOjYaXD/+zzV+psit+lfp1N5I2Kjbf48Zdhn/N6kSFVBzMXOciKHi02Y7pj179qpPprMC+aA9zb8pqFpWEfcC7n6/s1Xj1hUyATR5l1jHJR4F/LDOdIOlX0c8CuCoFA5DqLXU+p61/3uHTwqfrTwSr/YxFVC+zov/vxf2JsHXXVdVF9Rsmu6Ttc5Be0CMDzRxj2IrImB0159Ydh33vmQDKMPg29FV5Dzda82ZQQ0LXAdh/NIS2uWoRqIFx5lexYfwTXlu6yF5B0huNYz+QwZjim/VRSm7ZhYFlryfqVt7+22wmXcTd2wI830cB+RRfW81pEjwKPxUXJyUO2Y2frqsbeG9Alz0cWRZ9msyL8Ds5iSrKSaqnDf4nBOqpHx8hlzQaIyGXn6lKBrQ82LfBh7zm+zzuNY1aPj1n7Vs8Qt3GPpzEEfpD1CPCyg5L456QyCYsG86NjNOi4J8rqiP8pvOlN+j2yNSlqB9Xa/1tCtQAwW1koTOxYEFD6kaU0FnxRBE1wkofnxTJMCgGyADbzCrB5ITKaE3kaEGLm0yp/qK50W8t4Q1Q8/RUoZZWh1GIfe3gW6lmTWy0niPI0JHvAcFfDqS/4WFGCHGscKm3S7f6fUqHg31hJn3ynnpcpqUxpM7L0GIqTDZpSNGFms8g9fW51n1PnnVNFOM1nSsnLBLSW74FudhbSS5dIKZURtmzLJW04nTZbuARkAfouKryNgRBE4+X4utDe0kIvRRnnqZ61F1Z6J7D92q2zDZwRDvKhSanP43BU7HFeBt5/VI9khFBii02KX2Tc4HHp7LM5Qd0Zk51SZYk0z1wNZ7NxJpLzhZAKZs6u/EFc22qeEYcatQ7TQFeglct+l3NKlhDBZfkmVDmjB+GP0QvltlyKd04VJejLbhKMOOzyDkfHqP1AQGzeEmQ/kmlzNAqTt3fMyvqj9lebAM/DfP07KOi0Z0BodVCc7QWZTyXO73rG8c5Wa9CkQ1U0j64F+MqqVvHkHqsP2kxzw4Ui/b4XmqSAAu3OgUc4DJGQYAq0bFurj9zyCjlhMmqlTTXKHY2MZi35AGH8FPWo0xQTyh/Qufbo0s/KD1WT4qkMTvXyma5xkcgroo8NM04yYWHJG30VSqvYuC6PUSHprH/O89gr4YLbYknp8yyhftI92GXSTKBufKOkSrK7Xl3imYLvVnrJK5gpscjRxTGnR31NRNq1hUYgLxYzA2kiGFVmT8I+HdI0k6ogKgin/qRszXppAm2aOmY5Rr45J6xdv4o1hzSRQxWz5nwLuJmZZKW808pO1ghRtUNmAaO5zgAiuBP5duLW/p0glGr8oRHQ9wZSB3lb97i57DLsU0FytI3BYQZNUe2e1nt/reOGjQfUmwytoSnKx2Xu2NcXmNdNLRDV7WglnLvUC+p2MO6Nwulew4HQ/mkc0TXXFeFddhgEzEPT0IXGyuVgse5fmgTaRqIPtFHv/NlkfsxFxul99PG47ldosUiPXfGBrdAzS70/kJN7MlMXaXvKuF7ctOmhsUUp7Il6vphWg23IocU3gO2H0hqxyQC9NEc8QrQHzI2MsfeeUHXW80NiXecNRAYivgG57jcQsLANgm/yQjJmy3W7FscmaE1g5n1ldmAHF4s7LR7Jjt2Fsu3BmFktYzovdsC60hYsPPox1LkYNeL/uJq2eUYcc76tqpgwWoEMzmHk4IBEnmVsNb1itsw2r+1JC4LXgTkSD0t4sMgA5NaSnjRoW22nDsyHRb0ZjWk74e40zvDlyRYf+XGWDNVDvuSDNaoP1ok0ziXAxjxPMpFWWEfUlEAr71Kdxu738xDoWSfy9cuktIecDxSeMCkWkS5oCv3y1JZAXKvGT3JmUMbvcysdGOw0qNU2Ft2eUU5/Xd2xc1fIRZSNVPZoZXyOt3pzNK6SgKjrD0llDB54v2anmH14/K0eRXsoe5RpWR0zkxMoM0sPSg0A3KtP2NZ2JHzHgT6ya95uE4ZPfWb2XlPfomt9FNlrTOwQSpQOFyAtT0DN7ZcWj85KWg/7cGI+Iz9cyLGPR9G25yyyZzgAIOocn6PV85RQoN4zguOUclK4xhUHxQ+eI17GTkO3OPSA30yk8ejHNbgv72jWR9OHAmfQIHJpCIdrO51PjOzXMXMNp9Xpcb67BR9kOZ5098BsQBZN8uHyCrJniNGhdzTASazi9heZTjkFXAowOhyPerv8vP15uqE1t2V0aPQP69CWE9Mz8aDbd37DkyDtk2IukWXR/38qDRtsJ/iLgu+wzC9fymUuYED1cAS/Qu80IG/vayRKIrt+WR/sGsVDPPHEnqACv3epCHIrxTquPC9CHo7NuwIf5cbqY1QQ2ESVqcsb17AnromHaVbV3Da3dKL6Vu7XpjJstjR2Y7/LBLmtYYb2qq7d/7BKkKVHtt+mWFyskPHGMLkbyROf1V0cMHVmGaekWeGzytCh1GzshA5mWwrOcSxbTCyK6FHz640wlpFFeoS6GCBzm2WzADFPHPmQFNwlbPBZrvZZQaH8g/etzlib7INEGYuJuqVJkvgwnQ5HkK1oIVlZHR+fWbat1uszoaUyhSbOjC1VAE1y43d9/IeYpbKgf4OAbsb1CHmGphrGSk1NU0hO/IaQU/1H+UAADIV5xQ32VdqSUlu+hZYtHtIh1/w9boUxwFXmPNwCYoKm3FD3V5MTAsg+rrH8Rn/zKu/M6zCobs+LWyjBaelq4Ys4O0DYayqRrHbeng3azTv+frY4RXg2OcJ8F17pwi+0pwctqxsBEtjQA9BG6fw7/PQTaMqpiRbEq3VhOafkf8lOlOwOxyP87FkIKqmEJDqmyia/+qhBMmKIfkgP6/KlPndzkaSvXzXjlV+2NZn/cX6ztnQJqTMCKAfaBlxL53zvHowt/vdySiO+SsanZhcugwVBrLMYKPB7dMfbysr1ByKDiwu6zB/CMFyiPLTbsTKUFJtfKrf7BHPqX25+DNsUuYY2XPj0cluw/EQr20l7HKl/Dpd4KAbojIHckw3hImUfKzNWvgY19H/y5w/DLO5wPfj5nr1SXxuCLuaRkC29x4junYMMoSAR9Y0h65z83fQwkhaqcmYNgBSEz8HO92FG3nojrwW5yXOs7h17h9RLBMBenP8xEMULhSN9uJ9KgWXVKJ0Pw9U9pew2y/fQmCdzwbFqLpQO3jxAqKObLa1sf4BfPwbw1EFyfwQY5fCx/oFoGgshwUYs1T/dfw38XcL9fSEcR+2E4NvptKR9GMD9f01ZJXBP+mtlucxM3Zk741C/ysMQdw7efdAkUie3+d3mXgmt1ZVrZ2aG1j11Pr91F+s+JxiOjSRktoiPP3hXrzvUNCpvvnsIfDYKXrgKxdBqor9+xo41R1yUgjRHct1vIgHDG8NY6mR9ELd+zwsox2DjDMAnuP77x2z4I7rTv3g8XUyzdXaroC78EJCi5uPx3uZYtO5g6SofA9lIJ26C+ZYq4OgBDd36812hOGtIpGOR7RvoSXdt25yfkGY9J6ocQQ46IEq1on+PTZUPyPcMLgUZ2blkV4QBh15/XzvDSCaCXqbb0v0YeXjPKulUo2E6cQ3y2050b/BbjtX+GVlz6Ibodmq229nSabV6YtpCdPDNNIa2cI6k68rFqU8XWhOnQoHOcIOFBLSG+wU1ceLOjX0Ig0I/OSTbKdA071O3iYvJb/m2MzRz40afBxQoDC5msGjVFmD/V0sM7AMR/fRYCR3QAIeFkJ79R5XYravjntOcjBxu8I5HylSJtcPaUVNytynXSfF6gi5dLkz/+kbUr7Ya/a0WhiFK/Yn4uf4MmhnG/xY34yKMbfcMP3td6/g+2YEuBR9nljg1h72daA340+NtNeQnQR/65GwM+JGHb2PVSyURykb2x9Du9Oqms892gmcOmiiU1FcgzuzFV1WY33g4+uikxNgWZsRvnESTs6+zXMkPikHUd7xmPEAU7Gt688gjRYTdsxWcxqMyUi0m0zBJpy7l6jAQKaGM2GH6R4RiyB6Zaxkw516NjsK1IFiHjJ3343G2HbAN2Fwd1xqbNePxgoi/+nIkl7Jchqb2Y0W6mZYYZqkTNM6lVccwDBjNdsWMFE0E6eR19AelgwEn7a+1XQgh7tY7/TVMYhlrSWy82sZnL0kdD+aLCE8LgMvBKPekY8+xcLBVugApCOrNjLbisUIPooZ8m5p7UY+1dVsqL7orM9/yyiIQo+CQIZnK2aaXa75GNSfDRoZNgMVQX2kYEhlQQYOKTS2UTmbadxM0oxYEBXZKmPv9bafKprVxSvjo7/mzlXZKKe6v1dRPcZXsZnfrGFoMGxwwz0KQ/lgyu2zrqDLYUhRQh0i5AxfW5N6UI8EgPm0RzauZmEG9eNd6rRZf3OtMGxe1tbi8K3vTcCyUQMKHA5A2zuGCf6x7PZMhUVlChQI4WRBET/ZANAcr1o4mEecLhs7GntBkgKxNtMUauyvNvearroFjwN73Pek2Xcnh9xahYBi1s51jnP7L0q8JgKi7fp8siSSpwuhafsKmPqrfpgee0z4i7sMdU1xFN+R1QcljQ4zYCBPMjnZ9sIuxBl0LeDtfRHkc987EEk4O5/pGxJ4sBx1MdFYg1NN+GTuYQ7cIYs0si1ogWhCKx9daPkO+Y3yZu3uU3ciazIogOxJI4gRoseBOyr9Ldpn2NgIJzpDS4ReyMY4YWluFHPFNz7bdjNRI3rcLfGyjg0ljn8fabS8c5XBkTSkB5rMZdkJ9rm9uoN8zR8pxb2mqcUNV2n8L+vnsCMJWjWJ4UanBlQdAZX8O3iQ/EucWQVT/YMF8q4lB/dc5U8PSLE4eHoeo3AEvOAgXDz7F7S7v0MSRG15IKAYVqca3eVAieho5enogszrMOXstOPjLqjxR07Nblv1ybe8tB/7t5eFRQuB7VvgVRW7P4JXlshVPQQJKCLPIamAN4Vtidcw4I1HxV+QsR4uYWPYxqd+KQeTn09fQk5WtKKEywkA7i7z33Hs=
`pragma protect end_data_block
`pragma protect digest_block
827a0e92c76f5d211a45481966a558f8fa3c11d0af390cfa6fbb5160aa65e3da
`pragma protect end_digest_block
`pragma protect end_protected
