`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
Uth/vvpfYIsSw7WbLgkbSRdhDeYa60e3AXIfc/5u5CuqrmL6X2CJ7vmL2vFEhhfZKBEJdg+6JTr1358PhpBDufIM70Kr4TE1cjREdEL6OV7RBTPKL2GOmrtT39mUukzzUa4TtYp80aUBhELrdv9BnToiN8iujO1b5qRnt01qdowXHKJRLu8Z4rbxFeEaCj/4aPUAXEhqv3pV1hPMqQchjWRlulro+YIzzUf8mkjWHyMcShKCkp89Yx9dNQLn5ZbW0svtNGxFzzCKGBlybKEV+JWk2j0lALZmaEiIEfxAO8M1c5nlzB+MKMoqn6bm3CgjQoZ/CpUG260JHIRntIjFzbvsQdYDGcuacVG7UxcJvZ3nm47s7Cy/S/zsWArbxr2bbfe8ibDLTPpSfeRDYd865wJUQKjr/PitSA+2wITf3Adrr1PP1r92xNAI/iHyqL4PG363mqBAmLj+znMvjSUHTN2BdsLpwgJwR/W7URizLYZJvf4ZO4o2Lg8Ar5KanoHPNmAbnDit0ixJ1h42ZCPRx/FbjIfZ123pTFC4HHGXZ5RH3wpzHY+QPYEah8N9mtcYELY+UZI2BDuByW4r7I43ygCnfdBpiMiwWekOaRjLxCTVxTeNY9TPn39SKkNZLOhytrYer3Ak3Ui4pt+mBCYQNci4qJBYAVYdYyIhBQc+5zh7EV1M/eTcRYJ8e/wVH4MES4N4HKFNA2MI1SywHIXE8kzcB+bC2ni15l0gzmqUZLvXwVkFxHOe4BVsC3rE+I8a+UWUxUteougu8SwCiYhDVddzKDzoJvIZnHk9aokHBytSB7javoXpzbpA9sdr93cGnNuI2ZF0uV3eJyToYILROh/rNN6EcMZR+oqGSCfyXuigbcrdOWb3xaURyDz2RmOGVV4Hwt/nz1ekBAEsVlIB76BYn7pgR9HN+gXVhTtX7tVc1uj+QZcQuFf57RXZDWYZEiMbEWdaFDf3Qb1cP7DJhvIcjz/YdSrv2nPvL+yP9StCusnVou4DKXOaHfsy2FircrHMFydz9lDGRIQp6Xs5iQbs3n3ZNAWqngC1JL/NtqcS135x0kh9Jjzo3FSOQBIzg2fjh50CJFwQn1I0mGCA2h10deE1jAPyx2BiIupEgCzzeh+jW8LRMTj/XkCA9NUFeX5nnaKvfSxejJjVMtKBo3ZMMEnCrdl1B3F+NUqkRJ3njgJHPT2xOZeWwSqmcDRCU0GWcUKF4xZVNuGUEEcsUzbv8MApR0o0QmJ0uN8I4fhiFFh8eJ9z4Ym59rovHDsemSlFxg8yuS4uehNJE3IZUC2dG0HxPfeyNd8NHmikN8WpIZIqOrnb2Fqqw9uGnm2jTdneNmFGs+KRyekKgQ8wLSIGtXL74f9hBrgpUhLDxwGC8TPbdKu11zp9wyo+Aw46jKGNzG7xhVapm/moRooXYdT7P8xOcCtYcaj0yN8HvmgF9UQ6jsxYKsMu4wFErmuRpzSggIqNb416/fMiUI1+GlESmK9rcU7Prtgr7lIsykgiLryeWOiqVtzFT20fzKD/qPzhJ/+BzcHbBkNAC4d3pHPTIPdBso2dgDjyDBV9rd3Tg10KXWOU4d6MakhI/GFLtJRyF2brprHqQt3U9YEROKoeCkSNeNphJf9yqYWYfXF+Wur5ouNDx2W7K4pHbPOFKzvAHR4xynXI39zdXs54Iz7ugxxKedlIXQ/kleADMMxC0xLLjZh9RbwuK+2L+Ddsxh5Lu8Ez7XPLeG1krWJoqunBBSt51MT32DiQVJlT8QBucKSlqPK1vLhg5wcWdCPzwRnVbMSYGpbL+3ZBRKAQSZqwXTveM+dOdxxZdwQsA4hg3pxLDcR1MecfHUJX0+zTF6CRRxd7MNroOFL5Uimgutwi6Pr8ddkc5VYBzaiLQ0VvEpSnAY51UQM5m4+CmQja1jvYsrh19oFLqLRHzCd84jO7mAF7t6/8iYXJCD+Y7185fU+7xpImPxJF+Fwi41JMsfN5Z0f7rg8sHmzGml9XxZyPgdZZh1UH69Kp3ixx3Oet20AVo4Ot0KYXuMPquBS+pDchRUvI6lORFll9fDbg6HBKz4mAhQV+K+ikcemwCco0qtKLpxTXiPBwD3v+YMjVSTA1SfQ3S32XD5uxAywUII69HcExRMQMufUD9zZNkYBdkGbTDF+TGlNXticMDt4Qd6wADvpALRTNH39DvTKFZ0f3xFybxjypYfgpa9QRKvafcdVmQbmczxQT1gDDMDlIVpaLEhm6xBfQs0GB635Em+H0mOKruHQaOmz8GtK40U4SdgwOiOTVF6+BA09afIm2Q4/Ao65z4P+bXS3vk0ZrnLmBg8tC1mynjxH4iUT3NqvJeJ7HE5Cx0OM4u8bwpf/16VGekG/XgskottN1w03ax10JaWUosGs77rDSxfjX5KMbkpS5YwiNA/TFeLFFY8C1J7BsL0LXJrax3jqNeoEHrBjWz1cOaCvLCF11IKv5CM5SD0y0zQqiaf8lYiP4YWYz6GS76KfcMhpFKzVXQKAkBbn3yZVTZY9VHnhqWpUiAsOiDzJEosW8N5BjI6P0setJpgDjUGZH5Ra5EcVSjr76dfrxYHBmm+A9s92DS4ZhLhGQtsFTaVtqXFmw1rCAiSH1AwrikC4CIXnP7c092RJv/4+3R8GQiCVL8qWjDUqG1ZtWj7x36+UBVbWJcdWo10jt8ocRPcBXboE0xQP8de+njfWvlgwR6KKzVRkkdbVGpU0urkn+TRlFFR2zzjq++1ZbYr9qjaTNq3p4cUscXevzT1ibe0C+hyTERpeX+9Yu4j7cLBOnl7sAakW5kVdN2CERfx1qcIl+P1/9eiWjNGaqAaZz/xxLd1k4jnbMosB/Y+s9G3bxRCILBkNjidmoYE7LqUzLaPLadRyrnulX3pVBT8zuDraalm+3qm3B1hiwbEjRmcocE4T41WoWppuNStPnC2eVT+3TbwpNM2q/HF9hRg2i3TKKJitcPM2Q6JF6nkrqP23zGmMlbGDlHI9mYXr3ki2C8zDoAG9ZFRYDjJhLGO//NMP+fonF50UKmUxsvjPlVRfI3LQQzRhHfHjv3eznCl7scMJ/l2SuiuwhGRkcP3NzL7DFsSq63bbmCUMvherUOAc1s1JGOSh3AuwMfMd1BYamv9A4tVPPau4qFoWsWeIJoXiN64saZQUrm4iezLdipws6EubjMew/wQ+Y0mRka3y5Hv5/z+Ubd6MVs0g/O1+G6EmP6zJeZcHtsXP0QwyQJMP1+gm84uR9T1PGKw0j3KV4h24QyWbgOHfCyOBs/0/yMTPZxXL6vxknqmmbN9dc9LWa/Z1BCbg6qtCprDRaZPLJadz7C6YtS4tciDNtWPuFM3JcJPOvuHqm4ON0tcpULGYn2M2L3D/ZCzR2N1b6ICX94BnJnf70wsXL5W4NtB7W8KRCQZNh8FKLrfQZctbboSnebWzDesqnF8j2l+jDMaVrzQUBL7ca1w//BqTAdVfkqoMrtCD+NptAgo7QWBI/d/qYtRQA+Blin6LrPKTp1GGfPswyQ12tgwXTdLSC89sYYQhOqvWe2zXORBbywCFi15JypWAsoE+1L03wrvNJWUaCjzytzoIRIzhth1m2OfR3oBOsQdDyh8oPbDX0id0oQZqW0ugLfg4CWOOTd/yj4uQagLOwFquL8QHLZ4wEcN/e/5aLUoUrOltcne7tVc5HhA9A/S28NLGuFaOgDg1uvaj1aLNuwN7XjJUdsJ5SysNniVt0tKB6lFu+U+V5XzFaHBKzvUViwKG/pF9rMLr89m/hjo642TCLN4uq98LmumWoeHixxZnfnRjpjtR8crGMKMXJkyXY3uNseFqM54RHlzpnuMtcBnxE1NMv3cnQa8Cr5dPKoVCPl5UXTRtK6cuSH4du6JyRVRVA9U5uTHsGVRLprIKedJwqUb7Dc/atJ4U8b4qdr1sK9svi+gIFcrw/k/mahLBr545P8wsWt7Gf0yjTZMnLPohecR6a7kmyzDgaiHVyuvrpI+VMuXmhMo0Q20D3hIoGCIs292RU6Q8+j0632OzMz3dTckeXwWCvRAB7u3hmL+t2tHhXqPvxV9zvOiurF3HNaEkYtj+hmy1hgJ79gKS64HexqN1vvYP2KEe27udQLJjXjVhAdhoxoKy3VvJk8ENmJ/+A6f92VJfP+btjvF1mRbSSoDmJMZB0Wd0MY2V8l1n4G9xzM1TBP098xDJ6lEzwdZrtkxDe6iC1/FxHYAaDfH1lbVFhvi4qQ2Y9dqK/7HWx4dsjdOWffi5DPA4XAV6zmxOREeLfDQ+v2ce8R8pfVkM8IF40WtYV+sNJ9VpCEJroqGRoTaHRmkfxsqAxft4livUmb1TNJsJSE9s6iucFh9vjkypNIAOqoUFk23dn+VgM+u2elNEOUSEFuFaKRaNMQA44uu2IFzSpnhXRIkaNvpVHQiCzdShizCipH4+ZDdS2yBiT8j82cZlcZTwSZRe/9T6x9pma71wq5XilYVhf8HKvScTKzrp3nY/KQUD5vrb+lnFWsBRZs7TnvsFRJxyh4vmAt2xrec8uucyNUw/nOwm21mNidSwO5coXLp+bvuUoKyjrA18RFjDj3v/gE9m45AhCOzY0YgwlwaRBBPeH6wPbgRAPIrbC4Tsr26BrOcGEDEhp1nhI7rR7VqkYhdNow2ZB7qSZ6gongRWqQk4YceFVODQjZUtqJ5qvosSVV4f+PUOPpSXPpBKUHQzGQqz5no5lHNVQCTeuzHJPjqSFN0jf7QrkHx0l30Xv+fkuHfFkxTOyARBpisDHUU4Z7rQDYWdoTb7AuunAzO4ZbIVmoYg7CVO+a2F2vUpJw0HoUh2ncTJG+sae6TCWQkHjEnkg5RerW0VKw4k60kuoOqy/vzTsFmF027ZP5k+LbNd9FqPSc+wcP2S5Y3ZxvY3Rv7/EVtAoeXl7QhLx1IFp/yJOzhDBdoT58x7ADoPyzaUBf1HlmQUstob6tjKfnfaR/nJ5NnkfYHGO/TDx3i4OdasmKTwklta91TmrMLNXqRvRx45UgigcPtijF4ATzhxT8PAffjbL5JxJ8Oh9mrPt9oYYejSiDuhNEAT6HIWOF/84eUVsCnqa3xw72kO8zquNWnvuD1uAKZgLPzCX9owqdQE7Wtgu3xMIX/AcFVbStGJg85OYZwPdDHicZTikrPoxprpSIb9bR7tdYygMFaqfTjprVN+a13V8M4e1OxylMxBc6k4kD1Wf4apSkSMQPKsxYc6Rg8joX2uLQ7I2PUP/st7QJe7lrUR0GhGsLErNBkfPe7ipzk1ICfXepySzxI3uRi2LM+V6UUOip/Px+n9FgIbsh5XEL16O+WLfEwUWEijY8kxHMGuAu4HSYT/Z2lsYqrPLHDwKH/gcOOvzaGvHQGUSHF4mbCbAcdFTQ4TAXoYyvBew+JpD6uULI2XCIGMeKaF1djQfwE/+QbtzUUKMQEHFSITZWweyzMWaQzcXDFTUCmrJ4v4ixv0mhJNk5s/jYLA2ykq9uyG5/WIDyFLIX2iCu0KsQWgdILsBVM+GVT8/ZDC608A66pWa4ILSOceXrtiH5w7DBVZgKChgTweRDx39vKJErNV/uior15GWquPwieviRlJ2CmEnJvtO4wVa5GJYhq/xb+atB4T0gg1Af9Zm5Qc71bh4mRm4wsswbacW36Dehzv1D4xg+qjmFjCoqhLGUxYUWVY23OT1dQ2ePRjVGb7uNb6nRscaXL+468D+UqRz0UtR6oOUClcv6RABjAZ71Z2kl3qmce99/YjtibRXc/PJvcf9SUoGHd+fXchwjJESFiQZNPB1D30G5ds7PPgA7VShkArONtdA2fGgmNRceDy2SiwIFiscQjTAwhwi0zKj7NAuzgOW+DyUzPVOy3qeRf4YP3CSqQwjxtrhqp1tbvhAQ/KRE8rSMXfEhnKRYCEyEU//INgL2tkXFjxY8qIESB3wWIiPmZzEO+RYWzqeMSGbLpqgTp6dGa31q/yiatsy2w/xZ9dErgl6Hvz2b+ho+C+PmNA10F7gfJkw6ckt86hvVm50PCOgKwNGIDYDgSR+z+TZGKZyRRjDIDhNqh/wxAJNVT1RxbpKjQCXfpRBOQo4E9ikpQE+2Zx3PIPxEMemhppwJw231hNTi1pg96XAIXHaVjF2EOzgMEMOhtE4h4jovpoORUcsTW9ZjE7QlPZDEuxFvgBKxQ0tnmWxHq3r7JUIaRuzTiyJZoOXWYhV/c2kOouNNbCR5bb9641m3Tx9n7mDAxyTjd1OX3w4taPOleEaCG+WTp4993uwaVRpCnQWn6RK5phJWMHUjEb9z8OduZUPQjmnRcfc9Esfv/5If1Zm2ZgeEF1Glich9MmGpwIgx3ESKbF7dB0hPq3zjlXFVxrTT7J4lh9G3tD/9+QxGGLRzfCsZfjuxeg1MWhKROCEYwT85gdppHvOATcstoxdkdySDNVTh5OvMMFn1DHGDh4N1BnimhC6LpLmC8r+wN2TY5iS96aH5SaOIX55O2jQWWTKIGDmKKuuLzrdJhXiauSpQDQmfasXeyoOSlJJU6fXoxFhl0vsMiGMJrWYhVk2ZpM0fE44WAT/o7WihO0IWMQy19FBQASDTV6eByMY+MFuaR7LXHF/zT1FdhltwUvaHGCNWX6Bu5zh08h19lh+E9uB73D5Iexle6D75XSFi4F1i5GyS+My94rjKEXVbOd3TLxOGVeyN31R6T5fxkmktNPsYeIE/lZElQ1yPPEaMNl9+fVjOU1XBBGR9yy4pKepdcz6kGVb8k4PJQ1oMPxvvdYARLrrEvgCd+cpAj312VvHISUOVmSEnG1m0HJvEcbdUskmzw/jnPSh4YDEQ+OjgTW0/2Fg35wDpBymE/9DMEC5yXOvsPqO9CmVm0/3vJ+vESUgedvPAVk+PcD5xS17D4xP/ZGYyKVPdbxmXYenmqkXLi8zGnY090YVGNUCaPR8UKD12CR5KJ1q+gzDDVaBCMGFMrtNH21bCe1OTi/RmMBmgWp81PHve1k7cXoZHMNywox7CU78gH+nZl27/tX2C+hi7xTLUWNfpYmgD8B7f+24cODl7+9oXJ28uGmoDoruwF5T3SiOp99QowX1K0zZxERhCTbJPYaLrGA1ARIZdkMP+SNG4eYgzZDMit5ZlwlscwPl4a6lzHQ+8r8FYBZxd9BseYUwscO92T3NYKeUOma41fJo++QBk+FjZYcRtm9iaqgTS7Tu2kYmE5Nz03vY5sFu5+p3N3rnd/Ow5CNnY7RmhMBPg+oNZZAjPzjGCF+ZaAQSSPtEHPqbCQKiTvc0x2V+VcqHAJFVPAdD4jE1CA4JCBC2S/GYRPwr4p3Ixdu1pP31rRdIHDCMI5gHsFI/HBKRBdyTp/15/8whjzTb1S4g0lcsurSmb+AJbGi/fPsrlQkdMNAlimgyDKeSIAO1HCQVz6SEP2aQxM9UDi76/uQb8YggnrV8tiSY5ci4/E772Jfx3OY7Mu9B0TUOeo7Klx8cPMwkNnxqSekglVDeK1KzHI/W2UgYBjlHHCGDwx13jzYjz4l1B+Z3f/I/qosIzHMuy3+HMr1uojuHmfIvLaKu1+0BJGJJP7IGgeNWsulonlwz3PWrN/u4Uc8iMBhej3N4fT/R+FEDC3zDZWEw2gD44onaWHyNIZnbaOk6OnTc4c7DsUUUWHFvyA6p1EISs/wmekkUx+zqupmG0welLV39vjk2rYaH8zhQljr7JLPM1MlVJleTf71MTGJZVQexou3SKOIaO7rXRecDlxfL2BbtxmyO5CwDzDA97JVchGeYurm7QEw6nJ4XVCZBx+Cpwo6CFYk7Uw4xPd/tCoUVXlEbLQgy9PyXhphSV2iRLB87kUALW2DL2x79Bzn6di0x0qDszN6zIdk+DEztT/qPg3D+rqmLmKYF8mdk/do2mJiPFD3IowlYtKs0wtAbVWdUW0S6r7uWsz+PsTnqrsboigznSqoSXtdEgnA4KjyMBeb842q5kwZ80w/p9czuYo8xwl0jUjn4QEhMbMHcKd0e6gbVt+tDjuQIRvWNfSTDsikCtux9WVc8Blsl0UFnmxkGTteVUaJJtYyv9XBsbzBlfBDR/Jynr9EM+zJpkS3F+vJTHbPwhVwhJ2XM+4PMpRLs68VRjfoftgW7sJGCAkbMfmeC3KvcApbLzxwJfCTbfOLBCRPTqf76dJUgqiUiwJmOwTHbdr8MhlgagIZmyd+w5yieEUeBibnxVeKw4wsQxshAOUXWGcXjs96yZ7JJI25ZJccwGjLy2PqCAmMmh0f3MJeuBWSvfuEA3n2LtrWy1V9UcHIqWLfSovnthQY5bcF1uxajs8Byh62VVq3q9v7o+guXUJCzgpvsaZCC3gGvzclP/v735S7wGo9IYQkXQuerw/Gbpwo5QzW2PlldBde9WBRxfjKKMp/FaAFb2MR3SoBkf2UnlHMVFZCz0h3G1tJ5fALYS6fh6cbhioMrOKWsFBNFfipxxUmKsPWU0CmJbyjW+IZz35EdMmRkwmlSXL6I0bE8j9a7J4d5sX7Ry4v8fT5XVSe73xnnumvJ5CuBuRUfk6kUxPMFR0JZqGWKnrJshA8HWaAulEAs246AwfgjArINzSj26rNisxDHEnt13IjRSTEd8b+FDnA9iQuG0yIoYSfLrE5zCNOeP+AkmPf39PKylF5p/Rdv14AwnkfIa5jNDMsLe4VPEOUy0diOBKN2hdux0RafhGCy4t/kD2Cejiln+RQoCQ9BalIWqRgJ7QjsnOcFzAluBB4J/z5bXTLKRxQkVL4ozNiRldIHAxUY6UdXFByvalaeaztwijkXlF3W8fNcNKPARZAO+GDlQpEE27vMToT3YDLxuX5LD7oE4WA0xuqjauX7rF4q+DzcNLCtMlUvOnMtZMNmL3mXRCHsYEINFr00mT9p2q1uwJMeAHkpohkoHSxb2NOFACGIXWQXXc0GRsMC5ZerLjxqD7avqfiCnyADgfQjbVF5d95d5wCkUrNVHeN6MrXmLPm5TqOWm2m3NgxW0+MWpf5x3zDxNsi7T8A5+5dE8mD/Yql4zp2YZgW03Swadgurd1qJEBYQk6cpCHPoDiQUcn80FpiAQA65Z47eCmhYSJrin7ZN76kBBqz3pN9u3ij2NdVUa8dcMrG3s6rYtTJ7G21/s8NMQVrLjI71gz890jKxmxp3cvX1XGBnxuzfKZda0648rZ2cmUBh3ibwz7u9iEizAbSCuCMztO/I2wxXqP4Y9SHxVgZzjhsd36w96nIx/MY5QDQnxXnuZQGfozr2E8j3i7jw/dOUaMLHPaN1LkTbDqslsIN7kP4CEHnHi+YBCNf4U/SidG9+r+iRkP+hSlHHYlg2KFxBzv/1CNhC3wpsxUBPE0SikHmPqRkC+p5RU8S+vTM2LNTJUD86ycy9ofszvcXCnplNGUHhFXOh3iV4AREAZqkXi5JySAAGYrlYDt+NT3NH04OKiMknrUW8kWZ2JiKh1x9KlVKNDIheIXm/tjwkUtf4Ue9wePw8xXhWMXXJ3e3ut7EcsgG3cfPpqL+KqxlNliucj4cSYmfEFWkalnGmU4yjflyzFyXfHCakV9PSQOY7yjGnUbyfx7RSkH2D4RJzfSqmpzZZwrfaznO2SjT5d7hO3S/PI7KZnrsDn9eZbVnFgPLUTwNkzy5jyEKUkYwyvJImdlz6oqhAxVJjeZU6gy6XAKjNj4HMfinR/VEXlt65a+fXHzLDSQ/5Fh1ThZcwsb69EaBsTdO0IRg3yJYbOisaIAJQtXc/VquosnegHQ5jdhgEX2+1zdIUkZYYr+TXSXqyHztdfmTOEMtPbOkCqlyXwcJfP9NLGbW7Jlmpi2uTaJZlsw1ZMfxUnCVuDg45/db2BkoTzyOkSWYfsKnKe5FfmqKS3376m0fM44GNQ6dT0keSMLrcRJGfjoIX67NXSSD+8IRB1kcVPz8fb9re7oEaQm1l3jsDGkSuxYwOqfMRhtt9xm5Gi8UaTLTqyvD5MsXEEy8BpKjQhqt/EDUE8/7nV4FMwqXSJi5WFTU0WPHE0uQMMw5cDXPYD9YCTPzJhxyXhR4FF6vmINHPbSpJrIhlI747oc7r7I9RnJsTM+/vbIyBKFDSPb6g8bqSechn6jNS8wP6UvaeJ8WwRQMsG2pxTsCdL9rY5Z9Jvq5femKOovJzbyAu/ZikT9ZX5IeqYpEjtQ28RBkKAaHMVEQRIky5FpgvLBg9yxC4kmpqH33eWx45h9pBIapslf7tOjWWRUNxKbUEArm88NbSK1aL+f/7OcAvrg3RC0MPqspLRA+RxcxETTpf+ATpcVCgdljQzFvoypz/46Zvf3Ea6TsczT3cp2Wgf9NJ9nAVH/vrmA34VEeMBHhisj8S3f0eiFmB9YHVawzuJ5uglpOCStYBKhAOCQOmc5blV2trLNtxuLrRwmJb8+QGl2R9VmGlWenlr5Nv0Ok41LOH+VDJ5grOYtVVhtfBAAoiBNqLqdmNl1AzuHBeC1RI6pirO1tmwM6ulgcLZ9/hdzCe6D3HoAbd/ndZa4q0wOlAejFfo63FGqAX6apR7oOMNdUWr83jyii0q01rt1AYGbrBkdCLBzImKNEaxecx5V0nfxLQRTnhd8cydjoNomh9ftquoTrObmLXQkbSl11CuHITodN88nOBiQa5ddY2mrZLsrZx7031mnsMBXLo5/NtuIzNaQTeN4NymxZmsN1aPF6kc8ytYUQXSi42OHuDEEa57dh13uJtYFTvBUP2/NbhQq4mY7rkbSX3yag5jm2TBnyzydd2WqRFyEkDk4dvSu+S6q4wLJT76o38vUSG3ID03b1bIxyIRL3bRemUYBOTUuolHo1rdKOp+ABEesSYR/ICW2RwdnlVoXd347rIxPgVtH4HFVIqMcRcUuEIRa0J1FF1G0tTQBbWQqKcVDDdjrRzCZK5Z5My48Qt0NbQ2XoMOF81duH+w9Ky3bbkDqO0usQlqbngFEpICLuhD1jfP4Tj/sHZWLWYSOwyWBo6jgOVInrsNjRKiWllgRqvED6jAnYU5upsAHfzBQJmLnMmUIcS13EcPuXjjSMBasu4fuwH13xqQglewHi/3OXKPFSuI2NHI7zRQDE0bcUtXKE9ov9K+Rnw8OZwtSXZeZUFRHNIOCvKOVlfldatV4+Iq08d1DBCdW1BeaW/hWpTzk30i2RX3xkepg4gK+U/semW7ANGRRkfBlQRpAf+EPbpormkDKiyIX5RlnJQtt0qJyLeqt0jbeW4etP00jH4PwZOz5NHMCKbcYPUVJ4jB2dRqBWoIjtIKfluTtq0tNHnkyT7HpQFSOlbiETMdVMpI+xWt542sl6QjOb+206wFZx5TKM8mT73LL4MJkdXKfCo75ogXSi4LclrXAnvPQfaZ8GMSA3eAxcgPTCmCeesIs487OusXzS5Uy1ATlkSwGyRBJrhhrVhB/OyLqlX4ZKTYxNRGSRXxpQSgE3YihgVeJToThEIP33TXaeY6tNpyJXKQiNstjUyI8QVxG/YYCowcCVD5j0UinL1n1Q22WMlcuRt9Gy/PwzI8twQUFpwji2Yuw+ynNtDci5RJhaLL0L/7N07ET+krSulXBt1IKykRFjOznFdNnsa20CnbZYSghyMHvhCUkAdaxMgUcQ5hEjb6YEvJkaw+tmInSGIeoSSzRQMCfv45yeLGmdYWxxQ7vGrp4Cx0zF86fwZvUupk9bRbiuU9zf2tHsi3b41yA7decEptZYNFO1N2R4Asuu90FuKn+8JYsBhpkZuYlCneFpC5jr8aIu9APItXMaP1+at9JgLUjR/4xPTT0BCh2uQjpfp+z7iBLSYzqpVUIovsA+52ipDVSrKEazQ0UUXEgLo0A1fCwxvRYPFO1T2vWgz73jPGCzNj7003QIsMaeYvgpVpjLouI4Zt4Jq/ON3aDi3jL9Xp5ALOOWGJXtxl3CZtkxZ2+OftjDMnP86tfIqT74aCjpbkwyTCf1GUY24StgDRuJ/jI/ZR3XjTQ3UekjD3AvMp7xrJWg+nugOoyI39hgzzjRmkZu/UpDsYIL8xd6aj0ATAhKyajPTmjMcO4bh0uZ1U9sdMcNz24z95QIBbWKF/b2UwqTWJRqnFxUczSOGt9WGwTURNaMQb4vBw6IiJ9QHDGBazUGSf3IbxDJMT6wT2se6mPFJ1OqC/z0Cg8YTQvjDPtLiHx/1Rl0ZCSkJQE8lYhMMDTI+E6JSJl2lYSNfzqYBii2DWVy70LhRRczAVvhgLZBrNozZb1FPjMZZm1PcBppO3hlWNqHDlH5WPgNp6xjk0MCbccniwNDMSSrw2Nm90sYT2tqv99pB9bty3aLYPMBrZ7szhOjdkKC/3UroxAzPWcLy1n2hZ0gcYF2fX2fyl8p/fjJ2tGAe5qpQWsi4cUpAOPQNGMuLFj5PHOaU4D/XjdBYyY0jX3JPDCxlL1kKJblYhmGMBD6qJolqXoLKI3IerzX4gsE8J/WaD4Li1aW8u15dCriq6M5cbVBYFbIf71SY0HLdn3TVHmONna77mKoGb+V1Y8SIIkTITuy/l2lXyFKT1NwAVMjgG9+woARcf6u6lf5tVXL9qY+G5z607UKdYA6jM7fh21wCZHkG/5FWQ+QFGNXG40M9rNud4EZ/GJ0tF11lAUtj1EpMH8a1UqxL+WgESuTK/aTYITT7IeeFVOn06DmzS/L6XakiMVKRWHYjowzBV7HsOzrnwk3dGUp5N9tHWwkAYvKynJ2GyGVSYrkP9zAMl0SZ3IAGqvtkxmdZW9ORB9ReCufB2W0AjJAC9g9p6zjQyJMes9f72EwD/TagZXSS0kXvyzzoaKHg2iL7cvQ5vc5DZdJPg7jAUwbboDkD3sWUxz664rx/mN/envJ7zjaOIcZRddcoOGy5L/lnCk5/hb82frSvadkRIIXBzLzT77XrwKVSw3d1YlYqp+tVVEHaG6BemQ4LVVDRJTOARUV3ap+LhaU7ppTbTs0vsM7kAFg5bc272I0uaatm4sOIXIoqTxVfK75EVCvWGe8m7ro4ifcQ0lvyD5Ix/BfMumbJZVoJf+AmEnViG2wdTuRRBPSIEm4F/wU/L31uv4eeY7PdR+lCFUIPLD+qQRyHfF3zZmXmstaib2trQXi82CpykIDDMhm6WeDDrQEIBZr3mVjqrJKQHWdsEBb78KYevlLS7HLIoPc9qi/6hzeKnbpfDUkH+JQZ7Fop1yjXH37sk4DdEjCAh8LBYIXIKgKDpLncTiK65QvLtwHiVaKfuLfbh9vOOfke9yaEBcD0S0a5bQRzAIePMi9BoDDjYCZZRmkVfCfXa32ColkC8AgJSShH+hEBWuxWxhOPErCyGo+Agx5PTzPO0yawICX2XWyqL7Jn4NGuPoIvXHFrndhAVlEMTlLkc71riKViwY/ll3/mjv7mDEULk+K8pOHhHWhiIDs0hOoWSOfTK4fnxjyBiZZCZRjkBGih1hiPUKizEw7rqA3+4SynUIJP6xbywfrxxzkFSPXl32hAE4L/vrhdAf2DmjfcTyfqW6xTwWjNvgBbPmBpm4pSzgrAvUrI7XdoQ4cpdjQGCjvLOupUjvg3JgWOgZTLUbBsjLnap7DxYH4WOhrIIsqIaIr3k0pkMJDRgPzcHFPCtYlkxZpUByR6+j8poxkHG24DLUyXnqDs1urok+8Bn6Ypv3OVw758pVJ7U97b276gfvCxjv4UjYpyi9EL4u006BivnRsB3s2tKpdag35acmY/4zz9DletfC2PFEpv1DYueZK8GHodRku/6rgHm5b6MJ/XG0ODbcRSt00P+PzRWITfybXZLjuZXK4tVHgaTg5JmwU6hUTAziP1cl+v2YAjntjOVYRKe9u4T2xTCDR+gVCYXUlfM4rgw4NNuwkMZou6dmpPLGEFXWEO+LdmhlZNclMc0d1hjlbogxWu1XEJhiZH5ovmIBDqFYpThLnkR/MMPYFoc7balworRfGWTcWN1zF7A0s1VXqHUg9AqZ4WHP+Ne4bdp51BMDTykzWfn5wMZX9ws/jb7zh8uZ+sDhBhaCQ7rhxoS5y9P4tH3W2pjy3ZHH/mIQzCaLNwgQDIU0mqJIf2zOGdgL6d6G5wD7YyjWADLQoAawGPj8N/Df3XqE+HtZ26rCsnKKLQSy/yTtQE/YR2/QuM2FpdRI7IA80J5OLetrGtHslrGMCRQwfIzmlXa82OU6eCx9g0OxdK/AGu/GZDRduEJyVdUJdUSXZqn754oMD4GMTVxIS6lISqFfOX9QEBtE/ioi2qgcTXsd5YzWUpoEwTX1PVvfQOzn9SM7kIZSoBdM3WDO4TD/1igQT9cMbVLCYoIVahUxVyr91Dk3x35E8XVGiKx/jdMEueCZK76LMZ06G5516VbTq3iW8+TLLUclT4YnH1vcw82AObAHgjTzOlCBOyZS2Jj5fqamkTevVphEyzC2VKumPnjssw9fa9qC4+izmdB+iTuXKgJ+crX4OZRO4/ogxYQ9F2mQOk/rMpKNxO7TSS4b5EflML8dgTi7qluvECxnjkbnE8GqggBtEcgupLyVMupYdIWA+vcbADKF4/0i+zm11AL61xJ/Ak840edMQz4pwpRUYYnfktRhR+U5M1E21OamI6mpQSM9+dIhZQD5uvq1awicPRKG3FTh0LZLR/hkYQ/5Shi8L/awkUhBxorqlub/PP+1xkfwRQptIqtqyqqXvJDJWoi5BzJ3IoepEWB2WHeaPJE8Cyk0yeWxfCkVT6MQV9qCtFcl2wQSDmlMq/8huYbRWb309CHxT1SPUWTRhTJYMM0JkOcxeG+0R/fRMPxbptD6aak9NiNyL5ciu2/9EkBz/A6T+Dag337affCXjnc9TzK5CXxZBmNTe8dTKHzzXHMHPUOldR/2l+31y/b7hlY+UL4mcCgNV6d8zqZs4iVOJtn4KhFsXaADdcqipX5bdzE3PgxAw/xrNQ+WwN7UE0kVkgCsKoK1Gc2vHdvD+bjDEdzhyZFVkzNB9JyUj5eXTez8ddAhieNX4GFHt7iAvrLax2LU5UMxjqpRW/Py2x7bcd2QrKkZdgQxWzoC1wOz48pEQ9cFHuSh1ngr58ByLdr/ToJ3bbFhiS6aYuwjXcnX7Yt5NrbwcRFI+/9b2o2Dh7T9YwRKzkBCRQEes50gXYH2VapJE51D3kgzTfiqsfpTp9Gp6Y0dq4N+OuLjP1tiL3CjMQq+ZpiK1d1cJ6OvH6sUViZr6Nyy2+EUbNM1sRXfq7l1n/3ND4njjevE6ehZxkbjbUBiDSkmXiTzZxLBmhIj1Q3P3cEL1X2c1xUjQw9ZpT4zYSfDPy+ERDV7zaVBUjeRUn0Zbcm8eBzIE85EQw8Fnq3dRM2pVTWTuGqs/cbr4eKg9IixNzoHKR/Ny1WrcnX5aVWaDfUr3EP5LbOEGfizZ9DoDGbyZ6xZn6n9yn8hnm5H/OgcRVOZh4Wut9fw8N7jStvTsnkqO71QSdmTrJqcVnZoMJ+ct91sPH5ALLRNjd+nnMTezEf4r66k7P5r37YK5Hfobcw6hZ4KuJ6S+35qALiNUkjbvala/9knauIiwMhegOT8PhDfl4uh7A3bGwB4AQTiBxWzUDBfQJNcRG9epV450iG9aew6OcOIYleo7jef4i4F00JwizVHOXblwSjVgvncUtvSZuEV+AEOZyIaQdGZ5xU188TYJMpeUU86EHy89YvBl5YXD2S9qHAsJECkTQh6Su+NGOn4i3/hk30uxkYU4KuAIAHylptQYFtPjTrEIHITGxM2q5N5Y3EJVfEHm8aFPY4PpM/XKNHPEgoh+fyAaZ3QJsAtQ0o9i5fMocPmLBRoUuvPCN8nTa0YwCK25WVS4JyBxsEN9LqAUOKCRptZ+mPeMItxDEFmb/G+lpti0hKgv93jKuG7XFdAFk1pB5VMZ1aiAnc3vlUip/O88d+ezQd2VLcdMALsFX3fghV/oMgFatBHC1IYNLfhmVUnLc8s/8GkyeiTkro6VXNiaOctlT3CW5UO7hVM7or/ox8yDGcv9DKznDdj/ZPKCXzjXZkJuVXNM6AON+VLiB0Jlu4VPHa+OVTrgYUuW1qdMrIbDMFFSg+F152oHaGS+2ECGD31De5WCr4w1RKWMQy57EeTdcKS8wLV3UlF1kgFLi99oLy8fz2TWGP0rYFbiMKLfQ2oB5g5hwAyYeYLjgX+VxwF+Pb8bi7UVpK2gGmkJPKorLHo4yazVqc5l1nTwOyj+M28wFALiZ/dnMVVWwL6lemOi2jOqO+o2WEBFv3pe5DA4YRNJwBH/kwt0ynNhyi5wZqk1eHRE4Fg62M4NGrq1ITU71iGB3kn5xtwytPPxYKLLDH8dasTis2MQNMgqKbH1kmJQbjMACrNLgl4omijNLMynkhVE7EDp+jotJHos0/WyDg/6UY1RoEqnIYDuoxxufow/Eb9TSa+T9C4t2gznw2xWMgfxjMxDLIiC80sOYBjMgL5grDW9oZix0jpPkXYENaWg6BrolMxBCdlL/GXP9RMXa5kYfZ1ko0SIfW1o/1CuSbOs6uxuDmXaBvWXyAmi6IfwD8v03emKTOEOpt6yUjUe6m93rWQQnpDRXIpxgvafqW1xXbtiorQK5WxfMEQo0NNFfTmOwnP7s0g30p83KtNRfkZNE2Qfz9jyEaNcD6A1qK+bqUyI6kTBZHOhWrvOufZnToUkMZ+Dv3BKs60KwOr6QlQ8gIXct2oShOC4CgfA5SQj3yXyLDZF5o1odFSpnK0ES9oRYzcX5v+Jov6WQ91MXSaVsRZKn8HqRza+/S63w7zb1LM1CeY66Z6078W3VG+XpFCGWy7h94ljylvF7X4oZMOp+BOEuHmeqBeS4/j6ykJq0CcYAEzzQpEAWner370LpHeDQuiNH0n9tKRqnB4x2+eQgoVz8tYY5clQxAU7Po7fY9pLOfX/C89TCD7NwTgab8/rGlwZG3n40A+C2QeTyyGFUPSPmw+8LbBEpV74hoD7gA4CLznNV3QqwztXcSXZmE6UiNHg0VB2l6q6dTTNz6uxBSzCTt5BGC5TqqZSoJaGvK9M5D0Aq5rejlSjJNQRfm198erSapxvO73iCtbXAG362wjDOzVTQn/wQSwzcOWZq7QMCt+SNB37oNk3Bt2UicvBByhlNaHchF8U8C1ZRoaIHtdKPqfE5xdwFLzgtu3ZjcRiPyqhr8bGzLMdzl+UPLxMcseryMWyPnv8n5rPK7Fw7TlbIuM6MQhkdFN4kHqa4gOpCYRUw9TWAnmyqO/Bzc1ZFHKjN01xnow68Dp+LOv0vsRpFVKOZAAvhOsmCB3K7wvufk89wzW2GxDIBTX/ieXY1uifo+B27Brht53MnnLDBxQyguy1GaQsK/Ulj9eQaDNtVa7uhlXSWJP6gizn9f18ZR+VnIM6NVY/xVBhWOHr1IvzZqzl8bsADEKZ4a/ifwjw3K/NWz9BZQr7EmlvXWUzNDWQ3MYNb2A0TcTWOjg0IrnDy2z1Ev+IBnn5bZERutob19sTzMTYgPE9rhk45hGVvQDott6t5XwvLtVzuj9oaixR+xlZsUw417tQJd0Vuhr3LFUXSSea9FNbrjbqApdfEx3PM4hKx/UKEpAM+uzczjV6Pxdr8BcwPtzJ+7WhDlXOWXYtPNIo80b+9z+iFnR5qqL1eAOfT6UWkXHT8ZSUaqWfiLkXB/hcimc7SK+CGX9lzrdIE95iAvWbkh/96sU5JweU0I1FEkUGz3lDw+nLW33V7K456t22/SI2tHr1vvnicq7U4gvIr+ijOakoGt7TJw1ywYgu2avfhcLXmkpntLHTAPbuf7sXHF1gt4cq/KG8CdibIDGmV3EtfLxZcVpniBQU6/n17ytnJuMXSzzMyPUPXoImR/0tUIisBvqlPdILebLfOITyWQfjVa/yBG5CxWprOThqBHPDKbo89B6RyqVLPbDUhQlFADlLsGMb0HnV699QoMBlM0kwadEWfhTbacNgpAj+yvQqCBprjItrUQIBJSPicdsJ6jfLghUmAIqK3nAvWJiX+Oy2cWz0GAwaPOjLmjK/xkFnsn0bFrMFznb+rylceWMQjavEdixcW+jZ64Ck94Ua2wPNWBiPDVsA2izo0zVMw7vWFAfinfBOqVKBfCA/c+5bS/+NlU4zyD/a1MnAyN+f+0iE+51mUiXrlhnz/qe9+7LB6zW4CVvcNaMwqhdDdDYVaopU2KR9LDZQn4Rf0e1N24mVnfPZQNSAEQ2fF3qmAmx75n4k9nL/xW4xM98eZi8JzVKHXdeprE9J5Cj0lezLt4IfWE9p8vCEM3vRzXf1v9zC78c3oFQySf7juaP5LDkgevoPscY2iqVmgklT604WX0wYf/8joVm1hFlVPFhEFnMmIso9Jy+bYZneg5FuxcrXNBGVLZ/LnnEPCDUeJ9pxgpepQujkc60wxhuCak0JpRzurAWn5eNnWOwjbLUndMcMR5VsZiZEKBpqTqjCVuXCc2GWdjlYNGiYYwoPsUp9BSJxcndNjRwVADo+zuhRULdx7zd1rwKYlBtKWCGIFVsURUWGbfFKTlY+4cMdlXKCr/a/UNlvz+qfok4/DpZajT62EPeXlVavs/HLGUxJR1OHg69GldqvU7zRw94ctfq7KNuhd5hLaMhndUkjIKsWQIzXvWczs2AG/KGU3zpqQbcF0j6KG0zwLdXBFWL9DHa34a1/MhCiJqiY4pw/aGFkpQs3oD1mQaatMGb3VQCd4LETuArpA1TK7alixSnkSGWfGe5DWmBkCHCcvu5JZWtSJN0KBMG9kJwe7LG6riOCYFwaKGfXpOB/Ab0uORpWLsBA88l+Bf36iG6riHyp2LmiPgLRBWRh0dtOUdYCsznCv0wCs52FOlPex6nDZIcXz+cOzEdUm86LRV9w4P6t73vBEpCCbhS25KMPfyDyaQ3eHQgqpXdAO1DYu0T6xQPjs86fU8/aANKSeb9LpeFFWRLO1+x0cC9/cxbiHgG5xhNcyXXJOGgRphCYC7o2KNc9yUNOzKlw+WUYpHMfrbh0/5onTh5JAo07UNkfDORgfeasce9qvlyuxBOJNScGgIEyv8CWjd646aSH2FsAj5LKcO1topCTcAUoaeFMCF5SPa37Qhg+RppRDZJwYjjJIG31ix0WggK/nGRQI2tTCNfhyQnXYRsD0N8vEInLYeb0/+tv65e72v6Zm09mF7KSRwrJF8ZhfQvBDlzES+3WfMmcujKUMMRcNLwx6rilwI7krFWUlc6aCyKD/KDVqpJBYK76v5HVmoayoTuPovXp8oDGvn5Ry6cRqHxpfMiBVt6qHA8PJQ/XjOlKg9r4zYBATGhGxspc8f2DmPSB+GbgHnj/B0hle1IEfxXcmmTsB2ZOHM+YshMEAr09CFBpLZygpYZopXWCimuJZEa9NcMH9WbFXN8B6kGB5c5BXBN3jbaF5e7QRmIplHihAQWZ5KhQJWywXsJj+eJlJW73FnhUDhFklUwg5jpHMESwbCeyHs17WQiCyNW3bbzaDdL8gjtHOEleNYc3o6fn+DHIS1BrAsGQjUl5CsWybBeP9frYuFiiCqQotnJAhkb4Ew8M7r1zWyT+kb2wBtfgjrySCdE/iv5368p7ZM7RIBWn7kEQ7avNrI5OaWIPxJfePSCKa0dLX9gTKVMI6XtsEBhBQW9k4/RnoxaFTkcTR/QThlVkRvqi8yGkmLXptEEOkFI3jh/HN0FmQUSDBwOromv9bt+EDztEhyOkd32ckap7PJWRroVYDkoJfrcv0zFRP31X6LR9LzNtC8YhaFqV/NDbEQdk2q2lPbWeSYHDiRkbDNoZuuG0+pABlJ5zVf+ftGDnzNMIGBg2eOCQ9OgMpcw5Lx6gW2oVttZEWRbKYNAHaiqpUWlWWgcCbCdugb2YWTLZ6gwzLXCurbsOktFDnRxb6RlQSnECEUcy2cSXFxQt54yuZXFuF6eVHBIiJ4YvGDjNMIF7S2k9iNGu+sytWXzxtkK2yGWGo9iVvH3MUjrJWpYQYae/VTWTLojpeUw+b/di7/fnXY4iOLm0rO6jhjZthLd+D+Fk6uVWERpKy3TB+lmFl7kWwamVvO+MbV03VOR6IYEDCbosS59/cQG9MIZSTvFdmXXvRYxTnMC0RFgZHRetqDNDdEqGVCBXRh62dWIcRx87F7lsM/suBrRt6e1MVtMCrEXBd4FEzdHSWAw8rvmJYvGOccbXt1WtsFxjX15SCSWJFCxQrhWj/C0eSInuQ1RzgmT1PUAs9gmp07j9ACHF18kMuqruwyes3QRcClm/4cGF8gBr2FG0tV0jir1Wjgrh+YCBdOu0ws68yMeefKf9/BFIP5hEfaOPnnNOf303zi+g/7b1dOlrorWpxSLkVT5pVKUxXOsrc92VD13PwzW8brHZQ+CT7HAgS+c05QWJtXV4IIJiiXzJu912LwOfxmrDodj9psc8bjaxtxXyY00K4PmZa1BvBcjre1QgCdokHBnc5qc2owe/ci96rw4HfTmAsxj1CYVHKrLgN7enlgO2yhqRSk3nvEV4byDWdwu6M2kEd1og226N8UYbPSZjKwPnbSB4QJTyFl5LIPKZqVds+ZqY6QVKs4E1p1uwVj9AFM4CUW9JT4w+xHSXibBbLe7QJiJTGdvRSi5eB6CJBaTRdpTbgPu5+UyI9gmWOQ94IqSB6H2fYJzsdN91aBlkJXqNRPBKKledt/bMBol15cgtuhPL7CffTg25OicbjchWbxaR+L6amb7VeaDRKjKa5y/rF8AJ5+0su5MLchHLtXS01mAxbjOMXW+ol5fIaM5qPERlnk/WD6ZbQq6VNxuSx7kaQFdwIDCQmnIdyQNDodPGwS4RDvRdWurQLc4EQTSpzkRBSiJd5WmliwCrcL93H6TLj5aW4dSHGpL7Q8GEmMTH3a2uPpYpb9wZKugqrtN2p3UNVtgbcZVvr8mGH6FVJMsgI9ZR9g/YD5yQhjLJIv/lqMaz8O4tO6FpxWL1BTbwBFVUjKRHY9ijPYNqGFdaDhl/zk9jTIwjNJF6k48fuKpIAFVVNr3d3d99H2c1i6dN0QcIsmTsQhsOCKQlNQVWN0kNnD7Zk59XWLMNIXS2UoS+WePXy+gm2lm53Gj9BnqvpAmGVLe1fQEQ2J696opOujTLCcHwdUcE5fw1nKkYWsB71pQbn8E9v5Kkkd2oUowTj9bCCFVX+Hy1vfklgOtgCmYD73Zd3TaZ36vQxuj7Z0URRMEGRvIlgBi1KzPCCAHR/s3VFMbEBGiJ4vP9G0TrNod4RyBLcFv6DFYd8WZdl8rtySnhUPz5nl4lS3+ZfetH6bOzgXxJAjxUHOLVHJVTdKO+IYRxKRW2Th9sSvIRJdLmaWWdHsY74S3n9LNSm8A7APRCzeeMBZOqORi8/xxOjPTW4Rpn/vrpk/V9tp4PHOSMcXmXWQ8qzrCqklHLC3fFK5AGYpfvcZLU6g+Ds2H9hvHpR+MxxnCVT3+ajwU9qVIdmvHvv3aAKPvkUsZ0QOJusVZBovo8UK7sSn5ukyWitS5Dos7w0lZQ7kSMx2lSVddLXWpgTyCFsWyg/QV33AY1EzynIxXmc1zTLAPCYbtGXE8zFvmCTSc6ijEhblL4B6yXQabEuNkJ8FFd0FYyEzkzPwF6nT43La1ZaxCwUoI50plo+z6w5fV7rctFH0k1S1bGvFWgKvW7fK/3kgqFSuoMPJkgunHjPN1OuFdy4MtsbAZxaLZQ7cnUGhGub30kXPe1PzWSflsMyamCQ9t+Dn/mSkU7UR1A7VF2wXcbJyNpSr9Cl0kE801A8c7tctwT5Rm8/h7DgLrbC2xLkEswr8cSzc7GmkO64PEKEwkxAgTpfyDjC5FsbJ4ZoGkaQ+w1Q4/CwjUUhvuguCIxnuq+kjVfkAm5DAQW19Wnj9vFy1Zlp4Sx3/KmiiEmA13KWVcGks2vqHT7Wg4ctWHHNhJ3okxnjjr/nCsSBLcsmpF2J8waE/RT/ouBzEox2zbcKMSspvtev24NS+fS8Zq37TlP4ICAgD0HjIZ7m0WDKZXwQbli3YquRipyAeCg3SIXPWZXb7NCs1DFgaQKLIjS3nxTJNxV3p8ppLHh0J8ORwitkpo62Hy00954GAhnTZz9DEYevHmHj0BwE9U1KHrvPcXqu4NKKEMJjwPP+u7FEvDxFmfgYS93gpu2vUcqv1jlVnofYMRzUKCQ98YBqd50wxOQQUmcN9wqQpkHEuY4BwamQs+8/eH5ab8zzuxeaIPGAjUS5xGLlitMSO0RArHFWr6cZXdc1vF7x7RVthx/KDkYTYV9Pl5WUVFHckubedqa6WpAa9mscUQUyLkfL3teEATAGwI5CLWUlk3/kFNU3Ni1ECCKVh9gv0Y/lZzO2nY7kF/0RQ6B45mEjkToXSmQrDBpLQ2mhlv5FJ/8lTO3jO1CE5NlrvaggPjNrvMbEme5iSlmGr2anmrpi+F7WH2CfrwcvLLSDHDJYCNMRr9gR5Rd3OnrRWX7fCfgn45Zgw0yor4MzlHii1l3g0vACigWWRHOdIMxnj04kiyK9i+AELwzFvwZIrk17QaGYgL5AhCA9vnZcUUhhiWNZupXidb4SoGhqGNtLxMUV5RPmLKmz0PbWBnDO6t1cfWMzPFg90rrAonk8RJiZqIAw3x43x7iBDfJfQJJuuLj8bZgbdgavF1dQckrwWzxR2YYzcOIBFTpF4hpFiTHvSeMZ92fOyrJqWHqnV9uvz9OwICmEh27FiJSAY2MjEhCawVO3pop1+SbfdMZM9xTM4FvXiVHY+RdllydHBkQl5AYPskg3ASIIyEkTdJI0+NWu0CAlHjKKzSwkwSHKYbQK90t3aVWioWpHDVl62nm1Uai51bu+rQTOx7Oov+aKJfxWdLEvvszdxvNV8WSAAjUUoP5KFKsN7A4w8kAWUzot3Ml0/ZkLXlUAA29m+3dhAbWtNAbV++8LuP64XUDKqUT2VveyL+3o2zh5OMuVP9ObG4LcsQC8qtGv/1DkrPQnWxTvXvZd3vPXpgB2+U7wMXAm3WIP1PH7wKceUjZvJsLsknwvz89pMDiTEmmozSCvL8svq1+8Q9pYz2sY65xdFNkV1npRVBxiV/1v6mHTMm/hFX88hUtULrH65d3oca/MVWF2lqhnyJLpr4kBQYhM1/iC+iI6vAP+gLTeIJbjmFo94wgNCLwmqziyiFf6mU/jcvvObdww8mCb//na12pdqvl8qbAsan/SlE2mAABhvKwEG2z/CVoX79j1ra41hZZCqYxil47dzgrv/vNGZ/LsO5Z7xk9mtkQyV57TqZ6+hu+uIiojY4IUsg2S94GOPvSZYD5UZF8CiRWDDTR8LOKwtB6byM63cZ9S4F+R9abGzeegko02tBPxp/o7rPAT8kkrabV639b/YpWcD4mq9U7DmC9AlEbgDDSroh90VySkRi3t2W0peUqQQWWKn+5HhrMJ0rbEDrHj6x/mCl7E4EBtCWHPznRSzgo3CGEF1b/kjTEoMA+FgtzLz4qTOXuTCa8fwUwmKBxFVHFF8TM++dRrFysupzhSdUmJA7B2QwHlpiY5Guksn+Yxy2FYxFHYpbB/OnzTVq4DEo/JLtCYYTt0nuoKGGzLe8HUqeecfsybFBkhqxd8HfDAVtgt4vTMzGK50R4SImBJOCUdtadtP3oJQO4koZc2ijcXJ6iukM3PW9Z8da9qiGqqpW8wvkQcPc4WeMnBu7c99AacqIHZk3wDi3cZw5lnqTtX1OVryDR7vzSeaf2v1PTR45+uGWEegtvGXp8w0ihpTZ6puWASt2Hkbk34bRoGJ6WWAGqdzr6OppGa+3CComVabPIYArUs6vgrgITyzjwXZ/XL7jM2w4VggQr0+6hZGkfiDn1+tlVJTSrS+kRCgj4QTiZXzZfVSkg9RGoE7UHGuC15/BLv/6lZ0eSQsQujdfdkRXk17WX2MVTcJsTSRM7zIyprauW6/nzid0LU4vbuzyv2q2AItqIr/dINcjy6C9/fantzLg5rW9kSvbG8jQKgpbfztJuHJajAkWJgzAhiZWBcboAPmMWBjWl8qkXtcXJQsoXVZGSpepCxLxfIPD5EMbiHRprPGct8CSfVtgAsQSIY+GB7MBBPsYBBu66rJ0ZWCRmT+2pHx7n9kxKPIQc11X/Sr3sOGU4rLr7dGV3OZ/AtSiY6zSfrUU+6lFyXxPQ2lWTB/Ni8tf/0k6vQCMCB/BTtBtYWOwsjTr2RwFJ/Y5qkD19EMs3Hghhm61y5VnSdbRW7+jFXynJfnO85umf2+q9LFUengOB3BivFmhaxv9L9gG67KKSOh1GYtDptHAYQMaL/AZhWlCZ6yuqv7Hzi+rZf6ujpz/uIgguVbQqSKlGf5K8j2JxMk5I1n7/sHf98/qstsfVXHTDaiQpeDWbZq4aYY9+oyDXLQJgx/gAuS+SNxKzkwmq3CXX01VJG3qtE2M5oIjdKttOYyYJA7KTMHETmuLGiMA5TNSFPYBi2UVvsQx1yNfA84Nm/iQXz16T+usXMOdMmP7TDGFHl36KM3SYh5st6Pt0zqrV/G5gD1xlNrDmcLi7G6SsE4IZ9hveuidMa6hvfBXxpdwBLktOwnxCrhyMEGmNTa4s1z3WrFvn9X04N/EtGfL127t6IOggG6zWO4dKy+EirMwqCbE7ZTgzot3SWpeC/zBDpKLaTToVktXcCOUSpig+v8FyBj5vj9sMjylRlMETzgQKA9yY+9/AmrICx4uV8RiFRAqZr3AyBL10zWaMiZTkFkVA3vksT5aihDadjTkbHInunjlsrzGRlRDWp1wWrw0sD0cZjL6PEW+ObCeVTzrr1+IO+uwn1njM5pPrvNAdx3rlX5/WSVftVWp6f9WjvxfJJjdc8ElpY6+22Kjb65uUGvoGWLi3HenIv3j2IcKb4De2TUMrR9QtXdBexw2+bZY1A0Vt4OQu13yluDBVRN7vU7+Hr6QA4wP1JEQS69E4uyWZeEjaf67u4s+a4MJQr/ByQ0TjCJ7+ozxFQBr1UlB4HBOg3q16vfwf25c+CX2L/Dg8gCUmtCrZg2IQzIxaPK3X+ZKbwU29MZJJqLZV/O2UhBin3YrR93ly/MMvPfbzY8FKzW4rcfN9m6/tkDFMupWJEqTqt6RAPKfPyHKrIHHlSFiiwwaAvZAShp981y/1BLAQw2hB/IEBTeEZo8o6pMUFRiCWz94hWSj2+gTC1bblyLQ0mrb0zm9QGlyKEaaLgzCY8OLeA6N2jkA//AuTHoTwomAdKFiZHKY1Bp31jeIwm1NyZKESZAFkXZu/wysTkGq+MNnP/lwMZfl2JtPqEYcy2bVofL5yDG55R0uxkqm/kTW2ssEtwc1tA6ttHkYWzC2ik2XqX96yqhTAz3rkU5MI6Tux7uxYefEaXMkLQc5SBGHS+/L4H9UVNOb295dX98p1KfyhxKNJYjchDbozODbBdlMghTSZq3HaVGzxwFvGzo3yaaG+iYKQf7vAJ4/6tRxqTGglU4L7Z4kFn52IsguM8Xk6RXzzXMFQm51AoePWmP3nqf/7GZIK5lU0z/zxQNFIUS2VL+XZopGZlfcv0xlohi6iGWqAbn9JSIlhuM7KHFBvWprTgFTZMIPOaztGQ3ixyA6QUjo/SSNwzDZIOmKiXwGgJc+rh/yqFQ6zd0grhnYvSq23ciIxTGAUtey0tp87uihzNTUqG990lyQNAqaCHG8Lj6/+44r1yqKr7uBinilE6U/6LqzUwVyO8h/xGdJeLxNt5rX3gAcamEO7SzFtgG+8xQo3U0TLnFb89Ge497TAGSH4rzbjmiq5D4JNcrJ+Kuw3UlO2GqwIWG+qn/LhtAks6Q1yhv63zNHoD62oGzmeev2jFOIuHNgOmPtacUuh9K6ZAl/Ip2GA5ZErYDX2kTbTPUnMvONSK46R9sWqCZKMoQUkC8ZbxE9rUSUxjkY0qCnBZDmzOfxmp7m433MkqRIuup/K6mfxQOiIZcI8r2j+NFrhv75C2XurhwVjReZB4CtT3ntoUCzGl3hFN+euOKVfkyT1B5zvnuQymWIaVtdcGOkMj4yotvyPyuPcci/OyPcYunLwozSN/KuX0bXmazwoXZAKT3hZarWqdMQg9SaiOHzzzmTJqkcAPZyCJow19Ivj9G64Lqj2Rt2K3w1GBDHgRyS4pDZ5KPAorBJh5B4QKWztYkwIEGiu/hm/JwxsXEMolTfNFnvdv0OaussSr3pRnik6uZovgViLCh+WDtkYRUEW2X+rSWRFxW7deACi6aA6vf5IN1dbpe3fSNwACC2LLAGIRxETQw8459hD0A5mmPAQR1DWC9qi4tVPCxCGvBTwFlD+g3/52Z8Oa2/OdorM6xy6d84M9Q80S/eHAyON8rtyH8P4udwwG/n+c5leUeKFqCi1ASwCx2deNW/CicRfSqGrmM07n0hndne0EtZvqHQcGIiQGWXIoxpQrJ+/r0zvIKQSHTY3LSLUmajhqpar2t4gA7MBjx9id/rbMVjwaRG87d95Csr+MCcHHIrOzazqn7AK2LW1iR9TpifQbD5ndBUX8q9GJ14Gd0LBF36op9hJ+0VRwRFPuBwYwFhkDuxvriTiiogpi85QcXTQ71nk8GHjneGsbJU/fr+BqgO+ELSf8QJTx3ty+G6uZ9UoDK3THuhYxA18dMvcvJhHTB7a8NUUD4aWR517PUvbv2ZPrDEMNkhUdeYqxcN/hC05NfsSKCYxLFOZj6w41NDZ6y8bpFpQtbzkOyN5NFEcBh/DJXRnOVe/orM001CjF+sA+jORwqF0k9GmLCpzP26A1Um5MpuY+ZxaOIiA3Iz4Khe3Tv2gGC3E4iqTwM0VkRag0vfdDzpXv6wQOfKh+9X5emr1/FNN/USQI2+dRdmnBiB1v0L/OGVi3NlsriMEJA5wpLsUb84CrUxXqllxa9Q5O1PVH1MxGrmBqbXbnR4S4+/P+Q6FuKlLKk/monLUlHMMge7bgXugaMqkG9JY+wLfrIKOJPHWU/JRmPO+2kzqxckH77gPHYUSdE++jdDPJu19K9u/eoAeIjywlGMed74nfkzblEgbMX+LUwsOWgkqOM/EmDEG40POq6du8b+Rp1LP12ey/p0tUqoDCqOk1Si5tF1poCpw/c1HEy/xHXU48KaGtvb30gXVvJlMM1UgYqg0vtVjYWChjaXs28Glxfd4jPqJ3Ohq+gYRx61N/p4JiGAzxFVAuTpFW1PYkup1jwXC80MlKr3WEn16q/sThMAK41p3n9PyMSIUKtxw5Fh5f0azlEEMPMaCR/l+o8zzfYXn95VzQyjTx8R5A3OEPpEqSdiQqSXKTpxCdoFDmb94l/Biz9kUDTtDkhfiJ73sC5DOIbx7MMv86vFpG58v/xKXgKKyka3lNOvrNHd9GDyKCTYo1Z66UyBRzhiCSKahvuJLhhFNZbLYtCXo5TMNFeSOlJ/g1Xa90QponKw77MQ3vFWXtlIcZWkUjHEXqB58sOmbGk2nmQ57m6uKyaBWUJnicWJFGq3vLDziwnX7O53jauve+2cP2dewhqguBJAL+K8UMYHjBFXf2vDbzR5cztWx4g/wK1n34ApK/xpPImEi0DGeWd4uWO/sCQATmkcujTqwGFMh+ru/rMlDfjsUu256aj1UYbAQ4y03uWhzxJcyB5UbSUnOdD3b8Q0xrrWKe+Shh/a7MPKIFjfMgziA51sAcfS7gWXH5i6/jwRrWujXec1Ryrz5kuE2Oi/1nvVesT26H5RgWMZ8tw1zFyavS19lVnFOEiGzbhw9w9eeatmbcTfzlZb5qxKZ6XExlZX4ftcXW2/cXwNsvntaPliX8YlVVGqB4JOCLGPUlKrq6Bnl8PMgX687fc8mcxLnZ1PDo2YUUIxdSHtIocXHKWLAjB93uSlmCIRSH3ew/+NdD4QKKAe9D4OmGcGCdBNXR6NdDBfQqDYiRVKNM3z/alpjLzjhY09r1crTbSxvHr2EoJGNFg0cQ3zOSEo6weAb7S1H4PiqsfuYBcAuvm/md4wslIkJdV5IqkAJXVgWE+CLSH3BofF+moR/WGt/wT9jSpvorggMGjQQtBlkd1ZS/HRvwK02xCS36sDjqW2REbmSXaOeZCL12KPIcOhOyQcINFMJ807aef7wu3cMUFfKgcHhHpcTAHprg3AKog1Mr4yk0Rk1j4TP7eQfNacaiYeo291RHolh6uGSsAfwTy1hsR1q3WTth6Y8Uyw3wOES1x6H8wKGjiBpoODMRufYKURMm1nFyzxAEnoikwSpen9E2mmd89+/1rNgr0yvZaOTMo36yOzkN6EG9YMahJltx20qGpnlnmBYT5MIsWYyVXRgNlsZeGp+XjaYM1syRDSVfUO8U9gDENxMVc2x5ZM6ACpo2nziX4bo0TKZP1oqfiOiM1uAZEn/d2tqEgGK3n0e9iyN/goWGX2I9Hgc+kzXVznO0XUUe8k7pwo/mK4C5ECZTXKlJBXTJjZC/AuQsbnHGlJD9iro2EYwfDEcUUpyEBEqFC2cT/7uT22GWWzXRD4Y+2RziSc0L39JJR5ZrZEop4J8J+fIntpEf/ISQCTWdTf/rZ6p0ikIEvtc2AmSJdOWWQBA7AMsczSeQVHd2jBwvQ2fPnSciYUWO/vYGSFwhvzKhcIUItS2HMTCIUhzTPfogc0PK3L2lQGTAG+ptpmjnUXxnygQ6VclNb7iAA3VDm50ECB7dHr2HK42vipiSnbnZbO7rxFFe21w0PKBO813ekiD0XQn/c9AwBWO53WdTX38IKnrmNcFPEXf5T7oy7rhFORAsFlcHBYCCwEEuYPEYyIUahud12MQuRRMam7MoSGZd7T0VSOBUfDlnYPq27E71dWcFDSvEij+JyUxVEw6Af+1yDD+XnffOT/7LHdr+FL7w8+cNJHgtf22XSf1zWb6hbYvEYl69dArH4uJ563GCrcgPB/8TnVqZ5leEVQdce4UoHEFdre0Wvy5/5YeLPcexEQq1AoUsxXieUFaHGE0Cgg3zH3bbegH4jYuonetIiNf2l8YoMS+MVcywortEGCGv+AZFNmlstVxmuCFElHJPotrlh4UFXMkGH/bYaahUA5LNunbB4PTSXByPTP3AOwNm1oOzcztnOqmaCeiuz0mYP58VB4lFN2lE5FaYoUz6IbEQph4vzFVo80mNDwD47bVTw7arbybaxDQ1285ugNFfGdrfkufYTc2wBXYEmaAdQfqAc0/VusQrt1DEVI+F+h27/hrg8Qy7+XqCZtqGFeH43BaErb6idVBphzdjJhyr9jc0siqb4ZavjhbTw7AvkOinRamRCDD1VrxnhLXz7BXx/vCpOhLt0YwmG8ISG2xSEFG4d4NGEKPP5jQ16/3RslYdLdmWXytF0Q0hqk9MNRyD58GSUXlPETRidi+PuLWQPfBMzRfwVeMdC4IGOjCi94ZEfGenV7ofm9bMPFCntxRPEwYwSMbHGW0ZLQIwfDTSioxcHgLfstSlwytiW31aRS9Ou5VU8oHgldgzcX8UCeFJVAF0wzgVTGwwUMhtoM42aF/wORGQfrNMd+qlfpYrF7qdoVtgrtwGIEVt0ek8SKro5dWFgRIcx0v3pn/CFTT4k7TgpIYBzP1Zx5vVPk53Twjcr4bkdtdjxaBoch/XRX1p1ZFjr1il1vPu2sd8O/uIOQ7o7K/JnY9Llf3+ZFAeKBPja2PIDLJVDio1vyu4bdFFzMLX9iQiSaI2EScPLwyF1LkjF9BSZAp9d0RcmN7p7yIE20dramGxrqR4itQkruy/ixSWG5rCX9a1GY65LWNPRumx/nZuxe9Ru0/9sR397He7R7YRfWuJN5tXcqPR3SiLnBP1MrBNId8fJkcRvevxv6ZsI7eqnZ+D42bQulSnYgYFbZv9re+9Io7QvVltIq5+6/A8AtjtCGBqJo+WWm3aLD1+Cqw0J/wrpDFGijLwZYm3LWbsvIdVl8j/1iZ1+FcuzjVqk71+FfWGqtv4R2p/FE5nhT+1E+0+Tav8iEoysOjyywhROYlLrqym/p0Vpk/YtGA1WjOeOo+IQibpKwcsrj+Pg1WDJG1mR5r1915D+FL0byp8tKzDKFmkJC/m+2qTYpD2530BPfcTDm4wWuklY5nJLPvkp130itj6kcWhpo1pmoZ0fuBh7NZtLtZqlyELzYubqTn067bsHdho4SXSIs2PPAZf5VmuKyC6nQtojRPOiwi+ThqSsUihyNp+VLnR2a39810AJEtwr0Um4LPlkVNbHpb/BxvO7tZMb07wdoSZ3xwLxet+a68/1vwVm8Gnt5eWi3ZxtcpZ1Fb9Eszi/FWjs9rNZd9hi5szlbkn07hgdWingN2SN58YeRcQuytfuaTs2388O6JjXGWEyo0gQi7N3zeipJoPHth4yCcQnX1sxdktxnalpInagafRIYZ6b6QWl54Hfv6+Sv9ZDoNEEqzvlasv8JDkJ8XiePQTu9AMmfR2dbgSmfIzlojvrfHc5EWjomGEVCdj55KvE8z1pgRGc6SXLCPFeP+q0YrV0iV4b4pya57POFnZC0hcGgeoEQS9Fgafnfpa4X/fUu1fjUVeoN0vV2PqWXkbAt5PndvwiCjeOTto51pyvrK5TKNp0RVraYEpYfSZJ3uBPD18wCuLDM+JTpFAu/+nIXsMPaojN2+9YWOH9fBts282A0/2MFhQ2j48sBU96CnZo0lYWtY7baGID04iiiIIzaE38iIMZMmu1RhcKSZZg2gXIV92MUhOtnZMDCFTN4F7XG+KjZqqkt2xQMx7AeEfbDBAngds+VARDidV02hmYCRzyf6I/2P5CHATTEYFGKfXzlx6cYhM7p3HCTZu0bBzfeSVxjs02EGq74hfxm3jH48F98xQxeKTdZQdVxOqbU3/dlrSDcSdr+OLqxRVTBGWYR+lPY2UDi/+r/WBon5epnPlNeBSHYj+1uHVVhWX7f0zGqdANGl5RcYBnWUnULaCto7HlcP2ylfn912xikgkVsBrJNftVDXsNAUbgRwaKBFNv/xmHo17TQhemvlrNmHJJZB9TBeepXghjggkz65riyWeKv4iDmHahSDqA+CELNTHKBTFyF/GOagTAPRTTlzwNlCgBEPHmP1FzMvzikK6fNTMEqKtjqfErCoVjRhaYM2EB38HPbkXkxViq8IfAFCJcLJzVThuAcLaYk1pxZkffjlgq4wQhuviU0MJaJfWEqZpQ+AO5MjZSbDbubE5oCRRHi1JMToFvF3IiIjpqHpNMDn687YL5YEAVDtabpSAorYfRXZYqGqvXVktQkvH0Pjcd6tsIvXFWh8cQSNdhk18s4N/hch5TZ0g9WxZKQacmbwOUF2xRFx0azl+GoSKb6v2rST99561lwilY/zSNeudCHo2pq1RFAWhMTNxziHsmSLAs7yci2aXKiJa0b8XBd8ZfG6dtKYaaZlAhwMzl0f9Y//U9k0CnG+v7cIBgxYNzOoRj3fyuA43+6DGqLYhgABBUZ2V3UEf7IJ1lIbdV7UI6LyFzea7L2T2XxGJnA0zpZ5yFu1TDOtrExXXGuX4ffi3nseevXIbqVi4jdatJ3lHLge3YNoe/uhoyrr1i+/UhizsZCZp6GcRi4ZRMj0m3ebwyh8bp6T2CFOn7Gd6np8cFuPAhWhU7KUbH3rlCOuQHx5eszYGk+sE/SGOfKMVgDE1jm5Krp40rrSkDkvSxi0vAnP4bENqSNWLJb8v87MLKAul0zTPF6Av8tLjyVIkMgmhXxiJiqZmonMNLZ1qlqaRdoke+H/29XyHhS8CXtibbktm8HvLZQ2kg6lWVwxcNRRkXOsIsHATtSfceEmZ4OawLAbn8Itq2Gch7Bcyk8MCZyMOOiD+BSuwEeHXLONdzB3oBBrVABx9nwFiqzdvB9TTLcsWcjsMywRFMCR4WSh/iSO53SSfhViy984exMOuqcJaKAekPJO2Cfp1eid+6GmOF/HHJwYpv+WG6cjoc+n688SeaPLAslUWFY1fvwbomNMq+HrrV5FvG8Pcwt0oS3dyBXlA24xqiIRlh8mlVe9cNYTTb0zC6omiSSLtMPqJzyqHyjKGboToSWaCjV9awoRh/xk14ihE/+4H8hv2/d0wgz5vgKwx5BNS5Ie7NPId/ZKdx8vGeRKd5xh0xp0QCc90aOGlp2qc7e2rEcU4HjXHMnqeLE/t36swLUBCRWhQt8aGec6lMMHxnODZUAee2No+dcYcYTZFrTFQFCdtEblaZZ7yloLHotU96bsI2EtwO7fkgoHS/zGd+2+DVWQhXEwtvyq/6pjSwFc89NzTgwYnoA/sFQfWjO6yPXmxk+9GURqTYRvWY/Fk9/UESHFQX5q1kKxz5MPhOXxmHWRXiAGh7NrUMkl+3nYM48oxTm+q5MVuoqqDSRbnphwR+lzx+uhd14ZpHIAD++P7cS3x8aIENun1vGTDaPXaZH+KhEIqPtb89XVbxhlZ6temDmvl/4p2ze/Muwhv9KvKfSQ1oYC8swbVAdMgBTj9dz7f/4iFq3ke/RdioEUNBSnZJI2N1w5LKiMZ7ZhRJGmg83eVVBw+g4H2ePnrwUM09iaGOYA+3yY/E1wN5V56rI55jab1BtNwyir/7wr13xN9IsLRMu5Nin/7ySj++veQ5+wAxTK+Itoa6mHwStpoVuTMqnvGDZ8c6eXfBh+t5rVClvg9IYKGw0BP2+GLiyJq8foyCx2yAuLzNSnMZSijWOmxlk0h/KLNyTBCcyxFYXpadejJC0JWd/4PrQnog+WmTjQmjbb6INVz1eOFsk1uUhSUlPHkR9jbOjDPyXd8aVMooOt5ntGd1kNod3rtjfK7tERyfIN8bBNJObgfLsN6XkN3LpfJ5BSooOXA+eNzrrW4E7kcCC5tYT1aiLOoabqX3bQne6uicse0t5CzFqCu1Q8K7OUA4diabNmXXS4vMEOJ52TanFKEwfqqMO7nyXEvgX5Wk7NuXsOwkXHeemt1zj8Q8aiy3v9ZUCHdLMBYqIQGb7ycMOEhBU/gL66Kzu054UGL81RvhAWRHIuztcdS2qath2JF9cu9wjGG9YXfiFdQo+EKpyIzbjFtMXxv84WwlT2PQRmi6uc3Tv1iVAjAs+FEu33vlFWYJggXMrvzpdT3H+kRZFBcmvyv0DcYJk872XMzkmookaFktthmDblVjq20URAbpDc4Jq0t5ZhAehsVyD2P/Tn6YDcmK8pDy9gpVaXTX4d4jjkFxYfOeUB5IynsHpw+yFIrqf5cX0dmkOgI0LNuuBZL640ZBd7CDTM9vyiA9ig48qjrNNcb8bZrx1KygwCSFkcCp3S8+EQXrP9AEfwRjbVmbp6x8CD2aJ0tOTr60v94S63WYQo11dimmGauH9OP+Z+SitIUGnLhV2rt5NzIRrNI0Nz09n3bWLq8pbh15IcLRlw0HdWKYMBf/+J1L4XFB31QfIBOnam1fuzuFGr7V5FBsFqEZy8FPdYNMfYMil3MDRPai6sV2IQkQ9I/15l3mHft22dT7LGvjR6ExVWEjaWtkE2uK9PBCh0YMZk6lIgeaq3saDrSVuUKsOolrf1LRV4Lx8IxmJIZNigIJdPkrSW1+dQ40AOgZsnSoEBwMVTaANB9T66cQrDBV6/E3Esmdb95egNadKtcRZZa92JxVFmWg/5gbkMxwX/95p26M68JpGfxLgYGnGfihR64ZuuzW1L8fGxJ261HTlzQMYTGS/0CFaVUsLDdmvvwviKZI3WrDsb6kZ4tQrFqb+bXkFH5iwQzl8S0L0xQaCHVqwxtJbFu7jxY659HSelVkMq/sSrgwDSTmZMzO6GJerBfXTc83VnWgk1EjUdr59eRqldtnIhhmnJz0yCtgGy2pwucZrjQOJV0x3dNNAWZR+Om7oBcFtfS6gZ3GmeKv2bCi6m95kl/g3pwfLFCSJVQUUqhEDMKCITZCVTLz7rKjFfJnE/gNPKAMZm92S1vd35WGwK4t0NaYQ1jPjWSMsN7QAbzsyVjwYtzbk3h+1HRed+lLWMbL/7td/1M8XiSYiwutFveoSqaNOSdLCk40LSgtQSbrQzVLPWHo2MGN0OfXYSr8xKYAGLMIk/eV3914Mir7khjXreMHGmqTvDUgrWKISsMdIMW51XL2UPUIcw6w8uZMKqo4Hi93bCT5XW//ZMHFPm9XR5H5sjmBvPB5ztvSRZBokJ09hUSQvfGa/8ffRVirpKvVz11OudAmTj+5Wm5RlW0Y/bOc7amq6bNKOIy07skZVllkgJvFIb3hIYqpYY8g5Ih+kgceKgL8pLGO1qRIgbawEz9lAzRBBLizCj2AF5V+TyzmN2g/3MtCfyBsQKLOLlxyI8uFrFdfYtIUx/sPWSIxoDOI1MMUh7WksLFoaL0L70LzK4LmD9Ny/Yd1hE97PsGg8kFhgU7naGnsWpdCE05cnbyQC4xb44jpVDUYSKF9O3xX6xPp6Oa7kVxnjmtZzMyB+HDwPcTrUoa4PVjpxB98LXFg4Pg2KfJJzhu0IdklLk2iA27+/PgZ2yKLk6jkHwUjH+rC3zya6nnEUL0NJ+IdGuGL4c2fWdq5030zLIOTpq6/mf/1WvrYLod3czm39BdqdIWkrDS8nkBtvabw9yDgJiys2wggt8h0Oo9JcbAuRn5RLH5940R3HwnDrJmt8l2AIBY5bA9kaCeJS0u2Z+n0lp1r1GJrbYisbDjAYc9P3SDrqYlZ5C33I+Lc5lKu6za/QUU1lBNBJ1cZqj9GvEV1Xt4EjUi/uT3bQtHdhs6CwSNlxQIDyx/+HXCUFZCdiAkndamW8SftygHo1/XvnxHHAZkqI3LCzhLChe1p/Yefeai8vEQc5xeZd1j0wH+/MEC2XRtd5I1hjdjf3Wv+GpHgU6GEItcKh0INA/aCJMvrZAO20HlZcdk8bPmikMUxSDtI2e2jkI5Gvm7MzUKApqWT3nCvWLSJ5XBOgnIiMs5XGiPKgwFfpr/oBPJovXn/x9t6oYFv5XCl/TJ1DOhu0O0GptVFmpGQlwVGkndXPKG9gxP+VwjfEcAGT3iCHiouR1+5w+jSqn3t/DbJgVFtncCSJNkcffD2VYf8H3cwIrQ3NqbGRUVqWV1o4iYfw0r7qVJtC2kxcXSbeojHt6DCf8/BU+KYYTKfK5+NkIeweiGjvxKWbiQp5jewiSIHTpz9Wtw49yv4mgLGi0lLHMRq32ZIrRa0Gk7uzmiDZ0tvzbMl2TR5XCV8x6SOahkiHkb3WZI3CEG6xiC8uyjN/LoDdIzRFR2bOWr1QfRHhCEj8VLASfVwvYaHkjBPNRMlsGVZcXkWEG+aV2n9p2g+bTfFfk9CdMHrJ+tTmrjB7Bp9QXX/zU61jwgwHl4+mVyObVjV7oOd71BNgV2zr9oEW43alG4hTDSe1Q3kZEZrg6chaNcI5oi9VWUKgrYLhJYmBq4avNKmkvln0Qe8XKLrFi+emljK/JJrKs7dgF6PNeqf8URTsh1RPlWRdlzecpaw5uIGix3TQS34kdu9+INA/91MUOpOFkH5lYIThCqpYzT4iMMEA1jHocvZWNxb4X1aUIhUJ8hgPVPtUOPKdOETGVCMzp37GTZmAyL25x08xPRfO44c50Q9BKEc2BUoZXypbF1VvWRSozza3hhqAjagJ2Upkt9ir6sexaDZP8y83xdwsYhaq5omh1TmyORlNdO24Lb9gvrbQ72mEDMjZT7BfkxtUz0j+Q+gkU179ldflIgD9FTi7m1ZLwCmNZN9jFbl8lAU+1nG1M0eI9JPdrBNbfMM1uoyxdkcLMyYVxG3jmHHKN3Cg33kAnsNYL5YkftAkH2b/vYZAeMkn66IjBROnN1Worjon2lJze2mMcSYT4QSNJ2fi2CHAsYXnXRSmZ2lbJVCS9jGr7SLUdo+TrClzqduZrQ16HL/Y3MCelu+ZdrdgUeG2sPrt4BHaNOid80rOR8Wp3W86UPqm3XUWxKt1e7fO/3EWLwr7rZlj0C6c/rmLi4vUtlZFmibzYuDfbq206n6EDmIFWOQyGqdW0u4VF7/jx2uzlrFtTcYH7q1uM5SECAgJbxh0WEpJGyEbWj1BH6ctZdl/efLS1ArdVpgmu6y03M+PCAl6Rt5C7nXclIHvaRwPlFDWI6HlxbHPcX52EWEOXPpreIoGkkqjhVaU4ZPtStfktD3cur9974Z55kI0669eCmDWH1ADwDTwjTC27B8FprnucO/604b3kc0nmjuNiG3Ggx1L6EiiUfYbkDYIN8pMW2sfVUroUf8DWQBVtGrCFuw0RwW490nAL4LH/lBEYMS4zFJi61dCNgkqREFGyUyPRmeSxKsDBfZEqKv843YK72BKaUj0fZ5f58uj30JJQ6avY0e3hFvKll8wNPFwMReqDDceI76tByuRXW7ZtRM3Nok7NwxbQ7LDvHzn849gKmK1qRX+LEKrCkWx2PdaezzQpGu/TdFw19QPm+mAO3lbJmhjFGfdTyjZdLYoBu6NwcRRB3OfvoocsOD0O6cwTORgfUrAGdlx4IOLhwyHm40lh6wtae7DsjgCbJoMOPIt0UBJg5Q0qJhhn9DLsBJGZmIuCuh54v7990Dw5LlZgJitaL+aK16iJ7BhQfiOgAaDGlPfmF2uKOjX+MirP4etFB0IxmjxCSbqo5OGlFbQ5ZZLN6RIFtgX5mkVUQLTYxu4DUZXXyaO7z6nYyHJ/R4KHprM0kM6Vis6T1nAqcdKC30xtVUcUd5obvrfIBizuD+4KXMiwPIi3kv76jhX1o5+DrBMjEFQVU0WLL3Et5IfGsh6E5Tq9qW004TH9NBz7etTJeZ9431Q9ICArzHPyK84adAQqc5+re6YYjVvdOCRHSB5KXh//XAndZt4jLq0E02g/HKhZCp+x6aqUvHH9SWutWZLqdTdWbupTOMf9OpKu5pVyujwbX+5k9cEYa/a0BZJaAoJvhvWQT2sbfmXYvjrOwojK/jmGcDBIStyk7a6xf4+qMpPzAKb90IRlOKemYFN4n+omWJkSOM+T74zDBE4ABhUXQef7+YTkN7EaqQSdS4m+VGSR/8ZdOnm01a4wdNRjtROyZD0ynY+RRkYrR9wVpgN0ewruqsDsxAOMU8EGfSzrjR5KDRleK81u3/uK4HucQ3BpuYw46dbW/MwhCqUGNo+Z+AL3Res0/UE82ze//B7nkZCBS6xRcdnHiVij41qaNOGje5XtyzY5kAONxbhlCLWBR4qYH7zmaFhQxb1cfnsdGMqrqSDP+5o+/iHU2K2IfAjmaMkrHf4dXhYHgpclmueW2yErwZyy/IucA7W04pzDloqYpnMGVcYQSZp/XEbAs/C7NUNQeoNcHt5l7CNLvBv+eUCm/UvwpNRsqOGIrEN5WJZoWQtBIcqwPLjg/fieBneGe8aAWBl75mx07yh8mnGbs/237baKFgtjzBExvvtCVyy+j/cvX7mHbJ9Uh6m2xWvEK5vNWGhpnID4vNJKSsHC3KJaRfXHzOGEEueXcIkYAtSWwjO0OdsmC+ulnC+29uTqL00gMzTokd2F7qFbaStcYB50XVR+i9nS5eWpQw93BlwX7eHcp/zEnLQPXMl8kX7fLGCNIzuSaZuRBw24KDGwUXCNFfZAI4CJkSya9sqTx9V3KYgmFf4aAnCsdM5vJxlwL9NbByGdwVei/DRKTyYBj9uH59JcbLTjN/UOVdPfTcxzONDDpNZ0UQrUjSgNzjyo7NLOneo/xHimw84/jpyjuKMotXxFGGUtoYINqMap0Jr2II2YecQHPHKRij1kAMNUZkz5zh2qDjKAyf1P0jUt1ZA5fVEogfULjUMom5zAToyJeOPDdL0JsD44YqVTGNMhyHmJ4xGr5wrdb89piSvvZb2L4GQ+MfIMdKoKpDsf3aimkdDykrnSBp2ru4NyksCrYke6iaHLjhis9PVxd4EN0WUin4P4S8M/PIWw7hFfKYMpjdtK6Ou9E5csDno+duiGMpNSsMLR+NZC3/PlRZ0Vbk+GWAgLEbk0qqO2CAo1glP5xsrK9Jck31dY8L/C4/wX1DwFzIqviQD98XQBnPUwR+031JctaQdZwaVA8KWyC+tZ7uIyKYcXCycHVi3rje0PR8WzbdXvpTNtg4TojPrx/XTK6tiNHoUiApHURbRTYdRNAjyox+scNoiA315htVTyNuDCcQxQ/rmyjIdc6DUUCY2zJquVDJQ1QQ5ALI5lSu2Qz+pZ8jzKabfbCan5MwwqGhXVp7nVmdMXqEQTXkMcfFRZXxXjVNPl6TK+zuqhIuo09F6AtTlr3tkWQB8aaO0sFVaVl2eeWge6bsp6MmW3QswLoEY/9TwediGfCbbGRTVDUVfOxz7RCM0zOKXrI+4L21a0MU41O9aTgFggbKx8HWtjdUQOYh8s6W3KhTTsbvSLtRwIUQBPUF1PYaNZ9XY8X0xqYDdubyCN/DvhAEIRiVh9rtNrYoh3lhKEQ0pEomNIccxjXkQwQYmBZNhO66MP2l3vkEBt1SWCryyNuNaLf1WwB6vu1OVX+th+xM+DWXxrY/9ofO9KmR/y1kg2Ib3NUgr2R5sq7B4cywxeGmh9MEwEiWAY7t2mvgRC336R8zP3USAiy5+AMC9ev2cAtbC1/I2LKNm0P/ZNsrw6rv1J0rv4yFdf0LaPxdA8XS9LoVrBO01ndW+2q/ZwB8vRI/cGJUK3Gv7a54eMBw6xJtouetTin4hNVYQdkuYG7xmdFaGBbKIolexc3oY1zeixJMN9mv4TVDY8u0qzRT6xO0j3RMwUt7d3hMAoqWBdnW19uYzBV3x1TvTjx3rbrpO+e0stofFvkyxbCYk2kv70WQZH3VoXU28fPpv3w0ljFE0G5Xt/Lux8cPCl1pjZCMxwRJn16SnDlbvoPKfMRbJdKxA+Od8JWjghVCMXBAyIHjA+trIe8xk7iH4BdF2ygBb+1xlu+/3POAUgX1s5LEQ46JwqXn7nKVc2JgYiUa39ualaPZ9sBJ5+L9tL3RxxVWI/4sIQsU9yr5nRXfm7gzk0D5gVq5v1vqsefReNxhRy6FCBakLUdOLtDmmpolKSaJx4VvjMTA1HwROaX3w992kaJ8C25POg3JLHdIQuzYm/vct9CtMA5gNhD7xIQcpA1Geni0xto0mdUSRHzpaxLAFVoOdpFIGGPpjgrFd4dXKhXEcBcRsSjbjDg4xKsS/Bqo78WtcKIqABKhzvYylj5g5rtZ8evHXoPf1ufsnkXMrB8OJV5br2quTLgDNrV5qqBFJ9DT6ERjj7clFbEJFWRTKJtNttgVSgf4FpJ6Xxxq1NrLXBqH5CtZQJX3K647vQPNn2SmShkjYgGyG8c5YFU6b7NE0Txjgwo0k4GAjqpi8RAclSCTpdVMqXKNcsZ7rm+bKyzFZ07u6CAPi9UcoRpdnktnd33fc0Nd9VhmoAp1CoMnANRBNdlCebZSO1F4EVNW64K7rOiAcyfrS2d6Y8/KUO98O/GRBSTcXeHme8+txqYWMn/1l0tpUx1L3O4k8z7ywP0vU1I6FytfgCQ25ZQ1vn2stRW/qlD017DQlYfmVarKICU6MkP+WlxIHDHHI54KfYFoBhfeGm2g5NS7qg/jH/VWjKqlX7oDm2754Jbe06crz8nGrcCLwdPNbwK+CXnGIpuYHfa5I5JIFb2xaDaji990mxFZSacYma+WEFaH1ix1C5st5rrb6fMyEH9ElZ/2qa7MIAfV5OsUgPHSpR3xQoJ/qVbPnQ6nUKUfNiluCb25hRBDPD9X54KlPGqHy6zMjUb1ziiFsQ4T6KM19k2cCXArCxQS+AX+zzvdcXIk9NxGkKX9zmkhi3+pkoHE7DvkMEMj4InBdMDXQlOUmTcRGqaeSOPfgIXLSsNTnrgjg8U/6LPwytHavXtABMn0iOYPmv2mWmYYlUmZLkM2sv85FxKASuzQGJw1D7xedqZj9huS83uG67wkxEsfFkouJRgHAuPVcymFsIz3oXvvPDhdZkHNw4QmkMHaIB1mVdq79UHjg/RT2kbxMEmKZ6TejmnEiVNIJhk0ixgS/uHaP8Ut/NhBBe85HrFEyts154ZUK3HhH7d2nfTsRR0/7fhsXmIgbgUTncxHZCRKyojQg1IjZrQezDeUnfbX33RAtqcKLwE6VKazhgGQjJOAwRZ7VjrKDqO+fpCmll8h49Fjn+lT9jH/6SU7VV/U4flyksGFAeURm/5E/rhrMdWEMgoGY/hO7wtg47OFITL0zkHA3ToBM6S5vKSvSRcCvZiXh2X5p1fdBMgkY+Azygyw+xXhU5eLr2AsBmThayXvxRh5KA1jLj+wjodcFLKhHDnOe7A0W3zFjLFcgysjHTUiXbcLilp+mJrjL28+z0F1wDNy2QWuHn6SP+G+lrd8hnsfAVfZpK17kXtT+wV0yDj43xK7xQMG2uF57ytS0v4ZNmWtOpAirAfWDMFzAfPkgQiumToyLhw7bBFgsI2pH/aoqgyDkbOeLJReLBdfSj9D+mJQVPzi7CDCbSxuN1R6B4vaVVDBiSHEET7DDCbeYhL/OMWhEYcd01BwDtQ55TziQjerPyQdigYa12EbJgrPeLNkVjqMOlYDVGueAqq3K4KHmX9l83HvYAaIS62lX8WtvAg38+VWVlZrv0hWtd2LRZ5frzihJ57ydo7Lw0h4LumT6HzkYpGRnPmk8DgVh79sMZbCPILL/EX7GfMKExIptscfwa01WMYkRnD1F4+2G64i9OXrn5L4DSRTUOuE1RY562Lqu9zrTcidCjfNmiqy9lo99FfhuG/25dibg1TsVjdOwnZ5+igQvMiLgxGS1YUf9n/gg4OD0NwPn0PFoPuA7ymk9YXoQO/wCK/q21yg8nB4AuBzvobbrsXMvsTltO9+MF/bVp6BydufgsJQ3y+ZTwy1p7gwGY1B4FBaPN1PpAzhbIPxluk526LQBrAHuSqT5g+RW15yZSD3nqwEPiQ2IspTTDz+sHjasDSZEyhR1VOxD1P6zX6JJCt2YUZvdCZ4+A7A3MZ57fTdRH5jd7oBhMaMGCmJQzi63dd8f+4k1MEP745gVOldq0Y4Xu/WvICDJYQwTbHpS02yo8XWAqaCmXCgMDy4+Hqq8ndgbklfDl7CWQS7M7nubtesxzfevtfkbxJXrSzsTKKStxeArz5PjCBGrhZXqjuaCCE89vOtvNlN+lDiVXsqUohJ3NihPMqN+cRBuVO6wnRv6ncgFOIdVFpAsgfL3rTmfQCMBszFF6mzodxVfn/hx7khrPnhLIRZyY3jH0TRYD4NarN0gKFFvQV8rOd6Sf2fnhNotgI+PJp0l+ACPAyP+6EZLNr8FNzvJqjim5F5ml9GY3+tWgiPJP4rBcCCK/2nh8Gb0YAG7h71ASjrdLWc80qGDyq0pfqUYic7UtO8FdNMqvQguYQ6fWcKhSqZMUGxbBu2aFw54qZmAIUUWaPKHitkbEP2wPhP3oLiqLD6gDhSiN0hbxj1I244Ryj9cNKLpD6LexzjhUb1tAo+rWIVOOj5LkfLt4uX70DoeuS1/OBvN4t3R2+pId4YRh08g0J4U7yZZ4Ievm8yN6F8pTC3FoR/0XyG3yGIGSDDsmyOYZXkOf1Wvy3y7z5GDwtcRasrujG3IAWELgEOq+FNyhowzwYnLr0WwTvuzXVcJ5Okm7DpTW/TJiPzWBqzWqhwbTR/esssbDYY0Hx+Bdbt0LpTK1rRI2/5AilmvJJpUfo1BF0yj53+zGmWTLE6JALHclICgjXnTDWN4zadcvNNGD/TQPjAWv2/hZ7nRcG9QfHlPrM1HMk+Q9nG0FTjZMusT/WXmWBWQlHn16+mcVQ0/rxcDs2SowUJF5TrHclocbNncI2ibACwD1zA/LAYeAGvYwRmGYzxUCSOoHC3pbwRdaDWblLBf/Sfm11RrCvLqFMO/efKMhobfJZi4wedsNJj7A/L3tyT9OY7HRMBUjoF0/CfnSSnAe0Da4Tvq/rN2YwwBE2l+RISEufVGSlDXPKtCHrSvFpuz9FwLX0Rf3wBm7dPph7ZbghlDDhl4xrOGqELBb94sLQ+Wowt3MCdBQ5myX4aCoQsAY3Tap9rpFZ7qCAJOSBWWYmmoXyWXGYaG1xXCQrYhne88AMJZf1HXndgl1MqRTEkkFovAQKxD8MmJNgnofVGEvsbNuilbCffsr5P78XS8SuBOKo/fMiZANtqD/PAtkDRxOyXs/Pe5kAurO2VacMUXXd+sW6EopL0tXrCFiRz5DwFVMG1H5oDkgN+NL8khZG4I0ROoy/A1VkDx+0XQof/TtbjXe0nP+XFj5CqQS1KbmsjsLOzMc82tWHO77iH3cG6uZuRyZB3rPzgJRtheBjT647nklA+lJoMgtkLHj0t0ZTzHq1OoAQ82pJ7jhdkv2iLloJINhYIXfN/Z2EJ1lTVXbxgY4RJfAWnloBQ9TB+BnbY/WaJRgDJs3hGpiki2HeDH3/LeTnz1lKxslJeBUQSDNQhuzHvsVqYYhyiurEf8/lewYwwNHkzMCQnN1R/DC+6SH09lzF+lYp4yNM8hCJi1xZLD3DvwrxAzDYPuGOanNa1nk93thagYfPlLo8y+IixOB7RcKVggN4g8PRe84YKRaeXqxXjdmp6eNBIGqA1sXraJ53ZU62PCcGBiltWfiOUloVgMoqFa2rKWlyr4kCVeDBnlloh6tLX5iHema9/cm7+2QQ+yM9pdprV6wBH/CRQUqRSU+2q9BWEtpacMc3tUEj4Yf0rzepgXsZFp3GKkFsH72aSie4VeDDDsipYfwkEeocd9t0Jnn+AHmghl9sCjPugT18FbTrnHTNxkzTZRgDASCSAE/IcDoT/pNpkX/kcvNhOIGccrd/xCKN0t/VMR3pqFcR8hwRAr9QXkODN5CdEUPifiQHwkVpigd+XVAImLGUwokaM/EtovF2Q48ZhscUZGO4Z+TSKhd+XE5QepI620y2MV+hbeVdQxeqv4GUp4TIeq8XzQUjgjhvo3EwSO1F9K2YuNp3S+BVCJb5aMLjteWBug5LtAvXsmZyv/tnCRNsDu+g3KD6oaVIn8DecNbh6HvA6qHHgtC2FDb3fGFQpObzfCsMK+wyvJYFJJdMkSEWthXi7CHxCU41Ie+tgGOX4cMs6ChwYik+Ge+miLivgeW/fu+uLayqJZBjNoHfqL/5e9P8/q43ixaZU9TmdMOb+fDgZsgHHOp8GEr4pgpPH1x1BhOqR1y4RlQbc5nQ8He+xkOmnySVKQbl0S6lCxqjFomIGn6C7gczK58xUyfHCSuLhjc/BoSW9LuUUZVSl9LDrhJiBGsn6luUoeQgE7I192rZfFlj96E279qvmG4Ja5ksXSwch21EoUi72/c4gCZZo5izTLnOe5W9N4MxCpN6kAK2yvw9JKL+oyotEj47ggeo+Y8jpnbI5RhPdrzl8ny0Qw7ZQCtwnM8a25bykT3xbBAsxxCeM0N9MEOeKcoUckq0TGkoOUmRDljwqWlXaRX8Egq1/4ryAAJzMUIKytXJVbn2hV8/FmV3K2Z5GbhY2SRNyF/WHZqO4hAvZAUKJXvmOQJafd12q8+QJRt+0MrQXNt+PEFMPCxSX9QRXq/jTZKjiYcniyukxtpoj37SZlZyLKkis0VHUTLktstJOHSuUbEi2vhN1M4Fg7RQdOrKI1I30G+BdJp+s51nKIrvU83AqpeCLHoEEeUmj7lZrB4fnkRT5BmhpZ/hktJr9Wv6Fnn+Rg8xQEm/ispDrRvbu6574/tl2Y+VZnWdNei2GuQngMA0rYzhux5VTVaM/AmcnFDrKeZYLyIoEZkyFkq0Qnyy+6mINcTzHbVTU0EqmeHhAz8gp7ieF9W70ijqurFQXdUiwAljfn7feWlQL4TrgkpZ68xdk9VbYY4A1B8aAri6jTA2FbeEQnr9rEU19ikhee87rGLOaEuHP2MXH12n1LBE6Kf92FJmedm0CXh97q4eGXQOxs5tkaYI8lBlKPtt3p95XJ6cNZWuKq1m4Dl1oDw/J4CTlbCiSVJEDd9jp/dIZwG0is4EUVCLF6HlPPDUa7IoMenxyIvqnzfJq1FzEarDzL5OIE7lpPAGD77MIvNAhyczC4YNztpxRb2ni6xCCSFF+sVWfxaF2wWYt+BT9c/W0LELzM2sgFmJu0dloEn6qPklbsGsz+pWglccV/11qf35G/y2xNd8tAWEDasMmmi6kcxujVug5zAp0TXUYkJ1hn//1XF9ihWX9tqVXZ1N7UD+/toyOH3XRlzZ6rhp4hajaHSfjUkmESzg60O7VXbURpRxamaHTXyXp/6YHZ5YoyNlizC7F0nr/JXp/a2iHxbTk3WY/S6PP9+v5Yu73FBiL9Ww0PWD45/bM54z8nTacspLi2MkpJmEshCwmfWnl3QYQhu5XTD3sMQXgc0Nu9kpebRJzpIFYg01I2BH26tQ3rVt0MTl3aX+VhjYqTHAfXdad1jQpnPwx7OEwrUPx7SBPU/ss2czGnAvNGTDJ86TqOgHWykAyGa+pmTzRhiJkDOfVH0e1crHOPtQ1kLJm6/zjN9enr43XKWuaRaxp4W++k35xLEF89Y3V4j9VV2jjAQTB/+0jjewlp4sdic7Skv8rtKrN/vskgny7XElmL+GxP6IANMzGhfCljgoSh/BmaWRrIrcgL6oe+Z69A5wZihDSXwgPlK/4m9y0a3YbhnEkmTGb17oZsBhhWZUEyplqfgX8gwokuEpxzu9cteQgn9dN6kAQso7jClzWIN/9ZGEHid/qvOyg+wwiix6qG3vmqmbU4pLhC5zw2UtOiYErw1Nq4c12MW8CI9IaeVS3PG3DFq6zgpZpj8+TdeRhvtXo7G8hm8eSACt3nejXFT73Z+XTBKrsSG1nn2KFv3hCh0atSMXT6wDojQSjIrrgmVAYjrXFM6ZuyHWnygLcDFk4gqavM08/ANF2bmgTpS4Ipf1xAQFsyEX3c74Oq7zqPtBdmWVWmJOsSdb8ca+3xXucDRnp5feY24s06gO8D1hk7Ldx0vN17p83LFC/5E2CXY/hwEQ4OjZAon8wgGTlU7nrwvAip8j9cjPO62msylWZFcWSjN4b+vvMIaF64IwJEWXk32TTUko7ymmraUzPMXqvMUJ7emXPh0AX2IPNNEfLt68oYLjeQyoETs0mukjtUym6L/yU/82nBsVGoGeZFqOnwTel9KZEBa5FNELAPwXXVU+0gGV3KbYF2SHwJyVKIspCMZBcnBfKic/9p85zE4tLBXx0V3v+rCx2rT46yHfv6xN+PyQTyMLxg4P9lYHepETo+LVbO+M6KEWsDwwNfcm5iGfeahImH07r27X79yBnn4ZABvMXXVTdtldHZ8rj7aJ6K2cmK2cT10O23uj7zQSwnoMpa+9S5nqm2UqKwYNki0PdPzfY5j1QcdL/PgpYE4rK+/576DkgONXUNRNq04oP5DbrYBnCgEZ4XxVyO0jxWuDzECeCyyzCCvEqjQt/YnLMutK7viUnTJQnu/NZHgC2ZVyvjdU/r/1DUw2hJ9giAFbyu3vzkeIANb86njCFPOTZ4iCnQPz4IT6zUC6LEKwW6fj5V5pjZ6MdorGZb+YtCx21SGM9d0GDLaE0FnoiEHpku7YKKGTnN/vfz/LeO/BF4Z9yST5aETCrO+gEEXet9sNXHj4O4GT6aaCuLNffqJS2h+TN9qao752TW2nIQGtiuJRnaFcV5nyklG3dVHFYpM6CoN/Z4tL2tnQ5O7mrv/S6Sq+b9bRDfasH3GUUxMAR55LzQg/fSFSaEr3V2t3i2Emw8rYukvQEtSm0dKdxvtfciReo0emwh+ZlQM2WIHde7eFi5y5wFz2Ubbyy/ZlvLGeKGawOZh9yVkzzSTSE17LgOuprzteklA1wl3KDB96KNl+pgzL6Rr643lII53Cejf57OpoYgJxIyZ30M2a30k22m+UOEyKqxVB/RgYJRpl2XPOb8LfxnMZEbdNNJmuf6V9VEhNBw3gmI4B13SQ9zYhjDpRRafnYYGs4UIV1ARYJCDZLvzxmq2dZ2LcSzW4y6nYOirZfot3G37076mKR3gNhstR6FLiNRfMLyzyj2UrHsjqPF4/NUl4aoo1MaH+O+hbuVArsdnyAvTHcuO1NQ14bcoJ2qNHVeuKo8+5L9gyWeqJJFJAHG9zxpVww7bEMIlS07IvsIt0SXN4mh5sptIru0VqB2kpdg2S6vqECSo9nMfYRPuuOat+IWlzOB348CxtFJbEgoC3xwiCu7+Xmcf60MR2BZ92sMRxs3uf8aAOOr25Dvp9qQqJPZMUSZGMSYsTq1SFmprikrj4RuRnfpzGZc6VnA1hn48hyLsC3JIUMJa9G6c9Me7y/XmNgj3yygOpfh28huxv6zwuA6xpslrO7T0GJZSL7YOywlD5ObfhxiXdxdpJ34Dmy7HyvaqaM55a0F52vqmp3QIfOH6mr1HUf0l8AHfXnvf6T1msZnaQBjAUkyXF0CNcLJe+1WciAt48Ytp4CIxtjMTeh/g6h8lMbQeFx9pT/97kQadQz7CarRj9hol4rD85M58GrqgOogAfviFpF5CrpPPno9tIILduQNQYX+8wBdPwPUq/4+1nDdVa0jTUatAsoqaqx1/LHq6If6c4uJG/yOqVo1RytqbFuMxrxnSIjawGJVXKj8T2W0tJNLUpJDbwTMx1cPNH7BvVhG62P9qDobVaMENSkxopNQ+U+VSxJjnBjrQcCfKBl0IiIme2s26TLAT+6F0NVdNPNoQjRck2wVkP6A6f3Ee9Ui+mlNn9sqcz/zNt2kYII4hatmki3SPJvSPcBDNF7zQODTtL8e1h7yD6RFG1r3RJ7BAt05hyfZ5R7T/iNqPLP2h4zyVrKInfuy7AYROR/8ilMy5KTmKys2mg/inS8CdVSRlEUD6voaRYqrGXPUcRv1Fabw+rokqOwWVYVwX7xdSCAaixZy+9MWIkgIHI/oSPrrQE6fSvbFh+sr03Qi+RuKOh3tdJED0akfQUOdKy97wFa0tlVHAo4JOevlxL59UWAftTdiA4tVhLzFt6vrSFO6aXY4pky7QZ++s/mm33ngvPyrQZcWR06TiDYU/TWjqFY0yfXr3sXVO9PkeYNgFlUrZn/QD+5pVBm/mNdDojs5zeMhQMemkN8X0vvPgg1SwAchhADAg0cxt2ihU2pb9UYvjgjfs+xJUqvu6f1QmA+XvPOF4nforPN2Dkf4czZo6xi7laXXSqFX6gfr0PC1LaiJPXTNB6GbKX4GidRVhqEUb1kGgV6pfjIfKRiJ00l8OYdmOYuZYDXoMDGHoIJSjNyfWbaM8fM1SPORmTrOk08m0g4VnNV6lDXIjMOa8bb+s2tTIVz8LFQb3wsu+3rXOgOup5KHRszmYol0wIPZU6VP7iYm/L5xvEYsEQXOF5481HtyvgG53oM1hnjS2cVgoytMVWTt67gmEe1LrqDVeLUz8xeFN8wxyhbInhKmeX+vC2Va3t6EZhcMiWirVrj7kaXCiVYyRmSpngsTyHhOMAvYjoP4B08ArC/kQV7oyVhrvx6gURakp04TLdhEaVCTAfKQdvpribMpJfmns2qNydeLfrCfEJUaLXPyXOWTDZkFOi2oyEm5QSbkIjM8kbVbe0u+0gS6zUxpirQ10CgJ+EA5NvTA+0ntOi5XXTBkIpKQRsjjA5ZuDCuekkxGjr+ZWv/7R8TAWLKCwcRFuqF8vXmKVVnDSDE7mmnLH4ntcC6GvZxXGjNnUth8Oz8AdvKsQxPZh9B8Gpu4Fxq9Dbijl+Htf5QA4ypFUV2O8cnkPRh1Z2bLQqT2WVLTR9KhPeEFCQozvKAbxXsybOwKQURPK7rophBs+azx2dJLmggHVh7ltC1ZtQ352MprjWdOLu+atWnlK0vNgVGrjGs9anp3SfFILPBH469xer83LZcPkycoF6fXnmsosrjtw8Agf5/xqCoMMbnicYn8S60gzfOlBg/Fsndq8ArACxKCay5u5NhneiyEg110ZYcDbzr+4XPTEYEBaE0fylSeKuHnWc56ynsFumyV4v+E7kUzI3KJYXPTgzkIZekSUm7FywPDnxlrOLcUB/yioKiyf0iEdrIC7EOr3jhWqY7iPkBt3MPDY6TVmY7JA3O4y4QWjxWEtJlcRjhoUyhMYEDfVQkx3mWfh3gXXSSqQchR0sQvsvYcLKdZZdqMVW6ohr7y8jk7FZ4yXscHD/cH6/c5FGNp0vqiQiRwdoQhyephPHJbpZw4uc/Ep6D1OHLf9A6qze7+Uv1Dcq7n0FuX8eQP2ifs7rE+nhNfh6BWNgFSlROsTWEl6hp4jt4c5OfGOFmQ2CGRzgdcOWXReqKToS+GKF8WjzRrvjiYFF3I4C3bjXfSaARdLZwpMhw2XYnBp4TV+tWJC0F+AsputaU6P79q6MqRtu1r+utKweLMMtDAn1m4nVUms5AIdEk/xFuTTtP61+AT5q06atLpRFBmvK9SM9JfiR5Lobf98NGYs8ml3uegj/hTyNJKIH8dUMaYdGbHfUbQB9LIg8K63Zy5eWRaVClmNMGrRnQ9GfvUarBr9q63nfJ9Uwre3JICrh4UmbpkEQ3FoARXVvKsXF8zg+MpRGPAgw8IlOrjeC9HsCZ289GC1SLRQNhS0YXxIV2RA2aS1wkVvaovbV+O4gsSsMeWax9LDOpY5L+N3w9plNjsmIdszWkQzEaggNUdKJz9QCQeaXwo1nSFvrzHUBqvwr/5nP8bp7hASsJXtW0JnHUN7jGL9Qt52i0teERmi1YBr8jW+vTppCpWhuwGJX2S8hZs1BUdTLj0KS5e1ixiHw+BM7DhgE3I0TDeaYjHcfifNxaPeRp/7ReOWZeo0PtdALJCkXJqpoxzX7yDCcfWPaufEckNqfB3iE6zwUR+G7hcrl3CQGsSlaDWPpmvWSulvnnDrynaac701QoSYz9MvERj5Ucn6GA7NWMP03trTfpUE6noyzNe5QHlN4uWIA1GXAhutV7pgua8ePyxjzrTTx7Nz920rfE0eK9eA0f5T3SjbHCgIz3jw5CU+FwEWGTqc1nkqeILR072Zdo0eAeR8zE57t1z0vuyLLcVjEJWTJsSbqbSjb5BtEJaANd3+il7Yayg7loJBTEJW3V8M4DAzSv2AeWeSBvKYosGNKj4I+UcheL7zSH9PCXaOnGcZcGMf2KanTwpp4QItLvsV8LSwyoMXcuVSUZ4DTjyxMpjDdIfx7gAyqC3ekrqhE55N7oUrfVr5SalJIwPHKd5wN9NwQ+m5Cdw4sB5fpdhndXPYSF1U48eSDN00cECtZUqXxrb5WlGFyjFL+mdJCfr0zIEXDvs0wEQ9PfMguP/15D+RGpfbiu4Ig8t1tdxiZV9TymQ/VP87XS6prJ3+Le1QzvQArMrQU53JQlXUFeNBVxQRbRRdjPw4mUXecwZmuhTJWS2t2rVUAt1UqplCFSWKQ00RT28JFlB9emt5/Vl3+a0WBfMBGKOM1WqJLtjBNiH9QJ22iEReSWke6GMv3totkdtS5hazWzcTawkxyqDhpvBNe4+HtrhAtYKYCoRd57nXPxtXNs51gDDOaIZFNyODwN4F04g6Tw5zcPb9/Po64DMylt/260Ovsd/0dMx07dP4/2pbPegJF4U8I16NiSgvHGmfQ7x9k4Ffdwxe7NDBUEZ+yxZJqAVi5570rGuhmpLyBtsCFLej0b9TbCXjuYBMvd9nS5lIpJt+20BbyWs6PxwovpR+sCB3ZMwxZJ4NlzFkphm7K9EVGRo70mQrDUtVeW2ieXnEHFMZeeueFxccR89u0qDLfmGr1eS3LiiW015xNoU4+9Pnj6hIcWNcfN7ZKTv7UJjuS40PS5c5/OYoH9DKZewecsVzhn+k7sCtLI+WtU5BfGKktUs43MnlqG2VSvbcMi+W1qBL+yOymNatFYD0Wq9ERG5L+RIY/cKO1uVlAMqCiycqiYozoPn1oPrWWKq21vXO1+ZCdC4VVQoE6EVkuX/DstJR4nrbgXA9M5uYK3+DlCEPrEc/1MHLkrPR2icMzSoxyAZpUJ0aZttHi5k/2vgNb7nkfaWZkLGrHFT7lJ9VrF8OGW+LovVdOcm8QhygR1XuZzxbhVITAod6e2yynLMQUc6JyRFQpoFGObP3ZlQF1TZ8Lk38hpiFZ0FEh65mw0uzWetPSYYr89802Kkl5H+IG49F0h+N6oHQMwROK0vuRHVEZZyakndBlaPqx8eWt+jzbmM7iiJVsyL7rMzND2fZGIM4G/2OsLSKdMrHEefz7mKiKQg0Nq7LLygEbyC5IOQ8dTVUZtRF1eQVFyJ1jEGU0jcE8oqmxk1TEoyVITzxfxywLITJT3DuJytUaxV8x7rHRlc49n3VP7RYv+uw43v2pVsH3xZqdI4KehpZHZ1fUTgpD/PjR2DWYCiRFSxZUPmaRlOPagKBtoVVK3abzG2EwF+MOIy/iu9k9W4vEZ4zDDUfMF/PibJfzpEjXCUyEK1QPub3BwNDzK19eV+C2NojIw62fg595rkMPsTpnHEPtM13DtdCUjYTdpYTSUeT1J+oweq+sDlHk4bKGjoPLN3HamWKrTatUhnOr1BZIgIPYuby326ExU1+5mEnlu/+byDE4QMgV6zN/PdNDqp7PHT9PjGm0KrBMZoVVP+KYyGu17uRpRfV+O501/7QiQKc63PbeEo++l1aLMWjgUOh7wcTy/8EE9cuG8UQR4DLrpIVRoAduHDNZwWe3jvAA/l/bxLxN/u3+UNKWeDaqjVivUMtC6cyL5AQyIbwPJbHiOBz6APBpQ0OkQ3NB3B/1JAifJEQWOkXDSLYAvPtreme1usgmA034kzu56T9uHw1UCu1S64BEY1jLebA+Ev5Fl97JVxJckQKlKmq8c6QAXAi8jMV4pBpnxp0bta1XNY/B3DZY3+2Z7ih7tK2hIMPLMsCfZjV4MATeCpwyAc1yJhcIsHyKihBo+snoxYuo+e8i9Tb5Fr4SpUt5Mhq8MFyMXcV9MMP9KyHmq8Up0czGQzgL14wARbBFkhkD3Cv3UgaYsZhFqf+TehhczalWxT/9Z+zd+QHYa0thw9RHrJcvEF8Hwulu2DPzKUdMwMbQs5FmnUo60qb/f1OrEeW9BtyxMD727g3yG19v1Sou1TbLuT2z928qwPGfqKIkJAtDzMdbxnHidDtEm3tPgKJitSFvhS9fay6rNbku/ax3qyfTIkxRP2X1cmYgh/tIcGI+ra1eTSgt0DmZsRqojbweiGYZYR1JYWg0vdWLiivdEu/WBk0wrQn/1aPHLsqa8YnmhRibz7vCxfPRHROgaha+VljTxmDI71dZhLqOYHDHLFYHJWiAg0efeiy6cSRhl9pZwLZLX3v6Hwd1KUJJnd1GrRn5HarRp9vkGbT5EOAT0X/hxfVtCvia6mpzVWQblJU6oIvXeYFm6WbkqSppW+pvMYjnrzzgCAOx6b8EXYWHj509pnd8qDRLoFLjJuJDILZEPtKKQMsIWwARkwW4Kw61cSrZzIc0tlDW1BqSn+G7w9qmxgMfJ6Gtmco4ZZBwbY4buJsRDBemLbbVNxp2FiCrLQa5qSzmJbM9OigiLto6UrKcWp7P4HORy7fQeZPtfZmGbNkvEIBvIQjbJMV1TrvWf2ouXaDvsfil9ijczMvcJ2XQ5VjFSDHNZMEKekzzLyoZY+GLl9iqaPAcOtfJzpPOgujZdICV3OiP87YQQ3s5LuvLcKAw5+sHiZLqKo2PuTSa/j0zvGWyrSxwhf9fweSfzB1I54DLQn3T/scGYYEkZlhnhqxww0FUhoWQVsqNvBhctMnIaXlF+DhQz5ZLgDRqulweTwzySbKwsa3HC+sNpOt6lngS5c/pwa2Ypj1wngIhR5Bee9jmILGA8qiiGqItvMeeinVr5J3LBv0pwp4LIw6ZeIdxbdiVFLBJS3OAoF49FQqqvXFSnXUqdHmWR92VXbwzfhEhm78J1G/9xqWD6AZ8fX3hhNkGW9K4T70y1KspK7Yr0x85x54GcTYnEAAVB0xklTch1F5Ncu7tTp5tOn0S0hZ+wJEzhrBcaP6uZ9YxXH9zMQzi9WNzRFKa6dGOIM1hY2fX+TCLoWN9FSvRFdG99AE3Z3h7rBefYyM4+24FJxO0JtiRrVKrP/vhP3knRRifRmgBqpFacD0HIqOix4N2njIP8lVcRXvoOCYu6i8yJ921/N2yCj46aI19hxUkSmPcnS0czgDvKJd+xpmZ2YfpxzM1bge0tVYhjSbLQSb079WZAexOxQG/4Q1/UgR0hIBEdaa/uVwGOiDInKho/PxEJkV27SIiJIWOZ8fvW/soQA+WmEJ2wlMXDeuTgyos3Bs5yJhgp/iojx2E5GkSbTOKRlHLxWBfy/lpoKrWqq7Njv+xcO1i1Mck2T90hQ5xa9NVR010+ml7H/lWVGahs0wB+WSDmpxsbgBLRAaPNfI6MwUiYEAwg1ggvzGuvksRS8qwI9hzw1JextWhR11BtcCHFoyPKe5aIP4adfmCty6tDhXi60pmhzUV0siMpeDSJEVxwVdYPQsk6f+0JrOZFpvrSzEXqh4To+WuFShHyVF7JCcYfG8LD3UWNSUlKdLN+b+hEuyqXt4wg5BZ4kv7ZvFfiiyVaTV0OL7IrYhGo+Dry4pEfYMg097IcbiMde9n85QYQdIcKBxC/smhkrlMAl0hqO5/HDnbRolMT31WYGvBMi7P1K+uUCxH70Fki305Z4NdUEOzMKUXYajmWD+NCz2zdnF2GG4+8/7vNM80lfCZD12o0qKr830uSwNihck2oC8p4zlCWRPF3G0AgokUdp04VJUh+QncQjsKo+EpFfEolRDQ970Zg0IiYD9bbKGT+qsf+7LM82KWeH9/z6IiiA6LgQjwgF2P1faZ2xCNed8fM1ZKQsfnzcqFbhF510gAtud89WxqmHI0QJCE+4P7blc+FnfQHEt78N4sP155+yq1bOCIzXJVh4sag0KAzvjGdAlLHM7cuItuOVKYHB0CIKzfczMqUjJXrXesla0AgX3J6193oNvAAibYwcPZMdV0b7R2BqZ6R+Un1RzTlM2+pFilf1VF0K2gSp9exSbDTGbTzhjotP8wJ8gpzWjLCjfNWjzq3sx/yQnXIPADIXBNuGEsM/5vS5aqJcpLLgY3573R0uE34ySebRVAjPljUS9kJtNykBkEXebHxtECK8dR1gvuMXhrSr0oaJJbMw7uwcxmy83VzKm/Uc9y2BCSNieuDhB/e6U5Km3Lu+oJbTUP1FKDWUsMYzu4XUn28bFAxdsUrK1OQJ5ADXyCApf229/5vwFVLW2hihXWJybSE6qfdz/ZziQLGxQzJ084qQUlVk0fIPSoEQ7L1OlYeM4HRyt/193r22jMrvPUDPWByhfQXmv4OLOHLjb5Mv3RMnDmXJGnr6MUNFHwfTdiLNtIIIsx3l3TmzZ9AI4eSH4ZASjSaUHmwNnvlvY+GDmsXBX2kiVKuWTDtcAI5OM22T3b08X1oB/pgWvVIfYt2F+HLWRRTxXTMsoETIwXmPfFMvWAPdB3KRlqo2nkdcbSbdzGmnAJwmnJG+PxsWV/HX52TmlMbpY9Ea9jEPPHiQbBKIE+8uvPeJXUi6uO+GFoaktuyAxfkThN5nkyuoWypP+aChO2w8cCHBNOHl0leg7S4B9JJtlAZixZTyq6Tl4FMrvSZE/VWNQIXiNpmFQtH8dPgY49YiG3SELhDsCYP+KHdBXJht331Z0ERSM62A+tKjLpqV4DMKcC2X4KUTju0/1u87e7YVNSrtHJKye3+v6pbqbDefJ5pnJUjmx4m3vBj+hDpR3wIm/zQXtAXHN3hhhBjJgq+K6KE/u4vuuDeIurVDbhuQbIH4Zwz3HPyYdv+XrmqGpG4TZpr4AHLuQoA6JvZsQltK34U6Wbb6xMMQ7ZYBdMdgklhJ5j7LjjovRl2OACjakx421h9SZCRuHbuLDOsmBxvZrGxjvzOJLNfTIdaWRpilTtn7EIYTDc/KnAgiG10QMLQWvOtpQePIHQrW+SI0lgusGHot8uHPq//+s5VotKLD+0Tj3mOwMKZvsKTlES45fBvD4mK7e5eqk+Iwn9o/T8Enl5tJxeAUC2/KTUlIi2Rj1WMG8FzxiYUEAQ+trVJrCqe7vNnOJHkQMWNSH/hDR6J1vyki4Fd+ejmMTNyLX/JZ/jY3yQ65+9eS25QDzlLdpCaOhEcwbjU9WWwxl/oS8xaBy4DVhYt/kESi2ueJtLv3SVyiQgBYlfzwDy7wuEP2DjMjhmhzZ6/ssTBscN70RsO8X8Qg9DobFZ2Fm2TMltp/ZLWg3EDfyRZe/OygavE1XDSf31DKERasP4Lr2L93KfmBkIGcZXS13vcYnAfJIderD+nfdoRlrXv/L0h+X/Vt6ze52yNzzNL1vvp+tkc9H1P1cJkiGBxB2KR06dWBDA2kmD+JDWMCfm+MgGT7/+OwD2Z4fFbHgDlG5WruQOmmqUJtoMIj6S819/ZG3iyBbdpYLBBEnOoBFXXpw=
`pragma protect end_data_block
`pragma protect digest_block
d968ef716ab8fd82c192aa9efc4d3b8687c811ac3b2a3c28f14dede844eb4859
`pragma protect end_digest_block
`pragma protect end_protected
