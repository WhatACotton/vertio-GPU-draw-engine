`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
FRancKIkG8HM0SJ6lRYHwhD4HL4tECQ+XPkSxkZeePMouHCnYucQB8VrRePgOacmTglqwLhPHNaIAVQ1nf9j/PdLWU+3sjysyFPvBeVULkXu8YRu9NFssq2bGgUFpy0w9rXTggYKaOD9ZJq80gzaYXXxMvtbZFSHE3lMw2fpsPCc8gr3p/jMRbi5KoBEBc2iTTORv1uhNhLO68RJ4xUw4uf769xjBquSuJ1tk7/5vPYTH54WcHJf9ryi5eXYwXJ1c/+h0Shu68Uar7A8623RUAcrSskJEqzK61QtGCUSTy6CxKPENFBT2oqVJWk3JEtFAPmt+k3Tjq+o0E/ClhWgr9CvxLC5pmvnzJn51IwmTEvthRZZJTtTFNJT1iLyYmpGZ+OczsUXSfZIdZ0BymdEIrp6Op4ns/Lf/tcjzH8RunBhlXNh3mWV1zLWZajAQ4HiYFs7NshFOF/0sGXFhSAXQwhg5cUkYvb8dhFXVUVDoXbtfYThzjV1x8FFQ68NP19hYec24K7FFNFfsTAGJieBbVCTmOhh/CbtV61qoNEhROLOdYCDFYUH0hrXhQqHyl39ZQZpsycjRQyi/w1zP0jRsjeLx8OtSvrLTS2iR6AoW5YaDt8FXTRS+aTv6XgzcrR5TobllMNXU+xxHzMG6ZtpYmkax9FfdXmaedgoJl/MH2RMDCl7aTM5lUPcsV+Wc8IADgeLDpv7VUivTl4vESphmR1vLdMw4ogzipT+rbQvSVa1fdmzLRzhkKYBSNPIcOnSJIv5SNBmR9OhXd+FQEBCZJ2Osw1KF0m/enCLjXKRTMhPLiSQMQlEDw6jmEQQShcp4I1M9Nc3XrHUrODfVGge3xfgpe3TVcEDcE68jVrIYrzZUHEoBWLToWV9s8gzqr5BnDpsw9gOUyAuTgqtZqPWqJpSSY8hlEaa8LyA3jpfrEKj1VXT5yyZ1FF8dZ4RnG/Z0GURwle/rWf5bStXOF8ZPAUkFWNkc3Nru/9bpfnu0ramXmUo1S7J9N/KehbHm83WWLZFToj3Wkudj2OtEKRDQ3DKFrbXvo50re+N5XTh5uITFjvSSVT8xM75eQS5NFVGRqr2wv3dwKncq1MrVNIGp+ji4N4qR2XMblvCfRWahQ69UVdWN5hZrBBswI2Z6AoshuEL8YRrr1lFy3utIXhVoF6vdOeUNoaTdFcqjjOdJR59SuJEM+sXq+vwTaP31zHwSX8wsTUxwdbwaVhp5F+cGaWoCnCykv7GX+qgVPTAiocP/+un9KcjsD4lsAIG1BKYlpM96yxleemtQRLDX0yQYIVBmKBxKPtpGsR+ga38+CxDlYSuHEQr5kuCxPeu/HIWDEwLOUAbypfa7fOzD8JHpcEg1TMc42pNg8dz2JGv3VhF3GT3hKolFjJPHjWmCWFnNkM6lt4ZhXU5xAG0rfBwEoYdpxN0VSQGpJfJfynaK0khhP3dsN1n4gKiqUzJDktXX82EAPHzBpq6MlOuinMkmY2jYEtOrRQTHXx3Ff5qFTdTbHi6zTTkCsuaOxVGB/IZchNyowoJ/+k5p0Tn5sD2mZ80CLn7JLaT3n6DObC1q95G3Ua4hkiNjLS+9jXVS4oAqnXDLQXR+NiCngpxWrHdLzcZpUxP/Jzd4nlM+68B9YOtC2TmoUuFcYG0jpWYl561g/qsP27RnxN0g45qyG/1EMPsFX+dGE5eTM34Rz7P7BNFg3d7FFgt5nxqA5gvhfwm6+7Wvgn7WVLjd0FQQmvI5GkK9jwamP51mpK7nSsVSLqIwFfa49Y5aW24Raz/nx+Ctdj+r9BzQKah6rW2vw9socpvFPYntHs/RzaTjjq1c0qUhqAv2dDLUJYC6ItcBRRS91a6O2hrJIQ99FuExk0B1x7w7jAIAR9IUZvYBEdwt21rXwgI5XCKI5Yj35XSv7bnXPB+tNzfYqWMBxTBylbJOmON9jFt07WnpMH/zlmTcKsEDrUKITohgFD/wxp54lmlm7j3+pWnEE9c8CRh76vr8VlW6VSCnjoUmHSUU9QZMNuL1INgAGp4aa4mPs3Qz/CFt70ByIYJ0wvGIFtp6ADGBfyngv0Vkf2YgjL0INOSR9PniL4W5GHat5bFHYSehFoOkEnVx3lsEV9h0LvHxMLS/WKpUeAX+sg3FN0vd8Jwdv0a42X0nEUY0aoxD8VYaHP9LD7Lnh2dmBIv2uEBXt7VpmJbYwe7nAOgD86W6cpftjVT1k7PwbUq7gSEw/wWgfumV4RzBTvipL3pncMXSSGeLhyQADryio4J1az77jjrPrvkKT6dNi98Pts93eVWEItqPOTXDXkjKi00fqR3lH6U2l3gVPhbGYxCJd2VeA0MwHxPGxI6eFKWXq46l//5fpWSi+Y+RZ8fqouW+32CCTuZ020jGVkzoOK4TzOqlXnxGKQ4b/GfoOhBjtc8hJJBBffhkNY4d35qoRYbcAiIVN8xmSkY43pluWK8w7J21czFrCd9cGX9tu+0AO2l3pzvHWfI9f14iI8UtHKKhl1z0Xgf9W1PzEwwCB0uLALOy+sk4mtWQWnnQP660bEXdALjjXy+mXMrQTNUm4SW2+6WQCh04dy6xvwg4jUPBBxBRAevMJCxMY+YjIzjrEDgI995+JOhl9bLHxFUCA9lgky1QgmM/2CRSmsq/y2VjR2jETsMh7kbD6fR1yox+pzWJRU7xWvaiLCk/n0rc+5SkvIj/m9uHDcIW06HJaM+cALGosIZpQC5Iie71+XAkfJgwNSVFJjpyKZMu1PCXbylcK6/DWZCNqONT2o+fERuJFKRAyRZHXRVyWTxcwzm4nsaOoytyLjsi+qejOYT+8XZBKsG6ZeSKQ1ALT4F/nv+9MKMTjcaNzOYds3b61Q65HNrx+htw0dsVpLFlJDhYxI6MeGzY3xzKch/ivKLs8etXj0c8lnBD+OpjwmpkPxvlRdFXaDk8nhHyyqNYIsLiD32NWKe4HXX7t63lt63id0ufN2t1ZiOOBcrUJ1RU7FwWSK8u+nntHG1cu76Cb2LJ+HGabP+ZhVygeKWzjc0s19Is6i7tHGvr7sRNnEykowIbYaq8Na9YUGrvfYXesLCglpwVVNHe0vL5d2Gl6XRFjyffyQSsgP/KCgi5/S504AgAhqz/Zr+/wnCrQ/x2NoY8pablox1Gm/pNSSNg7whHLHJWOMGKZwCno6jo6OzjtRk40hSY3MeBDNnPknz4lbE25GOIHWsfvPE76fq8d0OlOoCccX8dHWo2MHcKl5xNDRdWopZcs74ig7jVfgq4SK+KgkzbZpFPZak7Pfs/uNTk3Cj5JVrQeK3lI97RXp3CeIxHpZmygr1gFuGAJxlo8hqXtlMC4OoesHnRGlQ1dU1HjhbhGIciaW9N1098Cp0HDHECalJgwpOe8ntwJL37ZWv1R7svvxnIQK7Qpw9G8LA8IzetVrLb9hK6Ha4HeG+VqOcBgwMAyTRCJUFw+QJuw3wwIsRW+RWe+zXGgjmwoYqC6hrVIfCmTuK1zOTmzZu1VnsVrBES/K0vl8xO4xe+rOoqkDrWsQyQS3nwVRQTI8tU0Us7RDc0lNtDE44MjeD3JcTFOLoiPlK1BRl1l3aEjoOxCf0Tid3ALc9Z5F1ELumLA8cxnLx587qTpXFoKcqDIPA2c7qGDJpQX7rVGvBr6/oqAzl9W1BULKGF+f5ZQixkMsq1YE0ethLgPs0bCjdEyjshCTrrRyx8CeEFDToG+PPup4J4K78xSraRDB13he/rShgV/oKda/fR8YXqphrUeqE9LgLE41nemEEHcj0GvKYsKZizz43Z/+g+lZlbX1JfxYfmCGNnDedaXSlRwmvGpk0tqs4ghH6nUHWCmMe9ly6eMRf4ykUkOD7wObH/waRAqdaCcWYsUnPQQqEn8Y2kYSf6SE7vp8l6DpkEl881JawGBdZemyJVPSf0qI2+8owdFJCvr1qR+0d9rAEarICM/p1GHkzA4WIpZYubHONbS1EnIec4Rd6YoqfV3YtT2cY2fxvryRhrDMrC26gDS95ztYAN3YTmpS/S6p+bGOomcPyrJxL3hkzlSmxyPqa24ePOGtuf8kzd5sKZCgdOyvhsjdQV3GZzRmWdwuNcxqagjDp+Qh395Ttd851YMPfbqLXOPEtSnyoeykrG/NpITBnTRhtndRHoSBXHF4KpYH3DeMuWxRH92WkYGVd7cGhSt3OhKOJGV84JklMgiBDuX5GuNVyYYXk8+Dug2pDBMJHF7lW44qGpRt3ofwmqRL7qZf/yXeAXfdTvDj8K8aRWfTu0vxHHUaOy7csFijhVM7yq+lLwLQtgXGw8IdJrkp1qISE6TtIPXAF6kju7eDQG4vqwGfV/cZhQGEqZDBddzDyWHLbdI14kUGwhSuy/UOOEflwg0TTVsjKDsOxKiRKr7MeuSLiD/GIVNkkELpH4jm9hg1Dxz02EsmKq31/YBB4C3SEYfdfUO2uk3VLdLaacRE+B+aI+s8AmFWid5s6Gn5iba1yul0rNS+FuHyKct4E3stmKEAScrJ28Q3R6O1Nrnmz3duwcXpoIEem3ipH4znrYvFZaGUMYvjo4sjJUxwKUDyYIJANlRJx58rBn5v//TK7xWTu26x5A+2qiZyvew29IK+cMKSGYbMPRpm2Q5usJMkFwaPoAwdtwNW5RGZ5iT+KrPCo8MPLuDmYVfDSowTZHVjhTB7TmV82/8WDKgF5fPDh9P4him44fmh7Z48ZbLTlLFDL4HJDduA9rxGNwJJiJkbiEFHYPRBVp5jmwwaxvclpYboKNkDSfbNwRW64CQSJCxN0zB/hBdIbdSl19rVsoe6nxqxBQEy4jVS6BRDRyCQtBIgIeAMToQGFHUfHrcsglgFcFpuzXXa8tvXtGML/5iCaKy8xaCZlTJdkkXxr57H3Xs+E9qQAnJGsFpmeIpeVTEGsYKCU3R4XR3SVaaD5aRAVbfTJiVJARQTKPBr+7DV/nndpAyFiwg9/MtLkAaphICFcibhL17omweFqv4A1Bya24FKVrLQOQlAHCLKaxmMJNUVeQUN+oos7yfgJyca4PIN1ER4x1i3w7BkY91V/iqVg1yw2MSE4S7WrQhSa7Q3A0Nuwsl0n+0ZnVX1kU01cc7ySR9Srjux2mjy0iMo958K4ZDSt7uNZYI+0mCA/nxuwHSElX6i0oJv4ZHULD2Ol49lpa3wygkrF5NcGGAW2e6GdeHb8mJaaFNgFZm8puD4+HwV1CTDCTRs2Kpniq6+3/xxJus0e7zrj9zn+leYnIOPgoPOH8pLfywJ8AJ+gzuRR4G9W1ahwjWplRQCW1I5K3UBlPdxSYrlGxgTvDZH+eOXLl7w6YomB5QJVTbPqUBD1zR6zI2DEZ27RPsga268nbdU6KV7HhMVdppeOa/d1KhIK2ELU+w7tYwx/1D5KR5OJakUpWJqjEjoEI8lc+fRMALFg9i2QBJjB1KwGQnbNDjdweTLIvKCIaszXziFUySJ6BtLZpfxjMXgtd9WJ2DNnUOr5VqOtrddnz0J3hHweLspaJIWNGXObKbkZD1fNakdeRpFpc5F43IMZcalJIcK9L3xcEaFt1rG7JSgzdrgKTqexW68d5Eau2OIC/Y1EL7FFPzIUMqnDJ7xWVB1JhzE2v2mjjipXE2zw8woe2/MQm+zFYu3LzDL/fRxBlPhuLPE+tCeUbmUkUdWP9k1HsGq7d7vfh+n1DqA+RYFUGZcaFsb7JSCBZssh6eZUYs8jat199maAf48nCZqrqA3vi/QLlyjMjbtJipE99I9oIdbQuH8AUcrVaYyYcQ4944zI5Ycea5cAiuZ8OJMUDuJEShivfqfJvZe5Dop/Iwnh994G3yireFFaypa+5r2Ia9AhPjFpIlJVdJB+2t6GaTA5BKzWJKk/1UNpazIvNaHZNC+s3LTel6MGz4stzt43pfGKsvNnM2uPcb70WHysMqL9ywfrYsStBQ07NQKJpk0BatRwTUvjxBk0PW0sczpPBDHqHb+1lWDagD1MwHu8KC/HMCtr1ny1z1LxYchmSOn7hWZcmsaLo4KyXm92dE4NtNcAAHWVQM3BCmarmZc3VEJRxfLCOSIhiZN4Eca7aukfGovPfo4Xqh62YYB8yMH4EATjS2G1QXH065ZstT3vdeAiPPMSj41JAvO38N+UPFnaJHyuIGjtWPqD4CmOV4fticpABZE+kMcrVfVX83HV1vGG4E8shgDyKwxGuiXxPNMn/6vOoUQikDYlwjyb59F3jOTgIW3THu3Cw/0HBsYdQaMuCEa+pBqMBdhTN8WHWOT47EcJIDPVqgofDMS7qiuHANiMOyX38jo/KTImruNVkVPrlbHf1osOeHofzaDOScHK9fgziRGDk3VyjTFnHBYRJ5z6OCNq77TKLzaOlcYQ5mzWekU6tXhCoSVZs1QTOGS97Y7ye3nmEbUTi1o0haSlV0baV58r+2AJ523/I1sm9ZZWVdzVogYEkbet+/EnOL8RhM2PjcmOPcHgpCvTqdV6teuvOo4DRDaeT2UnrYwF08E1opy4lZ+GBX4LUmvAq0QOZq4P5On30nxmsxVyHeL2Ah1shmq3HQmv0BpOUgkmT28y3/PuF6XvgcAt38WTspGGH5HJDaQrGzQqronYXwv93CwTFkNyAzLO01XF5Y/AqriFM/2xYORcI6rbIG6IfTRz5w6BXHYZIbRTd4EowhJaFsiRWUylirbIEJl8rRfbcM12K1qZiAoY4PqBRQ+YZYqgKCXm3OBNzNtZG5DdJX90/f1wEk14wHvUeDnZAb4NByikF3CFmShOlLtiA0qgw/csRLC88qF2l1NoiEGu9xtU3L2Q0E/BEcBNOfvk9nkSd5B9a3JblrQTHvLMSst82J6aWTnQfKpJaaDeZdTfJOm6xeHsVvlQALzveaWuwxZe9rrb6Fb1afZxxGoWgb0IMcKHmW0mZTdW5IROqYzzAcpGxF+d0Nw9EG2udKhecZqOrKWNk8FyKvP3PlhQEDs9FfJKiOaGjlbkQfB6SJPohh23CG2L/D5GdSjU+rqCmdg9QRr403TPuSWd8WMd/KoRe00MekBHb7YqYJdxVl8Rghzo9dPdjzE7zu/v7TiySSQLGp8k5MidRvlkZ4PaW20WYC2KQ114eyS18zp4cpiLMT7IhMxiB9+wdQd0yeEYjHlg6+2uhS84TqhbVyGvOjzmmm72p+g7J2vtpBB/EUNCYue4UPwcwg9FHnXJFhzQSujV0BSmJvypqio9815t2eUm/sTP65wFYUJDPTuAxhuyMS55m9KbaCUcEggjZscItJwfoHjpgKUoLcR586HVTe5bHIVynw+Qht04bkqCFEGTmLQsqjxDkMENW/J3QASuX+ZvfTVPEYRruv5ZQlNwFQ2++hmOydvdUoIEB5ayR7rCjKKI6Dt/YXxvTAxxYo/exbwagV4WvrGBncJqV3r32dODgUk90VCF2nAFa0fwm60Xhy363m34WXdIAj+ripdKexbqI7BxZ2pWrMOKUffrC9anjbgtKUtK7EArXpXIeaLv6LmzfHtUfiB4J0znla5fPL1fQROIMaUR04ZC7IsGKqux+P5vgQpa08ojBom4QC9qKcCB/6s8gU5cvTJDtzRKwAcHWq0poqNQG4vxrHu80I9LMMdbukT5m76paUroSem2LQ78iU4cqzGrzp7+rWbdyP43laaRl5sgSZ+dN3Qy9+bEGp7JIzAorjtY/PbSxlXugrmIzkQi0hBsn2tvC2EsUTu31DwJXVLnjpcppBQ8QkZzr94otZlGw4kUTOuDUtj+u6BKVMesbBEYXBO0ewCsdwEWxG3jJY6YqVZsbLahCaF7EjbqysnNZYnTjeaGMlK2ZG+rczrrrphXdePUZeCndJnsDE2mVgRAZYx15uJ/4UjeSB78AInzAgq7ZcdRI0+9qqQuUryCmHWnlS0Wj3TvI3lZ1+ZXJseJCM06chBmBx0I5miQR38FEYbFLjdSPFi+15axE0raK3FmKzaVBE8fOToSQgU2N4CA+XbRxL70imC1SfQn/zZFlQ4uHsp4Axd2nH+DQRqvAiE+NBrFza+YTpZJvjYk2FjY3ZY8H/6IK14ioiLlcEgP8WbVl7X2lOaBmYI/kz+POEb1xFY+eRIxZDRIt8IRbyF8izGkYwmZGW0J8xa3x6aTLkTvuUEtRuEmnkT3jHJdRFo8ixP2KwmiuEae86+jZriUENMKBT+qRrydqlbZsOkbkhakXg4gnWlXAxVICQlE0oARN0P1HugLnYQpcHHEJHVC4fgogv4wYeliQZRbZGfYm6xL4mim0v1NUGiVHbul86BPltPEWnLNtlK8GTvoRO68zeFLCmpLk6BsAmembLbO0inUeYJWRD10SeTpxBQiACoJJ0Tpq4M8tdxt2tmXCaNxMfRdvtFDg28VTSzlv6hhEqEfBIiRwUusc2PWTAkJy7vuQJTlRVplQDLFKS/T0um1m0KG8NGAXXJQgygSlR4msDoXB9Lx20IIU9mFIeimTqh762eSYprlmW5JXrAMbbvgAeAwOVLfHVnUlOYQG8/zY2/pO1brL0lTHdj4k5M9UG9y/NUB2yBK6NRJfx7tOpI3qyRri9idEUdVevkjD47W79fyJ7Q1ZmCtAHbYvdJaLPB8i13tPUygC1ltAVMAHmFxJELOQKD4i5p8GTjEigmZ810NFSYM5S39iBaNIY7xWIQ7559stHR2YgqGf4q7spn7+Yu8BdH3LX27k4+q190HAm9Qx0IAw2BNEjUIxWpvrEo+01RzQj0qvWz1RDaMXEeWRL4iQ8xktbuBL7UaeffHK0EYTKhU0tFV04Qj6UkKZymOfnwIAWr604sYTfPxbVAHHlJ/6ldY7+cUvxvtZQkVAwo/FRXYnoouHqs2FPItWkrwN048gugsrBzyvU4JvKr5xLOdA8dCGM/m4eRK2E+HnpzucjpdnwqyhgGiekWambRlmdbERhdv/jzOXgupLcv+XpF4a6iSYH2iNVOJKxlp6YS7JlY3PcZYwHcHn76R73T9HtWETunaHULDKWPaw/Dzn9/28l9WPlDi97CElloVvza//NBbOfoagczDvilk8iJLe0UZ/09p5x5/fWcv976p0Xdtf3M1eYV4sZADoAB8PpNmJ/GZ0rxkNg/dLl82BO8xrBt72N6LOIF59NhpZl9zoQT2gikdvCPvXjLrlo96hoHt22WQsTTY/721iwwJhCQ1Usw0LIe9XeirpCP6EqAqwXxg+GM0iX1GNECrRVGdb5zfZWom0SrMCftsLEMKySUpP5D+qjVtCzvP5i/4Z87PKfcBnNHR68Jey84X5xhmvtzLHyRT0azbyOd8Gg3SiYVm2+qm+Ea4Y/zmuQlPpHJL37iXBLrEk+MIReXzF9Au74oHpIS8SSI+o/NPLyExbj0TjGjzbKrXPt6uceYKzkJvMKoEZjtXEDjV8ii8PpMWOV9hBiEwjI+Itgu9GrYSh4ItQw5GW7oLGNmw981KMkhXg6urx3r4WowIbp45Dg+YO0z/kTPhMvnHHH9HYu8RPti6OZ6B3CIxE9vFJv3qLpcUHkQaCHmHPIU1r5PI+Z0cjpcNH/gkrcbaajwzOx67Nq4hgisE8F3Bk1JJ+U4nGr+Wo1E1K+4oC9cke8QQ5a1iRU7SLdxaiMg7H2Qwgy5/M6JS/liMf8wEC/2WQf+7QztfgwT6noOobVbJMBqvg3OLUoPuaRZJdGQAehkIFKrYsV7ku0f1LQP/RdDPU8zQUT/EYnKmgbpEJEsyiNZVsmwa//H2BCwyiSqy6cdO7enr7CyfD0ogN264Bw/zW8nVKY7djLO/T8Qm8zEnLQXrlA9a/31Es3s/2O4duNlHoEOA7axlfpziNxToCRNV6vSy4NvZqRp1PPcfK+SSVqD9VoMLF/SfYQWpksgu0d9b8HuJ19gXLNeduI+1pu5rfNuZnUfxE4TgK3qOCVgVWPRQIJLt2muUOLaIiisVrjPbPLefOIlwe8yI/TWJ3Cmmj8aWjMpa7F9m8NgmYfs4lNLMfHiZHkvcU3E5irt9bBoTiYnIiRGVd1heCbqY2FxVIaJqMwLvr93p959jaUuhEOxHNH3U0fzPpO0YRXqI201JRuOfFNvugB+m0cGuwZ7griU+zTxV3q9+EZGlOhA+nwkfGaBYBlT9bhIh5brBHjxlplV/vjK5iHd0xH+zTkHjRif8d44n+CjswEG2VZrikk5TfEClooy5L1fGxw3EQ6eYW50hIh37FcOocHROrxZu6Ua5Ut35w5K9khG1LHqKBGotK1d2KpB+ivFzF4frAQ4xHDYZzIJDQ6sG8FeXEiCm3q0IZnHzkDnuNwc1vO9ENBpoGJPyhLWaOWCkr5ywFwtq+PtGVK0shx3uIqR6VwpbJHw+WtGW3xudjm92ehbwibIkVqa+Prc4hwl063wNZxXHY10iCgGGo7dW+4ztsv4uireBhtp2HLqNDeNXAb1znTEy6XYa6jJRrry6+t4+PHGtLQPPWx4gKQSU9wqqYYPtEeZ+0YwoA9Pc0tlyrk32wwpgVFBGoW0eLvoxadsOHICHrfuVWHugD9XbiYGSkZ2vxQzcMdUEzp30e3COVX/o0zaj5pa0/wkrlE/eS8BXAoaD63v+6kRQttSjj9GNmH7f83DCMNS/AozzUAQJPUoABxmND4xq1eyELslKluytubAvAAJ0oBGJp2u1Ul5QG5V9YDXRovAGjzMdPFniv7mZVfhRwMp3LwYc/nmrEipaQVe7Zjsd/adIaPDXznmfUPgSfMOrfgVjqFglFw/kThGb0GqRd8fdLNxMmYYevLngDVu/yHJAgkgAwQwzW7Dy47ZM2i1e6FCj/bE5hFELzoRG1dPtLNADHeiTVb3MNudUZHhjSTCYK2CWtUT7laQubwtAjw+W6ROS7FHBL56HKLBRAGxE+OoiaytSavln7/58DfWltnlgEGyzTtPA0nws6Zp2cYdSHDwl7O5fEgIsRCY/guCsVABwge8LDKT772nLyyM1bxDqHrc8Wth0BVyhFNoMsFffiEvYCT5nYMT9ua53mpw13x4+yADgq5rIeOxBQOidgnWUgyjfJ2m4UNqa39vQCoBBp/wlkC548dQCnAVHKmRJZ/Co89X+KVn03a6qLnUUaGSy43HgNQlMiwUkzNXeBZDzABshmN25JyuhTOx0HXgCAC9vEedRgUmDBhAopxqGPsIj57275as5bEbsZwHCEv6KV3tCN4qR//eSfUsJk/xjjIpbg4t3QCgeZ59jtCM6MdnYby73fji3sTE7iJMaGnQm7NgI5pU4OaSgECaoKjTI6YkzN6tODx3N4aGfabodzCDtG2yRx6Ro26rS5zdCEswe8z0j3BTDPzGxzTHIETJw0EJydcwGk9MMR8a+AMJF9VIcN/Yq8aJx/ac8Et2YCBsnph1gcG0SM1ZqtQeAIwszQFXZS0bfpkVw4Pd0ZRQYbBYc1e/1Q6grZSEnu8RkKphcSYKJ1FaXLwSXXRWFs4R8j86p8icC5ZB/s8ONHZdhB8LirhvafqYxph5SSXt9TZdDmvS4nhF52VZeJoWw8oXzjXeX1/LgGcSEHYi6sSn0ZA5gRAybV3+bA/bSaDI2NhnTmiFwtIJS8Hm8RnrwrPS+3gCC5LRZcchD4Q3M1oUXitcW2woneIt05WakdmUn6MHZrFiDnbkyJ0MXsTliewfgWIyHME1KF3HY7n5dNzLaDQ/KU/9nqPlXS0eCr8GuWQBH7faHXuRR47geb9ebQBQ1t4KQEms5C8Jxke+zzDXchqSx4P4DA3y1n++PS3x87ZOV0Ww8QI6xUJEzQELNER4qL57NggrHd8za9moSnHHYje/kMvXC2YkyvzSVJxyOLhgxeLDQb/BF8c1pxuz/zB6gcTDQW9JnlvF1R5Y8i7CajOYeBwWzI20PfPBw33Z9zdRu+sodvZRV3Du5SlqHGDFPrCgVfI3AnmGNA5tLkZ4oir9SwIHC5X8n5ff2aimtdDF5Me1K2dCHkkXqB9aQVeKL7ikItPd2iG1Cm23qxhW5xIEPrOx+KsDgCAiSuZO2rQbPX+h4fR4HpG0by5RCiXISLMFntkCZr//39YHktZftJKQ4zLfalcbMpkMFkEsCmnUpqTH9D9kCS+nQdA/P5W0nf5a5LbUg+/vbz3Gh9/nkE795KuWto1SD/zHDwUTNigJuBIjvu63dDKPbUgGGKtusZcU1vWOEyef0WAPJJNnv9L2krtNWw76N899tJMsX3QaXN5URRi61wCPbntdt9tO5RvNtk8oSYeDH+Ey4V8k5P2+eqZwmmcNIPflLNZT/vUs7zxxJMqrnNdaPdED2ju2ohBNE1rQ3TyAQJjfNDmFjDNzlfnsGoahKMgCDbavUlRmXt8uYEfw/G5LrZk3IcFyQJ8iqeJdijDPmC6DqwO0ShH5BbZ+fBFNg41c4MkXTqFe2cpCFPr3GHAm0ZFU1u88VwybNwP317vISoJnDwTg/cAnLLAyfJ++vLFoK9FopSVQXw1M038t7AduY/ROcDbnQ54pVRVyjs8C2fpds5/BbiL47R41GbUXQWYecxsGsC1vkUvMFRY/4kVOdPMIqCKZ07zZFqA2emtmT/s5O8+7o8BzM6aaUOpb+uVVpQ8y27XR1Iz+TkJFGAn7QUmfYeiaBGxL985j/1IrILYNMm0EoCEvLFcjamkLFjlI6lgl0Lbhtxmun9TcwH8Xp01Wq68tF6NWFS3Na8GnC+ZB4Fu3fsRD8BhOBJ4YfRkXftxeCg/FSaiGhyX7NjXvPuSwA6uFy0Puewv42Jr8ArkFac6IoVm4TKpgw/4BaD1oiifhcO0XoydpkXC589OWNkw6QW+I+p+O/0mJDI5wi7/cADZS3mGztqwa5fZlXZIqAmahZxOs=
`pragma protect end_data_block
`pragma protect digest_block
2d388a2b7cfd7bb9f8165e71abe8edf7382b401860f6dac99f2282c5dea9aec2
`pragma protect end_digest_block
`pragma protect end_protected
