`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
byi2G+z7ywKs25ZDEs7BbH8W3llplFMCeaFcZ26mVhzTz7/fsIPxB1S8c9rn3BIUyRwtLk8xSqHXyC6lZOevDP2Flu+HYP+mOUXICYz1x7Cx54JDgTLyztmWp7ZJZ1JhY03HfB/d25pqY0DAg8ZYqaMR1lrgy8BdFgYCmijLFVNjq2z2ji3dygtSewdbT6czN8Tba47SLX+PH9kq34KW7Ao1qz4onhS0wbhqHDxPdknySuHp7nwcuNpFGQc30AcgvyCxaAVM5nRbyIr0Fu4GasV6iPbL20bDMyTNInzXq86MTKmuv4A19iz33zxPYwOTNb1fm7TlP4ZKlEI+jT+/4hn4XW2ckopIHrPCzQ581L9h/JMTx1LLJcbwlM8tOGefFPrtauEIuoAcV9i6/r4Pab9cqIZ359+OjBmZUBCG927C1uNRCXXXaP1wCh71O0NGXMxI9GY0UQZzWCFNFF5RDRrkqPw7G/PkOALCE+a0iAMBGASnpzpob2KAZnP7jqyRFNvtj42mP0wX7thGRTFh16t6MPAokzXE7oXUaVMwOhlLrbynxVMdqRY+RFNAt0uRVaarMFvRJskH2zrh+vcmBYDiOcb/shCVFA7x0XWjJGY63eDWNwM2oufxiDiQ9q/jIZqzO+2RoMUgyqrPLin49rfYJAdxrb7lmTgYpzI+eepQi6TmiJjiXRmaJmK+EMs9czcY4leM6vrn225UfM5yXqvHSaP3AOd0byNicgZkzYTZW5n4bcC2a1ofZLxdyyXniRMj6r9iQe+Gqkpr0l5KHzlsMYZnMQ+OgYClOjAj5a6yNsbVOBcTWrLx0bGMfKV14vcYaEI/b8Lkd7Zgu38LAdH+8T/mP56+72x6rEvrBmxnFfcQa2tCXl9lp41sQHLb8wzEoaltLL0xZPf2iUO58Dm3tIWgchf9xHSdVY9J373+3kgSXfekr14kGXxnxg3FSWQy4HRMWyxQ81xcIg8VA5x7ZhoH3pr9tLaEroNB9vXguczqGehSyjnGMy6onYN8xMoPHrxzGDwzzUZa6roBDImJrXF3UqHO1rhlK8bYhCc5bLJv+ZROKUvrVobDDno7yPb1w/xt2luv+BsoIem4r8FWv01AR/lvULYKzTApzfPOib+o1FefmRnOXbS34WNFyaSo0Iut9B1p2CTE10IU9Jc7w1J5VIzTN5+5mkjoFben7JGCJzgOUNTY8Eh6BSbl1ucqsk3U7NElEiV2NDxbd2cLp8H3oF5Ke/kQlpG6e6VOqRknTfkhYUgfDtk4DNY9ZaJWoqoWaW45RVaBlAl+ANgAGORVvzbw1K8pxDHVV30oXmPUgeUa82jLKeAvx7fBszZJkARhXMQKfoRX8qNRyvecMPy1ZZqdmwO5IUwzRLGLwOqm5ow14t4qGfbGPEIXhuff+XV1jhBty+S8L59PCidDoVZRRUhxxiwKSaU0dhluWFubFf5AAyPti4IkYPd4SaNIQQxwadauJirniwchLi3z3e2dD2A/qzPLMz46z7aZQ5BZiBFPX82y16UEwuc+j86a9fWqO3GP0XIXNismJKFs4zVZ0JpgXO2/5/0SqsytpjcSjK9TXmr3eR9dNA0HrDmt+3gsEmXZGOSZ6NPUenElA8CtnjaKlBTeF2S/Te9rjcqd8CYu6QeRSjigS8YMMV/jmr/W06eq7qYPB6Jd/NLSC0gzUtDJ2lj0xUxjp0iza4fTv5zPQCunSwiidUP2OhfVnlX9aMCCibZ0wW7Y1ENRDNljZQHwlZFO3f9p1BOIvhLRGm80JtH9+8t+qPx3iGhT9I+PayqsRwgqpUlCR0K+/eG+uV1yCxsjDkUYoPnwtIy8Nr0OxKiewOQY6s/96px08BC6eY3YQPSwPMjqRElGz9sfNSk0uYgaMP6M1S5W9YDJ9PfdvNMrn7NJurZbuvICODSF46c8IHc3hcAtT72IVI1U0G/xynx3L1imBRjywod+eDROYF+NwF6z4W4lqRsNe2v9gUcc69cD8RQpQ7TrUfZDkGyWilrOfmstLDaMjVDLJqzO/PdDHcbpZYpqOsEgthw5t7zReSnYC5LeZwR1eRgZmpQOTdgG99twXXlCERhvfYQOXGj6h3pn79U1uoFj3kPp5oFTraEEoDFCyqPYED8eGKWdVnHLl/g+AiO26L6fvxT7/5vnP9H+lNI+eZyDcSzQSsMlzEQel2Kx5d/ltWPAO9A9klnawk2w3vP1oyVq/mi+6g/l4JwP+dSX183x0m3oBFdtCw1rohk9Zr4d5EJTvNF8iOMzqgx7ZC/EHV4WG2TQb4Vv6Yiz3uGjDUbHJmqgKM/aRrGiy7UmwHEJJCcPLwoBgUfYUKlyVs+JigR+J/zqfci04yq12fKuyjy6vtlZzmzqKFNln7ucs09df7ScoLH/IqEWKCc3VvdhLxTdtxQfPeKheQYYLWg0//lpvTI/kzcFreXxTNSZ+a85Xiqzjk0zpsS/YVzp8c+/FVmfen8rusxssFeFpV4DhNk4xVXtezgUWH1tFEYD4BWGhejICX+ierMBg5ZnCJ6+2fTsR2S5fWxlP55wNoe2aQi8Get8ZPG1d6nrmeeP2G4AJRf1ykV/awDkwBOp7P5BSH/zDDPMAGlM8hlx0jcF+LnImti207XkvAmWSyJ+Rvx/Le9Uc2j0ZLrdKkoPehdUf8G386UlulFPsVpyQxROskxl3y7EPQp87mVK7vags8sm5uUi73BBXJCrq2/7yUJQ+yUY9Q6vqQuRQ6b2ENDBCWdUTg99A8JyZXquZ+aGOYk+Q6AiHDnrfU8qJ1lCV+Y9iEJ0l0vUyyrWEkJjbCnzCaLKUfgJJg997mQIR8jYpwb2uKNf7O97Q5+/srKvQOXBM7bn2hNNv/gbX+l9uFYHlrsRjHSsCxm2arvRCSAt6G9dGNm5fvD3yisfjKblfUeU89l44JsEUg9MCG8O3VVB95c9W8cnrXLiasxWPcEyU+vzoTAYQJyoTZ8AxntARyh7A/z6qCvDStP4C5SGWQr89VQRd84cotaQY4mkhwhGzp/wwBfpLxNDYUGZQd7cKuGqr/UCDzbeL3ze8ulB/S1n+Uvgm6YA4UQsKLIxaNKtKh+1kCnUaFtgXXb54fSGZGmA5lXkFg50YLm4xf4tHcMrLcPO0GiFODPExXxAPx/PyySbGwxk5FHxR3iJWUgyOaZQvZTAAGQ9UWKh2xI4zFWyhi/bdTRLroVrGJGmJd3lg25RxBb2jyoX41O4MM4caVb8p7sYd7dkXXoSbYlwWrJX1fvhXYvKm/e/OSK25Msh4wafDrKwH/nt+wJ22UF9RfIHddl1sucXl7NNnEuCyeUBzCs77UI0ooqE6b+15IAST9e+hFLNAkVUmtBlMze5/jxGVqSv8qIpVY+GF4TjWgq4r27k0j8bRem9VTpz+4j7pD1HTJvEmEFE7IAsJ5megXTfczebxAs4wKm7lbnvLz/MtqR/mvRxYmfZFf37T5kqBNqAA1XOkPlXYiWZedoyqHFV0Z0jXZe1Ouv73pck+UEAPkKH73YcslolUArGpxjh8ZdqjjsIEZDCG/JckDLEpovqh42ZTk6eWib1EhnCLUMhBq9jBXLXtf0ni6osh8RbB3G2/ZfrQn3tQcKgN/wu03vCFE7YG+lap6doU7KOIFuXB/JbPXdy2imIc6ObZTvbQMMj589Ergbn82EzkHxfersnQNLgpCUKxxlU5FctmMmtka30g5gcOYkbK0l7KN5UhFk9uJ+jBpqsMEXh1+UGNuXTaS7D2xfgXFiBU3ly/ncN0DUYA8KBbIBPbAR5N6N9t2jU749mVaYmpjj1jO3HRPk+icbLKAnfqzmfEi7UwZiyppeMCJquss6rRzke3iViDB9RcJPcS1WYe2Nvnf7WP/fjAIbkBiAVcGPVxXGJ+++5TDqUZ1h489S9l2XNoAdIt+5oh+IQni90Mxl39/7VTwVWt169K7rkruJ8OAh8vgkHwrudGJqNCuG9Ntbnxomrw/rgPE+I9aOPZGAdfZYCiRoByqtoi1mK24DvqQwd+TlwmNFy+kRLokhMkKpOm4kATPmbSJ4pgZgOdN6aRcazX+mMwxW/jBz5leVQGXTO/pwxH+658LGCU382oyplp/dgRsgc/k7ejS+i5kz6gAayW8Imcp6X3UoremYeTVjT4MnpBbRT5K+Ue4vsQ0+biY0uNWcjNTf6RnvttHdON1w8aZCzyrSnXdFPLRTmcsWJ25kpJZn7QktPOO8IhxER4ugPIRjGRSrc+FeVjp7q6R0w+13Se6nMBpYSLh6+qlebaZzeAf9CeFk3/4gSpw3j6ZgUv9LXXjoNmFoslv/kqgCZUC45mJuVsQc0biY2XpK39JrTO3OZEF0d1DLON/SgGvHh3Pmg8hGpeiKnHXRF049o/qMCXcxZBeyUXhDzbLoShzI/C/UZNTx5fh3R07GtJZ884KIgnYWNv2KmMFUEkp9r4Rjr0Ib7Vha7z7UVrGzBidRQB9Y8CghtHMPV3uN4+cwplxA5m2VdORBxZUzhzW3BtMYIwQhJ9lT1NZKJeeVIf8YH4HaVICQObieSHahb8oHKz0/TYnBTKg2W6zUhvB0sh7MJPR6lqLtsM5DPn3SK8L1KH5CBM1bA+lVQdUWzOW4a6cu35kBbpR9fwIEp6h2KAMjVKBFELpmcDL4EcgQC1sYXF8WJCrxEJ7qQ6YUFIipRvwnW5CbHTLj/AK8HHpfkoK47WJUWS023EnKgP+zWVvIChFeCvUswgK8C+K8AwNaNRpUW6SjL4j7KykxUjSG3jRYZuv12z1T0qpTHy2yOSW8nyIy9Q/km2PuEzqB6zhgJXkSBrqPebN+x+tMu31+fa1aUTfEi6YxOF2s2v0c+qzU5Ef1izOz+d6tAoMnQ+CrTlBvP2TaxECtMYLQ1PUw7eoB3CqaQoFbS32fiO8qz08JQ2BRFcCQJ3JgAXh3xpaRUfog4LeIBol1SkA+BVfluiVDjuvs4SGImtaSGnNzlmvelev1dDRPosh86QW3Ps+2zi+CtXa8IGm4VmE7ruWxtFGr4Uqfjs5d5D9fIQVaVcfXe4DvQJw2gx0sEI1JSdnDElLhisrx33kC0uHonrw9zTB6KwDOU+D9I2pav5J4CynwWa2bXEoyh516e8jq5MJeUzTMeVMSGPApga1nqtPmrFtnXRWzpH6uWJizcLAYiqmilyTzfLUG//R7zFTBYWV2nleLv0NqGB9KQbwT44ydb+lckrHcnPpYjpeQk2O93YEfPeQ8ANXYRUCFFUCUa39uklKVBDur7gGJB//PZMpCZ/Bx/yhMQo0lv0LGD1maBvW56pPglwJJ63bmwwTJK9w11mQXMo4t2H8PXRJbZmqr6WhLcTnda8xKOSFWZarNRTR3Rq0/bjNiRoQQxGzZmHmZ3m1j0oIvLPAqV2GlURCnZnNpABn/ZAbqPqoM6Ta/TcEu7r21JnFPXHKxG7p7ZjApOS6dlf+vzOtrGXHjI1U/tgxx2xvsjUv+x1XSrtK8K6HQOU+udzmJH9zEMwDbXmph8yc4NyV4gOSe/kJ2HM5h/rj/aXsurP3SuI6PsLYfCDxopVVlmytXVQcEZx+5h8o96Qr59gKowDAdsX+/wuIc6t3sR6px8YSZ9lOjejkXwQzJzv78knFcUlXrbEtnR3qjm5xgQBkDAG3mGsayqQ8Rl3wvKDmeD7wM6Fs0PFqxcvEMOOh87k11m/1ghQFZPnIZrCmB/L0kw4NiA0xCQpHuBKFCKIcDXkQ+lJqMRo2Eo0dBhvHaQSvW5a5aaGihmjvOIr90whvQ/zQaoNHJo3lUkcK+c55fx9ip/A728uumCwA6Z1LzMn+72iWK4dV9bQ1MNJ2WgO8k1QBJp4d7AGwbPYIgS0fl6sahs1BD31tfKRdc0GaUc+kKE7wntnY1dIto6W84+s/tC6InrGfsj3CxKxKpBmGwCray21tsmwBJSN32bH72temIoa+GrkH16MKK/VD3HWN8aoew2AZC9v/LZeFQdzZwviPo7M/m4vTgRc59EpycTFYl9VRny0EClsKs70u8OH1ko5fHgPnE1Na01cb+fRWvZbuSG9Sm0uiEuI/XNXcwZtCWCXAxpfBDXTaMB8bG8eJBCIvjpQeb5ODYEeaM+uHNaJW5AEbVsEjDzwf3ycaGWnz5RGknCZfMTJBeRG7sBLwFPKFdXPQ/A+T52AzS7hqcz3QKAMLSiLKoU+6wnp67sihzMvryQNYWF0TqWd6UqmtJqQIcxd6PMqb3HsO0NAk8sM8xKLpwj4txW26p93djXUoP0N9CjPi1X8LQ2ll5jUePqPkzEyM04dhy2qAg2jWfMk9jy7VPaEpxM+MeFjG2/C2kEEqlXg2j1F1Bg+al1n/it59hsCOHIrLWDTEuCC+rMXCPpjyfX32ssJLIC8guDzbmyJ8eGOjIR9luC5Jo0rdwqFU5AFDO/HiYfHfzVmXOq4GEBt7qnrkPqBUilHvC0HXh4njlE/zXtiUIm4Ax9j9VN55YM1JjLtaEfB2HZKhLi/eRfJhRGnu/P7ZmHgZt9UVhXZBd8ZmYbKJ2oJyyC4KYJnTJsN2pvInZJQRvaCDf4iHhapu65VvEkYyy3/JqP2CUdf0KQFBeGu/I4imaSZojROSqFkq7xOTbH+74IxDdRu/vJPOBqpMi7uFxMR3Yh2pseUVM69NEukn6x2yMhlX+SwOV58ykW6z20d27/Xa2TW+gu9D8T/i2N0pRRMIFMFm1Wy0DJnLzxSFsPhEd0xwOBimzFRRP25ZPCrL46j87Ld5vIbENiLW567291f8xjUFH6oLIhUdKqIeij200MQxjKG4rSN8H702BdtKqgBkyGpZkzYSVQDoBFxVVlcON2z5dmYv4kYZhiC+dVa1+EXy7TzJcmswB3kshAxvcVJqihW6BhavHm1Lt2mgq2wRqifyr/Ts/QeJzIjMy1vSvHl6B0ORGL89gZ6jR0ubTajkZHfK2fqRd5C0zs8qqRoogyfa00t/h4DEDjyiEyEiaD9nTvFrWlSPlEUWiXm5fF7eQd7DZmu5mn7YiMg1zPGVDwEde2OYwz7nfFWcs4HwexonoQS7oVzI2m8aFfoySeBPWF+Qoo4VBqIw7RJAI1PrALaJj9sp17DGwPW91544Cjn/ZYrFG/UG4t2Owo/Dupfxmp8NVUHRzkx34OX9ecoUr+gGDxurEsrqDeqaPb8Dvy4TotJhElNmh4HYeAUs06R25ln2sPA929Pw6az3m/1/AyxZSU1FwngEyBsi4BbvFXQdTEzxSOE1vyOuQ8Q6Eb7uloS+omBLQVmKZotBZ4XKSBgXVGuhPBkP2eFBOAG+CrmUhbfU1wpp4m0gCFGf5XeohoB1Y2aFIa3aAGmDcffHXZ86+Nm46ffb5pAuD4MwbdJyGBcU4GOdqvvy5+DCL7V/bWg0nVJ3BvcnBRmwfkE8vyPQdHPWRzJCa/AWraGzT8lhz7uVL+OXqc0s3aXmfzzjyrvXWuuGAteEsBwh2xfpgQQsgG/3KfXw+j9uuXtxM9w97JRjmrH+kFs2RQXkyluxpyKJV96ZwY4v93YGMw+iyMhusYhPMxqSLNkZz2L0tVLjfKkxx+Uc+nsEhWc62TnSrFD327IV2Vf7VyEpDc57Cb/5nM+2vv5/PefYIM9WDTDp0o/ASFMRDTx6XkMdJ6ubGD+cSRoc3wA4vylyP+aIoqLzummNLCadoCdUm95Gg4y5htVLEqc5iwRVcfs6V/DCTKC52DENntvKgx2T7d2I8azDn190+LAFUP7RI/tUyytldJMbbjPFhBqqADFyZJdrULzHT2lWxwhAQ3/eo3JsWw1uAkShn2iay2Vxm767c4w3Yw4HofJvtltllqNkK9VvML3sv0cd0ztjk/ETi3mcxvUzrP8/2h5M0AwD4vt47Dr1y1EYRUJAajE60qvsJG0N91Zho12Sp/IE6UzLrOanzzUkJ8ObMwz6WZ/nI36ZIgIrtD9Qb585Z700TkW0jxHzb9xIUBqUet/YKfrTz9mFSd/6X2XS3T7P8Dc19wFKfzG7TSJurpGVbUNxxeNVXJGInQM1QMee3pn1Sak6oG59Guwczs163m2Frp59D3cWThqdQFjBZaFcQGNBDvd3XFQhb4jF6Pbcj1GmtFc6D/ZYc5v6a4Xz41Bykx0g3m8Wy9p8zuc5XcLA4k5aCannCWdJQpxfErECf73YULXdlkgRSbk3J+QJRgzZfGuQp1tlb8b1eFMjtx5TCeRwXKjX8pUhs1uMSCH9Vm5guYmsc1+90ZWY5wJZDZOsfxLAItiIuG/aQTD7YUmwZgaUxoXaUn6nOiRA/exc+At7eLQsrZPUUQ3sZWl1Y4ti8bwarP2Wb6XvBl4IpSdonAVGaeOPLpymMg1+0JXbM19WICB7s4KgXTPrSdPu3BAKfEhg216YgQ3kq/paMKexIqKsKwXf6UeSPP2XX7LMYC5Vzssph+eXJLD1MtL4kJ8lv1G/eSPlEkqWXe2kWL6NuqoW/qc95ZdyBf2dDxdLiWX9u5UqzGdQ9su4Gw8l9+/UwxN4B4m4xpBmKzzr2oNKgChMTrdYk1pMlGJXDhLiplRSoARyGjtdP6aWZIVqFp2FQ8LDhZw+r1L6Tpd3g6rCzywB+TNhZZOQbpbvLIsVP58D/ZNXe3yzsWx9gxqMBEzrmYce6UapZ+JjIDSiPsI781rrr+DOxDCIaHCnq6qfwCb0di6xm242SN3OymPMP004+EpLnNREz3DlqfVuDfOH00ktO1LHverOeksRRKVDFueyiHJhMoia+hWXbfwawcW0ItD6R6kLd9yfohCzfjS7NRh4npJTlpc55txuRZv7q5ObmPyI2z5xzp70RyqP7DOE5OMJfYOJaVXs8jx4t5igE/sIjwSTKbl/RB3Xatt2zTpaMKOnNboGK9dzkEjllrK04L1W0xlqqYjWXrJe8Ej2/8cZDKJ8HOl/TErSuqfndpjV0aUGREju3okj1pCqdWIaJ7kvMQlCcj0D9LYP1fHLJ5iJdMzi1RGAuUj2kyIT8m7Hf4eQ+OiCF+XAJBTwF06JQt9qUlbLPQHL46Ojs2HaGkhoMeaWSHjv3F6UFBNDD9cw/bHpsG9bTD6vdWds+WmL3m929Ao/3/5qachITMqe3qXQc0mQS/E3TsgKnyVYLMLszql89WuQ6afEMHjuo/NOgwh7T31BIUs11qixub8lG2qRw3p8/OHNFHVJbBrVEb1XQkbpJt/OnT8fBCC9ThTKsDgo0lDOd3JKWW9CKCjasUk5nPY/9iCRBD1boDImtHR5gGWRcfnj2mdRSV7Qq5ESyXMf6ea7c+iIOpYYAIUhdlIBzXPPQmE/lWXIqTBnVJ7Rjx6nchrXBceucGTxI3AsWJWPErsxy406rm2pmQ1nUvs5zZ45HZC9qQ3rCU5EQlUGwPOWkJr0qfoJR/WB/V2p2WcF3QrIK41+ai4UIADRTOnnM5k8XhEzuXPmG6kFUytuUjQOCrkw5nxJskpL4eJ2jrr4Z75ILgrzUoedm8JfIv1pmPupQRzJwMVE6NY6TcS/cBI8Q4p3iBqrNT30gwCLdYUXZt4vxO2NDiC6/ap17Pdb57PKS4jPaEkVMSIT3iRYknciFnG31/n9U95GqENquX2X2rUGp57f7WMzW0hlQWwWFySKQcQ3+I9kW6+HZwnklkEXf6YUWVDJmI38ye/4SHbD4ytuuaFLdsWpQG4FHxh6uFd6X4b+yCczNXrEqQmp6rNBwQH63FOvI8CW66h70HID7bEaVDEth15bKVbHt8m2YmWCHKNhSy+PTcYKKqAmtOpe4BvnWZfI1W6eu6k2z6D75NRwyNpTDQBsDFdtb1vDFZl4npbl4hoH/zCVUyljFiZRWGrWrVRhQRZhRsYKKsk3K+nOrUq6UDSEB7jkF3q4CA6qFdZrvr34z0XyF0qmrZHHVWuQtburQqOY7uJOVSkiTEYBgJxbgh52j6Ue+LmDUWNSZZ5W1KZx9Ymv4ECeQYkV/no3cEWN8KCNgHtvgLP7E5Z3XDIi2xn3gm3YaNXr7SljriggvBhbbX/ERr6iOAxzmCgJzNAGXI90JFTM9zcMmcF8Y9DFkvfSl7TSzNA4v0AMvD47YVJCMIePJ7sKm6z+d6QgYtF28NloeQwnRhGvShIESxgod+oKmnQoPkaRQs1mgLS+NkGrOlKpVhJlcokjE0uaTSzNzpogaE5mRgR4ltPHzF8gAMizfeCGkMqIzrOrzHJJtWb/zu18ILoFd2JO+k09V5kuZ5a+8MUC8sVUNzda5GIq8BqLppjh8P/FYfOPYUdNkGQcBSNqzs9guZkRgcSAC488JkiLfH7cHIIPerEj68fqz4Ietq92OUl56uUOAWaXTwZV+NDi2XOB4EhHGuNSA5A3dhtt9wEVsi/Vaq1gmE6Rpmr7OnQlIrKB9qKdamxzo1ONsIzL7gS1Dix1nSAlZpgkp5FT09B3y3d29b8KYF+MDGhJcduSIQesHh3nx2K61O5gPls6iVpuakfmFTPu4k7V/ldgvbLvMxpvA/+gQ0UJoCP70neO+/p7JzjnDB2c3Q2UYOtbSvbFV4kU2rGMlb1XCMnbnxs58+xibFkytXjS7OfmA77VhAEkv84C+0/4YPU2+tz5GWRYb3bYh8kRQ/2dCr5N6lvdTduDLelJVXv6gJ4dlRrUsiqh4+WjMdhYyuc+m6vP8AkJMnegkLUgw7BwpPAntS7HqwJBxQvUuze6eLj0eBpHmNoHrbBK5chYn2vmXbgYOGKmSIMISrKxlz40FOIfJWm71uzmX8ghJ2pW4AMAYFyitxhpk1cq5oFvNFcZ/nC2D+i4M2oeK+AHG8mqKDJoMOU3AwKlQHNHmCVohgDorgWZ1AUutPgZwHoZhgJgsv1En2Qu2mLm9MX6LY1kvBkQXYNhN3StwUiDzvldikFCzketlMVkSN5JA2QD8CZH8DAev3Un2X4DRUynQ5ee+8eJCtE2JIqIteoDShvqLupq3QbodWs4d2EwqNzCnZcN3Sc9p6l5BfUbk2uIWWlUaoikm4GlRYLw7AxWPupt+sT5PZq9iZAIEKP8ZfyBTP32sABdS36/vACpdTizesG+1lvSW6HzM1WctKwFA2Qn6qI62Q/TLluRbqz7pPKaJdWXx82cJgBzzV1R0i/Q0CMG+QRsXn46+4/DPM5NqLMif5sstKry2dJEt9LfhVVHRTctvrSeDNFFZOY5IM73lS6CXJWuKkj5n5rjPNtdIWsPkeMsczX8RaQfVqX0u3HMOZTstJIHsayVtJrhSuf8XEw7GV+Rr+C1Oq+ZV8yDBMCvxnRpwZMAJew1VVM7AiN6InBz2AxmikLT7mWB1i++zA3PsA2uUxM0Pa2tP92SHxv5gZxHFom7fhsQwDhy8QBGLQBspr4gL4jySo4xCOK3GM1jiAT9COYPPZaCzgE0q92/hx4Abyiwd+zpfBDhgq/ejSwO+Rc646EftwXH7rvq4eOI3/DlNzvc/Tx+D4Eq5GTWsG+Kx6uhOYOdWC8fRLNOzc5qratAezVFtZiHRmpw14Zr+OgXT1qxdooiuYWljrAmUEcsp0W202Yy7fZwDIj83M1rLpm40gJKk7mS8gSrASa2QOD3A8wYVUp2SIvrhpTPQH8WqL9WpSxa2fL4gAvb/hE4QnSBuP1ZPt1hY/HFaibJq8pemwgeITBXQ/SueMMKLhf12w0uzZBEuK94Tc8vnwNo697wLh0+CqOp/57uvQDr7bwwhMvGUHqtUbrVScpQD9G9XX2x8iWZO9M0h2TyTeJYrL6A1leG7TKtSRvULQrKvQanV3P57v/JLaLaF64lXv/R2G6CLWCNG4+AfynCPG7oSpZ5roB3CYWedAt3xo2TrREssqiwdCIoDBrWZddhNtNoQ6EmdHv2fm4V3s5Gq16ip0uxrG2jYP6gtQjEu2IBMksR+D4ukFw8xr3KoFgGj1TgbgMZb80Ovy4o/dHQpqEJhriurOZPOJUptKSZS66Wa0k47KuY2wPG/090D88aoRcQAsuuqGWI8c5gODUD8VkwkAFar6XGG7F2sRuxBKrQhAzA7FOgVLg1weRuVAQqAMayox4w6lIXrjVjs16c38hWoaHI+r/JaPfmC3X73GSV4HkyVPRNm2wg3P6B9yWX5AV/qI7SE7b9qPZJ8D6IzeYKnYT7tdxAFe2p+5OM8H3KkiLoX0v8J92+1Wrtj7640EhOsmO7e3KBaQySQVqGOEPqrzuHK/MtyqAl6mN17T9VCKThga8H1nu7JD83qTWNjUN64BYiYRPX3powZWOJLpXxg7TOKS9x1Qntl3IkQDybDyaAq+9lh0ld9U6HkQvgJe4QVRZqJp6qAEwMzaOgd85ZxXN+o2buk5CtXXPvuAEWgitk1TwAqCW7yrvKC3RLFipagENnRh+7x0F/n8AJNTN/gmu5hJw8szqZh6Tu4UheehCouGrWicxXTRr9Pow4fZ5VdiS6jiUp8/qK8HQ4vYvtnIKHhT23jG34od8SycO/991+pscPl76rrbcDHyqjmkK/h2PqQwLhY0Ljs0OGO51ZXyTY5PFNeuxYCN8fG4U5d+13fqc8k0ljke0KS1a9sOT+sXC6Q1C2v4zMOLFz7QVm5v350Qby9bMlTibjBeaywFm7xjN3tmXSsJazPueU/h5slking3Ujt4MFMmIlK/bE47aAGkx/U05OrKO8Qw3r5c5lBMbn//8eESgsQ9Io6i5kQnP8MYLlS/r08C2BqljUHZo69Q8wmf4+VENryKkMhAnoATwmWpduPHGBg6npLY+HS67k5fk/tA2P1BVV84j22KX9OnA7nocFdRfRK0T0pJ39RMVhZ33K92mLa5wWQc+HmH/tLRtNWjpyVHH0cHPDUxc7+z6SeMsG4Nu0+IgZ2e1wBPOapktkjfld3LZocsoN+SaCmA/5MqC0hFQXQriPy5Uv9NH4g6CD0UUFf+twHQjBlULNSIMnPigM3RVVVy7r/xauu2H3tguFx1zaOGFE2VcdjcdWnzI/u642k4XjfsEn4Pm88grEUUvlsHJPYV7so2cz43YAJhOKSw6NmlT42iCQpy9gIiNw/RDTDULCYaFrgGF/DK0D1/3hnbH69R6PKBYg7DTvENozAm9GrMm4vJj/abd1Ef4rWvPfi02BcTvAxdb0JdLiwirJbBsVYp5+gLqDLWyuC6UYF6LChlKCO4vngYCFJ/f2PT0HXNAwCqnKaPqA4IXMPMSHkNXOJy6CLL1clcVEOP02Kq2UByX7z3OQrMT7PCq0YsS6PrWz5Nc+JoZWPICdENILvO0qoL4SieZhmnIHgC4zbX8KM3PANsMM//MP17kahPvNCLBeCpB/jwI3+j5rre3H++L0NZab1ehVG0PyRcMmGnIr9y7REvA6YzgQdy1SqD5K+xjL8mCxtb3ZJN9GPBxCLNKiOdQhMOoYSEnffKwZQFUfDIO/ZUJgpjea/4nW674QOPas9xMr14tjLsB9iazy+jecANrqDpgsaUsTn5OdNc9chy4EHO3tC0saFBk4r5TRx2G7DoEmF1rQVScPxOuiAW55BVGmdZPjDlJtQ57A5RhdX4vjTn7ycH5MypRKlPCkm5htfZDqVobmPGcZIbjBDc1qrYXVri3URWx8UND77RWaFNlE2vdijh8ZExy9+mjWwJcD1Wj/pvojOGx31akko78FZmKfV2VV+IoosBoBHWcmwINVCHWy6Hqc0xyJ/3psPryYViXpoML9xRBs0mhxB9KTdzBBuh2cIGn2cft06iicUS1yYWcxiI4OznqTeVuvndbMtE6bZbcRz+LXIu78qvsorC6hZGUqgX5iJoBfXMT/7RQmP4APn4mB4kZkIaXWleqzBVWcmTjS22mXwXTsZm1vUv3SKExjUS+MdxiMo6u8543Vg6KcqJQMeia1fLDtAnror06fOyOGKQQaqDKqgfn1JJSJ/5Nulczudj4I7/g6vRZ0mvPHkw1O2j9nRdBLX9OGVWUg9hgAZX+fPYzOdfszM4c3Nh8muA0JN596U4SvScqdvcAbBsjGolPWx8jesq9hbRbY8WX5nGeBOHorUojHV4uy3dvaSOC0AjRvHSvCPTaaezcjUtZY4sBY7hBWu2gPRfp9qIYh/BcQnmjOShkXEsRykWmSluFPglN+ErO5Xd/wQIsyivjc9eMZX2vrbHlqq14J9Lf7Peg+ozjvOD1rh/2YKrRnAKlpPydZ+0AGjEe2IgbyHLXqrBsgAit0VbkgLVDnYm2HxCcuteu5qe3/qJY+QHfGJQ2wfSfUywYjsBfrbeLLgspKZ3U+qhwBXS6veD/BLgEid0F6sIAA6ZG/kwUDBm1XaNeNN3s0qF7rlUCcsta8ZCD7VkL+bww3pWtl4vFvT/1+XtYXY1q0N50qzdxXMa6db4VLq5YZm/NN2EMKC9qIKdSJqxYD10Tr2Iogg5dlEOm9eDbxxABL7uc1Hiwsl8gwn0tKLSDL76014xHzQ6odmqnqVrYBq0PuxBhcH1a5cya8U0z89p+2GNDg6LHjVQG5GVUyTHAeBg5ceEo7hgJe4Lhtqc0qLqF+Ju1jdVVPiAYSFiyQa9PbjFBbKN1Y+KpmQUuAGrCtZiJGxiTt7mYvWkFrfJjm+RI6MFjW8Ve9/0m20RyKCvHVb9OTmermOYS1T/2OGIc4ee0GnO546I3/kEZgDqUhhZGAyxl3pxIz42P+sTQrWYx8TlRrO5us8bb8WjM7YMOcuXOrvxOGoJGZ4VyHyoZoMlHku87B165MDdeP3OyOMytiZqmSyPax1rALiroRfXUqMcsvJdsp4etUWMR5LAn9b/HZicZAXZYwx8tpUIcxUhqgTmSUbEpmiodwFYpS8P5+hE9aodRxYUdN7hVOOjI9fVfgMhdVUN2Dq9ZqFGnYaUiIlIZoZznfRwao6ljanWiKCnNPwaIhDfkcvd7sLHWtxnUZe5Q9e/hDlCkMWdrXY0+6yYJKwWmWr0qQQAJr9Kiu4VIZTCbcuz4kOyyf5mO4WEOSJ834bWGic+IaQ1BuzJDvli9ikFfykXXCGZs1t5HIamnRHwQLs/bkAt/qQ/uS8FOvlV6roMv+NKK8ilpfHCE/zY+VebQ939GZDLBckJndKsEf16H49PJE1fXPoe7e59DXaqlGIdpcfsSFQBmez72dvVWtEMr89mnX0RuT3q7K2LMglCfPnU1/N8z0FAwsSOpzCaXNNqcoclUu6yU+4YLGKBbmfcRZLismtjAvbkY8uQwjwXy4hhQPB4pkIKGZxLfmcLMJPTOtsLDQ2bEbTEpJrHTusY3FJbSrxwR70ITv5Fc+lBGMhAQiTMYM6VmADpie81qSYbI33YuOaYyk10nYWirEmnGy38+bKAdCYjz4V1QjEbYAlya03HFtRGPUDvHJi7l1SR0ORu/iy4zEn+x6g+kumeVYbliEYwQsXV61XOhpXQbQ8kfuHWaNOnFh4KO/LdiF68KyPrRoeuCBZcO6tLCuBwJleITCkU5m96mfH7dj1woGjoO4EhyqdE3Wwexug7Un2VQM3Sh96GmUdpS4t43wJ4OI5OtLEa2IBLbY/9rl+RC7y9wzD2eVUgr7kK8Y23kxsllxgr7oVf7+uxVwIOqkojXtlALAOozXWpBoSXSEPF3VBmjTBjYHe8hlKPJpusuQclbJboUUksng6MzGs/RH4LgEkEQm06F0JfN8EmKmQRDdZpnCdrwJMNyFT/ScqkebLvA3Jwh7hfpdL8dLbsZboljshumyS5y8PyDDiXL5/AEguEkfuRLkWofCkRCvJhRhVxVDUfE89vSpaPjV9hUxVRMKTtf3n5qTk5xNxALLcl/q8Z0ZlnDcPCxkP9l1+iJSHJbo67BMy/3gU2+VEXc3Fhq9c0g3+sTyoW6ogtp/dveqrEHf1bHo/eYH+/YgCpCwRW6sed5LFktpvf+skMxoMmzrfkdjsW+i40J/YkOnvL1JvS2X2+EW5zErqgPudo9lNarStyG8prJkHy1CZHPmSksfAPp0g4FJ2dCsrM+Hl76nP4jAbOx/a6nOW7oKngZz0+g22Vd1oOZOGgaPFcHrbip2PWg1u4IbVsBcD2gaOI4ktRrdOsLNgrZObRNk/aIIrzcuqUpi1q9+bT7lFSJC38yc/HigYZYyE+MdFXKT2MzIrlrOBW3hnyN4AezrFIs+p4A0HL2EFlaoaRm8tTEvit8dN9N1sQ2OWzUr42SjzeS+FM8HO6dWMvQKz3idd0F9U/n+F7cbEZW/csVHl0hM+UuDC5D50Edcjca513TqNI4Lfd6lKTa2TRsGV/tvxaN4BOk5gk7Xsnxj12yBL/vUraLfwK81eWhwsyrSAZgVZtj70isilG3MXg3Kalg8bqpnnekuAAPdE1JeONJS6vssQNv0C/LoyjL0mnQDejGY5RH5VyRI2kpgoMRkp/6qzE5JiAkedFo0KEtHzULNIc8dIkMVCLn4PXcNEVGXtutFMP+7EH2RNq84UfKBIooMb9Qypj2hKqU4dq/nbHJdJuqUDgBNlQ4JGsRfTb99Mx/iRd9++F0NnHUaW/hD2za7UWkH6VM/04iWcGpbBX6pGtLf8rdmHCYaR9MNnFjjJI7PA2ytm90I/Q41FRfr7Lv6OvrKzQSUAYP5k/HbHsItyYzwiIMCwTbKyx78j3hciLBfEyF4kAGf3EmdGCOnm3+bSMlT9yon2q48/HrZRwFVptQQ3gh2EBGTfix+MehCjXruesy9RLZbuksoYzosiuFmwJffv+ivmqhYbK8uWmfAr/QqzTPxiy/4REuttPNnU6Q+If0wHJ2cS++VFW8Z30HBpODtAPQSnNreLcIKLSuGF6BaTDEzEVUPXS3NZxZHErBuxUCkfy9nzrCSvxJVitz06Vew3t9i8YKv/cJAcJWOHqAUt446pDVN9dKvtcbS2rIs6PqxZ9TgZARdxoOmyIyDhiAEQwT2gVPBfVKGyRRXatGWjjGccOkc7Vn2MCcNy4syz574H2Fvl1WFlGw0JHZPuJBSkF4dk0yC7KmWTNnonHMigqHvX3sMfnqu4cp59GWR8lh+lnrXr9OPj59qdhT0WGsK7cqm5gRez9vXScSphYUNCDyU8wtFqenk19coZf4FePBNXeN3RBhq3u/VgEhsBRlWXZe2FG5XMo2oCt7kz8fTMs4pGck0U/gEYXpdKQqMXmJcZCecTbZq9a7pRba+i7HvmwopisgDZ73V78q7JCeFkFnjLv5qSYMG4hXApHro0u2z8qWEGPktvsCp3k97oYo9+pHV20eVOL5uPq4dBOpbnQKq+cr5Vv/7cEOJOZeFkogc/h2TvvtFFaIPLHfaMRshoRRE1Mno5h89LjHkAgPF5l8NjupOQp280dMdeobPXu1bhLHcCbgQYYtEbIfr0ixu6YnWbXBBQqoAwzhNbrKQRdgwuiwweqwgc5s+M5jQvIKwhjyZEA/mNeGEsb8YpzbOECAX5VLDtHa1m13bxqD4fwuUOY6CUVq9w2WM9cxHaafcP0pMh2KweG9G/+owVR3g8bxFSXtb6MYFBWHwnhjCL28lPZQkch5pdei1yJyVWHC5NnJLl8BZqIkEhCfACE6trqBJlTrO/bi87wxR9MUBK9AY8VXCTVNXMJwPB+19IalfzPGGifkfmpUtujLm39giFUAN+4/AH0lJ34F0IPuSohM5oNmJpgJyXXGP7P84rW56kRcy9ePJZbIbKuIAJeTUHLC7OQDOcqBNZUAc0unkjd6pf2ohnT1l1aletW+RxQwLeGduO5lq0fzEPlv4ViFHR5vuMSYrP2P9UQHjG10ULYslfFVainVKxew1MCgxxdEeOJcqftpq7on40shg16WEd/NhECnOxU54eJ5hyfFU1qDhe+IN0+9jSJP+t/PHFQ4eOaF6trMDbK4Nqlc3n3ywjYm0m7PcAhoR5ChOEm6Mgy4RS+MXqKiYlB1UBOWqjmRc6EjdqD6AyTfOGQElfN0FikyIqnaRzJJfCA2SCe3sUR5QI4yZpqV1GU13tY6/ZyrFF4pvNN5tWgkhN5s1glP3VHxIr4hiStpe8s8PGyrGGwMvzIsfi/+zZGg3hBMd22DFdJ/MUsNpLOCr+n16r4M5JHdY13ZXzwsZGvqSvp7nliikCDT0tf/7kf8p9Nwd/UCHNb/3GKa7gOoHBFGToVGZ3phl22rpKu6Q3cBWRlUchPH2aG01vhoNV8onlqwF+4LI4iBAK6jH1965dSFT1u0w8CqfwwIqbQG91IHO8EXf5aCIsLCpyZ9JR8ZMDITDHTu5U5p92M/gDgBn2YkjDmzv/uGWsiO8alWPp/7M0ryhUepgJrbZuZzDd/h7mt6uB9NllH8FNpucOvXEhqGixclbnXeP28c2PvVP+7T0REF/2Hf0CyCmzUA+b1R/S7j7sret732bZFpbSqkCGHxGi5ffocDPG2qokyBgh64x1/cUb6Wi77khDdgCH87Wrjd+g5GbB9yw/iJjcxuZTDvL2dWFFWtTrdOvjYr8xrnjm1s7w835sYeb27aHGnGgfXA7TeiT+N7srDYFr/uHHRSPnoBt6OXVHE8UyrX0rSBsmqVowzYxoy4h1An4Svu3BYEJcbEnFKfITrZkrXHy5OvcRE54uomKWD/W5dyhzmRnOS3LbW4JMZ97SeHQUj2pyumKL7EEcnw8LOunRfPXJVpWNsCxYOM7WHZ0bs0J8t1q6a8r6QCND5do8ah3LcZXbXqNMI9wJuU+Ix3OW/rlvAnUAIAZJSmeoTzeRQC9/sf031kvGqiYCppzJrZZxa+V7r5n9uJKBAfKsv9xDno8jKRNq0IzLDtvPQUmESHaQK/Tw1pHhZjbhQJxM26GawRrZ6LJgC31GE+tsv7eCuy5eyCuUCoUJV7QSNPhv0XZi2n0kYONtknn0/dcgqSQg4utebGXCoHGsA7BKEVr4LKW9BgtHVAt8NEfi5HaWMUlAPpb1ZBPgLHyJJSiA+IUF8CJmuL/gufD2mbaWYDnRpGsLupUhg3fLeEtSbjOqPI2hq3IjWiz2QpLED7TOtCVWDOiPZWk8VAKIeeDaJPVB9jn3+t6I+sb0elkiBqW95C0f2Be4jnYYxFcINk2mX7a3yI5udsE952PF6novfVMbJkTYXmGgAX5X+MuvFYupdbpVigNDUapdfVpNAz4m9tPSdtrQfpnpLyOhlEWGZIp+dzPdjGw3D7AiWdlXN1gD2zccM36IzPgMiC+WQBdfPMgwRaEWql8enChPs/kvwo1DcfBVFRxKh7pteLvKkn9HeQ1zes9Kl/Q3LN4QCdudXeHOjtiSNuK8f/icehGi1mQz8FXShGQgiSIROdjczx8nBw37pCYzvUdTrAsZs0L10zbVxC0aa+algnvt3QN+F7SKHI+ABCjnwpyUUf1/ZDeRzMRJhUXs+cTejnLT+MWIf2XqCE50BfwnGp992kZvKlRfVUPPceuRBVKVsrh65Kk11Pgs2ZJHZXYc7NB1EbUcCwKQp3cHSD0sjl7zT9XkmN3Dec746cT4epf4d7JZe83sRWVxHeIK0ijJO/S9/FTx0ncbNvZzRwR0N03y5M5f4jpWY+uLnpbmJHerlEqlClWlJSHfhdHNL6DNk1C2EHMphNAtoNnC31wzx2wEq3Kdfw4A2ZGM6ZZ1m16PIQAoA3GG9R2ucaL/308fHJszeoEQcDU80DtFSycI9j+ZJbUAiEhfEyl1NhWsI1vACRza7Ju8YHAcoHKfzgB6IpA+g87mlyVUg9v9EppjJ93HjotXWtdUt6tp7QLJzAPO+6ekGPVF565aWxkybpFdIpTt9QINGktkbhrW/GgRDD0OMQ67/9JpmQX0Ryqvh1d/y3l1xGd2MpagF9RJc+SGVEWli/lRy+2v0dfWKiKNpPtCPFfuWAiP6GibslG+4VOfCCDsCPzVSZguaOhQORPbbAtvyypnKbCwkWj5LdeB1ZhtAMOuMnhvYpreDCdjS+jrreotbtFWSqoEsVwFy76C9c7yXr0ux1vf3P2vDS52bdWCkF3vhpuYL8MLSlG9dI6bPezUGc5HoI7a+uZSGqZBvzOL1BYqawcxwZi9nvKucDNq48cBVXIF77JrLQdNGxRKp7YS4uPMQrQW5jxguhXVSX1jQVAYmnAXYykn1NHsVV9GP40xNSzaVK9ygzktCOwI54FR7J9DQYixZymvnOdE/D1GU83ajSfIt1vpEmWzGTFPcdMlRRKm9+Shi0f0jiNWVaXcUHcT0tK8bVY2tNmUWNiocJjgytirZpTusRzkQzz6tW5OOT+TRFrajQNnmXbaIQli1Y0VAVhHy9QUwY3TW5zWU1xo9gZkh7sjyS0DYKrmpF+nYdDYi5ddev6zKYYF+LNb5sljiBygzUqJRlOp2iGSNb13Wl4JWzpKEJ+1zxBrFAPLL2FBm5GI8fq3CEA4Rry//YdPmP7aD3+cT3xw97SHofWi5xQzsTA8kAhQdgRlNR8ockyYOxt19gnmRAGlTIhqSX5Rh2L3u5IhQgjdOjRysCyCftR/BcmGwF/Tezbdna1d4GujCz8LdKg0XYhNvdi7y5AEnikPmIu/mkBv+nSkkINZab/COdjkbURxRdcCpbP7uQw/xBoeJL4+EVmokvnaZAQ0T7483cH4pBhQ6XEVUwCN0SaqWVZW1xUsrJZCPkcrCLXtcp1g3nrEr+PEfDQc8vwLrpMAxxCITUhgJOFdP76Ig8ar7uXcz7mZze7n8qQ3USeWS/LdcAzbyawI8f0UHt2Bft3uCVMhctvYaECnI8/Ze6R9AnslYrRtNZg5W7Q1B7lSt9rHIM3QqwIVj6X5EZUSieZttEJHvIH7x/cRTue/CcyFryPpUzErq9FsuMhl7EUFRPVpBXBJ75D96c8uTx6hYyTup4qLr65XE9jrspz0OPrMp8QPj5LrMldr89gCN0a8dx3Pf0+3r/n0fYhu7i5MHefowkj6/y5lYR48jkqbQj/tpwa26fKjNCf1bikr8rcpJ+65sziurPAwwd45SJDWYIosR6uI4QcVoPkK9AmX4sqGQ5tuTPCHiZ6r4GgFwzksWOaLtGXw7j1OYVMnsClJGPiJJzNxfFKKAB93SVR714RN0Q/7LlxszYAgtT2J1BywXPFLuVbaOYB9Hj93wscv5l9tyI7vfN8EdL2w0HEfq/HE4ce72NGrnQW898b5hW/zu/V2/6JdnTzPFhqFVQj0fsf73ssqHf3+e7R994H06RSQiP3iXFGUvdOvkBstL8a3BEATVw8v4tX1mMvSCqQr8jgmN7TNVbbFqJXNWVNATcEzAuqGeD+Ke1E0MnCkJfmWJ+dNb9gk961b7MXMYW5V9FjLXvva+AOUA6Jf+BXj8K21UrLB0v9f/9lBt7wm7ht6IBLrol272U94cPT+1BQp1tcqYtGAW+bpOxe7lZbQsyczSLKTS0lqnveNGNwiEWy5BbBHoYKFOkCkS+neF7w+6ipYhTh597J9bjoJBJJH/2zgxo+Icf+qkNBGKu8nZEnWdPrb3bSjzoNwsWrmdwoo8kTqU+9Ke94ROn9h0DcqXdctVCha0DVK+QrvpAPS0SrVFvIx8vwCJOXLJC574xrBqGp+n+Gji0Kbqa40Lp6UX2DSkzppYRMzcViYM5nRxYD4RvO1hNVZRVUNR0sQI/TGF5vs65evxQqovk7Y8YlR7DgyLue8ysFzGzTfhIjhsWCfbHKLiqyO2FLMYiAZsYtiA0W6W0QWPu5/xnG7ZK0dY/mmsm091LIynRaCdUWz3jY0d/+a7aIyZC9z73r9lf4KVa/i1Z1AN6Qi0Au9VBapqoVmckRy1dwuxWeOombH8I7hDRrpkPJUf4DDyP195D1VE7YFrAV77OTvCMKeNFI6Jpbx9gVqb3zdkzNeA0OapII2IWfwEgxFxeUwZZ0fQk8FUw00l8IYvvFvcATYZsVGiLeC6/r1Or0+pjKOdi5K23qS4R15JWnV/Meb9BiYkNu87nniB9DtRuyPsne4iBppeIpSiS3OGLNGImViOJ6tXwCcPNyjy5yhkrNDhg7+rgprl5YYAKsSGYS2mDkmRqrBedr5Vm744hPBY8CvyyK+qTZY07pOHkHw+07H99XsD5InH/vax3T5TaPg8i1Req8xN5Yr5XScrFIyekLQ5avBorw2PgQ44EG/L9KdERIzFmvl6LuzO0uj5nIk5Qjgpa6aBlpg1ZsNt/i01SF1Ojmo7xkb1q1UZG7ZEcqKlJTbxL8cGOGVEY+GxDjFKDq54mDxvM7cY0pTH3xCbgCfKO0EfdjIA7g4rMNQBS/NbT69mGoZ1FWBOtiUz6ezMIdhCpS9zM1WbON2+lB5Dbc41/Yni2B8hVRid3YpQU4T9y/u4+SYZUXMQnqgsLbdBJik8cQRF6rEP1MS6ETf9UhhJ9Lh7P51Z3hg+00mxFOg32F6AjTXBnp+sUqS7E+trICXkQv6W3WzWfBRnoR+s+2fJZBiW8YsJ+UqooOaR7qjBuE8vCjvvjqa4kE34hoic/UylwmJ8/v9ia2FOzolKbYOMe0eRRzECAURIvlqISrxnP0UV18lNgeLg2HLobH0y/jJkdf7lWp7q7xFf9QzM6QhE+RBNLU7x2FzCNozVqw4xlj0FzDdcQU+yOTHTgFdscUHaFstIODLckPO+B0PhSZIFZgGUAw1IFNaPJe5e84ohniizahHB3b1V2wv89ocvqwop+J/OEomb6WGb8RPp1z4/rKe67aGTScu+mRtRtj+JIQsrz98kdoRzEe7Oe/C2lXGYxRyObl1s+yhkA71E0Qq2hqirG5iPEY+HNKXHeh+yQE/bdsl5XCjnkOP9dOkQKPZGGMNNZKEPnpdTMEn6mWL5dsnJViRe12qrc0KilB0s+5n0l4uMF299waaSfvJHsU9PxF4A95adW1uECYuW/sEhY7BhDD9cM7b5i+T6WwTcx++adjVmQzI6fORZ598wsxyUblaAeHYCdLoe4u4PjAYRJ4R4P5lhtiolcvN+8X5pOr6pU9mzH+224AF9Hp3Foun3OfWj6qP5wV3VNLwAfBVVJIIMU/ckfxK3pIFF1JDRgztS3FXxI6rj3zJd/zo9Y//hOhDHKCRaU1KCv13SB1DMzQ8peiGggYyF7T60Z6Rw7a8Wh2fakISRAt0Ob8AQDVwuftI3h3bZoph5N0Vv9No6FJZDRLELLqrLIDv+KzwS1nJP2da1c4FbyLjP0CLqth22Pz1AWSK4r3qNN/R0Y7xZRTqc6z31nCLNV27TYrAvztFuf/HHPEGr17EkVuxKRx7yVZwtV6PGfj1RhnNz4lQss4NDogAG8D8Ur4fsmk5kRB07KMR79WVTmh2AaWuCr1unCFZfFyuR6IpgaS1z3Y0p3U1jZpW4mJ9rLl7+malJ84SpHO5nTbt73Lp7h+UUlOKUWQYp9v/d8lNLf3ZWqtPc8d8Kro/7Va1xwa5ndRepY5Tl8rZH9eej0LLneXYI6K41sqrtbRxKoHyhOywBxwllwu0MYdQaGbQgs+6Z20YZWRzbwEA2AS4cbFR0gL66+bc1WWLNjnbzzhcRG3xR+7gGNDGbRGY3QWroEQB/hb89sJ3erXjmrwr/MOZemPYCkcoIEx/Tg9wu1m65utRrD5Je5DVFMUL2iNjqSwWj8ERuQ87fKuJjmAgGXo7Oabf4uja8HdwkMTXXxb3FShvi/Wx1YKJsfEvYsTk0gVla3DOzlDwz2s8CKnM/e54Sf7Ittl+LlN7tCGtLDzNAWx6oLmfSp6XGt+lg6XAqor8xJRbMnnrMBVuc1ABLVnHlcdiPbXkxzkgqGijkPVmFzsRt38iQsicmAw16UDgsmmuXiD1i83kXnemRt8iY1XZNfJl8pqLHxoSsgPGNedRakQpN5FpIAEibfMauV6oXjkKFizFiQg14OGET6ICsYHR+7HngwHiILkzqOdpdudvR9B1EAeUMFJK0GxaY8VcJCntnnRl2Ed8OBqDKFcr7FgKdLvhkMbxqqoUQA3DrMn8Cpozfc++SHZtEtg+2OyyhegyICr6aiouApLHSaqGD1sXC6DTOt9s+dOakFwD/GCEHeFxc/Lc81o8kA40Cf4+yVt4LFrR7f463eJvmRFFBHVjYvJJeJhQIUKs+2AJh5JWkcbWk8l9tiidk4qyA07EO3C0mHFCtxrr1jGiXJYt1sTS5MsifLhE7Sv0FTIR19tlU/JkyAGgy+Tion+k+xKK+ywBVsxHCWh4jitLV9Wna/rycog/OJJTDPBKOLc98eo/Na3nW35ADqJ3owxIdPkLLYbq0d6jyxfp7+zdg8D8edz1sZAHhFJgSyb5xVv9u4zM6cs6myux3SfO6JerSAjCgjB7ImezYcZyWCe+/t5cW18cLfndsWXm+82fkh6JycMFD4CSdmQgr2csEKTHXTMk17r/XvWuskFg2fF3ckUzlVHFHyczdDNZxjkllWNUhwbmdwKw9Zt3K43C8+jycUXwEo44stODf6ho22/Grx8uZO+DNOtrTVjqHS8Nd/rlMUNttvs9j4pJQ88+bNizc1zBwC3sX6/rL4RIUUlM053Qt0iKfAKe/rkZLjEHyLZusKaOF9X/d68vIlEpvUUeJNHxX91wm7LHbI8EWRsCCC9delEZcEvdGRYhisp7fvGzS50fBN34XFtcNLp3LypaZZBcC6DNmN5kGZvRmzIGy6Peh2H4QNdfLuWGiQt9EPrYbT9F3hZIIBe8gwRQ7mV12So29QARKkDmFcksO7HOZOXb3BxhubQ62Pd6FdHyC3+DQpCeBCXckVm/AEIo86jdDlHi+/HtZ79HedPEgwsl/xHksu9ANQO+RUvQMui9FeD8A4cLsdy/sDQ8khAR0nCC9zgwgUk0hgRDFcJsqWT81+PxErylkXt8UesO0J+CXeN/8D3YQXEeZhaTnMI38L0Dn3BgYbRAEHoKbhqIcFMrpjHy3Tj18AcoG+MWYe5pmryvr597zfVm844rOr2by0cl5PkAHYWqngp6uQb3s0ncZaAxc+kyk8oFtIzHTCRjfhlj4HktVFDkXqUpxy2OWGNKcfxST9xNMl+L1s6ik6HyTP8MTenvvwsySXVCNtce13VeKGSAMkjKYB9bH7BEbCgRvRIy3WRdk4eHf+OM7lSnRECTkhHOqI8qiZkyhScNrhTRSRT14wnBSdqketBUQjsQOTIhyoXYKXOHPk4oULFchbsMRxgWDddTqxrylUVziZKIJwQ9hZSG9QvmcR/VG0VSQs41TOFQU4Cmwed9L69rpeF5F6LRdPSr4izRkMVsHPokeSWFLW8LM1VwTkK3V2atGT2fE+Xc5L0g0ykeUetAoqRixkeX4CrwL0puZoAfBpugi5vbw3GeRop2THCX0jbyocQbIy6aPZjX0/ugVpjJlvJirMxHhJ1BedI3eF/JjaimaLtEySoWFX9sE7cc6/NKmcerlb0M7NwfhYXEs/rE1nteHEeRVx/HzxRSIZPAdqYssAzjmQoJcMluBerkOzwUSYs4kBANezd8Sjs3+Coz9f6hWGm9j+et1Qx5tIW3TKE4kbvFlh0md4bsO79v2myAwlMXQPaQ5RGbF9ilpIxkPIEvuds7WFoM1a0KaHKny86ziXGmjeVn/4E7CB0vuzO9ELNrzM+l/6X76BhPxmYkVY03shXuc4o1BbGNzpteAc8psbYe0m5xkvy4IbP4fsBwyXnBN8bywG9lZucbSyVt9QZ0MiKBxideS8v+QKuDwuum69qtE/wRrwL/S77CVIEy+EcY75fn9fLwiUdAsVSC10sAOqBpKQ7zYxFw8kgJTllazHBu5kscgs9Z7oMGTjK3CQGfPH+pRjcV2bCB4s9UZej4mwqZivhALIq4Pl1sCubSfIviF4xXSk+X3kM4tjsodSxQiRhGQxTP2W+fK4HzQ7jJBrNKvGS+lkosOle7Bt9F1zJfH5bTz062yrc93ein0/7kXFW0f8N4YwBjxMgeYagMUHxW5t/lbipRam5g6oa2OHf8OvpoRiRbBFw9xiEWMJfN4Iv0RAQ0jF/H6vzIVRrazCwXF+bx4ujkJd9T3Sj7yRmH8QAwBBhF14hrpFfcdaGhIF4Ejdb9wwIbUVUOjawn1d4LrB9y9DGJ8kyJMPDnUJJYJYfICS5ToN1XrlT8SBCjIlKCayTIbdB4dlUkENJ8TfXb+FkGZ65XDey7YV4yP1MVT/k4u8vDiW+gPrPnBLZs2J9PlcQIfy8LhGloJg4Ftgiug7wNICFApD1Vg6BXXSlFSklnM4iEDJTUh58GnJvUMz97KPDJYy8lkOpzkfvViHHdXLhk7AGEmSDLsmgqR3ZYGjvu2AE5Kaf74jObDXS5/KsPJdnTvPg6TKEJdt7zncFoFjtNjQRGdVe2bidltVABwxsKi2L/FgFVC921e8GRlsnnl+y3U1C1VVQoIssl9O4RpofswqrBg+raEgH/KogkPC1Yr24jXuUsrNZGYpwJZxBodT38WrNuSotR74BCCN4Tv5zN31wPdYnzpi20gGtgAqjtKTXSbmFOn+Ic47nB9emUggnvNmq9qsg15/u8HE9eSJQJIZSU7SbboZyxj7HIvz7POSXQoo/xeR55T20YnWsbCqOPSZLqtSqN9bSdWEqb24DzQToqCmTOL4KxynzvYpfNlFlrKcA3B2KlN5IpTSjpAmz8rc/V2bPctvcrGxA+lh12EJwBnt50xEZDL8pWBFVvA+awewZb6GzjqRK221O09fF4/XWZbfSnHC5h1RovZZxgrZ6zZRcMBxQ6I1ASxReetiWEHggeyYowjgWndQccipQiBWV41LmUT1jHPGQExCjh+0RTPxnkAwY5jRmDFfLU2B1DZN7Z/wzvtSOIP2ZCH/1iOH985w6xYFEaUyDRsbYzQIaKsVh92fsFNdV7qnMEt0vBE4pqFTHQOXxlH64vmP+NBGPN52kaNhm5XJy7Qb3GpLrFksQ3+kDyYEeFLNmnMwzl0z3u0rrGNvQjRheRQd2RqzQdUpPUxeAKkzcze8XJiSNvlFvlbKaIk+a47+iqaEj2MwuxZr++StBtLCGaVRmKfgQL5bNGa1J9/kuLaLaUuOqe1m8vVdOSuBGQE9PpVnYclIJcfaAq7FxdtCCFLSHeGhLGwEzaTm36bMZofd6GWnOTcNXJMpstJDgU3YAPdIi3Fv+CdBbUGamivhnv1trqNmDfjDKxYgATtE6/B88JqUUc0fJEQLmcpgx4rwyNRqiWhffZHbLZH6e/KsY6Ved7FbUccVNoW8383eQ5i+KP1hFGZqA74FPfehEtgR4o6XZIZwG4yCQg5jd+zD2rBuvw4PNyH0WeyEYi1Jeq+ryYYC++jTgPtaCZPhYEVppwLzwsUj2KeylL7S9VisCeaMy6m+jPOhA16wuOXiFeNG3j2+hfeDoGc/xSdlm3EFFx+x8tIrZ/7HQITuCPCo8yDZy3PQs++udyb95704wSz1vKWq4SnP81zpp2Ou2MGpXckFMm8Kr6K0PDlHMDH/HlEEc4+sDH7v8REPcAfgK86sQEv1DNN5H3tt6mI+EjTLgD/01iR5E+dcsyrUAowbhpgmXFOv4EWEd5imCfPqKxlfzenKWl+vJ8ak8LeQiHs25NwvPyCsbpAGEPXfqlxwKMNuGTrBaumCRh8JeA5xuNCI9RM2JaogvBSGeUucyA4SK8z+0PMPW46xB2NPWIhOEVRn85RCh8QtcMnUbWCLKQkI48x5dXuXnGMC/6LlclD+pzo5Lcq1X/rl+s/ZQ4Sc9tIvZ9tNze/3FHeO6hP3/e84KUKQpIdO+vbASi/LDwy9uEUkeCQA2yupYb6p0ALD4KEIh23pJ/bnpQN2v6/AcEA2sU7uDNz23RJxyeRK1dw3LzzJiOqcG9KWNkzkterTv9f5iau/thQTdWjjqexU49a9bjmpmGuhpIZXSi2KM6rUzTLp84HCmYPB+uwwfvp9vlshg4cIbLa5c35mbpOAKQkQZXaNI870ARSoQbgXJ6Zl7/kuTGavSobxXNPxw9ODx2uHYZDQLmo3osbCBpqBh4Xy+AZo8Oz5OmlTBHJtciqg5gFZnTBRKfSsIIu5wDlTwx4MivNpB9bxUeQVYbzqxA30N1ly9l1R7lcSVMuJYB9Hq3yiOm9AIDtufiYKP+bOO0f+fwkFyKoNpoBTN2BWRIsZP+7tL775ldWmh2fdYZdHIVg0oUm7TS4xm3vzrFAbw3BnrRhMF6JJrdB0z8tVCCi9ZcVDLQicStwyj71GCfPCTJYPBIRwwgrwPEGWVAOFhHVI97Wrp9KkmozlSUA6RgqB14l/yqnh9vP3Gf6CkzP+juyloCA96KpObfNmrbEWBDnupqmgW+gJTEykhkH7E8tFKTqoSSZ4XdZi6NKW3fC0VdMMWs4wN0RHmr2QLoJeINWBvvwjNptFLvboACMPnZBPtJxSDp6KDVrGb3+SjVjBM2H4zEqR8YEDhoy3EceTPzIqBgTKergYiOlCIlTj08XUOb2vclcuDOeuSGDlwY+BLEUmn343sM+/Qnvi0zO723kiYELbOgjN6Ybfeiu3cceswyKFFG+OSNQ3jRPtbldvh1ma83H1lCCSm11jP7gtI4NEepqkEQecOP0SWn6+5/jHRAHvXjSpNq26uhIq+xivYSmi7swrz/mdUGVRaT98pR0rXZnhHLt8v/WN4Q2cuOFvVsre34tx/boI8tjUPuEqvhK1W5xTgKdp9Yk8lthvxHRexReYkVtfP4+lK+ZcMrXky8UsoUMs0NAdbGmg9+Ri6n8fMgywr4vRhyT3ASnZaTt5uxpe8kw3mzieOw02w3EcbXuP07+qBpey2S4fjNk6miGY9BxxlVZFlZr5z1XVzadoJdkRncL36lPT8DWY7K3486BYx6kku9m3/erkFXbw8iTz/jRWKLX2sHjzw2dqV0cYRBU4tMyxxpJWAi6u9X9imqgSFlC55GHxSsoMK3Bj0bVbkQdHh3yCmPC+O1e/PoUVfA72rFND3OK0kxcDI/lTOeV+S0EcbzjZDfhpq3hCXNbOF345Q8q6aC/Z+RUVa5mibMZCFocC1/tRun4Q+tAk+xXTLDbLr8+W6CgCgQSOqxN0KeuR2VGl55jMdGTGG8wjYEecvDDv5CH7bcxR82Ogr8bRMnThcll9lq+IAlcMdMWmxOfzrPprP+uObjuqX2bSUlvk7CBld7ACuzs8ev05150qkYsvavsVkHhPUWCN9SOgurW/ys/5MN22IiLqbHx9Am+zpNyccHwiC2rky128iDoPRMN/xOEtdcPoDyX0WQr400guJHi+ra920QYZUHqcGxyIz7MCgBWR8x8ztMhLqwAcQ2BvBvAjl9aR+uuaxyOkJBWrdatrxixQrNtVzZvoBMiAnhuqDOgLu97X5a4zCZuMXrlH7ZFgweJkQRMGAmgkDvTT4o1bQ/sbVXDve4AllxR245EiPEPPxvR3JJU/ktG+SMt+zvPaXWBePl7OrE2MNMfuxm16SCbVoN7th6IWABbltkpeJ4cLys9AvDeh30mj6ybJ1WC96ZfRuXhkvsgS2MfMuLXhSwrbcLUmQor/hK0Thmbe8uO5Kf3OHYro+kwr6COiXynn7+ENxs1xmwLTdcYgg7ZqLmGx581xtn/Ks5ulaz7u+21nQqbf7194sJDyGmef7I8VRPXIkq2cPFrhWhyK/nWRiHgSOSZIMtn8/QIwaeTx+9IA/OsgSsboURnPVbWgNOJVTeCm//dgCKUt5RjrIvOV3Wj8jO6wZobTBk8nGVmrsC2na/5l9qTmgZ9mWvXg7kXHG+HdDVmGbOyy5sxDurXPP4xr05xezgpDN4P1gAojAcijqIKwIYnInfaxg+ppguAT/bPjQarT2FdHLeHhyKk9elOzX93dUgKxINItKYuZBcO9GAXAKw4mckkKkmg7bXMewT1OMU1oB8YCfyaEm8qJHSjLRBZnqbS3uYKWsBQ0eZt3DgJNEvq9v4eVFiboP5OhY6pRaboCe1zjXWvaCDxeYevxUbP5G32ntrKgfmv248qUXgK7HE02RACZlOGbbn4weJRI4OqX8Jis1YUJfMPe7HLOQvl4IL1bHUX5vfjcOX73ouyyFLPdpqDTq9JNlsQLYBuQXF7ZCECSLwflXKlztALtph2mYgmiM12ZqW/TZ4SE05cZsE8Etsiz4Cuw3h9wS8Q3bSU/pB34vDWWwfcymQxP6xMVQZZdBj+5b67R365aref3r+LFMgWF7SPxr5gRrLcbnesucHJ3q5qh1BP6VOj3a8Tnq2c8cal6WebmVHlISq148VAFN8R2UrG4Dsxjp7qSgOVhQE0A0Hc3qAMf/JWZ0vGvoB2KsxMI77pTw4JBuDWcCfjr/Ya/pbcnhhy9ODwoRDIl78QHV4VTBelTo1U6cEB+VNVm3wgPJZPJtW1WajZiZof39RjWK+tv/I+NF54V6Y0l8RKpJANyIK3lWP5vyi0k/LB1y4UoDE+OA0juhl13pLsnoIeptnn/jr30ZvZIlX3DlzOAHffE1HBwRjTU3OgSvxwbsFrRfFz3D4DuvBWSLZmUjX4YSEiUwWnV4RJPtckJD5KgjH6G5JXzy5+5QWuWIq6bnKifqi4TGRl0Zuw3sPDBZT79O3bIb+cOQBtaaI0XwpInuUVvqGhAJpJD4397MCKANmreKiPEf/QN+7JV1cw7OtVdHsLzbAJIEey7+ddfymXUz/9o1iCYelB277G6M7tRIKHxRyYUMG16QVsuKh2V+CbrExj5NqNPZYB58wBomci98PB+AAcNFdm6sQFJj6GklsHRTxudP2RC8con/1I44gK/G6E2nLWRAypGMAYDygQu1/CbeUefu5buzXMj6wCket0Aypf+/sE2dEBkc3OZArt/J9lnPtfY+0TFX+AeLWp7DGVQL6HigELbTeLDEsveYmWDtFKR9OOD8B0jiWLeZ0IDEi+8OKxIrnXwkeHUlNlQcnrhJrOYgBJnqkme/5BRlOjbpdrw2zO64hJIYCDIYnBhIbQqrHyHb+gJBUhkEFrInTSxc40kCFtuvGBBOrRYC63EwNIofJRtM5wLAInivINLWearYrsaBQtwxz3pG83Kj9CGLefUp7NknMa+s7QSfaVjn+N2y+vLqIzgT/5h8HlD3NOh15yak23eeiDB6LmNIGjsf8qrjp3IChxuViOClgUogdvoxRStnFPPl9030zLaCilR6nDjJ92FS5nyw5jSkDoxevDqgwghpRLY83mzM9jnsGWM0qkYEVV4Qs9/k2feCQoI3/5QJF/PYlW6Chaa6ZiCMQSHTz9US4iFo6URAxRdlkELa8BzO1ayQPKKqcGU9yd4CV8pUPZyoSoc/V5N13k7mzXuY/YwsRNzxSn1KY64AM9/L9A4wSlBVGD+LGFYuoR6tpzU7cw1on7aEsxywXs+GWntc3lfPclCgvXLef5RM7t6bE1Bl9v9gLF7AasVYPJog2yOeOHlHszBwbb/29GlW2zdZgl5PEUhtmJJaXWRKK8mk3++5WrVSTP5Cvfbru2xPnhF+ayPHhMyOSAY/r0owHOoX8mjtOIMWOq4zOcPwxrIq+xUpSbw7Ou/q1CPx/GZZS2r+Qn84k7OhCG3uWYVnwBuzlSnzlpLyU6L3njpEebMReI4dT8YNAYMO5Gr9ww2GGs8T3NBvdqaNncG+m2K/BF1FprbyFGvnkYiHJORkvYfYQkmifVdQHk41MXzb8XqA97rTsJxFYHq/R63cfu2p8dKdcHTw827rerEhisVEixoyU6swGJV4MmXustsg3jm/TN3zIHTNX/DKjhgnp4X4mYRT3SXS8fvsDCQjWGqKqT5Di8Br+oHzawvEc56AhVMyfOeu1Tfd6hhOAkBL8ocKj1NPuj+ofiuMSmLBMtWUGGhl10DlBXhS2almyRK0TlFkToe+ZDl8wKZzcvODGaj4isKRzYBSRyaIBI4+nmx1ai4kHbTTDlUdetOn85JjAqmQX10xbTTdUdy0m2QNLoeGGV3QbAeKc68QIfnG0whQDwzt+QrMxGJWKDknKqAxuaH7DqDOdxbFayYgReA9hekf8XgUEo9hQioZ4e61QtA7/fe1x5APCYabW7vMrpesoOXk4QdNsVWkPCEAKiCBAH32rLpOStsFJ+x0U+ZrPFEHLDwkaPo8iGvP+NSIBpyEWDNLyT5FgbYnQFog/7BpbwqC/yjEbDyHOgWLp3J2s0rBoTy5YrwWlUwQenYlPumnDSETBvKhjD7LrJogdjK3Hfw5Dn2jiwNHx0rk/TddRMy2BoDwER/v3OBulk8c15ws238rdT3w1BC4imfsd991rvUySP83Dl8P2BjA8Ky6SgEc5JZztsRDZu8E/ahHP3R9xL9Z9XujTCbSbdCloDYnh3sHg+bSDyXOHPGVe0tH8FlRo9JvQQb3gZmGKjjmM5n8hKgDr3yWIjsDuOlz/p1IkgVx+Iu9RMASUKt39nO0pz6P9hhpN4PAc6doNkfu2oylMj3sAqeYYueUXJ91oTGm04O0C0tlNgSxqjqrrD1Ju76adrf8l45ej8F96nn7C4qCXGxi7517B5b2zFUjW+qKLn1XgRIPorevLkFa33Rh2Uo4g1HHigLotOpd/XscwjdAt3/071Zf+WRPcnb0YaaZ0oH2/7ZJ03d5NEvplm4r0QNBsnvwFtGe1OsLJAIIyH3Y2+e3dvt5aS9Z8euFOT5ayGtAmLUohfAK/MW6FPvscMY4IKOtQdhwsftxnV7JiiaOmtHhRnoIokdCMpXiJR7or3V2mWIqCXvEjBa0p9lbBRHT0Y6nVxgs5MGqUDITFkZLlRQLdpg4eEWVnIFeqSVnqV+9jOwVlqP3W5cJra2aFsMO+YT9uAGD7SuXpyoifvAFjc5v/vWTrASluUK+C19DsFb5Jsg9PUcmNiO2dh03DDWpgIZ7b1wd35cLM4PC+FUvSE+QmeqiaEww2TkpgzN/2VJ93Ho1E9b2QRDcVf+dfC+gspVqsaeRjliihJGihfXnGyemXUG31Wj/435PYn6cXz4NxUKtXSkgHZwRQmgGQ5UrslQPbZsVHINJAjSNe9HSYeDI96dsclA6fGDV6PHMm/XSP0LyNGfLXIuVdWbjUPDe+Pr/Mmg5fYnOHyslUEannqeGbz9vB9k34l4XRnxfQs8f6Lvk2fu7Vdbk0Shr9soA90TkzNDdqYFXhvBxdS/JvcxMU6f9T74DiCWpmX3bQzWx2yW73CYXSZihMQPR3CZYEitXu2jfuMxBQPtY5w90an+FiZJMLZG2rTsjKJkWO/53ok69yqgy3Wrr3C89GjeofesPWBGOhWac4HQk5sHuV4mfRr3sY9ARtWP0diD5BiAhZcHnEY2g4462W/MN1Erh9KVqCWOvYVTnXjvoL8mcWAQyqdPmeRNTYFXecLo+bVWfy9nQWIKBMWLeNGshAi/ro+C30CkNkJK5byA48Sux5GIA6yXclkoiuRLPiKKtXHpIKnIoC+SjE+LAM0ZKaUijsuGozwfo0bUfvxYspAZSiaJVdpTKNdiNB+W1oDYx6S23RpSkJ2vTw7pgMJtrvp7FcuosCaiZjmEiPMKCM3kMjbgKs+jzgQ/+T0dYorcybWAtxtkwtKpvR9DFrLvfHd6Jm7ccKMzehhMUaMJZLHahf6vlB5H1hiUY+1Qj8q9vU3l6oZ8fgoI6VobsaySjlgwCUFYrPzWe15M11/5+a87KJzP2/jFRb9W25VyH3lO/DhkSEO2coQG/3eeyTazhb56QPIJdvGdg2137Jr60UHpS4n34WDYHju2B8/QEb4scU4kUVGqUj19pflnyu5CX1vJbNrdvbfayOHM7Fx8PiTOfUqs+ScwE10MlaeQuXj50LYg8kOGkGb4a+XWu6PDomvgQegE/yVZJ7uU0jycVWJP/fAEujBD6wvZsr1FMrunnkYe1Lmawd4XwvxJqLnonritmaCg28JvfrI+ptZOQamfmG9qJxJU96932yyBn96Ee9UtaLgkgyBem7++uYEOE8M60UNwK7NSrxOIZzt5QC9vYnMuKCtPlMF4JhY28/KPLYMyFLJq5HYAPVYW1fFhJ3jnjUkbuNfto27U3H7VGuwKRed5qahErwtfCpiw8vTljCdV/SPLYqwmD+by8m2Qrk/5aZ+KkP8JrkxP0XmmuTIBKdWGY6eVBbMSvsHlwzJxgqqdOWnL8eVruPhCTc6II7ijAYLGL83T/fMGcCmi1YE4wGLeh8GcpHSxW8f6+GGOXF0RanAc48CnikcBbRQ42O4FH5ytniFg5ew59d5zeaZ1jgspCHUTFwGu+/+fg0nOeRFsxcIoZxuRBdzNqD35Gn+b8A3G7eBU4/fkfODNn4/X/j4CR8spL+4BXrrczxcYyb7cv5ZUGQH0lupQ0axwfxulen0UfsVsMloXXDgT6R8WAdO4NFv4Ox/jYRScDJl0UPxzw5p58F97J8L4d2EjIwLT36zI50p0xLEq1a6JPAp+Hm8W51D2g6WXdRrIEeoz7j7z3SSqaVJkSoVZMKpvy9MpChUHJruOV8JTzeVptziQ/0rqbLTlBAzq6tzCQzme6u6mjEGSwji5NdC4K1MubnwZhpQr9Bsneb7Lb5OMnuKQycPmsr8VcoHe5W0orY2VE8uz8tmLBP6iQJCeSw8KkYgQiC+0x2iOgJxNeVsV5VfMZnr6SlPcgcoL0dH9PtGtZkKm4DJMpx3/zjyRdjfzf9R6AEgQ3B1R4wkIn9iob36hVqfiaDD66NbQat/rsNSGAyG6Iy2FX7Hmd5d8sOKV5L8x0pyGrf84+CS/rC/1DZjNrGM3qVamEbFXj5CNANbL7Syy39iOPTYyfnK2wIyOGpC1gExeiUc1GkbJ48JL94Mov7N8mZYzpNrCpBf3dFcg6Yp1ApGmwxt+nowQUyS7XbpNIRiuPkJiMf8vCKsu4kmcWqU9ItHx6qw4UMq8D5/g7lwUPogk7rV+AAq11vhQ40+qjY4RhrCHvxdRgPEcXR5EI2HIYuvah4Rn0q0JVI54F0kr8omgGcIzsjG0jrQMdRm0JECLVN8CXYow2h9b+7cojIvgjFE/uOPuBxrEtXr1c9Q+bIo1rqMaqknSgl6btfgkRbDB5OqJRPZ6EW7CGNk7C8413iamFetWGfiqgG0onoz4wg8YOZ9jsXhiJX28gDobaQwpBUqQwKvdmbUEjjeVZ6/Aqyi2vLfZzcLknDqPEm1F0EiMMXb5+XNdiPVdRkgfMEa8SOLk5QqBKXWGGI8jE/lAIVbDreLX0wUxOfIgMIToltRF/Kr35a9zkvNtWN3sIph26aI382buCvTfb34n7uvYglGCe/mJ/AWrYwEgpP0nmBqRb+W4IXygr8Wq8AMJdg6SAUBulV53QCaMw6VP8cszCBJGt5V13xW6t/JV+lvrcHKyWP8zI5lBEmfas2OCp5vA2vgZ21PlobPi6HhPwbCcCUTzIdTBFJzNcwzVfQrfAjHIFSWb5Vmtg4wq1JrEY7AczNi7tacjKBOowTQ2LsGxOCRm+tWhA0iRxC3F9dMDij0oQ+VBdeoWLr6aPCnhWvcTRX/C6BDjp9fjKgd47NzT57z3UqXluCWB8nRREe1f205EAlKAAluusS3QQaH6MMoEWW8Cpjkmjb4aTuCHGszQJSH9TMlA5SJjTQCBWJvM+SXaAhyMPMUFZWicOjHcydVPlNRqPEFuBNinnfKwH/Ft9e4BbYUPkwf14J45DK5d+YXCJ5FfID8EFkDgHSRh033cl2lI4SYrgjJ3i+k0WzlGhTjp/t9Pj+TK75SjjAyINwp1hNN0O7JdkpfPqmn3+nV6c5EFmNI4hat/ach8cDUVoTycNk14MHFJH32eUm8zOdfs9jh7z2FzfSdd3DimhEZiMA7+xcM7cPiPdMGhuobARDPRauQkJ2FEvKhkMwZBo+E54C/FGDA3Wi1qO35GOgA/eNnMte8vtYUOXRUAQAzyd/hkqrp44r4WOzVm3mi+bWZ6kG4s55dPUi/xxfndl8NuAbNJyzY4+lHQDikxqRlpar4kdGcJ9JJXdXp0KxhbD2FDVlRjNJdoM2xi/J3M6FxfBbPF12FTjdGG00RRxJ41xYdigl3XRbZrP92L6oiNuW2A8/HXqORnmMMfpdm4J5k6tZRL5ZkHzZfs1HMdHuXhjwA5t2b4c1CW57yizBryFjX3anWzVLitt37daMbTNnl7PWBYgquVLepRLoTkaYXYze/TUBUnsQICdrvO82Dj0TqIyFHPsmJmDnSzDLqk6JbocW48lDh0iTOSUJDROVXHG6mZTzZyANFO479rjzj7xzv8yTOgfzqHeO03xAxsS0CiDhIwOTqLywnpS5RRcveWauv5y3M4eHAPHmTy6Iy2LYy+WAJIHdqWufBWzA+P/u53WC6a5s1q1XlI7DV0/5WUwI2F6izs0QOqCOQbqzA3uPFpDMVMAEpTOkJZV9BFt3lNcj5skGuBJB8eAZUVeqND9ZWUnVy/haNvLqE4CuDbfVfU83GtU8PfX9+VliUpk9C4j8Bl+ERr1EpEknrHMq81QlL7Oa/d3Y8tj9kIEhXxpV+ifDyphP5YPofQR5Tp09W8rw8zxWzMV7jdszXiMg/0F/2FBRxoDxUDmnDRY1bouyCEecT3eJ3rNeru9UarvS/sCkp2Qksvpb1aaMZgjyl9dGw7ustRcsKIiTtWuOVCF8xIY136SRuI9OJHc151MM6O6NvorC4YG8+Qtgw5+Yh7EO9IeGKpXdW3GHCp1R+jmVdQB7MKdoiN6FcwFhqoBJt6M5Kxv/lWLsyXsbjZsmtlZAaNyYFMjDOeuQurGq9kCYvfrm7OouCp0HTDN/3e/l7DkOZri+ns/rMC6rrxM9fMzZzyxWbNWG3GJO8NBk9ShpMcjcFuZhcFn1aR5LvxkdWEqW2zrY/UaR4lhMROnSdvO3zIOWxwle2ZL933T385upld0qrkedaXGT7w6PeGQMIK6tBnUp/1I9YH6a0Xw6mmeI4c3vIOiWpeH5R3tpWGhHdkB7eqErbSJRCSQYWYkwhzwIsOLJOo0W2ElkFMrnhbMEFUFj2tvt+I//ZOdrVtjjkXVBUQ6YHKZnqyAK5YqrhqnQOcLrz3rhKZZU6dPheUBa63T2ggEyJpCocsmn0ct+s5jQ6Abv9wTeumMaoTVuGjk1oBPn5bz4+2o/V1XgrkNRswfpJgSwqZNiGRjUqeBie2r9giWMCV3N9h+7xaQLvZMe7D9755QytWnIDp4zxMeomL8jGSnFP5UCr2qFTDmyQ2H5zZp7BScwj5/apx0gLIVPDbuO8u5T0XknMkcrR6x16ivJjEW92zFziHWQ8+3//Ir8Q8h9lirkC73/1MWWQm0oc7+lIUekUtaCfGtvC29nxVA/f7YDvcz7EFDVzuWLrXC9WRoRF56nsU75LVO95BKUrTY9qpUj55n7Rnn+XYQF+K6IO+lC7v9QvS3HjsiqnW0Oc8PAD5CcP1sMylaelVE7seVKoDFj9tnch94fMNufemDbDSINCSii94Tqz0YVfXIGKimLqIexrbdqymI1NVFU2PK5Rm4Fp/N7U4bV9jSHl/RETQbDjXbLmEZqPBazad6cr+ljJmrYcyFSyvkOU0EiE1jH3cy95/o/0lyEEDpX08HJzJoYlDAvEJmY53SQYyL69Lr9O4RJVf2CWIfVFWXxu5b49OHKU8xAdEObHOj8XYTQdGGdm75OnZuRVzdj28SpHWQBM9ynbENTNRLxQfvI04BYrnlNXKtFiZX9fId1rtI5N2IkAalU43jJoqicSgnAjCmbzJdxZEFTBMp13qFuodlZg3IJgqnpWconjqx7TpnOuKmEQt+35S2SywZ3XvdjIU7wTCCbvvAWnd9H1kJuwF4Ga2NoBfvwQWLJupIllTV5m3nR97OcMVa3yeu1Z/MycbjFYJcKbv4+1vxWriNBGaXRSfjVcz3IZh+lOCGhXF5BAnLrcxc8me/4JvUOH2IizmF/AqD5toualiCal1bC2xAADKXkDI1Kb4+RRwSktMCYpjDJLfCHiHppBpt5ywdD9FRLbIaQgRTccBXf9LKE3v72DF7bbg0LO+9mAPJ5o4VvgG5MCZ5+Ctu2bVoT9CHFu5svqd0TQfkn9BFOQda+QL0yVMwfv1Qh0ZYXQQS2a++f5AzdVENnkkIpZogLJnCxfX/JitRlWdF4XeZl9QP6lCusyRfpwktM/Y8wxs7XSOcbM3Psvmixegsn+uvuWeOqyhd3ctmsXedbg6D21xOboHFLhdWTJVNaIJoZH0e+J0+C5ZECLTR3OjPO8tX7UaKOxiNrL5qQfzrzKKbuOd2N1TCDvzhZfJXttZuw9Xi05VytLm+2rwqglOzXbRPRCA1WfApvRJPCB39e3WPh0r+5yJg9yvoFcua2AjvInh6ExvlnHeAmjkI2ZtXOk2W302IbfRliJdYXU3VvkkMWs5KICB8rv/WQxQ6lB1bh95JdhB4ghvwC5foaeicWqcCKEwi7PeBeUsVmTv6MwmeaSsf1C5v0blSjipLclLEzIhRtVHLygn4xwbHZZ/j8trkDlKIGGBzG9XUTV9+iJdAoy6c581xpOJn3ujqgs/XA0RIjqZHeVxv4Bf/bvAe4IH97j9fuONd77EcteL7o/N8+5lWDaij3xUWd2qsNrPbOhw8UnXAs0ysYGpxFVL5mbUylE3HXtxa3+xEwUydqU2lECLZbKFl37aZ2Q3eV+DiaHi3kDnEOZroE6CzGiS5XIZmYAtB11jAMcvBPJHTmrUuIAHakG3yW+cBvI+nTL5aBWojCDTGXiUfCIyweOXbpgMXzkR7HLCZSKXG7M727hYbC6TPsGKG8g8oMdKxt18M/Jn+xtvBgq6L184cIQ+KhOnVcrU96M/xUeIVEeh6X4wA/+wDrDvuLhZNnJ0e0QE2Ig0shYO7mADjGp5OBJ8qCuxrcB7wGnZUhACZVJRg4HrafOeQNiqORCSkKdljn/Zo4qZzBqOi6c4d6iD4/9PT6T83AuUhmnPqEK5RCLma0EYEXxGbfjtvlLwdSLWsvug/60H7KNUnCc72YFKC9AypiRGVqcloH6xuIQ0CNy409tIb4NOKa979hjf8Bi4V1IEEmAPVcbsrL1rvBGblcjRhKo2lNJ0nAsqAJJSv9rhMOiEOJSjZGLnOOUESEWjQxP7w78zUlL7Z/xZlx5uTw+S3HpdTzWiq6IIWvz48hG3IqprliSa+6CkyYZiLBSxHyOZ/x+HVzNQALgik5+ll+QUUDd5U1gCI5iRgkNPGCyUfIuy+tx7vVW7ig8pJKNPXfgG9iNW32WLlMJwqAnk+SvamxDd/RZ5nQhfYlfAH/VJcwsYaP8qY9/UjCcIEYHFi9pKHY0kCiN3czcNSwwtnbWpJ/b2RHJ8ZI1lOvxUgLBwhuQmXFw/1GJhj6UrV9dcnswsDwPpGOmO+8JZEueiBMLYRjrewfX0P1WU/Hj+RiQSTP8J343hH24f+S6e5U06b+cXFhEyqUquqZGRyHCqIInDBvSS6cQ1MbI5HsV7gjZzKYeEh3ejYr+qBmCg8HC3nuxl0vh5fE0HhupfJPqfck6WkA+c/rERL3r5uPE3l8NBHKPwVy1FFZZbS2lkplkCQKnSPgdSX6KYV08BG2x1fQzdc1VZQeKPfkmgT9P8YEXmb57wFuRFJwa56z3w4TFaqEr9088JqcHl8+15GeDRIhEDxRA/cOF/crIHL5ipYF/tcllyEdr1Nt1vZmwBshO0cGFgzMgA0HEkyah116OYWr5ABmviDhWnK0DEuSwnn7YZXZJEsyRnihfu9VlHK+/xk95Ik7Mp4lHHyTYzd9jeNNaUBTz2wNsoT5HmOJVMdwMoKEEKlIqHcsISY1UudTgDIl57X0ouYibPrQ5NGwBsrQ7XO8ho8fpeYF6SlmeYx1fsxFi9NCzI3UEQS5Z5tjv00fvBPMdcTs4D34ex+tpULAYDQA4b6MywhpexxzHUWhi6iy7PtohS9e0d3zfy1WLHCSg+HbsMFTh8HUIKKQJWe1jnO8OWta42auyKUocfbHD+EY+/DaqDHi2rw2bNkxaPxRQgfw0jlKwsEOoqQOmsX1zPCmhJ75q+Q+dsG86ytkSz+Uz64EP0CnRfZWwCMCR1EMJ+nUAycerZ490T9BKhXsV4TkGFy+D9qlihyscUihp+8GAkZk2uUysfaHuVWAMIg6zBR3DO+KLoFZNbNBfAoRqPGqBmvJgbThvdwc3xTB4LBZCnFWYxCfu+yBMK5WxG/5JegsEfHNxE//MQnI8bZhIyt2BOtXCbEcZbUbf9JKPVLovMQRay2o7f3AxQb4Y6ju7XI/RqOjxt3KL2NYr/AJ9eKjMiosGEL+8yLr0TH+D1qMqgigw2xwEoyOTRQ3C+dD3vdaUZudm4lVRBXUlmwlV/v9W+C1f+t2tNUdkek0FfKsWrj1J26lwI83VMiD4fqf0+VoSBtMEZ6y+SO6EVt27SWR2aGOnmZsCOyiZr2KylOfMWHXH7E2hFIuWCsfJYdOgpzoPn0HtKyuUyIncYb2rsOtrqvD6EUHsfE1uaqCBeRu9droPhWznk9rHLnd8qNrgwhwjkxRs8w4IjJK5+D6+g4OcSthARbv0rZLY670Hb3CHQ2DMKo4OPKG+ysFWpCeaDmER/xtZuoYpPzhPUNCMVEakDh/RdjoWaSelV+6YS4MQBMf2mT3YAYsDV7zvSDP+SL9dCK8aI+rzghU9z8IXQfBjTQlBoEbRwJilGOHKrrCtG3IVuubW0yXIHBYN6KRCpQT0PhIRoq7xyvm+P2RRXeEOvaaQ2vlTCfrw7IBhdnNPAD3hVFY9NA+Q8Lk+RaGP89zOAOxe0vEV5kY=
`pragma protect end_data_block
`pragma protect digest_block
67a960102431d9ceba06be5b136ab5825e438a8b8a4a89820c78f5a29b059050
`pragma protect end_digest_block
`pragma protect end_protected
