`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
h4HDeC0mHk4P5VD+ljxf9sMM7BMBz7GoWcb+6Y+M3L+XzB6erYfofK0GQqX0YFheNvMBA+hb6cXZJpbAq34mgwtbslIrHQY2fQWtLILV4MivF9qBor5tL22537MfaKiIREcffVnz3pfxlvsc53YSEUMjSqeX5NF2cUWuU9niMxqMJgzPkHz0lMOfjazyp5QaZWNplTR8a3jEYEPfYQ5dddNZeq5sKyEn8oehrT00qJEnCaAIc32rZlJZk6mor84pQlNNMVlSb6osrxHnUF3+blrQ+nrpF30laA5D73aoeuK1O3Q2ehP+QGRk3ExJANCHYm7SHHzKw47kne8LWCm41A9VafDqwo6eC5SDHLfmUrIdURZrJXGTxa8RHE96dgmI/IHLv7HywbA1eis+OAotK9Kc91ULoejiXaD8tiKMkfTqBw5Gic/XX7F+faXSMhU6yjTP2MYPd1QRjEYMrrnhq6/4MQRCe+pdbgswUaVWCpZsDMmTg9vf2z2vg2RVjt0ZHyl0SnJKJDKqqcGiGIRpf1Fj3rY8zzsrxYMt4Z2O9M3EAWZTSGWSvvTzdrBrqkAkPCpXRalOOjNOfPCUsfi4Pwahw13RBZ8PyJOBZGYtJh8YiMPcfoeuWBhl3Jk72N8Y1NkNgsBnW+jvbQ1fXAnqZmtx2KsJ001tYI7Qw+Ji6lqbTfH2iStR+sQ+/stm4DZ4CKYCQ05MznLCgH7raDvmoEDcKrs+F23hm8EiU38uzRDgc1V0ZQVxqxBTMBUmx82lYv9RZOdaasj8Q0OawYRWNvgAzG67IpEYM4TO/uH4YzyKSgv6a3hetaUi2n0M+C6DHy4I7sJy/58SlYR4sS0ViII8Ydijmne5VhHUmQH2PH6eEbISrJ8zmSWoHcZoivgIJbJ63GfOpWFY754NIIzDQNyA6V/j9U2kX650qif58Z+6TEozqIhdazNcDbrKn0i8+mFlfJqhU1eTkeRpZ1qVGF7Yh6PzjV8/Z8PKEBPN7mu5eD0TVaPBJiVYm5gyh+/6NDtBzrGxJb/4ois8JMlBmpMz2I0DQuLQ3D2H3kPB5+mrqzaLTEn0NKrGUF7dgLMMz71jSIZgbzb4GRMT27oss66BIDlbu5Z/Q4u+VO1Cb40SRNhGc9lIVVEwFAxF1m7sB3AiURsMBLiNljrqgCsyNMASZA/iq3LmlLaxYTtZwQm9la88kOC5e2F/BA6c3FafepzP6ETHEitr+cCNcXPuUFcF4Fo/pCx+j1+QGosbtX8RTAAeZUFulousioX26lwH8v56hpzojHAOG/W/YoOwCv5JcoC78j/7sOiLm0/9Z6XbL9ymVouOmGyjTBvngq6V4ch1k8Lumx8CAgHL73I2ACyfPAenfnH1D4ET8BdwiDi3LNFDyhl8zvHRto0/tX3VO2SOeph2/MIfk9O5dx9hNj00tJC2oDT3Rqoexv/ly4gEkNhOcrdeM4SW6wmYdtgyTNo6GchyQRrJQO+GDV/rjOdOgXPnj8MI6pYTX6G27Eo175Hi2Pbd5C3QhJWwSXovNVyoArQbclVl1LzEtB5oie4P+9cXrjgCDYkWsgquDbi4tjqSUd5hbmaku5S5DVGBPEipc7El5DnMsgMOZEwpnpxyPA0a25EWYd+A7EBv+W5sjSh3+DlKS/NatG7WpD4ZAnT/uvXh8n+5HhQhzJvvGTnAAxcVR65jjUVbBYdIxgwx0o8IJUDCMMbYofwKxWgS7LEt9Kx87JqrhehKo5L0hADePp40XsPlN+u5wiNTdiCjF+SGHp9I0bTe4joqg265f3Kr9Dl0JEF6k0TfcxevSEKSa1G1DLlPRxqurlZoM+uVMtq0q0brrflul2LszeYCbt4PNL3oatoeOjA1wasVLKMClzx9996S8jZFjL9snZ2Gs9eGmpih2yPOZqszq44ps+gPwu/tkacQYbIAFfIXubCyj+asJ+a/Mm4WY4o/5sisKMnqpdgCBLv+Pt7u4IFTLtrPhrwMmmmd5nVbjElveVEgr31a0+FMKQLxpSnPUCWBMSb+yPZEeCF2cPrGBruB/ptpHsJFKo7QYHbgVZBu06gjpUULZzGd4ADfZtDtdkbicW8x5BBFKmepVKR/PGoWdf46CwuQ+3k68UHXfJH8qWWLyaPSNodHdSk5Wg8pVdYhcbmIkQU9t+Zw540938fOvHfs+s6mn015tB2Pt9RGG4/H1STXELJxX6XnqMXUZbtF3BG7/0SZdibcvEvqRfS6mnowVH4bty+M8izovJYectRelU11W0Hd4/0H7+O8XSPEpXrWZ6Tl6spnkYIERWhRQIRLVZN72weC8tK/khp7KldmKXa/AowwKs523KpXwPVa4TVnWoRsxzjjQHW46y8ZYV9Dyg7yNTxlrtCok+ipYGz47qA9GWog9pQzqHSpe7apncf8RGVjyzUd94w3Up6uc5x95PhsTTHAKpKwEwz2Mmf0Z3GeX9ZeCsScPmDQTKv8M7i5F4y7tVwCZkC1mkuy732d5wJyH6R/1bBkTudra8QV6od58h321d7YniW9oB2n5o3B3Ri+cTe8W3NbYufB9qjSDVRJ9I9oia658C1VoCTjSEVTGG7JWE12lr0BV5OgpITKOiVgfdqIWSG8wZhvQvIdEYQ0NtBjwozbrn4PF9grdlBItXB2vlMKEL3zmCOtCYn3Hpev0hA2/HaeLUAD7PSt3N6/D7WsMHUMCx9g9jsQOWdfiY1SFdCiVJB6B/HeVgxeHsIZo15KAfEHHy369zTpxEoP1HDk879QGUhKGY92/4vUY7P7D5873SaIJBvHAI5N7yEp2qH4WPxN/5jqgfzdQ2rc4KZM37t8QjzDrsUDfaVzbwQXldi0vfbmLufC1C0dY50Tt8gygWymK4veHQy9aq2hgpyv3kpWzDXU9DdXkMC7OWTc7jsqfClpuA5o8PzgMYFTEF3c9o7rzOeALb+TeiWhVpFJ6WMG4+ueJAWCDKY+s3I9ICCcF8ODgjsSUvCDgO//Ck/jY3EDwb1M7c3p0uhcQgYsaS+6v2kqSO0dGJDMe2lNRXx2sEGu+m3bYjC9iRn6dQkp8q5X1R0ProgKMAKf1T4rETJoOcvwuWkPMPz38cmahEac5hW8Q1Rrnhi7cuMQwKz1A4eb1soiK9i4PcZOOVe29toJ0z1UeINWJtLwKQX9XvDsJAQYJ0uUl7KRh8OOP29Tmy9Csf644AzPaKW8ro6cYIw0Eov0rrA3QdljMHq0ncJ9nqBZUh3l+6KaYtpnA3iAuIRShZ3jTMx/arzyCZm0JF9siW5vz+0UVEb2UYO9uh5ilkuZUBF53M243B3W6+LOqy9uDNcfqbgQoDcDx6B8/3Yt3qH22AFvy3gS8Ny3Iw47PJ05lH/bm4B3by7dqx7Mt8qT9DJ11pq3mWyc9F3izZd68OPTj+6nWTU9MUF+qfj8f0mTogj2q+oUzT9mMkB2ba9RyMKtBQwO0buZbGu+MQ8Izz5aX3U8tMvCNTPLvFFw8urB+T03WGmTuFit3u9YSZaws2xlNF5Xkx/VS70qKauhObissfsmRwsgwEHok8hAc7RzmDimMU5BdbR6KHEoW85bmCL32zqE9swf27wcteeGt3sFYYka+h9k/9LhAE8flxa29aGR2T6w+7h0IosCDadoOxhzFRs6o7SPrJ07nJ+Q8qw7LMcszqSrIRru1O0yenUhKVhOBou0PpKwkPRzWXhAhsTScm4ix5tTnJE4WibdFmuqdOGoQk2xKn6O+5ALP+C75eST4Fs1Pw6Xd8MNRE1OXJHfnecXdtK8FidXOVstUQL8fOGOj5PptwXJgHwUcJoYGEUWajf0qTvBpLfVufdtRLCTD0rVgEvvGF70fJVa5ExDJozAtC+P1N/VqA+H5BW0PMM+s+3YpmZ4VSrMpbhKgl2Y2I6pIBNT/fqO0tW1JYhfcYgHvr8txKBhjTqE9ycp4Y3Wqx7TUz6s8W4NwxD/1+FAeFa/z2zHAfwwTRfw3zLng5qxtjQlme1ZSEobgZkwXaZdEFw+xGGJNeQkJBvKBDUJElP5oXIqdLpJI7eY+oz65F+40WmUsHEva1IZQHBFnJxsMdZP0oVrFJopfBt1w4C7kKojx6tUHlPk5H0yRKWYxgfYLrjH+xaZRzyr50vwsWPQ9yjnmJ7fdRZyfEr0XcDEmdNQKQJSTg2nns0dZQ4EK9J0pfRQn+xjcHSdhHx0juwtdlxWA/UlPCJe96WsyJjB2fgbV+Yt9j8WHQpSYYZBDIWmK3AW1D4qIjJzyK8oqkOokjIdv656pf2GA9QQXlfxWniI2ikiVHmwZwouXANEIXyjdNw4m93M8pn14aSrhtx/mkSvnqcyHRID7jdt2mjGkhO4fvwUoeJW+SecN2GKDMVryMj21W3EpVfm6v1uxumUETLlNipVz3yOvP9mLNa4svFsycdueEDmcW2xIt3HI/qr2xJ1/xiquYhSzEvENHFHJPFcT9fDW5lCPG9KBmWiD/jVlHRa54gCQtNcRSrLvVisdEFzm0n58H7DEQjlcB05s+q/fapAnKXIPKgnjpwJjbNn1BdoaHHMKEJQNwobiJLUgOZOvQk7IcDq9FsF2Hx2R8p+Xzb82ygR2TzXWrAKwII+wJ0uLYxJZXczLUMW9NJFPmBcBM9Ky3JvqFD/yTn+PgjuC2QFU3fle9t9gVBNfoU2rWNCqs0GuVYy8jJSwy7K9yoMnaPgGOul2S7UI0Wi9LeFHOzR6v0F7bKiMc4emHWJO9v4C+39Dkzgqyp4oQQnVqOF9afnzOrwZ0bv8SR2rhX0pxZIu2819xk1lkVQxixglwjMyT3i5ZXWyNUCcvY51i8xB73LzF3T+JQAoSyyxipL6e4uzcC8JATpUcrGjhcNaiWV8bA4VN/H6gk7ora1szQeyGnZHS8FaitDq/gMs3+1iIWZdlV0QrIBAx2jmnpdIOIJZ1PoyQ9m6UvgS2Ns4+MeFPSCcMmmwfnKTIJart+eXGTVazvx18/HIU7u/p27+w9gNUs+iI65XZ52TjTWonEaFT7xJs04Ba+t6Wf1ttKb4jC2drft03P8L+DHM2uO2OK9Xnbe5m5SBUi4Y/AlZ3Gb6q4dOvH+oQ2MXw955V94AqtDt9HPmatr6JALT5ZuBRN79MDvoJjl7Yh3d/E8Q95tpz5C3qhTjwoGI88GdOkgM34m4+IO9P9m0Dt/GfYI7NoNPpI2Di47hz9YRyd9QyKEXQep9ys+SCGa6/ndxf2hhynFy91pYyM/jvVy1Q5ZFt/3bBcUugRAPJ/lPpFYs378n8LVvRhgCCNIkiB+JMJF4/Pvu2W+R0AQp61jj+/18Igikl47KCtMfiENeGPYxhBJbhWrQfKvOqgypZa/6bL1PNG/UhhX00bTWMWjtEy+uQaHX++1tRlMyGx/ZNPaFyywqGCKwPiF5OeaRJ6PoHdUic9ujY0Ej2lEH/MPSgAWnVnHGA0OHYsipAteNFyD54jXB7ll891QABrWLftBeiyDmS6gf0kwJc3rrurMUW2VNeGM0xnhvaobZQdntjJh3cujQvXgSWjs1RIlqwkVc+7US117qoU6cYNbgVxn6TJRlD0HpPbC/Hyxto5AH08KgghfowdRx+HlFdKklabvKwuvjU8EF1lyHcsY7orWLuywqt78mKak6Q/BFUoxOguydyKUXOwSILNWnarrdwTo+s+WiFUG636D+hYyFLf/kZ/egi5DJVZj188KlgRW1AHFRkC4npcCnxtoVFVtnMpxr+Fi8tE7jK8TKpjD48KMSJYZlsyZsN30JSl1b5ZxLF5YiJEgtet2KSVNEtE/At5eW67tlbtF4aEl3m1XnQ+Hn+IjU9TQYZZEvSJAU5CV8pok8uKJOn30Wc9HgtsMmr+nqycZTQhHDIy695Jzwj30KiFj8J2pz252AWtSkzynvvYeE/wN7l5BF0Wct9gB+vrhlAOR3Kh1oOYGtuWQKrreNiKbdz3+qa149kC3fbIODe+NnOxjLLe+3uZnr/YFGU77PLwKggd92w8bVLSFjNoxnmsI6H8ohfj77Kkbi4jC0kSqUGdPD1DCbZAPX0N9kwO17uUr+8RMsXrunzRndP0GoYXnTGwo7pUyK/xTXuUpk0v2/95LOkZkft/jySvh0WV/F416yieULa0wx1hlhGPZmHW0p+kukWNcTI9Ppx0XjfAHmz7ShtosATV0mqRObQ1nj3vmjm7zyWXlH90FFZhDOa16t3P/UOIAevNRW31dY/GTQa2q2cdqF1x1dQg7jOemovxMZwcguq3S59tLEd+59Ftqpe2Mj9wAZwuWXcxtq80KLkmVchVu/firnT6+dxemGo5XUz8zNKDJm99HxcY0etyiN0g3qFc6rdwtgBV/xTDgYamcp1ZVEOoEXr1wPB3HawtZ3Tu2Skpgub7+nVwTY3D0NGMAbG1x4Z+eVQ19fVZ0G59vtHKtOBH+LZPWpifWUCJuUDYYrU3lxOJKS5Om79VBt9e2qgdZPeUhPb7DqTwkkbYAz1surQJBblMHYyqXjjt3I9OD7gDRM6IQIQo6GpF4XN/klNj26T1dWFIw+V+uJ0A1iEqDFpItShWEkTD7dbmRlnuAwJDXZUcpa+DoXicc5ZnCZrgzhlDA7o5GogXhUkg7rZQ30VEQmGJmGcxY7nWB426mte17vBpS9/TOsXxOa2ybY4d+ZXnPRTebhIOlZA5azvnrLPxBc9V5/QUmyMJziWO6klr+Lx+7RCmmpfEGyJxcSHRkJqLgLt43WGgQQTfG9TGYxIRtYeVZAFmtg11BQtG9/HioDy9y8O2ji+UJzZubAGRkNd3nW+FWH9/5oPjXDMyf1uWyxS0m0/HcDOo7607mJuPWQCGaN+E2OL9q5E/MY6qrKfr91w4Im26J2Ww2NOTa5XJ4Jn/TfZura81tTobajlpDUbEREHW8FQ1tIMwEGKunEgvtoP1/qShK+IGXOjlvhZw6FDIWKgCtbDPpb3pNnaNF1DFiqzJUrYMQ3/legXQPYxTacIjpCtyululNU9eF5lyI9GhvtAz3HKRmGwxgd1qFCEU9+eh33z9nCYPnRajRJV8nLj7HJ1uwzEVTeSC7IwIjwum1SdQVcJ/ZQnz8uF+MecUqxdPB/Ro5tlbSXH508dz9dCf9Holr1D5GqCfSBuGeB4dNbAIVRSN4tpB/0voDqvgP58lRJZkXVhNN/e+q9D3qA2bRMXGCmgONp0SQQAIKhQK5polYomv3YwtL6iAsqWPuWuBTSRXxSSbRLU/fse+MMYnu4JbtQy5TLNPPPXzPJR5CieroAT/W78VlBA+NsG2FwMKbILMt9cFgmCQRMYb7Ai8C7Al+2snF4AogCmUB3n2/uo1Iw4BQLubwps/9ksxro19EzgPqqQ59lD3c2+0rAdIw4n6wyzOJvDsVg2eeGW65huhBR9e9ZsrUB71ESRQz+GnEwa1aZ7OV/xI0f3l3PU4PFt+CHAiCQDxi56V53CLByAGgftw7IX/g7Gp57606Bswwrk2F0vWJDqo1YzWX18R7koomo1yiy++v0FCq/N7GRFHhOYlStXMeL2oWajP26RMbujg1ISPXRT3gG5ZnoZpj+JyQuu6xHkmC9A1exWcAkh5zWG/zL1QOl1rfogkv7q+1Wg8IZ6KgD/dPx48GIM9E1kmx4IDW16WuKdZsy+eX9XcYDtb+l1jCTnVk0yNQ6pS0jPkaTjDlfPzZA+WAMWA7o/aFnuHgln0E2JeflqR0wO8LYGe1QQiniqX8011CdtAj7lN2Fbrp6h7zWIOxBSJ/CVTaWEmnL17bF50xsLITDRAMRdgMV5X363V2YUikl0dCaZ0bKfXx6LAe7kkHO4XqEp0MTI9rnXGAU9SINfdCa1RNDGxaS0Owse2BN0lz/4xQg+XZh5fnBC5qXpMxcVg61kshi+TZ+MK28NJ2hojGgF9JvszOc40H0xhNx8XM1Cd97ePc/S5Rqx+JW1dZ0Z2Y7AbxNmQeOZpvfRSAQYqI4R92rggN5KwDU6pcdCZqWMZKnGLeKTcFIDy4ec9655TwKg88ixo+coktuk0NayF1kL8CIMl5G5ulZ+xl5O3A8YvX7TuyHlPDBgTCsXasIxb3xWhiIt6CVQMH3tDoNhmp6vcaO5HW8FoZFxQoJgSCuFUbaGjyhcDmhcBZrbtpRHJxUHA8j389f0kt0sE/jsm2fge/fBYU8eKxQclpByNBnEl+OV4YU6CA2RfmdH9+QNcYwGDwWw0CBkcxFThau5vG1CiiQt2rCFE7TtIQHtNVsPNnWcCysJtoJYnGEp3LJX/33MCoDoGqaFGvGow8IBo3krrZDR1CQthl11PmpphffSvNTls60AxbHX73LwJhFxJWsUTzyb8fAk8rMlqZR46+x9T5otKhhFWFUQpfsX1RXa+1myYWrIyYj/pUC0WGittEDvW6NQw1Exxi4Tto7UjKTowTslWAdyyE6v8Mb3cUGQ4880Pb2f4shG5yHtHSW5CiCoYG7r/+a/lp8XvByy/vx3Qw4V80OqFMJrGApAKX4EgU6KMmqg2/wXLdZlR8eexv9yRPLt092NK2OBU42zSppEetTvM2qD+SKy+zYg3WRVF+uhGu9c6VBQU08vS3tM7YsysRMunGVQ1ZPRryizFDpiQYuvwLq0Gyj+RU/P/CME64VrhPcfGBzIwEXmESChooDNVmIme9ArO7oUofS2dWacAe+bWKHd6aUWqH/BSMA/i9W1yn1T1KQUXboDPzCK1QmjdA+zq9c8+lV15bE+s/zoFLIKOYKiQ0ftyZExy0PoEViGsQmD5wc7YQHUfjUyTKp3qT15rY1YP/atZXb7iWVt/ZJUtYEq83WOGtJM1FXOrcfKvaplUzLReJ6RXUvq4nMDfgnjaEPJpFx3P/PE3dpcQKiwq2L6O4LdRS3imfHZwzWqixfUSOjiWtETq/SUD7T5jCbtGkt404dDNHkD4HnhxQepl3HIAGEl6gAyCHMr1mQuepKG/02zEu5diJ0W4keDxRzvAdc0P+ss5mMIr4Cv6Ixde0zT0t8RV0gvudt5PuHWPxczLbzplqmbiZus3CpAmmQwm/1RAmhGXIf/EVaYXSeq2QP+8QDCW9nT+6Eon9AW6HrnZHNLU90e5nqs0uUMf6gvX0A3y2icwuU57K3sM3oNrnGpwNAdYprXAAb0SXP1LvgQ1o1M7h/vkk102tTNCt8nBjV66lAjiiJBfIAa6UWHQD/2B8bDMFYED73Be8RrcZOszUISt5q6PuVYGAO2O4jBhl05sx1dyhW+bLcMMzz3ZjRpxVD30OQu66L0BbL7Ea9iGEDN6+dX3I3YaJsjEvGy3SxsIUbydBp4Km4TKKlrp+6wMEXtl5GiCU2BZFd9eTItO3SH57IpcKjLRsNI5X/DLg5nJFYaORW7DqazaeHqdOFNn0SMT4+4b4uM9vvp7k2JEGBnjBbAmRjDZpmh92tIrWVn0UEWGn6DeFC68OGR6oqvgoXwzDs6R/MIks1GX6LXoYy1omIQyh8jQktm3gkvIUSvybwBCGmXhJ55QQkInIqXBHeTf6YhGI1QY826Z6feXsK8DqAO1NrBejn9oaYKgcJzMhkS4GRWanAbw5jtVBU7RJnx05vijE0ooM7yP3pMxfY+Yu7HM6OnCdeGQZ4yJRWJtUyZ3xofuwQJYbGLZ5Iye3zCgrsminRvJtChPmnCvXfx1/S/ATy8jyXvJ8iqOISUfqpQY2RCXB/uqUY5M7vMo0WW6xHuukFZWt43QWON15DBTJ/zFB9vJzvFcyuZ98QKtr/6z/M0j1oAXYeq8hNMAk6D99NYq2vSKbMnjFDFs3naTmHnp72n/pxrYg2fuXN55KZwfYe7PQ3DIyhWNvcx1yy95AYKr3YykJR+xPGkcIxn3+KxtAEgvFIfgOnpou7V8+1upIIYgqlo2AyFDFY2XVZmfQNoVkmuea2/9IXSopZe8zI2hRb7S41oynjvD8q6U9vLPoy3aUO7aOIxIJf4v3aAEHFEuSGylzsPjv9RWF8bbqnfhUCQuumoEnX7NaPygfClfBccVVFZCrE5vnmmYkE193jTyUGRlZz7Z0VuNGWxUXVifCNeYl0ng/yQ06ZMlPyI3ZmAK3YUlQ9kJy4hbLzCxHP+pdQFZU/5c9l9imfUdHWCvGzLoA5Ca+j2DTbntJSAZXh3UaXH/rjEZDljj7qVp0geMvA1x1tqE6BoVWKpuBtFgPdoUjz8OqZDO6xDX25ue56UHOPuNt8wekdCSFrokRShxHml20KaT3Z0j9y4+IXLuW/qHS7Y2slmF/4ZJcgjiNzRJL2WCUyMbKCQvIvVZOwbumrA/9S18oVz4HQF8uwsPECt8sVsiCgfObbTQp6uXw1lR5ecimkCIO2j6sBXcsJdqQYGWJx6AITVvisn/XrfN5dXy/3o6SAPausS+sXWbpMEnyFzGuho+eppObLX+7gyvysbjnEKesO63e6yLu01jRPNQwpos63Ojsuaii4lTaFKs/vsTfYZYEQqOIjYA1lo4gMX9gBcBliGkZnbUu0Euez2tL8NGcMrYbvNETw/pVqd7fgS8ysAzkZyvjUYy2fbfqsBUb66cM0Eyxv+rUdYCEevnsvASvujMI+rw7dwHtVf8TthjFWa8NLSllWXITGc3r+lXko+iU3kjDyW6ETR86PCsAjc2z5tav8l1besik3d4uLLTHwXugtfj/NbI2ba5qh+spn4RbW641MOQm8OP2zmGctUJ6bzmRgHi6QcGWooayrDHeBe6e81u+kdzlYXl23NfODeGsB3pJlLbfSOQkEv//u21B9Vv3dOcxqCLx1PtRe5ukkmroNHVsH5NjVslduyj7gd4hgMcEWtNeNOCdD4/S5rgI984f3CKjFQY2IFddNklHM4JGSLmAtIn2TcZMR3qHF/Nj523zJ6xLDFUFcaS3coe5paz39RhymaCKA0G/NpdP0seUsu/bpG7xfn/FwpYTL1Cvh3DQkZznAkT4ik/xc/UMrkAxFnOUnFJ+sArSp+pQ0UoRIPcSV4oFiuOoCzbAYOg92eyeGYf2T//9FPvc2NMQ/sXmoH2HuEGCSgefsCIkWsoYb6f4O2jyvJAxVXg3/QEpL17P/9F/7/8P7RMOgaOvSj70JK62zbAWbsrIEprM2o8rpENUM9F3uZit3cIpXvBoenXDAUhu2ZWWkjx0MkSPaJD2OhE8dpB5qOTgyQ5hkqucz+r908+lYf3DlF+wkU5czkrDg5V+SK7ON59PD8CQOOoIUZs/1xFbiCT38Dg18xUeNxgfwKg0tlKABrKxmA6LnGnPDV5zyufH9aalbKcUGj//KsytrtphJ7ZEzzjGnmxqlB9E7gAMnxWwwvsCICdu9jJR9YXQM6LKGf+FPVK2+OHiCvIgiVvi/LreAG9Gm7sYdMlLjOmheXJkVwRnBjjj+ur4KiXQNS86eolXNcLnEKeuOTNCfKhevvmEzoVQaWNXZUpX1A+21RlmIRSwn0gVx9vYBguqBFZD3OBZma4HY+fLqFmhZJVo3JUz1PFzLccE6375VzNth4UWWE7Q6JH4/vE0H+1vgd3XtSjgxZI4wWiSf2agEMZigs9oqZyw2OFnXDWSKSiZaubsq1rZ1fteyWxxIs95sf2ANOwRtWO86jKgl9FKne2ofAa9F3xGKcNwB9AleXbM9YkhcmBM+q7ajyxnOoBCxFyvPp0Im+tgz+eUVbTtt/7lF3qL2+EtFthDayTnpSaZFk7dOlYpllicIJl9FLfs5rYkzL50v5/zJ72e9MlutmqVyq3IbalFSmVAcrPzs5pxLpx/rykd93hHtFGXnxvlCFXzwpiy79VonB/Gx/ldWwovmJHBha+47AX/GSAD3NCEm5avMEmy5j69p4EEDFij/8UdE5GbyqfyDnkdSEYUxIphu31Vw8P30Vomu0Kjww4PgXAvqzUSi9Yk+DMNwsaaL4BJRuA/DqYLvxnXLWd8P24m4PbS3WzfG68HULVkGWJ8yVjQacwT1eXQXTlIn41WEw1hsjfVQk+jtj9q7xvxY2JKLeMUKXr9EHSID/Pgm1DD905WlZTi8qKyCjL1PazgO4pdsIDG8z+fqsj/Y9BYK+spQG8HmBFGGFJr/tBcv7caNTc3jMKd6cmaY3PNiLgVygyux6AQnvlqo9fhQqqjakX9DGIA39FiTz4IVe0Xw28SzGj6zv8KsUi/5jHu+IqcpIdX4+SGM3ZN8NsqwhwmORLgO4IVGdoU81DwEsHzobRAt0431CqXcm/Gu/GnM8Ecq6qAzUOnD6qeLnBeGcfOl2KaPtECLbTQNB1rCoL5IY4mzCWAwAiFppjL/kc358IunZJGOgsRhiouFWyz//VWFTfTQF8t4ELHcQi55mIwBUnoxjMBDoooBywR7z4MWAPfeJYDB4BNPAwvgZz/qj5LTguEdxB2XR5PTt94OksUUJv+E55GSmCejicZxIWaf2um/qJb+RHMDllYVthMTK2DdC5sW203Y4iRirOoKikS0zDM3jJZOv3f7TSJkV5vA4YkNZKHTHjGMFRtKwJinmrcFoExoLUGPwUw/SkyjG/uCITHio5EXonNvdyIKEBgtz20PLXft4aEZFr9Nn7yVl3Eh8C6J963Sk1fHJk8j8oh3nWguOieTAZYCV9jsyEIx8urNzYA1AzSwbk0a1Njm14EdHOej2DhfbyfT7raIZA//+nMblOGx3CuGR5UkBNQ2CSBpG2tVNaUc0hNpjvBwTF+FHxTAqFzQ2O8MPMPS9W6yRfhH2KcfLTRagrFLnNbbA4CjYJlYYYl4P4r7Bcl+TNnbllXiwL+4kd1wIETqYAq2GuZiGcYNJuyl6//VojjxI24ohQTh/XEPkjqt261/eydkH5XJAYTxZ42JdJofUv/7L9AeFOCcL/A58woainqQKvS/AjCf6LXQYr7z4F+b45h3Yc26895Me+YWFhkju7k8Ey1mSuhtYUwx6t7fw5lvsI0ieI4HRrZgBcAJEhAFYSgBMKzioKSYjjIEjrmAfTrMwbI+KmqtqW7Jz2ewyL4wk1TL/j/A7nCIGSYz1Ld8zznJOW+YRk1pBRBl+DLOlfn7evl08IHAXyQDH4yp9cU3JY4jFnrMkRE4W2xZg5DuF3ifr8k0GF9osjs486PyeYE1atvwcO7Lwg/b8UkE21ufc7HvYflZNd6PI+XRRvaASNTYHy31W2zK2re8fgSh6U/STCPoj6zvSnQKlymzXMdqvT6wpLzdme7yysFTgsOLxn7tYqrhDYy6lJcoUYQfFvqbL2ucNt6i45VvXLVIcGDlO+Mw0ydizVNhkrEBvWlWZQfEUh1vFC2fSwG+YP8GnQ8iihNwf1CmFyqNp5p9h/YkioOYti64hzRX+EhE/Si2Bzt0WZ7Dkn28tKKfu5e1LqXr9YODogREC92Z+0KQEATX2HkRl+2HNdLNbUI/Ca1CJwy6tpdhVSR4HNFsQNeWXe+gMyTfTLhekO2jnElYzRQN4A0gw+dZEgWr0H/JrGshiAuF+cWJCxdcVvnXti03DNQ2soiOD0viu//mwFnrV2RgYbAMhfR6+AVBTUIlQ9uXBxVgEfQVeYVurBnAn6gczSGsibHQY2EtZs/8sgGwLYac0EgXgbPHTPNlwedQJQI3a6qc4x17ohuFlhVIQ/MI4RTow5aZAUWRWUj15394yV4GQmg6loGp0LvQDxqZL3dEB/6aTYYjfI0tCzic+SGSOZe6y9AzcyKbtTbb3KuKr7sS7hDGVC8Qj06/v4OW5VrpheheISJ7Ihjgc7IlpJF1TP5/dWaiHOqjULABBiUTOKuUDhkjdhEEbT1bbuz4EwEEam5UAWy6vERkP+p9alPV28PIr/mO2im+mX8KJuaXgM63t5D7PkScix3mKjOr/EcWDgxhhc+dq+wLhZpxRq5QI86naGDD8dCDzKjbuZRAGRp0Xo56w6lljdvPT4wZ434G6Z0WCVFGy7ue9oOhJmNdViwVTYey2zj5Ld7oZHTKzSnOPJNQOibZKAkzQ4hB0jEpAkSUTykr4MnNEAaZDhhgv2xFk6W7Oym7aCLAMpmKX7Ejyg4BtdX6ukNmluEpVHGqKHs2ecStCIbjLOlYthFqhhXFvXuq+caeg+hcSOqdj6f5p/vfcM9Ek+I6mDSFJnx9w0xFWTVWyVeH84BMy+OwxvdCmjw/So830TsG9TrFKgW2RuTQbK5r5jYb4wv2mm3TXRARHbX+cyn1oJ0tMnNu+qs91M1yRV/ivX3PkPc64Yy6gRXF8FfZcfc3eUfRPd2f41IYWrnzt8p56yNLwX0gaNzi9OxdSq4CoTYVuWWUgDe/8Wku0ZQ65zWsvZywjK0dqg1sV8unk33fkkQfzQjwo87Nnm68IMn665JDOAfcU9b5jaXf/YGdslvXhnTyqalftLQ6M2+aPaBCUyJbt4LS9jAqZ7lep04JknlomZL9PUgmyPlCo5DngC85fpzVAMexnsnfXY8V2HiRR089yNIMtjS4Hjf9BGFlphQDEpeVzpDNjpHn7WlKoD57TKanmalTEq/tElR4eRFs5I+Zibcky4rPO91oCOYss6UaZnBBNqTr90OTa3kfbjYqdrmTIOpZNoT8mG0kgBWTF92daoI77HhcpXziuWONC7RR1q/rDa+MCt3rdVqAsEeZ7xHBJ2DxxhMcYeZcMSXvj2ffLt2L+cWR12qrmKeIcu5q/ok89uiFds6aQa+fye4B+BMqJBQPHlTklgXC9peZGwivjCq7vSeNgICwQd0JgoFuVobhKroczEGd2vEpLr2uyFtwS0ObFcA/JVQkL5G7kY3iliRpOyjzFXxc0nSwjh6Y+A+WmL4iqQsfdjck16XE6XoWxkmN9OZQtvTxTQGPOfS8knJ+pCVy7+rXB64VCKJAkbVMfLZDIgUpGc6kcEk3RZR9b7rdhxWdsi1n8bsGJZTIrP+HM9kG9fOZsQdgCKJMtanXF5iM1xuGMiwrLJg+2g1qC0X7dt90oRuFppyoBxo3kYQH/sJMVHwKZ74+hktxOgDmaasb2GxYtc64qDzB93QP6orJoe18AtomIe1vccvlxQzvGsrViuRRNbgy/+ziXC60z1aIPy76Rham/+yL1mSh5vaPnMZWgRCjpFuI2zT1SgXLm53fBZiZYLFcxf3l2UacRn4v9oV3gALRPmtfds9BO/+BmPq15/0N11J50WmuNNah2t+RNBVdISv8oa+U9IwODcghzUCVlma3dkc93bhbOmi8tbwPbNfjIQN1qfBgeI/jasrBfp8h7tLQLhPZdcfm5BnK67IBfcomquCu4kzIrHxJ8FHZ+WpUffGa6dOw58xdm4JGbFb9bwV9ZtREW0FO6CGk0M7r2P1F16+tHWIVxIZpzVVtEEXlw5MkqDydd4yRjH+xYD9Vc6te4o4B1ClDZB1ft+mf0YkGl29xRJAodYCdCDrH0Ll3QPNK5TPrN9m5ap4ioiFvbriHT9ycJZzxiOsZP9lKwPpqhPsZhdoGRBgJU+PEhkInsMonI7Q+L2btKDPsSc6FGX+Ha/Fk+u3GDvwbgBp+q1CmQrmtMVmiijBcdJRG9EjDdd8XI8HBevNIGoMUzncw6D7MqM5UTpl7e5AOLQiIRBmfBR3cOmI67cuBMhppnchz6idGroeusMv0wbWmeopMDB48omjrRrK7bMBO/MIw3zuYIjw+j7HNY7StqmGLtKRlF81LuUA016nPR7UxCtHzGOFs+ihesHY8Ur6Zx1nfJEMGfEuAItKh6CO4bJx6e1gQG8VO+KiFzuCtK2GRWmnZf49j+KPErj8AZo8CsuMyCEiwNUvrGSld8MBhI1dMsDABvake0/uNZzrRhomvqVVOmNQSE9hUjvJ70C6fWCho1+ERf8fKr6R4O2IxK5zXuMMqdhcNdBMQwmf1uS+8Bz+WrWMKC/7tnuW/YUFHZpeXjy7p26oJlyec9/fLWQighSXFZ2cNFqAztpWfx5ahD/BM9q6Xr2ocloczIaf4Oxz6abvmUn/4hh9XZyDMMVrzH0JGCPVqU60FJNvMSVH351Ug6ofqiJYIsthWTVqHvl4pqVAt0227T9xB9N3gE+Xi4j3J+V0BXwYO4nsVmg0o+3J9E8Dtz0O36slZ/BwKbzsoj6Gma8AlIdePD6y4nVqW5HtGUWIR1Wl/0fj4O9pTkVUI6k3ZBsDg5CInB5kLAz8o40SjdlTbiMdOAN3JheNByPsmxPCNSdeVbcJrEPiGDCPi1KODlfNN4GsZ1pS4jkl6ozypoanUEXOmWvSIBUPMTfNCklfYdOZRWgS7JXVsaeo0CRugrJVmHT1jxdYSRaEdLB+y0AI2cDtCIDsfPwic5FK5q4Ht+c2s+OhfRaPzYgKSP4mZqbnYlENmuaL3I3/KUoxaralwW3n1K1sG5v1owh4jKluKPpc+d6Mfxpv2txMTK6JLFdMERPv7/yUz8ivREuQBN+GZkLWwNDoD4IORyaTrn4ACCPynmGxl348ONZ6WmsEUpUqEGTkdhvZ9e0xtHiuuSnd1rvneNtBo7kVec1kKzpgp8iu45D4A+Kl1uq4Hsbfyc3oYzWnoFbaARhuAjnGfhaoYNdwbsqZM3eELxnP4I7maVGABa+NnKvDaQ+fGsFk8HIMfraLfJlbTsTa12kJBY0rDauNzwIDQM+e6SjFApC20VUJGb72SG/C0uP1f0FzBhBQJHzDA2HZfLMxHPIW5odYIs7DpDnulPhVdhgOUlv3Q3o/ifWCLVR1w9cWmt5xW3qKUYo4PEF48Gy3NE9AeBekVP2MCyzrTJVrkirFQfDiQtuC+vpN25plbn/cZJUhqlfIZq40yR8nNVuC/7TLW657hu23JDp80uAL6nsdgD5+PcAU6Qyj3mI3oMLuQVIzA4T8cg7oiY6MKw+obJ9O/3M1j4Qrv8tQj7sinMxGSCzuQ4iNVZ0a7PiXghwTVDk1gK0mwMxO97LR+3Xwd5Xn02JBcvjT71lMotsnp31xWSwfDWXNN3g2YvziWNt+Dk8F8GP2FipcXCjR9tcGW+iFf43hfz0dZ3FjNKQIkc6e6VdeiE7/wqKHbbs5RHC3uK0ciKr2IkwBxDLhwD6+cEbQBIsHYRAYoMoDbPeSvi7+djMMJ8wnYb8c7CBxPdmK2wnXiwotZU2VRyGJ3Xb/ydpq1fcOOHnWc7E6zHt9666B6vaGAeqA7Bov4G2cUxbterp+et4CoEc4pbTy0C1kRdsTkq57AlIZSGq8RGOUxYxWsvlL348TrnBxvB9lRWFZsght/8xxcEmq1FeBAzGmA67NUPrd4e+y06q5FjhC7cmtMzlLu6AqD+Ot7lh89MUgWWx/L+Ie1RY6fnBuJr3M2Ca1G1B2rrUFRTfTyZ/kZq86nK7pBfnmrU/jGHaaECzjEyV0V6TFmqSzPEMQwQT2WOUAfXyhqzRbUHyknO2FkIA3u4RESbM717PEjizGGCptmxYSs9UC2JsB/azTfWbnWSdELvIu6vr9qPTytj6azVSOXevlcnegh7I8WdtwAo7g8Bu3iisexza6/3EdFhD22zb6Bv5HZPDwtZ8Tk3QadvDSTcmcidj00unBtta/iE8SKE0Xx/MZi4h+sK6YNZekr3sdEETI3ACXr8VI2m3PPiMTMRUjhJkjtaCGKikj2jhuIRNGlnaON5ZLWrwcSpIz+N2RlwQpBSZBgJ6V0AZizrpRQSl7wC7vy/t+ZX5m5QIdounBdb4iUXk37TILVQydJcAXdfqX2SJJW536jOfLG3xPyuTIV4lcvjzXZqRqru849VPBLqD0ytVXY70WASdpfDmBeRBcTHqnDBW817ZRCWuiVgJ6V351T2IwuZlpLjOdUvs0r60ncdmTDj8hiHQHOWXGgwGt3ruvlmeIle8BmxoFsEMDGqi6JP4xW+rVVBEXuuemEWWjCFtHl0ttRAymv4iIyQoK/hPYI6RzsrbSoAcyyus6g5YMq5rF+KZs/9zknUg6JYM33iMQtiDaclOfjvhVm0DfiJu3mEAlyLfdw6vO8o8lc3Ely6h2IiiqLuWKQqTzxftBfmFyYZeeWnq7m8HZ7/QRAIV3sFxkec0pSm6xvq06nBfUfj6PaYPxeErqe7n6P1z1CcwpEb9yDjgUiMjxz7jKnpDK7QVvI1Pmd5qKdMIAZmzrLEHcu9B5tIku0rrCBpQ21ezl938M65OXiyyMW3kEzoUgb5q6BBYRbRFislhevULbPHNZEBEpWqoXV/pBY+IUEiafRgVieEiHSXXdfy5r8gWcuikCYjKPFg9qAbqwDrxPC5ENyHCT1IsG+8XqfaOgiPCLHqvQZrGJbsaMhj7SAikzQDd8xCaQtBOIvBJiLHUQa7b1PStKCfmYmLr1QFZ7REVkv/Q+w/bGX9/ne6dDsoQ93NON7if2oWigynnsLBR5UCv6jcb3IroHVhY4P4P0l+2Ne6DS4EEYEeXJiLn08AM/HjCzNF0OxuiAsCNvn/LVUvWujF96aSaQL92I9g8u4qxI97nfMO9rXUjbTU2ZFMMaz3LhNO/6qhgnrce1Zn10Uu/I/Q4+VY25zqPXtIWNPolPjJ4NJyt7qz+5iRU6pcEH4V93lRcNI38pv5cCKao1aT+kUkqt883oFGzWJR3fTPSxQyeih0L0Ovo7P7S54GsPh4QzlgZZTxYI/ejQxbwY4jGuozAcoKKjSOxyZBAV/IUDABL0Y1wxU8DEtqXsFnK+f/IB/TMWiZ7FCL/2yMVtKQgsY9BJofRavHcuq5G8tmw8H9vtrrHk7bRSG1iz4Jb0XrnQywae2UrYNn4W7NTaxD7b9ODSVkiUOP1JByl7RKfreKp7iMHDB0sPxPvu80QY1iDMR7ghVpxkZ7KmZw0WP35gFZgCoMKpZIzD1mBISnZU/VA0G0f++vVOpwZMpHgqgC8M6EvOrpPjEzY93IjeKVjv0vEYcqI+p5DS6Wm/pLvTgWo+WANNHF45oxIkHgZjVZXoBftz/GQ7op34TDw8JnST0Uj3lsGKz3ZQyAxBun1JEaNSOo+Zifh2A4R/LMWvXwKy66OgEYK4ETgQGzi58lWskfY/Wq+TYPnwBYrt5P5P4e10kaZWw0WTc4IYg4YX59X56yJDS9aI1NfGGeuXbaMS2asZYJ4BrLHMtiMHupvnyW6I4Yp9EZO9H837qKW2bLC9eZZbO2auKnItu64UTwudB9QHBcS9fJkbtuUEPeUnqw6bY+vHgWRclcR7Q9cSSgAOPg9mPkPYLVWeEaRar506oWYn50yBfOU/+jAauLRgHT/wU0E/+AYDba9++niHL89mRrn/1xw9MiySSUdYyn9tzkj1H4nHtECDFq9IMKQnpDf9k6G17oIJ4rJ5dhNINofP5KbPL1L+bidu2iQehUf9GjLjQ2MvG2i9ODYf/zMeB8WaCnbN2YXbmem7xffidh6BBXvZkf5SR8GWun7TOlneDCrVdnPOAdiJMPHLzUod2llDOBBDrPHNmmctnq5oomoq4SepSOJTCBmcui4qIdZ/oXFNBKnZt5QEzAodkdRacN34jmUh6JVTbFnqRm+PwiZCujDT/cZ8z0MDCpmVuHd9DzUNYCw2/jntyrAH64/OXv4J8HBfCEsmd/YHGMWN1j+RNXx/ZGxFF8/V7Cw7f0Ur8SfPzCcAUcGcY+R/rXTbJZBEL6KpbxZuH4Th888R6qi2+pvoFaRk78Rnso/cW/rGEbanLxDziSwXtTYkWSudk92mH8q6yZauaaRNACPFqhNRmAgLR3sPT04rHaDDaKQZDv6K2o7qNbnLDWlEG8XMKEWinMh+FwPEHY8DJOseMUuVBgHivDjo0A02E58PpoWnomyIQbsP17W44s9Y/fo245e3xTmPWmKhi8auUlZWk+SZMjwnlpnJobCy99Cw0k79WriYrOnQmnWI6fFyo1BNWNeH2d6FVvcjWTp+n8opY+GpHrMSwSJGU2fA1JutkZ6suj0RxwWI8IDL/IhdTQzvLBgLwXTnBInRuhmWjZxoZT9B/pEYFQ29zR+o8t+YgqsVM8H5ZTGLrh3PQFnpALQeS/fhPH4TK6z/ISI//KkmIRgA6SXZeKfylhWxEI026P54uaXE9XALhRf6dICmdMUNnGrXnMGCa+yHuLZhVciS+KUrhKc5/Tmpr29GNQ5kIHxURxM4SjTjIWgg+jEstUkfHTF6imWqns4yqb1PUPDmR9VWFrLOODRiVWoJ968yhryzNxiBr4rubkQ+Q8XZq4u0CsoMtYE/CRmktMOCrxt34x4U5tJD+jP36uhBCOe8luvrxIV53q70Yg4eHBshnIM0XusTNrcQRT5mLQgNN6iBFIZxB3uALzDJl+FHsAGAO4Xzf9HI4anmVqxeyvqS3yEO2Ag/VyLvMTxSbPumkgD7OXiUMv/SUu90lNqQwEwS4J/qtJcPaWUAZ+6x1VTRSr07rypL5Lqpj3UowRW1TqGF1MK4tWXtYjqUdqGPvweI9hXd6oRT9wRu4VPF4b41Kw9x6LYpn1qouUpjwDN/pdkBnAEFk+aIowUVNJTBEVCVSmJN4+nU2LY156sg87ZzOtiR2wyDJLzZ5WOWGoK38Zg/z8P1x/gJUpF+HjQJfL9ePpxfPa5Axutxz6No6YbDXrHiM7Os74SqptKi74Y21gfHWVeSM3kVekGKxENonIU=
`pragma protect end_data_block
`pragma protect digest_block
463c4a8358d4847005bdaa5467e96bb0d4b2dcc422d7fdb9b761553e90480d2a
`pragma protect end_digest_block
`pragma protect end_protected
