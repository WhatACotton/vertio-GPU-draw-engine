`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
bBeiShnePt9IJWsXpW5Bij0AssrJq9hG9lDzTi5wt+Gghw+DmZnKHi35mzo9ExOFhMhFqK5GN5u239hAeGAueEzndrZUOi8ijPPx866g1GINr7L283VVgnj+pA4mWzo69x9Hl2JaW6JFWvI+TFsLzCgXpOG2Qg3pgfK134XuELHHxyJOJCuYWzAu++M0Q0QM+E9oY8ieWQ7S0xNGfUYXfovDwG8VhWDO2MDO8sEBExITlE1re2yOmAs3AM5nW+DCYq/UPhdwLHOBleVoJFxDtaz0/rj8DjK4iozbNuRYbqY99GHOlCqYRBkstXkf2bsYlfp2yOQ5UNn0VqeGFfyCyVChZ7fjK8r27sbWdOLMAvmgKwq3eMik8I3LdllbJo/a7EGngRAVCafPcH46JFl2SoEfUPyOEZux0gq7Vb4TsOwNJsBoM57EHBM8yF/fVbVZDV7biy6fZN5OmDRmiFcTu36831vUM3IF68PZOmr5tXO205Rn66Nqzqbg4+gWRTZxsSK/6gXgIbZnVi+7P4/oEagr+cn1WtqayJvc0tmERPCGuY2hX8X543nuM6W+PyWMGAOf2FRxbZw/CWQvS3dsa1hX/RCNWDaMF0ppQw9GjVq8fB7t5M+yI6pbhOpBzd0RkXfNUXGjVRCTJQPb5mo9JvI5/T8ltk9oOZzPLpnme3IcwUClVmpo6bBpiDd7p3ApStWuOlv9dEtqzyAhVgU28sQYEaPRv8cCleog/jx2lnhO/EFiIgLu21soj1Cer8v1dTp/6z9+XHZWXCKbe3BiBIxbXvAdV33yhpeoWGMuAeYgqo6SUVZSiN4HuuKb0/Ra2FIFBFCLSWeMhz7h7NAySVUP7ZK1DULXAbExPRwXHU3C04j4rVkLrHsM8f4CCqr+pTVNXvVZpOYtnqqiSPMXE8R9PDwalLeWokn8DpEl13OBbYawxYeTY3irZXvJ3KJllqPQFB75atLwC7ChsKAVT6avo98kWy88VJ1zizqJHNQeFvS+JJvnMqrhZb/WtrEEZR/3atQYjgy7JhSRr/HtzwCVolaKaNE21ioOGeFlSoukPwUsEtA3CPuV0E1iIFtwl21V4XV3k183b4FNxXYg8OehTnAQiILJcI2FkUnX6XgA4Z1WhpRjuUCsZbrDbMozMLJP1xwUynwK2nPmlKDyShWbeCyQag26pPGG+v7DhpsP1BtY76mS2uFtFQ45vifCEXQsg2Z/H4nKhiPkBRN0uUnHPUik/nwkZRdaM/84FdGqWhSWkgYi+R4GtNi1zfVKHDMDKk1kjpnBwZX+afb1nMea1VYFZvyBuVSM4Tyy2r5sIuKmR6onS6utcsYTMOMUGmLvPL3EzAYDAKUhPkL70Cafn8R+TwEBgi7pf1SEx37k9Hp2y4BiJpNC52Bu28+5UJl/PKUWwCi95iJcrT6laUsxHwQBbHhyX3e2LQ6n940mojlSrDpY9QqyM2VJzlqNO3d+zetezA7uPn+8WDvuI7OuDnKkHmnyvbQS1dEWIUOrddfYkwR3aXzpUZRhQL67IwBj98Sg/lDqOiPfW/wp4l/MoebXpYC5XjLi6AGT28+DncxYF/NtV29iQ09aX61X2s8ZUZjlRHeXk8O5Pmjm7vXyXvG0o5pzRRPSUOl8ljsR6kmdSeufT8O93CVRrfnCVLvN+vsxfD3NvzywI26JrcPsTxAy8T4IAZWhzIdInwdm9lWygHhW9iVvJ/E2O7UsupLY2v8xpRoa5SIXuUOGtRTzjpap5d+xgHoztQPZnKQIdxc0eWquBmY5yTRUVRofX8zOEj02C/wfOjjoAMP/xhpg0jvMBAtU/EKyafSMIvuJk+rYSnCgzAdjE4g3mwGrC8wnI2Ysba0XJp3HpXBEXNac0f+puvG4ChtNwHXCUo217WAOcXn99v3Mb/MVacHascPc9szfRXRa1ZLtCTICGN7OCcVucRznLGK6qYKgv4P9BqJW6ltJTzJPrW1MiepyNr0UMX3gjPigEG0BFBjRfT3EewMrlw1N/YxkXj/c6rq6pRC88Oh2j5xxX8BpO1B0x2MYTvRFwDDDHk6DSqG0R35WH4LH34RuftRZ30n1UDO1t4y37Rk322vmZuAcABD0tDC2+pE9ZVC4HiNeQG1h5wTrx7OlPmo+aBhfUhom9jr0ho0WPUPhuNWx9w+Rv6g0pnt9twi4Q3OX/n2WjtPuHa3MEz3T06VYk4X3E+lmQXu2plYu3KqrLqaMpXCB+D3B65U0QkbiNplr+0ssuy0v7LK6dkVcqm/aSGYhHkebu3EsbaIul0hPjAgFNbC1ieBYj2BG7FPClaNv5PMACoejgKQSheBekby/Dt1OAQ1CD4CSs0DPB4KJEfDstsMrjWXL8P40tAwNrkAGqmBLzUF0kW4ZS9OcALZQ5+pTFWJAmg9SVm+9FJ2L5n8EK+iRWhj2wuOqP5YXUDBT8bhuTGvaTttpsMRg6ilALIITnSDbOqeydWAPCxj7BkgO9LHYShMZKzWSiaFOBwEXBweUxCqgGUbQVGDwdSBmblBDiQ2yMg0zFgZvVKH697mo1OxEbp3LYbychQOuhJ2JEoNJbvMCBmRy3BuhS83W7PuJyAF6yVpc5r7CVTTew4l6r9WrvKdnYEUeiMm1SN4qsT8FRlyfqxO+rGeSY0tG28zuS7jCUiynP+YVw8kKe3JGJn+DCXfj98XazI0j0Q3hR9Yl36w9KDqaDfXv49K7njfGBH/qY6+LqONh/U9Hv0UC4zcln9r8q+6KS3/MTbx4jayJBgHadJQTD9XfzL++9jG0R95G/JIUukxzuSpA/sQpdu8j7fp7Ly264WI+fhJ7enwasv+u91PZSZl1eL72WmxCP2+xoyx36sySkD1iJ163jiuUP/t6fau5/uIgVlOQmpMHeXUmRGzeTKgnK4vi+kvJimulgqS/n48GhbMEJORVzSae0QPRON4DM0ZRkBZQN4SZLn+bV3bD+Vn8FBvx7a7Hb3oYXCa9mpHS3hRR3HsbVjWQb8Rirbr8pu3iKTfdSW47uI0O9kOFEQExDoaOTP/sb51hvt6MOdie74sqblQwFcEyvpsAQddH03ER3bPAnB1iZC/ygrmGMfVrC5/TDa9hOmFIpbUlUbF7UWO/zUewgn/Qfibtpt3gqfgn90JO5y9BSUrpVm29FZxX3iPbjv4e5FJWCXXws+rI2ZuSaSEvt+lhdUZExgTpQt5Njeg6dZApziwPqiujqpIaVNsYsyoA0SIRD8eI0umAcP9gFHHEVDRA8uviYOCHhQpQIpNS9d9FjhWeNr+0I1bFvOcMCTNVu2irbUh9oZB9k3qpxjEkaLN9zLkwBNK75PONuQgySmY7c0THem06HtOgYAG/EYfYnus/hURAOduZyLcWfgO3m8F9kVinpdlnOJXjP+eS+tFO23D62N8pya+VTKJ5CjDIX4B3ibQsaBLT5Be8ux1uv/Ks9KvD+em0O4lLhwB/VH1S9KLywqjqdIpxrpVW2Cm8ECmKzLFbkgyhnBGCXlf6idwFAOko/yMfU4LcxlCEWFs5XhjA04VG68AF13wfdCKlXW1fG2AbCRGyUS8zJfBobOO65KXHmHPrcO6OqwUtnOAsTqhp8C1Qc+pQoSQTV8qn8urDljSku6u+KaNr5kt7vhtT1Fnmqhy+FwfDJazaHtnWQvW3D0hnbNjFtDuVm7Fq1O0IDhEVJbch3/5CO/6ISvn7PCGFhswRqGymV4Pgga0NHnSWpiM5Vb5TE3bkYEoCyK288ijJjgelQRTXEXxI+Bl1oZEjAzFHMSF506IE6vKYWacS11z17aWFcx22k2ldVWli3jZwJfHc/HdMwvPnQnox75hrb9j7Br8MbQF24gjxnsgLio/FSVB/5f+8is0ViHmFWqa6ZQvA2MWeHKDvZG7Kdgpa5Aerq0GJOA7lCDgVNJ5wNi34hbafAD9GxpHo/8sjQ+I9rkjRAnJWqS+yFp/84uQiE3YuOMQCxxZgDm3RD5J3js2tViVeDfjFcyIRA48EJfF3aMV10BLSMMw/9OGB1zer+T87sCAo+q1PDAp90U9D4Kc2FVcFp4MKxAq005b6UjlkcUHy2kCBEGEvcjMnuvzVqxq/i3JoPTjlVQrMM6/C77V8DmcNwE6sy21kGmo/Sy/n5bKKarITk7DxwyT8kziD5rDd+8lVqnpdpocniA4dhXOVIJrQ5ntubO9NWZGB2J0StCOWD8z+RgcYhDyIBLpyiWvXGFGAK4s9J/FXvuFCNXd6bDHaeUGxFxbWWa27+IPQlEFG+LZ4Bcr4ZzAQFQyNDOIR8/XRWfEgZQUZPSuR421cJRC1TDZKI5SdwIeq98RpLal+24+gp2st1UyKkmR99IXMUG0BKUiXowthv+OwmrKXuVpHw+l+ZKVMp4v/AqSwEAr8votNq3DcsmrLE6U9YJS/YFNjbla8IhLp7ZGbniPht8aTcg0iB50uif4T/cdOcZWglSK37jlJQLu39W81YKyuHrzcuDijQLzFZjFCj5qyQ9tX+sOy3rURQNKXkWzvi9Mvqn8UePhIZho2LPYWBWXZ1mi1skPVLO5GlaWOzm+tuO/MW9Tr4qivcg5gsQtd2pd+rypFh5UApw2mrI58NAxMdRX625weHUTscI0nGJiS6f2QGdItGrJEj+m8YMgS2G06GHx2IGU8HKICp1mDzcc/fqNP/8TJNKXIju4XB+2VkAjexGHjr/cbCyHftWZf72M9wLSG8DTyuJ3AhWFB48oSLLiWaPOaruguu/klIqRC7LMbaI94mOIOuNp9/HLnqNgtT52eH4AZbZB+1eqJn0XG9uj+xXyinCwxwfF4CBz3sU8RPpIY8hLhCOxkqA/VNl5R1Kg63glrjYjGA+ogs4ndD/yy9Wa+KeL6uKsb4T2cUD15I4G1GMKswgi3hdAZuoeVVDzD8VtEH2OdsnkZ1M8+yejvWTCrxst1vvvLt3/nCakMQ4JbLrCD3YKDBxlbWEDiLkOM9nqslH9AC9tGvN1D52SUN65g6zNlyxmCwWI2oYpTKAVcs50nQ5RaGgsjSRi9dGxoHi4+x5KoLFs7edX4F76BY3WYo5DA+Pz9h49mNQdW/FIn78GMCK+qEirjf6MeRzG1S9PqwnNN5Q1zwIEK3OBtDK4E15XWH7O9FA4Xdh+LJ9SCTq2POei/RWfULx3pWW54P5ZjsascxbdfBl+N6UOyXR5J9wQdKjaWQwGqskL3nDmR2Pl522YogyEIfbCuUNxtOlfvf5HnHrFRSYwSrn32P+TMxnCBvm0TARjNGwH4gSUBADbH392lPgjF3y9uxrw/bhNcwKWRclWGc9DTeL2t3SZ2OPd9TVOgvQFUsqIcVm3UXdo+SkRHskjEjGCteM7TbsDhXsHQThvmPqAsmsi4TcAeykyNDBFtHIZlNwbgUbGnBn0pr1lZM1ZUcqOeXpCLW4F6L84jBXWzA7F1HnS2APdg/xwdMOH5009ptbB1Gv173/rt+ITHmgau3wozAQq6HcrU99JTndu6PvZFYtgmG8lAFdhloyn0b3rsLwGP6/JIYgfr6MufGwSq1gO9jsN6u+vZ+mBUX0VAtSrz4/WtTynhNsHM2fp/30Sjx08vq5uUURtcNyNH0/i2HK6TAATCVYUKEItUutUSDt2MN3bLkp//aAbdx8Y7AUnY74GESJaL3Ftuuci591vGO13O5clYF6wAAO5p4j4Ir1+rvDpZ09/ipZUgLxKb2sYmQniLjmu4L4hoUs4/kKTFG0NNF0Urriox1d6w91tpIBE4WrC/4T3kf5/YRVxzN8za3cy1crU7MV4nmWFRAaVOghf0oybgNBuwU7ThHCHk0xbHmht90BPNx4FQG4oct+nkbcWj0Twsg7LfdwR3xgvcYT6iYr16If+W1kOF5Xq6LBVnslGdY9Tr5cE1jWsqmacb5fpvjO42i6eukHMUFAhR9jIz8gPiwmb7YbO7LzPOzJgI6VpuwSbaIUsHeSBuT+huSk6GxNQIYqFmhYmVXCTD6q56nMX5+gaMUWBUSZ7SB9LLRRtyOGzam/99qjMiLhhlxUUrs56IscOyr+BsdQgo+JfngW1G3n4snfHWjhlFOQw1TgaoEpOuzsT/e6lrapkknBDMF732rhRsQKIKNDBQk83q4CKwm+j3DQB5hU/T0qbN6JfFsQClkjgelQtijPUunmpZEzBX5Zg15gBUYUsZcm43SHyMJ7W4FkBFu4lxG+6Af4IFp+tQ5FRsJ2288vQ0FRFJKSfwAxOOZczFJV9SE7lkxicZrLWm1hbLiHc46o8TrcoHDoCsQcBCjc9DBylITKxTx3eQC9mgIEydc3a9ZLnXNfiaCTQCMGYx3ZHhgOBsU0GCTN8Vyreo1pSVPf7psBNUpDywRj8s90tuiI3CnMqGiyzNoUdbiQIMoLgIlD/dDjOlXYlerit80v0Ep7L6Hd9yx1DLmhrwUQWZ2WNJsBpr9Z4WUBwnqUn/+sdcLQSO75juizZ4T0IUnDoF4y521Irc1sjNQS8zUdtgUjnc2CRbmLpCco8SfBMHQP2DpqyrlMTE1Bd3KHey/Lx1czG72I6pzT/3e83LOaRAC3Suxa8Lslc70G9v2Aq+D8g2yd8QEtZKsU4vhtRlI5CS3rHRkjaTmcd7xZMbSGPR4N/xXGNfVODGgsCXJWHWi77oFNIvhK6F5xHPf2y4rliLIPXnxprlFQzl5FHfkP85UxbT011RCfoBOb4Rn9UUVLdiVGLAyyRIcJkbMcTa11wF6M//d3MgKAT2MOIQk/mwSo8sqSrukHl3JBmubmwjzCJiOi4B+6UFrQbyOwHaIGLZ1em53mCSEtOl3/M9Pyu6uo+8/+kED5QryA8q4B3SaaX2Osgop+zrlp3SzBlexogl8jeiALFkX8a9ClCMRtpgiVs+0ZIuWu+gUtF6XeA6RNhol+71NeTdha52Ctej4EffOHPcpFDdP+Sa1j+8AoT2XeytKinggeuU4Rq6De4CWGaECbXMINuHDdAi16EWASzOgpGs6v42MY4dNvf4aNoLqje6xqjmW8xQXMGYVVRJnuT02TNSsrAvLDi4JTrwWH5WN201KnXuUknfOpkvVt+IW+o/LYASwIsz1vKO7TFIWgzxzjJpERSlBFoVFVQyqFtutXKLaAIlxoBeukNtCXQTTxACdd42BKjinEN7ZgWM1OnF0LbZNXaBahIGfhigfCV7eDR0wNS34xKSobRLA/DhnJgPb0ZMOag1yxR6/KU2P/UB1Z88gQMZhThTmG+PUAyXSCPGYW/GzD2PnnRPURy8GiV+WJye66/DKhXnU4i6zlJ+MojTecx66Z0YJXviPUbjAK6d9LAPopYfo7xH6Mdq9dhLrjcMFsHMT25VdXT1YAYCqFGUXzdcVkW0kgiwnpZURYeuJg1m2n2EQg4Ole1Ulq85BuOlqHVqOThLZKMaNwLABZ5P/2+7ddsJfvXtwVN6Qq7HL9/j8oKRkTlm9tRruyH3TVQLLhUFfGENjjzc7IK5QQ7wgiDu34HYVhlZuwaI/IhX7iM3LtBfGATRfrOF16oxqsjGrM14nBZB5pU+eYkh24qLdtlJTlczPqGuh/DvAUgwg7S8bUeRAUbAAPDDXHGA/OgbKDsFMKJeHR3kUBd3jwuYZcNqp9imbL9hLTBBjIQA+L3qhjEQNKfZvgDEe9sr3MzhYLB6q0NFV6e+GnNIHTVH39lWvZF6D40+gvPuA8nNY3Rnuaz3+NpBqA8qmRWYtliGwGR9XN8B9Q0niF+5N5bb4FKQDBl4KG8ClU36BBK8s0zMnEpOW5TMrRmMxR+iIlzpuP3fv4Xupbkse5O3AFRDyqjggcI7Gry5vf3NgcmU/V17cBxovAZR8JjAAoCfjeQTgTHlwsupsxP1f1EMUWIhkrtEECR+Y8XLaQA0DWTHDpmrKFbwHxRqTlJTRtdG08S+kBISqMDpnoSeNXtYV3vH61Pmms0S3a/2DmRh91jkqLmQgJYK/g9ewciwW/x4IKHH8bcnE6g/9uZDDhghzncy+CutyG+FJr4XrjznE/3PZNL4Gw0SX8qCzg3QkgLwgwxmB9V2Vrqp7GKiBv+PD2I8a14KOQk8b5+7k2IClG5b5xy6Iv9tqBgbGUbkLBfEFCJfSkx6tpdqj9K3oDsMrY7HHbRbgwQYFP9b/HzdwBMXuiLdUKBmBB+QLDNIeBeu/00lcV9nyMZo0FDFPyh8NnUwmV36VWj4V6RvtXrLMvzBvr54pc72LpNIzeh9zm2bqOLiD27yaX/Cf9Z4SS2DbPXRVVTw3/sfoRSb2YqKZMpHsGa2yUjZyFlUuwqV97cHEeZ+phNleyUJsWyYrWOb8d1Vax5aGfIMBJ6c0MHDVp6S7q1pvYwJ2YsdxEU/1Em+YJyJHfUKdgpzqAO6kCorQAlH9a11izOVBmmBTnNTUZLc2+AiOtKPNBEN+pTxaLp14b5wNTFkwCezGugPzIscdrgT5d6QVZ6yPvI9mtTPC2C5Uu/q/gQyB1sdBWe+vtQWKm/4qXiVagklVd5E9mjTBQUK4sD5d+gM1LDhkIZyMw5Ic7FbJz+WUaiQWvF+i6+1h/pGFM7YGWT5uzuLzrVTeX4EbuwGGQZ2G5kXYwYhabfReNYHWfZzse0u8GD+qf1Zy71qnt9zX1f2tcQKyDyVDgfrI2ujbPeWdWTnSEqnKCAV41nBGeKUZOC3xUTfmFn9DdGtg6RlYAbEK0oVzBaHmDehgmukNlaBvOdjrI2AYTehpeCkuTyNx1NlAqOJQ08EP9vltvUJpNIA/IDGNXcwAAN5lZ9W+uRO2z8JMOmrkkPhy2NFU73PoJd+nawRTkDvcHpmAD7r5H1ZUeQeYLiaSJScrDCo6ZYIoQEv/8ONb4U5vGS2tuWpvB3NWK6aiP7cy8y1spUFCs3GYnAQUOvrh4tJdL06JvBgLf/vhcs9/QTfcD6z3Jj3wGeBazj8/Slf++ekA96hlnTxXfOzR8bu7I8xQb5teG5botNt2ymD2GXQ+mvd2ugCmKWtVMqvBxznsywwneGGmfpRwHo7RTvoKyNU1bssiCag+T8slMII0nBP/mfgTYL+ZTojUyjrm3FsVe3r2NxrCpJ82yUwkA2Dkqnf6TITDm1Zx3oHW9+02XaEq/XXpewoGNQUYbEAAfoNZb4HeGSxJL/g0jIj/ZVJ5FM1hDDVhd4riDyvqaaxh4c9WcVRbQ1B0sJ2jf0D32AhYHaZCG7fTUrrKAMhmPzp/tbc65VRXisSgOsLtea+KLa9LReES4VYJcwYF4Ne5jvB6lu0u8LOH+q981zhXhA7w25d3LhfzSKem03a1CNmp03747PDn+/1pG9BoTX4UBLYSzVkXafHdecgUzKPUitAE2Ha3e8a9iHuI3dTrlJqLGGGtG8YrWToNEbkJglNiO4mEqo+KAESC3yQfb3nv8svRsdlzKSyUZ2ZtAOscwFswECKTeRgZB9OvF1/FcpWP9ycXRQ0WMxTFerbl5UZ07+IhqTID2eCXLwbCwnt0b1Aj15gJbir3OrVx9FyqA5bFta9EN1Wb7NA/WH5nDvSS7G0LHUaFjawg6x8pz79NCYmL6G/PtmqkJ9USer8RUuCLrKXaGCBvUGmmPJpLalzk079fH2C3FqjuZTM/lZ7poLO5XNpx7TqPOloazls2OwRSexoHfdVSHf6muSHFOQCn7qgZV9xU2PhySNalo9pxw1JGeVedVZ/vD8G5Vwl5vDYEOurZDauiSAKN2qOH0bPa27NcL6HK/vdBBTpd5XqK3Qimn4tmwd25sBNIDx6X5r2GetSD0Bliio6NJ1QjUmjb1Qr6ViDj/Tj8ahMKptp71a/cYjoKHvAJ1Xi568l3l1XkfFRvHlCE2WlAktoOBGCNtSzMZCXUtUhCx2rBBcZaNoCBhMf/WoVZhj1Qbv+umA+MGAvYpi4X4eu9YNgVp+9udM465DzoT+Vd86eC1gQXOl8ocx0vZf8rZHmReYBtxjbJCscBZr3jwi1zU+UBBlrzE/T0m3f29dCum91kVlCXeduyeIrs4LbGpCfqslGdYuNMjQ9N1pDv36Vav3eMfnj/3X4Oi+3dwDTHITF0c9FUR3BWpb9SsxzQd7C6oEoF3Jvw0f5Ov40KrXvyfJ5XFxtt3allp4Q3We4Hg4IG1m2i2+rtN5nJv8jUqHmFzZqaBkWFIvvUilMEB+y0UlZ2lVHg7TQLlK4WqExJtXaxNzirzxGMA7+NS9eKKXQoPBwpEPIOFcp4mq8onYKyTRerfrHp3IGKl8/n7BObSY0TKyY2L95MiE75Go0W5OYV+G5QnnFyxCzWMuiJOm/DgqVvN+SA+2KOwGAdcvJd0skRjJWOMWkozN7MxlTJ9Ud5i/DLBV74cwlgqPPUyTRwlHCPLj5PXQWeiG7eQYpLx3Ap7sysG+hVscY23ioDSd9pssuvOUikClRTlZ1+dVLYDCIYkw3T+LmeNknx5G667JQpQMEM9uPmWmiR6Cevkkp7HQrmvTVTQHbVvoEiLxA3/9fg0J4KoZ4u34xhGMjUiJRYpBXfUAyIL8YaKiJp79OUnIJm8wQiKooqM9zwj5hctaCxIPjWM3Iy69j2phLV1UTs2028a8m3fF7k39gTexwY8LEnIevmc/FVzid5sLQkKdgyMS7fz3MYbLJaVFREHSA6WaPkoRTpI9Bjqfnw99GJ3Tlm4u3njbM3BCoWEB0KxElbQPKa9jAbMvDk/44AW2pAhLHNOzWB4VrKpRHv4VKaNT5GU8na1ZYG5uwBitbl1htDlA0cPSQK6HMxv/cwE7/Nu7SxZEi65z/hLzNn+93nw6uivQh5LnnfYdtTd/oh/YATsQocpXZbbv7tu+euZ9xCs2JmsCF5BwN3V51qfcfVJCLy3/n9sC250JwLXpco0iSxJHFG53/YFW1A+S7NqzoI3p4YREsrMbUz52hw9KPBDCKCBJnprjokZMIS8ANq7hNbD7E1l+BxfR+8ZVlgpUhvNdS51HbWJ5mLXOsUlO9H3JjYuKZHgRhXqJLqOMSnAcKYo/fBFrVSQqCbigqH7O+k/KhQUCDM3vEkdtPPOg923hm9jOJdlP+SA+U//XNKkUbe4gaeH3TnhUpj75RhcLmwCcFQbodVgy2wBdTawREb738w9IeTzBRjgY2R7AmLlTWLEHWp46OEByxhYy1EbFPlcjZoCyJzGhZ7aFpk8mDzVM8leNGq+GUYX0XZ8mFDtPatC5Jhx2mHZBUWooXJ1zbyN66p4pYwNIOBwm9jsNWnUJfA7t02aIADH4PQWz4Opc8cUvSHrvZMjUzKg/DA30eRPOPrhrGRW+ERw8DJCbWcbPkz+WZkrvPoHeuV4t4rK/a2Rt5i/ckyL4J4Ag/9boNdfi+TlQfPkqDH3dNxvKr3VuFEnbSMaqxcr2xJz2gi4MF9+Pq3xngsmYtG7kfH5hQM/Mk6iTDjiVlihALSvpQtDixhZ7GFbZeEhKZIJvSQEqp708puKBoZ3Wb0ikj4iOLPR1Q5wWmMEp08qrBIcQZw+2R0LGaFzvR5IlOyJLT98g8wD5VIPAfRiFuYaxRlDGwo+ntwulIdI1dk9bSrCmVJ76CqxvnNQ3iLDNRRElOOm017O7raDLs/fRwxnKov2ofShZyJCYnRoQmS4AzUgYBwtLCmcdu5dFhfD0zAzmEJ8D0ERYVOqKntr1NP923MiTgsqdfTAQIAcSkuzWgo+WtmHqQDEK0DdvNAcZJFxIzHTTXXXFTwb4kw6LWExjS3ywCmD0vZxpIyfVBwmswCVUzmHEgkRqGQ46h3EaJ9KY6ySSR1JV1ut2luuthzIkAu8seDZkiPRHRbXcdg6NN+BJ2UIGa7I3Up592n6pTjOAOwrTQVfUI9LieGa1aqE63aEcFbymdcTC+m5ytaFVrWUMfu92uWQC5XGGwzi17Sqmuk2RexY+MAMwTnvNcUPWvUOycmgRxZJZ2FyNvMTBSpINglRJBcGeFvcnfeAQViC/WX2nomle+8Y1vLTmnERKgIl9KEkMggCwZo/cxL4HAUSq/0lyPfN9GiOi3uhphTO+OgT26jC+3UDzYcjGi1cZ37TSW7QotYAgczIpWRgXjrd2jvG59um7s64nTkAo8Pfa7qR0DbxOBP0I88gTnIEXQ4QZmEz84JEXzXa4i2lPQhRuo9faCCbSuFlk5/i1g1p3He/dWYkiAYTF4zdq1Ny5ijmhpW9J09UuMXsOho933fvklcPSMLKtznEgbocI7O+dauXHPh6l2WlPtwf+TvI7nDOL7ezZvt/spaVQKK0VNKKKow/02yD07TNHWKRfKXOOJ6IarTeEA2S6/bjkJEPGFdsv+pD/BEduuZ5N+rb52Wd9ncimYrjLYzxagdPoadd4jVegBIm3UceT/SEhXHKmHKbCf7hSsf5zRbJbE3RLp+KiuNCDLiwhjXjV3GwGycGkzJfa48UZ0o7xJnD6AD1hVQEkKSUoxpvo8VWsiiD6ORe0A/U06AvlfyV+ks40nnkYFyCxlSvzGSyVz6FE2mQ7e5HtYmjbKI9hecwn8sK/AWYUW5ylw7fxCoM/7mOlrt+mg4YRXxGy2fkVWpLu8UvhDy8Id/q8fFwczk+SOZTmfMPwgKuL5jNlnWuBaO+76bSL8U6nhjJp7KlAWaLl8re7xG0gjUXXmcmKb0Pg/aM6zF/0MTW6Ht/5zFiIvFS6TJZr+FoYbQOdL6/SPQy5vVYcemQB1drqtOY7kmhxepHuvUISetC3KsTw3iK/d+jPh/RBNz7+N0Xv+l1GPiurpfwBC12YlG4FbdS1YpUEvnEqOi6vnmsEkbEN20R2ipN5nwzT8F2XNiSmbwcJkw0k9WPLqrgK8D8fL2Cw5uwtiKkMXtVs3E9Rc6tdUoFr2RvAW7FTXeoxg5T8hpBlxMdYL3HYGUnltjgtaaOgbdHtDInRyELQsiHYWc7yoDa0WWO8SLWQBNq+u6QiN4GEJCfrH+Ci6nTbLQRGQeSZ0uMyEGEEQ5p4pVo5conEzrZi+ts459+X4MhuH0CuOxEzWdtFhDh0plLHDH7NVGgNUpGg+01B1de54uDMnbctTEpxN7pMFi+SwaYwWyN+15yUiGiMl5uUhwt208ytmnmwJLtZpSBJioMcqQkQiD+wmoIVigBSc8CbQyX0FaynxWXSBnd7StnxTx/KvfFPmWV0YFVYdNOI20FJLNS3Mf48+9yyoYSh8i4HLNV7VTTnwFrGI0wMO1kkXVWhVYYHkQLiG6RmQPq5EWM3Jnqy3J18bbDwkIOsxVSj8i0i5zkr4u2PBEGa6P10D+9Pn1kfgcb6KvVatAWnBZN8EVOgtp2eFrc3jhB6zVs+T83tV6VQbQ+iPWVM2KGklH7xvrFSNYLaZHsxg3uM2BJNR+5zPgP5JpifFnvKcCBrM1Meoho9BI4YVh96272KGSDB6Yv9RyCSgmcrdjH/jFkXs04W8e2M5pLsZBzFmN44KNhnWUi7pLLJNAQ7LOoWvwj2TqV9BVQ3WIV0YLXTu3EZVbRS5HU3pZ48zLDCyOpICxuExGWgmranrua6pIErVVxyDac1rbpHtNwDGaAP6+EJlWMqn4Rnm4Yt4sLKSvlkOih8BYEk0jGI9H7T1PTRY+rpFaVQR8gcJdUDEf+6jGB0Jr7PAbZysPQpRKqc3dd1tUa74c1nxTmQY4aV/uVSUevab9UAL6cSKLAK9T8VagLVGplZWaVIpn2W3HphoL55P2SMGC6JB4uW1uJnVY1UdwYeS7OkIrbOVkNrJ1gtnoLajsSitnufLHJgqYwOc1GwE2oou8d0AbCTBDVChNCzKDIge1QRLFb/MrDpez1pRfwMWV6NXjfHZ1uCbEFq8ufRliY1XYE87u5yOWWIbFOwJe0CLSR9VdDVHSF9+O6/zTQFZtCRQVYaFQ3rZp1mG299xScqJg8ih5aZkLmKJmRQAHpqNs5DWVPwZYbIBzPkc3mZDphwG6Cjy6tVZgQTMSN5FydIAe5lw2qWZO8ovwJHWIo68JUNRB/yA46bBv9c0/UvMTqNT0SwxWINYFkM0nnGV9g5tqIxCWGXqo8UB7Yp0eSq1luuMkSQJjCSMDPLkl3tBs8Ms/JwRb/CQ9GQgiDT/l3Druf35FYkAjjDpotJ0fD2UFVJDAsvlt2Atkmed1tZvpglBvTFTei+FemO2JxfNU3/aaMbOGk7kj+V2a7ug264gUBeF8QZYpnqVA6AaJWXWAanepDYdyxYFFBO7mMkkAETaNQ8UKOQfjerCsEwR2TSFKBsknaaUSxyjUkI+D612N1w+Pk5AKGOWFoK7IEYol1n0A6o9I2tMyNdt5GV9g8Hgq566u+1SfwUm4BGlxtuKhIlKaRL95SF+A8vlF+Hhi/QOnASdosqhDjIE/Q0ZY61a8CL4d2PY7nfgBRmAOeopI7KP4ugCT9vxYCJw2p/wAeinBHqBNIHgPhwgmTSthv1jpLxaMmRTnTNA7N8XYRqMTCu5f1zHkHg2tlqf+zZrs3hLD7bWc+qwlVJptHX/HvPP/ELjlK6z5S/E/lXSJ09n+Tosnvm4K40FXvZjunn7EPHaLhYI4+pn/SkjG63ESzDLFrb07AMlVMTyfuAOczKhgfSAXVV6dbq2cY/unPvJ1dsxWL3ckDiQiHasbXcSxxwSdKzy9O9c/9zg0uVHLyXfED5Om/50S8a+cVYdvS08a0Yl5iw2nUvRfon5ipfQ7brNXwPo5sjwjXKnCxeeuClc+Gh8HwPlSOBu/CC2F9JkH+SV1TstX/rQyEn/YSCUvdG7PI/LNkz2Nd3CupHa0YWZ8oBbYNBRuGyXkcoj9Jfi2q4N/uiHGKB1I/qsYDlOdviTZ5N29iBLB4kOZoXPDCAc4TB0jskeGM/dPszbA/9zIMZY7A1loaB8HPLZzFiZCHtGaMK/j7MQKKPizkdxB58tC6r2+l3YJBFp+o+P/DPa4ZhpOOw4a3vxdEDXf5nnmX/axVsAcqoj7TB4D9fwC+I7PkoH2PI3qPzRbsUf7wuMlL8tQVpf1x1l5siuZraO4JoH4aEzqW1m68XaplGCJt4YvuIvjdPNmlR+WYau/RTinz6/aN/W9q0oGlq/09ebGUMEfRDGpNe/z3NA0kn3D7MtyHmae1pXQrUS7gR/6AJ/qGkPS6f8UC9DlBvf6ufY8beY1kMQujkOjWwG/zKYfqkv6AG3jCCfUVlmrAqhLGU6JouWH5Gt5IoxVZdh7zN3gU8cVxJIuu7j6Lwx2V8oxbYVmzDi1HpZBqAY0d2giHn7eLSHKC8mpGf3TWDPpVL4NJ8Xb3M7PJi4zrPuN+1ailFN30wM9eU1NOGw5hStEB1HT1ZHn01Xz6X5OIt4D1VSn+Zhs1txDOHOzcoFpmF4nkulsQ8+wC9u7uXwNe7Y6uLejyJR+6mGfKOM7b6hUQYoMOYGBbHup7OH4k+WDf0y2XiFpDcsAhlobPN1lkUQP6ZMIGV0QXmGDkxwCjh92kOwJ7yt700dXE0oSD6V5s434hm8TeTnmxtXdS/hTsMQZ+DekbWhJebkEBPuaWS6FFvYhPlhvG29HPQrBKArC9yYONJ3Fo00N7OAMyPKv7TS4Ei6YLf9iEXPHOzVsZLltIciPo0Uwm4VpNgsCDMegoNVfSKgq89fm/vy4kAGsr9JYrcVm469g8MC060mHnqUvy9dl2k2oeFy+g8IeEm4F7OPe1XKlaCe8XPu4WNo/cCJyZzb4QZGo70k5P2qE6uIK97ulITmH/cqQRlG/qhlaU+8nraR1CPH8EElVSk3YhzCST5wTkO35lG636KhRos2GNJvuynJnoIFTLWJMbBrKdwhEAhYmlIhMJMcIns+lBMs6VZxZC9agqh6kp2LPinK1/ZUhXjuyCSHpKYhKacxd/tOIvzK+HzFzkZLw9h2BXWDN/mzVJh50S/5TNIFTO+ZK40r7vpZItOWDt91RyCEcT7XDL3+0d5soqZJYHavR7XJ32yHLPppC1ZCx3KL1ipqP399lVwmy1USqAwWV25JpVv2wYue4WoDZSkS8nMhmRX7nwcdfmS6cE/CtepcVHvVpDtlSwD9LrqrUSr+KbXOCIlNARY916Ek5V6loyex909HBFSlZrqWlZkEVecVt5I5VScMLRjdJO/pWLejgtN0MnPkpQaCZMEeFfwUXGio+8XFERjES7BcmKZE4EN1+2DPFtvFCVoOgj0WVSTooFR7/EyVuTTYU/dv1wrBAJVshtzHzYal2Q1ML05V3FlZY7o+cSPyjKhsGZrxZHQ+m16z/wLyRQS0nEaY29WYTVeCtrK00xtae2BosQENhhHjTU7byzMF5888LOIRnh00BCfKWHouYONCHPm9BXPXRbSgJkVA6t/LQhAOAsCVDLXF4H8Nm21TrEzdj5tWkjK4M9phhYKPGHcJI4k1kOARVNw4dGJ8GO+rTQc5LHiGrFQWJakWTbWBAZd154d4d5uT6h3AloPAjEC3zMa/RXNQRWZz3JQHZ1BSXTd3iqE1aZnG3Hav9Ymp1kroMLYTTLc5SKpEiqxavt5J5iHLXH/KOV5e5MsH4MaZOs06eTblV9eY4ZRQwYz6DU4ELk2CoUT/A9WC8F0UBGKQFsVWuQMOoYCAqXQwm/ncBYsrTHcUraYKMy5lWVE275oh6RlXj/8M+PYrAJB6CLoWuggXXwgxDWm/169LGaQefxBqp/QON+jms6xmjIS7mdJWDfaR96fPH52oBul2LmomszLXYHWOs3lI6uCLllelG56hDXsh8/XmACsyqb1JGH2pDT0FW6rSpT7FKxGWP2pLHS5BgelhF9en3+yL3Oz907u/AY1ipPfTQTBfrIpQxl4+OeiRhBCSme/RGwbDu7oknqSQRZ9cg9oe0GKpAo8I8DhJu+y/9qVdFiPR1Sc0JUxTQvcA4DWrO9CeuQve+cvAYJxabtLcV7O8ZLLbvMHI+xCZsgwH9vhqTj/X0pTy5cMbyeDty1EI9Fkrh1Kv8poQLNu8qLxRbym0ON8PgiipLA66PCCpEbbB2T9Tg60CKCC38kJdOAGAkI+Gx9nYtrJtQCPxFQ0bUXH4Md1BYhx2HLU0gIpTWu8q+cz1lsFuWhWT5vEjBQI28fVpw+1mhw0pxkhrKz8p6QSqWIyHeeM4pHl6FTE5Za8/bUBru/1RgeTlkwBMFyIj/sGw2+j9ItsPRRH0LmeQ7MunIoyXQn0bbBZ05U93X2U9/BbSwpXBKRyWEblD/Jkh5xdZnnujmVwjPm+z6R1fmWzVfw+yGpLtX6+6iG4Tyz2WwM+ry2mneY6/RT4XRpJujydIMmb9uaJvyuklbY9k6RePWIAj3kWHi9ISAE9Mgj56aHRtO9h0GHzP16eV4zEImOAqmnGhjlwRzA3510+hndiX+csrNZA1czU6cKZNTzWARbby6LqQn5hSXrVqlk+BALjrC4dKnYmECjwQCuVCjcj/+JvlPlvsB+Jk1ahMq1Jo+4Qw7xqJRzF7Nlu7psiIDMBOzMHGIV9hii2PPzXBtNMNC9uXHUHlj4nQjIPgGO4tjGLuleb/wS8Jpi5DvRGxORxYFHT1tQYprEnAV1hzNu/aIexNhyq2W3ciwrYTtvna+kgduHLVJoMacJtne1gV/ggX1eTeKjQP3UXQLdvIUUx7hNhjojKOAOEBxWk+UiGLDEYRnpwzs2rSgWq3Mc09uowWyl7o3KrVmwnUa13h8EJ/M8aLFvk3IPs67eB8vXu0iMbbSAQ878oie5ch7iwYAfgTYqZixIcC5A0jBBp6wfzp6UpkEKSNKDcv+Khm9kN4GcHvFpDrizD+p3qF+1xNU8DkDPYt2maFvDLutYtKPF0/Z6aNhIXESU/ILkEvudcq3DiXKxBMQYkgsJPK2dQy7G5NDpvfRCaM+aak6obYieFitt4f916g0ee/7R85oN8ql/pCnJiuaUINqjXAnGgERPhpnoNGetmXhgaPlkAxiM5USeCKWbHB+RRcuRP7e5uNgtyGz+Sg/x0dac7s7y2Y7dw860UfjBvo2ReNQFwGulzY4mSaMIPmhgdKOTzndxA43iAUg/t9rRFZUJzOkZ79XAZznt+KxjIVsySCmZOM8QLCRQrSHJk5n7zaHoMz4khAIH35dPc20wffHqLn3T7LqFtTsi4ZPb8vRFMC4wlLkKBMbLwqiRABW8rDbcuBQD5a7NbKQvWk2AWY0WU/VGBcyKeyiops2TYqbNDfulPkW/Q4w0MdhyyOERIIvJ+fqJaRrSyo9O6OTfx+PuEvMJz9OIxvOOb4RmM7fZVhbBrVZxpbsjr+HGO1xAJapTNcF9k+FhrbPbs4TsUDuxSjN+jEnEKk3RCVmYgxy0fMqxtLKwXvp1b4mz6Ws+bJp85lYlExJujnNPNU2N5uVF30cA2KJ9uPpqTrRSLZXW1Uf2i/5qgfG5wQErmwpRyPXRA/psI1Hmun9ZVFx7hHVccDfdewIXp/hDFEVsAoqmpEhgVk+ndCaTXWoV3Wwbd7+Kz2CM0ugFuCHbu/pbSEAv/DzUcwvca8a/eQIA8zZWPw58IU+bPz+kchoLmLHZ2jVA6m1OvcsOdxFBf9iIfsqyIW/aXw4FslaYk2GHeb26z0NlG6SnqiPJKxWwVjNcfEWwkQQZngP5BCLoRPvLH5d64TKKxjgnFBxMkIc3vPlFQnyet596pnMZSxyRiqklv/50j+R5+F3rzdHHcFVCkQNeKxyFyRJSMjQUyM0zf0fgd2zlyazqln9uuKjnIZByoi2lC5f5jgMldEz8EWGbA1Wht33CUntS8tD4C40dBOGz2RISE5xyBGI83xyN2DDLOKEtmOm8tKW5H2QPvRvrOC9YEJRHya9nWpWcgrczvdE1d5xAOnrxiSZrEXmIomqnFLNp1tsorn+zI0aAYbVJesM9FDOZxSSvx4iaQ4Iw4wPafoWU+hgyxnIhJtZemVJ5HmoDQr2XxTZLWVNRUJ9nJ9dtVl6i3S+eN4XP8wZD2vbJxbHA0KfvO6cMlnLrwYOcFEIYYzX+Ft49n4aR9BIfXWGMDgboZEHEXzAhz46wVRWyitUoCHpxH9yxhJrY5SRe7nuklcLP9lTJ6E0CQeZEzy/AXXAfPrjiIPAMZNnpBki2YRWhZmg+4KdYClhFW7aoPDor8ORMiDf+kakpecHDDdo54EK/7x5e/NCjsdpAxCu8fuXwUIrhnTH8tOurqv8Di0VDYfkW25H+KGJWLzDj/saCHA7YYo1TVQZcKdmbG5wWaZALgem/YtA6/p7XKp0IzpztXBPdJth/1Ys2RlCvGT2KV0YUfhdyK93uf8UGDRwYeAi8bNeNkyz/DF2OiB9oQJaLvuM7NMCAdQdi1m0fmxdCSD6q1mKTzM/MYbdnT7gYSj/hOz8R5uGPORJFPDQgsnrgKJAAxzHsAZzOxM8XjgE+xl7fuLicTwv5VOtprZC3FdMt8Q3FfMNvIRAK8+bRS5vTGo7/nPb/vmXYksxdMM27pXWpBB5gaNniDqw4PfLDcKphLng21xlQaiJpyzh/+U8DtKBscz3OOGL35ozp+9YIwqQdzqq9Z5PEQ+BRa15xrpLGlEppO14Mtg2NdvKsrKYcW8bRWGtahzAqmLA8Unj1CTuvsqG0p0lDdC+i4MYYWhsc5NlMc3+JR7r9vAmtOGASWJ3Z58kP0dny6Y4lZhj1sX2wncv2aeHMHXmMSZ5scuhwdd4ZWTAZgBvfMi98cGXjdG386WVYJ1iKapyogFzm+BYP7VHOe76mjQVD8wZQnYF8TTdaaCbodz9CAaqO7ihAdaBp+jZ4kjZJ3zGx2FVcFhirgUcPdPG6BH+i7HSP5OH6PBBz6RwUWzh7V4o4ZQdyHXV9pRWu5Xw0aDSQ8jBlC7tMOdyX2Fg4FtlSFV0XW9hNIts+nTzcz6+IqswEnLC58vNfMgBD/RBkktptgQDgZPVVMK4pPhuGX6s9O0Mj6TYYPHLCCXecR9wekhtTO15jgz41vDSIu49uTqizfw/176kStzD+kwEFSICPGweidt8klSx8jdts04kWKjNPpM7P0gFiFvqZIOheu0TdnfJyG8qiQgNrj1a5Ld8kDJOBFKN5IjerhtVzUvp3i9l6J7o0kCRmsMUOhCcC1+LzAiZEIjqR7lV2R7xGVzmTEo+FksdWNl/I4y1y8taksXqMd/euAgwhr+cp6YuXFcXH5MRmrTBVUHCb3Sz0CKO72Z7ceNiZrxqQ5VXmn5uqA/6Pmz8VEfnRTRJ8KZlQ3PRE6knLl2qk+NptuYXV00d49h+jguPEZCfD76zYdHbh3xgva7gFsQPq67GR9kLaBPMJwrHfxXIZWcRYcJ1DuNJrc4+N0eP6qEjmBCNw1XzJ4WnHjOeNUts6POSaS8INZURrlqzejSByYp+DRyTL7ih/nZEiSQ1Cfhfp76XoMjsfdg/hjhvS8/oRct7hV9gi2Kw+sGGwwrxOQXj2UpgDhsVFan3OJMgbl0mT99O9IFvSlUxBLjjkuK5G3cjray3EUu+r8UEq6AtJjcBedJZJZ3GEjHm8+Exib/oIlG/Fl++eX23flyGjMJumdr3PUwK0ulj9Gpg5oFF4xmSZI5hGIbxF274cW4ova0pdwC+56M5TYa+Ll0GJx7+YdtPa3A2UcqBjbp8hIdk0jhwFseU1U1sime613WwOjFscQEYWcdqbGbUlO2Gyc7sXWcZE4yp9ovLhjQcEMu6fL85Iz8RsKJMJTEkhvvzaE4jafE/fj0u3vev7OTfGkoH0/qQRQM6pNZzjKzQoaiEj9io2oI1yeeD9pN0rlwIKo8Crw74KB1uQCxC/+njQan7A+vEoSD/BCXURR38bVl3fwOHVt4mbNz008jY6a4ESWY4hpLroNVUInIeE31TwoXE8VuiQP91ioZZitPjo5qe+tIOyLOImlwegn9nGCfZV7jHQIm+LLUGDEr7OB+9MupwdjqbLofJdTjH0TOXI5mMvmPaHjTMDXwS3X08nWuHqLnw3mf0uIwpv5XBr44vdwRbFtfd2N7KkprC7/egQNsz/k5qYfTW+lZfEJVjn5tggj4YhrxfO0CYFB71P+8vTja3tZCJfsjGVwEKSCnsRuHAWaJ5LxhGa4oCTrl4j1r2fsIqoHP1LlVa72QEoThrnXjqN+Pi30WGd6/gsSJqx9GWgANVerjhTU593tNz0da/3jOPCtlynk5j8KLOQfA+vIj5srEGssyVu4t6s40LMQdrspht5/1/eUq2NUvpMo/8YRyU9hPLFcXI5HMmaQpDbB8px3zXWId0D1AW/QA/9KIg+/87c5lXSE6JSboPto/UKcXAM6JAX93FLZXXDgzoC9rI2UbGJphxaO62f1APzeuNJQAcAn17TYWIUeW7IqYJskTXakuQ3Rfjzq/aDnpuDY6bINzA+dqWThY2q5NE8i6F1iV3Ss3D3d67EsR/pjJFnfKXgcYZb4ipgYSWKkNZ1SvYhSxB7FZfPsyVF7+WeMz9Y5v32YF23D6+CAqCPBH3pgVJT7GTnsPEPQlQhBI23MAmcdDGZfg5iHR016Yz3dBmaaRKDIgcYgl/XSWuLdShcuUHeRXK42dKroSngtF/BCqu+bAchMmta6QCVHnrFI12N9k/PN9xm1AHKp6b8wTKtGwhazaon/65O0GBv2moiXcHQd6Zg7lXaFfFsj91xGad4jVC4Pv6XfwqpQcI9Gcb8ATLw7cyQtk5edyCaOvvxm2woi0K80rQ8braodsUPj5NquwYDWrd1NFkVBy6NkVQv41neE61JI5xMCYAVvz+vOOQYmzmVaAs3Tokqju1SHGP5WfKSMwIbs2e/T2OAMt+bTOnuibncuGhvyryXTvWEpOJNXvods4w2Ms6blaBaJglPe7SLF0OI2lsEJPETN6xyz5u8pOhYlqJukq3GDz+l5mgClvgRHYhDxBQLYGsaYw/DYfVvhbf0JlQElPwmyqR3rT9WSuu1GzSETzkIAMzRYVXkyRqBrkx+Ph6+Wi8zbrg4mIjrZCz9V00JhwSA6lZ5gE9/40VUSKW2uOx0UJZuPfCKUIv22nEaVWnXeb52/yO+D9Lq1WQCXUQS3oXdvbFIwDeiIZjCwxbA/3GDDi7ScVa6mnBWaUcpSqvVtqc1g7K8ydAUZSzcNj3/em6X8O7MVD+YiYDHA4ig02F6cxJnbzrXB1BptdjQy0qwkDlsSVGHbRBXk6eJ7CXBpoyNpiWo7gD/xZGD/nyR1dVxnrWsZHoFLhSu6JZcgbwiMF1V7vd86BYSjos0iL3inz9WsW3zMUpEnS+J0S+PSvEK4NEJHv8OS0eNsQ9rlfCik1JrKF6leTRBPIzTNK0w/EkE+7zetuph1K9xs+U1K29cqtjenLLlGFsvCNoyy9ujVgkP/DFwYOfVAl540+Dz2q0MeD6O5mmafW4FT5XFUsa6uebo0xGN7cIUOGO63kpVNkBhKqVyOoPoZJHeDUeX2yPed1yqQyBfKHGkZx7j0dETg7IJWLtEfkbf0G3wMtbaZZrLQFIAyPDutiXh9SiI7Bt352876o4yE8J3gKsWuI0+8izM35ANJaKim6Bdr/8QU++ZPWox/Nw4VE4kzOtTrh+iWShi7haI9Ycv/+8Mm9W82WpBlBzOH7gZaAmJ7JHHS+C/Hwj9P3u1she85+BTrS4SJqh97OTfGlRvYJI2CMskLHyAz/A9FgeaihE/E8C1CRcdCuA2M4fkkdTBvekrsXSHN8wAEGVy7vY3eBGYBLmxPa3b7US9IqUVP7Cdhc6yr3+pd5lD63U+015mNG1Hk43NwUpT8pUvERcZJwcs6C5oj7GpuuHUhcPT0P9284z86xC4YRCHxETGcZyDHdUROFoEqraYlplb/4ZaZDkGx3Om4ecCzZXHYz9HVV8o0sZhHR9qhP/OIWVgBSVdVFhX07xMfrUMSkn5oRTCP4Isykmwsj75RSB+apV4OATpsJct90ylQdSK3N6fAO1hYqoKja0OTjmfRQPPRidwzcWnmgYgyO4Wpbg4qhkITlBrv33pERSb1JquP1ZrXsEAHFIt7xeJiVmEef+eZjEEZTBvyQr0u2K7/4ORi6n265gFJ2C6G4h1RX9wAK8Ctq6BizcslHdYyFIRFZwAUUabmmBKq8jGMPkysyydp2KCXgIAqMDZLiGMWmlsbnO2IzNBWzaIuzOSIhQnuruF6gUPp/QoEdH2qRHcpwsPkmXxMBSs9YEDco+YJyfxXgMd80FrUYZps8JlVlid0iWR1JcuLi4Q/NJwitaM+TyG2s7SSJltsl25tB/AkXqVNupTSx2WkdDNJYMp5OzaANM54eX+0g8gTudSzbWRKdwUBEKUdjOudao6LJhQHM69WZ7KZyv1S0Hu1BmBBhYM54q9dqNwMPDO6QK4ySF2h6o8PEkpXJc98r3IaNkQIhMBXTFodiEGFKZRu1Lh5DXppKayODbqVJnGJgMIcxVIxwKVi3NAhut9/nauWQLgSE11giKR6D6EXFcZ4s2OaHqzJ9CtjNDrx2djtMXYnPcG5K8Tt87pK4vCKDvyLFSuYNtn1X+USHBPHcUvrRNeGQhH5mWlEdwDR2noIRjxP0hRZScTZ3RmzyMX0zO8bx5gbwzsfTtVfGjaQvW5kEoxiwWrMCYPn0CLbtGUvZnAE/60gaeU5FHIEcO75X48d93B+92VtJrIo308/srkAa7s18kJ2+gw3UCmO/UeBthpTkKJ030r95nPakbOGs3JZke5WAoSFVFEUI+zFssW2bYCtHqnZHTXuy7ttU0UYoO6x2UFbMbYTsMS01Y8/333jKvr5lLu7AUs9Fugea9fTAD3KqGyOc7JPO6HGn7khwhMZIhZz82SYRARU/ZSdFmNQAeD1oGJ6mINSHD1W14aJyDddUzEjq2bJkfFfCKBsGheoZimh9JT/hw2018kCOTnZXdmVPLa7Kd5SlmDB/spv3OMljDoxgM3o8kQAZ56Mk6Lu8uDu0aOA09RF2J9E97YbtCMYRVdo0UR5yXHoJieIPwdeE7L2avHgyXwX5hqO1eZfUEeIUc+LAaZx8bPnusGmolMAm/sRxXG0sWYS1UwrDZDRTsXg40tr0tNHstsOG1FL26dolrnOAA8Bs3SZUm7jiYGCO9W2GzFsdVhy3/mL0lQwA281faQHm4x6ai0i6aMZ5xHEabChnJnaSWQ3B7LdWbap7ORWQB5GUQaHwCfn9wQGVEz29ATv6rAeHZAwcUI6VmkD+lwM+o0MrmaUqT9u+hmAEfuVx8oEEOogpRxy759bCPpiDt4JRsunQxeKvTI+7WKo4RNdzd8o+wQh6nQR6Lv15bejW5Rxnet7PpLJV3uZGC5UnVZwl3ZQzPm3Sj2LSe+nOnWVItKesFGzQMEuCNCMaiCJ/MFqfX8V5fLQ9BhDf4asvI7gqfNXUo7VFQva1P49bO4M1D2ELNmhxVEchowjYYLKGkqC8MAFIyNQnCh67Z8792D99/sumElG8yigV0YqVb9725O/NduUGc5snO5sEbUFzhzQC02oQW72JCB0Sz2fDLI5IgKfSxMrF1ITk550toTnwzlFZLYqb8fsGRGtLgRE5McKXVcKV9axLyy/STuL8ZM+e3Z8++MRLIiNDPplDRJe6fpHqvVIc8EJCV2tm9mv5luYKEEvYdYK4qyLSggpICt9emMvGrAYTXPXnZctUu5/HG6Nf7vtZQ52LqQL6Z/AQ8u/A1fpBgTbxT+kIBTb98GbRflkvk8iO9yxEuY4bro6tE/kAjN6kjon4oMHVcw7E0+fIEw60bID3kKptoauGS7IMws95KGJphiUur24WAP/s25Enu5v/4UAaOkaO0QMi27EhcCAmdFLekEv7UHgUC1PovlioqZrdAnaXyXhadloLAAhFaItMNEjfY/eUciR/uOhdHn0EwPFRHZkNltyJiuNtwVFqkKXsIXNvtWgglbAeh5btMtoAqi8KGjS5fQ5ZBZi5J8LYbckVg6z/xOQaS7I5EayvPXMbs7d6Ma8WOY2SCDIdpcp4ISTfvMOiTIf4GuRJfK9Ns5loKIp/GF/8N9SfY5mgzGKHHX2zpUxxnE+Izb/n/iS/uuBCYL3uD8PKa49RIVpkRYsWx1fWEea+xBsVreJErLAq92s47BK74Sw3WPtr6Z3SJ5YIIKXsJ7F19HetBtprLk7I4yTMRWG+iU0MFz0UgboYmxW5hVGrx7jq1IhriB3UtrwWg6Q6n0U5x0+WEGDtXuFHK4YxIs9DZRv2xzIa84sICPfpniWmwe8EMK5PQqDSjqNxor+nFMGiR6A1GxMdXGlQZPyC13QwUP/WKLiOtXYE1Rps0M8Sl4FS+di8z4Am8P467UiGcsr3RjmIOjnpgM0CnDvu5I9yPMuEQxkn0Hqr7U0BBb9u/0b2Chya8LrxEBk0eDIif6Bt8BmekLPv0xZll8QWREA5E3crWvyuDZwGSGdO0RWky73HGP6RgTvaTtz1pgB02Zb+nFxrMstxyFTSDE54TRPk2o6vOxZXiAkeSQzum7kuyx2PzA2EsdwI4ZJTYTyLbu9DCZ4/bBbvsQC/IHgDFU1CM7zqvaMKcfMDaHdEtlU5+cTF9Zz5Bnlt9FaWBcZDIcaAGyK8rczbSfba70WgI4amKBGkEPtcpJn57qyDDHWrq3FLrz2eIqLmR8VxfCDrEjLPp4gnw+MEH8bZvInAr9P470+MNF2UKYT4i1MnztUEnqir/s01wIb2wRu6BicyB88wzZKeyLQH9SXzVDv5pVrSmaF9NbnAB6G3ikHJAzPu5nbfqie4C/uc5QlsC3Qu3oObreMH2FHxIxKyn0JLu2NyHE3KYIp7RojLoPidQQFW1H7xk42SZ00IAE46/89R0iGs105YReme2eQ2p4voovjXBDc+gjZLGQZUHs/KQCQ1vNTzCCSNYOj/cV5eOEK8wizTwkGRtcz4ssNJ8z1GDbdEGu9xAnElrPedhWmAcBbUUcj2yk7cQP1aaE6ia7LPB0KDIiXy3YqQQlUd0KF54lHdHRxs9VUkCSJT13jQw4Dg3cfk7UP144izBLcZsUC/ImeOdztTIC06KpqeFDzEeRssuuFALODP7jaAVP9kyJqGoLfg30FCWjwT4a/R+/Go7gNGW/ktFUXZhqzeGOf/FifSeA8VlfmZ58urftN+v5hstFFVmwj9VrQTNGvnvbrwNoF9ytcdAW4/URo8tzFxEsRAGNpCQPA2nyG4sTpLpdP4Z3OlwqhhBh4NpUcsyNwlIYliFnjfn5rxi5tiWze84YLYPgVq2YFlmHztMnIYYDumZlC+5NlUsiDYm/GrjMAKH/7NP1TpV+YgX9eUKPGb/7E7cptiCQGDaVLt42TDK1oLOJqs+p3JEQ+ipot5ygBgdAL2VcLR3QH1hzKsVbLeKtnVGQpUc/eSCiksdJYsDnYNTm43LhLuR+KPh5iT8xfDDkfdXNcYIvIKLP+jrYL7w41A4lmDbr6RtM1eC24DPOQpw6EEoUJuzMsbMhMnSI39TzRYJpLHv+clm72h/hy4ZhhnYsMfX4ljyFXIofLxXGcTf9tWpLtCH7u8uWkkrC1YyKQfkXfnFg4hpkw6V3baoELGu/QLNZmZ4I44J0wSkgdN44aB93+wY5G73FvyA12jje/KNgzVsplnUiovzzjR713/8FDAx3WA5H+058lPvh4r2upW2E+rDD0ncsyWsOQ21XVAS0b74foUqvwSVITkP77pmXB+tQSmxW+lMQayt4uC5ZaUFxPYSY9QU3nslkLh8UFnjavxeg51AQ0MOb/8x7/iK5GpW7QhE1rbhDeBeZkPOhl4M4K5xN59OtxLTlG4JmHvg6xTWeeHvBQx8raAxxuD9Y7dlwiZdnvFKDA9/MQk/8yjKWyTtzbc5CJRiSJ8MCcs/tNkupBuXeoiIb+w72v8WjJilP5p8WEivQfpT0gcW/E3dp0/0PXsMtCBB+n46yCUs1NZK/riH5Smh4+eE5JgIk+Se8qrtVxTtH49fGqsTaJZtEMZl4FcFUoHagfltGEprL+5pG9GV25Mm/YpJOhkF8hZDcb6VYtSfvsIYiKqm5rtuc6kVBKpSoKhXgPPLZlhpaCp2nWtdeoNEijwPich5r8nCi3wSZvlYgDhU9jbi4KE1IYgSKXnA7fy8blNn13kyrN4CpXWSGCY+OKTiCT677Z6lZTd7XVrXeJk9cuFM6dp6lXdPl/RVBsWr3qtlZEDO4/dBGWB9oTAUPgzhMAAnf7Gt43XgWPNEa1b6ye8S2fJToxuPwUxPbnWvcBvbF5L7FDw0eqUbOyfXJdnapFzSlkn8B802Yn3Q0RMYsYm7scK33I1hOurGEDvPGh9r7Q9Yatixe007GRv/ECh7Kltso36KfZDT0ik4HHRzWBjXzbjoZcc+HnYIqmc3mRKf1MbqDjluEOC3b47uciwFsFh4XDqnUwPxRSxBp4Afl9iVcp+C7rpypSmzXTd0ATUix0l9WzHdUGMy5tLmugoZ/baDpjVo136MMp6A1asFJfDDRHNW/5zPChLldeAes6ZY2RLFPoX4WZLFMbqqqzpoKr1htYeBELLMJQmY2GgT/jjZN0Zg0m8guSV3BoZ1qEofUh67HPhIj/ji8HqbTMHQ2MHOqf4rE3RRp82ejfTYbMoKEqoecnw4TL+FVPKxIT4cSkq8nmOyA3dEVSn7DujP8kuGWbF6+AVYT9mOePGxAhEeEK4uxF5AaXtA2SS16fos5zt0s0lOCf9i90SmwiZkHOz1DpKQIU/SWha5W6chAywxjmBForDEq0+GxkhuILNpoCvsleWgezYztJ9eG9FHPM5aP15iLmC4vv5YbokWdMPHPHmEeJBTcjC+CVgZ0P3Y60B7X254ouA71Lsogy4Czn4OdaMv1yplbPrXZokIgOdlFYIIyLpvg10j4t4lvJUchEMm3MUxdE5TqdxeWt6YXesVaBb68AgRcHRqgib9gjI/W1+0YT7DfX+JncsV0KJAp6cX8I+X2Sov7JBKgbA0BZXcNQR9j1EISwtUmGWjR1CcEXmSnUOKp0Dm/4QkZl3YW4Bw9n1GEzSMkhCNHRNsTb8/GIYbjTmaeW/P90ATLdmDP7s6rcpWNG+U12Y23Pv66miyhlUf3wFSCnbLgx8bMZhok3sNQLu/6R3Gu+usrDjmZbUoDPaVlvOkFlRnHBdJSVST4EIur1pu0h3Fcwg+Uq1rdct5Wnr6H6cWl3RQE6muRstSJgRDQOmLYDcZIHPoPODaoOMhbAmsuWnGMYauLMUGKfwuOWH2MNKdhAnLRgKr/PNeYLijvfjAva20N6A7R6WxQeDPBc3BSzHvu0pJ2lUAVpuistieBEa6NuXLH1t5hyaSrax8ihq40DszQVu3mqqgs8EtqYkGDlekr++HoMP4Uj7x7YxPKhI0Xk9efTYjIDR9wxrdZwxO6tsztICWNHh97/uXa5lY7AYUn/tBQuOGmMAozfm0o9+UfLznrtPFwraVbxKz1KtH6ziCy3nVpYRIGtFIvqHTtHs6zXCcYlElKpS/jcEWefdsu3UBb0fTZLVWAzrM1MceY+02L+eiCLxYW9wIbbSoRO3ggZwUOg6spSR6qR+mXTkkiQQhTQ/8HJK4Lze3CcGTNfbkoQ0mbUPU5U28Ea7aHy+Q/mjSVR6qc7h7510LHQ0KIgDW/8Oin79LbAD90ZqWAUjzWAVC/1jo4148ixt/ity66HfKWsGsDSG93vV/1RZRGn65yDXZfrZCJrB/pZ3Q+qw8ksqSqOy7eD2o+/xW58idgslbTiKCi+7dMY0alVUs+hOgM8EEco3DKrppjo0hX4Kba/ctABcEo/4ZM1RxaokzBMmoEi84jP805powZvyv0qO/xDZn9aVYgu0V3FMnXh3IDKux4stP3gS2UQ1njshIJ7FYQQ2hm8ov+EPyIpbg9ll/+Cu3cPD9SnHNvGSWhIjubbfGtavsZWU5Xm0u5/a8kqQBrq8iyZ/no7dsb6+X4L4EahklqSmV02NDSZj03GF6yi7pamb6xN88tAeE162nHJRYkQsBCeYlzXzbtBBnH+vhx1DrDEDvPSfjLWXeMLtVPbNt2tmSSjSxtfHjWVcmK1Y+GHEnEUbskeBLAdtY09Ehse3ENVFhYuYHX7NBO0l3KJPgrScgPk3j88GuUi5C0j6JaKbzG/TObJxFK7yKRSr79SBZaUbEMnEhQaKlxQ8shIpU+zLouOFKc8jD949R0kCmKJMvAsKRoQMaRZrrFNSRCvZ1q5oHifpdxvYLRPNOua2/9IF5T+s074jmK0GMNeV/L5+SLhX7leR8+qRYcbSsbBr2MbaGg9DSm3HBm71UUGkSivhkFHYC4hBVl30RPD60SsHsAeX+ILQWwqL4agyJYIrtw2V4zbFJsK2FvitzLVMZDxFGbjY51Hm588sSOzNtR2FEFlww2Fwf6Ye85Db6Q1ctT6IIXJFRau7DMG7QjSGOdcjoxp4eYEyyAxgJtbccfHs6AjUtUBqOF4rJj7UxQ7vtTSWEm55KQbXIRX9L8mnsCnk1d11/abMFIo1FM8aR++8AGBRxm6zcPLtFH7mv93gnLhyD3/2DXJiaXN/MQDTWxEEe8BALZwFJRfqHEZ9/awTCgycase36fhw9fadEtLCWGoRdwOeqmS2Ndp+ttWVC/dMNJeSJXHs/t8BtDu0kVjMv7+gEqrlpF5LywDSVIIsmFrcwampJGhquOGMjh97tzJH8P6cSbUq8K7ZkaFTH/AhVmld3eFRC/VE/v16eAW3zFkr/a4w0rVLlCnttgjyUan8VySJfHVbqaA7TJrMhGxJWVhxh8A5IvcjaWFg0BT48P35bTjR5i7zBnQh4927MAk+tQBb8hgUYCBffT9nPs3thaxXF4cYDirrY/rwQNZYpHS+eOdX2d2JPbYh3SVdb4VhZZGT6wc8as2ctB/M2+QULkCPQiMM6ZIvcRNHwROLvemvuW9X9gz/nz4SckPPsSr2F3pWennyPlrZGu3eVYeJ3AHQzbu5m9phv8km5pEjJwBZmd2fWDEoIe5lkD+uTknYBxNjUGmP5ecwYJCSR9pf7fm+c169o3K+CI/akdG6oi4HfR8h5jIJDRCKkTP38Vhteml0RlG7Z2F++sZ5TIxPdk7ZVx7P0odmEVuebBSXMIP6bFv92fEkELGWnPsVdGrPXeraSrKm/rjOQ/K7QIkJ6JBVj7dV8JECf/ka6OxUUH70X7+Fpf3NxttVBQrTFRIV39TTkXTZFRb3o9lp2Z6pe5N48oVNgsTmenCmbtpd7bcHM5nbb5xLsTVNCswdz3BGE1ZeKRpTJwP9fBf4BCKzfAkaO4EILarJrj/ZafNIr7dbUIK5e/U2q8b6OEMG/Usf6t+p83lWC5AV/mcrc7ZgLMs6pVkFi4Nse6PU1UI2QHXfk+5jryX54/MScMjYeojkOjvfth73ecQF0RLV1pDUL7eoZlpLFJD8tnQ73hze1Riq5s7fF1qYzRaVxKMuz+KsoaIordUmCIU8JpBS2Oq65eoj37cENHenxVl1+g61/lmp66xxNHiB2a3db9Q3AGDhOO9vHHY4DoMbr9eYxS5adsbVnQGlnhwFcB/gXLKR8Yf3Gy+UqPNhWFZMzOyMMjqnOnHT/4hTFPQ4SOcEfXWv/GPp5R+nIrVqWP/LpYh3WBIbGYCocU3nAcO04KwV5SY0npHp3b5dE3ioDAUxVp7YZS+pVFBrABt2Vix9BnLUdReiBMmDt95hvK6cddp/wzPartyYCQliT/xiBPNeOUnCA/mPkZoTbz+p+wrlzNWvhmu9XaW6diaCWqNxtelhA+y3LjsJmsnhzGDTaB885YMB/+811WJ+3pL5ju4axlK3zt0jcm9z8+cDYdADxSVwTrlwp4BsYjxnmI0/Mo/O7izYbj3ozAXWq7YmuGYyxUZKGj7ynVnTyiXnAkPHA84bddI/OMyNzXhd1bLp2/m4NS42VjxTX+k3RykL0jch+ZkZNa1Q04qevEG1jCXGPEStcHPJAKykfpiBBpRb53F7wDzKSQvcDdxkWSXEaxaWcRwHWqZrwIQ/fdEgm9weUxLWNaP0YOWSAU7uPG0489kcwrz3H1vWlWiESMEqD4suyn79ltRbS1VkYoSK3l7L+VxI+8+A6tWtk0Ss374eQIHUZ4PanilSLItMrZEpV767KL+NpZUfyCTIAHmW/QOy7V4Um9J6Rr9FP9EBDik7j8Ogo7nEeIiFUPBJXF9QJ/bfQuwyHGvmzWHfM3CbYM4FUb5uMB8Ovl7C3INVa/KyXNm8HJnkJUPOpRLEMbCDnFjiYK4gIcT7BEgEFbWC7raqkVqv8+LVgKwyZrV1CLsGuqKu87cIP9TYrCbczyCbgC9lyZSZ8Nyg5TLOtK4z4Fb3d/fzeRfrM1MHHKuOtggcDMHOx898CSZOHI59HkB4KfvraEA0RpgKcWf+z3tmnV1OHdfVJt9E4p6wiS2CYE6UOX0G4icvNL3NVBX5cteqgXbk6ykv3zn3oFzIVf61PwySnsK59l+Z2xta1PJMoszzI6dp0k0cB4ANDTj4YtuDmq6ChCBX51zwMoxAu+K5b9ScdbWT2oj8OyyVcokvZLvYeZfihjWpWgWd07G69rUxHX6xQmJPtxiRtWySN+RwV9Gnwv/Sd0g0m6bJ53PeS0QktKNv/osN6WgkfwUi7PGopuiNKz/f+10PL6qVjaH0eeKkaAkU689jOMEGhQnON3trKNTYPNNhi2XA5ldeAVTX6ou2T/p9F21GcWBtYb07S2UcUWUyG9ya/ywOvw7OMalJ1xPHYuKpfph9rq6hJRiBkPO9FNIQP9jIrJxMoLnL4VoCv4K3CNhOtQEJufS6HQhghcC8G+1pow+rCqyKJNUdNpMxwL/BEvLn+9f8N8nLBSEvwR/XE4D9gAg4T0fJSrYHQtLX8Z1qc9UcTOeqE0bnQ9Z16Tf5QzWNhYtY2TCCCAO9EnEBKgMRKc6Kr8fQcr5Q5sr0STl1KSHqEkc9NwgieKN4FF0sYz8jw88TuU1cm9xb1f91PBni5Br6PXitClSTEe9Tfibxpx1qkR4dVqgMWtoG4owv+pRXj8Ut7yU8nN5sVihto0vF1pAXmfq8AFcUeyihz9xaf95ShvyvKtDkfoC8dZChBhgu2M8gLMHHjks6ZfTKbNL04E7Bej5OeVeuTCuxIGLELvuaC0TTvTjVzxrvvYy/HMX8fIaReO7G6m/SpNwHWHub57Z7gSO1l2fvjN7IREWajfQozsG+HovRUheAhFL7k7Qg6IZPYLXs5uJhFCH8MLhkMn0N8/krspmM8AJTtKd0Lf+Smeq39H8XMeJtxPe7Qm1dFVPka0C5cTWxIMVnUbXQ4BGdVA0fSFYmEAU+QHS1/UzsNCtBqIayIF4EVXgVOVTG4TJO73TG638b6IWIZb1Orja7ofFGEPMnKcXICYtfVj7Ca9Qoc+5Z6ISi6BCmgT4RsZGzIQDNJypYPyzs8C460r/e9Pxkku1aeX8eN9UjtoUFEeXlExC7Ut+H/6mGkrKbGU/relxaskFUctfUM06QQbfyS7NIa3v/cWwB3H/ZbH44xQHNQeTY+3MKtL6M/2ptpIHLwFYLx9Pc6jCcH8xyuPE7a3y0BY9erQs5if6pBWg7Jfr4GwBb+cCkx5ooM+OD6NHs9lakdzLtujVG6uWsbb8QTRJFIhPlxRklZozM61U2RxRwQjEnAfVSga5SS8b9DVm3kNuxmi1ht5kP3IyXvLP/2H49RgYg8ngAyLOPSE5mkE/Ex2Xi88UFy7skG3U/cE/yIjUbcspza9BwnWyG/mteL46W//sAqKFpogHCZesQPWiZyLnMfkp/mBlp3f6AOBA/f1hgKgexubaPCTqAFca0W8HrzeOmsqwE7SbJqvhO1x1zau4gWkPPrsUgzwvpY2Qq9iTJcv0nnQh4e1zOPVDXeNbZcfoxnI45HWQwPsQ1zjqHNTBBjmVHoOgi20rKX640fRDHBaRCHgJF+TYljAjUN7E3HaDhDeII0GSiDSegvDsqKpWDT+LQyD/7ErNkwpyw/ADGbTuluo96hRTLF4qmBlDGGrZR1L+WRqe7e6ph1GGqrSQDbAOGJwuOeHZIO5eGlDIP9tMlov19Hs/sKE0zDhj1rrVrtLnd2qzun4OnngozbzLkgMlWeybv+TOWYrGPEpJGPzDzhWthSOxrnFWfj41BMKyqvfW26ZPnFVGwUzy7L8L71RnbgG18BQRL7NJm1iPvUwNVZK5hQWR0xrHXHfH18JmcnDpX7D/zM0JMRCbCX/ZP8rN+xG9zfje0S5R/0b2Q2HLa7qFVXZRHvwjEeI0jEhvs9CwQ5Ad1XniP02uvWBZ8B8NTKdnUju/q+cdC5N+F7dtQt2IfbPR9h7SYSL8iescLvWTH9QhAFrMMyHNOSwjrYKdQejWH7COa8dkf9ZR2WTEXtNC3cL/hk+YX3RCtj4NTonc4ruDZZT/O7iL/k41zW/tFd7V5zNvy311sXh4fcy5LxaxENLXWT7BM+MrxI39PY85PiSQ5GrIibVw6sJkVjCGiMwY4q8bXw0cpLvQ7CfplE5pAVYLKyf/fs9Z2EpAI9ZmIFpf4ySTtPvVAlcrigVxvvlH35bQrUC22509M4vAzZui1C2qcC2tki3s8QCWHu0qI37igoVkIeJXCzzlvFaJ+/wllUxzLZcQZM+/Xie4PtAgdVu1SbD1ZRPnDBAbSEcrHhT+BbJ/MyhR6DtZ7LbfUtVgKg1b4jIhYtaa95rRnbimWJz8SXfmxdZwQjYZ0buCqYO06dpng15gdwrMvJjVLPNUzI0fNwCvkIufOaZ82n3pVLUmWALnN/y8saWXHFzvpHymX0x8K3Xm/h0s1NIUng1/vTa2d8o+YeN7HIAfa4OL8gL3MRkHMeJgTXdeO/kiF2xEqXepjEBigETMgLpYm7ynOS+WtZLelH9968oBex+FsTZ99aTIzjp7wHrVBaPuKsPIujQ5afK24cCHafMFVdKqUwy0BA8+of/dkbJau7vNObj2mtshXYvowWN7lYhRBMMQ+BfKDv1ah8pFsfN+180bzqz8IelHQiO3Ied3cL6QuGwaEmgtUi4QhhgzPw2UV/kzuTnWzi1eZIKfu7AtQp3BQrV7Q8SNeaazGRUOOyGZvuc44l+GPbMJxBELyr9DKypbI46OWC5ElyPDXwNEV9hlVndkzkE42Z+7Li6fo8MJB9SWw2Zrt1kRmBQ2cjWZiSWu1DBBcVGzWGdumj3JKw0XO3N8JwBqw4QqMvbmmz9GdDJ7V9/Uzjd+OISa1TWFtKs9w6U/lj5WyQ/W1a7+7lDFEIreiMpDdonhRRCZ4ioF96EVxmbbWodvCRSi3L8sxq5QlAyjhvSrh7sTSakQ4vH52D9K6YgqoHkLQSQdXVfA2aSmd5frrsnvGm2uWMqrMXqgJ+V3OsE/AZIVe8VG3H8MzHZJ2jhWIWg2Zp9B3EveJ86R6WSs1Jt5l+sGBsElvia4mkPUId4vVLdqmtDKQddy+GSQh1vMXTXJLywREYG9tKYOVtSJjjBXO4iy0UFmRlf/bPGAv7qaSzW2e2BJd4smxkPQ3wsmkUJiTe7G2hV0zdOmo0OmTG2J/jeJ/rAfJtYi/Z6ulJ0IYtpd1G/LKqKLnqXKdmVEsLrF1g5nifJZXA+Bh6J9yYq+5K1nmBa6eqq0BQ5fhI8euQb3sHNQ8vdO2E2mnXsKMfrJxvUQnyqFCMGaUMxPPkPan7bpGWGXvQrV+YMhxF9vzSXb5tzWfd1qeb5Ezi+k8ISO54JXGF43sFTbN97EVOxFbn9UYqxj41I0LeRUaH+0/qKIqWXNcT3g1w3ulPLb7Tmrp/jTjezhjH2JnrTKrD0roEY39bMjqiECXVt94tqQ0eYA50qWvWvqQ2CKtq498eIdproCficOi/d4C66gCdlw0Ca9ugtYNA5GtCZdFJols0vt6V5N0RxdFyBZM4TviYw1tG9USF4Bg8JrQybTucWO1qrhpADaev/5fRbJzJDkGMshj4kZQNgKAudpOtBBjTj2/xvzMAMz7oXHbA+wF9ulIxaGtnb7htcwQ0j1dbctc3aOsTFc4lHM1WYUcOMqETc9JxqODraIpRDLX0THytHwqTyg0K16tjg62/hytgoJp6uztc/x0TM+zQSsyHCY43wriF7u0y9cGuPJiz9KNIBpX/1oCvV3ZYTtRlXToBtt+0aSfJVhHVEkRiz1ZGvJqfQ0tOIySQnIEdbKOOimOylBl/fe/GTak83ksEgAzL92Qk0wrWptAAzzSn//VQIMPZfyORg/BmDk+LnnpxRSRaiTWiQQnhDQaxtQQihV99+yRCy0OWhHz/S1pp0B/XAURgn1YnzhgqyNECygaNf+2q8+u8zyWPaXNH8Ub7+Aa1Pb3GwHHU6OI0146Vv4f1RacWBF7CR19w0cNzYbs/N/1iJMxJTNZ+Sb8vIPNBLsipyA42WxxssMtJD0DHAxQSrN9C22hN4AN3S0PQ9CTUMc+BJfVsTRWFt7l3Eg3p0UV5rzA91HWe9Ae4DVV2UUbcFObPdl2IzPHJNxTF4t3Iy59TXxBzq7SPuycxrc958kjw+geYprVt3svMRophzhrABgzMSQ0f3Z9yi/35JNIMQwCSZrUB1xaXNwvzsTNbu/j9NvQiMG3Q9BNHjUV3JeXR/Pma7bWm7hfpEi9U6go1gKGFdu9VE/j00HftN12N6gfQ6AoZuraKA/wxw8MCD0AnAtpaxHZDTACJyuTGoje61l7KU9nyfSsFlI9ZkVkKK4wUNWV+7C2wPP5ur0vLFi90UuAvLVzmBe+6p6N2XA7JILZ193669lxnR/F0XEoUfdAbgDk4QcHxxSZ9FklrRs35QbcVNJwEgM1jpnsMNW9ivkkLs2wL1HmP2Rytk2XUvxtQRpVEtNOFTJijRLBp3ibjAx1Hpn3nq4tjKzDaH6CKzHtfimmLKo/jyijFh76EUObIONCO/4xPhE/CtUQ90i3kKy4/mJffwD7ubFlh8SQuaVH67mTt52xzKzXLaVJrbgFgMXAu4CAiGusYis8oDoyqLsylNNExujuC8iM86ObNuFFvhgzYgjb3CR2KX/RG8/WJ054hQjfdioX8mvKrqSvrCNMZGi4uIprDxqneVKoYaVE7xxbUkzPWJSFTcoM2Oebn08Ojjn4OUwR+DLV3j5YUD7M/Nd4K8+XSDwy9Iwm3Hxw7VKSoFJE6wT6Oz8wERwfIOK30/DpCNw+ObMYMs0JzWlY7SWdkWHgpN/2fd6vPgyvxgaQty92bHT009H5vXWNTYWMZN1M1fkb3/UJtxJSi/dx+VVA6flOYVrnjFOFqsiIiWkq3caAhRhYFJr1S3NIkWXHZFYH4fvhyldiufKn5TDpl2uHu7sh3B3CKDDXIKi3bWljCdhQyy2o66+6UJS34hM6SN9jwMSPzBoIUR0w3yd19kxz56PAqOhwcwiBlwI6/4MqecPTPd3BWOYlK6JgqDUgcN/1wtmnFbswRRz6DVb7zpZ1FXFIouTlU+1GLdUBA0Fs932Abf0aqouWo9nGADOfSf7pam7Y6YURUb6dYpYgbCIyW/gHY7xPgtKpxlKohEVZA+zuyD7TNOxXsPhTRCSOETAeYLQY0WepOCFUFRBbL7Flfg+fSp+Tyi9YVej3KcrmePyxUI3+zzOBNWJ0QuNQvhDGC2tbkU2dy7ymIHkbzbAhD1WIAkx0jg7A14ACta3ZGqQDPmYAnETz70wT/7fxmJlYOWKBJlm3ie6cyGdy+TX0/DJgRLieBc/hAZMQSBVt8f8mOQeUhr88h3i4zQ5IPK07bZ2ZnvCVFFhy6SNEQxvYT+B4END4DiyUlMZxvKWcd+DVArKrDuENK2sExeq3a+Hc39y2FyOhABT0kubjOL4PcqtzF7CQTsBURbNR5PqlvoDsgTWqLc2uYF88y4Z8Zf5qHCrMltGqvGlrR7EY3dxcbJcFvrlMfCEzWEUstQ9dGocLa1h/1tJausMPAniL1CevA6Y8759sgiK6sOYWxZsEjrvfnuyKjAgxPAsLGZXFe5nTXA2wOiCHx/Rt/7BHFwBpev9pGoqGQLleh09eFyU9xbuVHHY3LFpfbiSAvibesMDXGrBiE26oJKwIVagBjq6LoJlzeigXMj4RQuuftujYSmSOfgcMuYAVzfCJqJyyqfL1Xw1T88jORktW1FSsMogaAy7fphvKd/F5CA5XpmKdyw2xFWm2qRbGf91tzmHACm5cYuB6+R1ic/+SsW/b5v5DzibBPJhae45CzVdoUtaxZ9qyO9uZoFBC1j9gWb0eiZrA2B9vHGfP+YOQILp0mCebmWj155KE6D/zyU4L2uScl3+ygHbcyoqB2h/Y1+NKqdjh9zy48a92kSaK5opH1YxV1c5b2Uar/tRETixZ9I8PjwvuSuMSAI2U9ebNMpvZu/ntYTWoodPXAxIYfUbhgWgdsjtBcC8m1wk/w0Fgde+vixpemPsJexxK2wgGidbOyifidVf3BLW64PU/2zyEoSTDpSkeYin63e3T+V5WGfrl6hBiGXkM2eCUlp2diY4iOo+Mf+63CVE+3NYyiQjyLRbASU0C+pW4AfuR4owcykWvln9aiMJI+68kdebQfcJiBQEj0Gc/Z0i6EEPxPGi8TAvFZrsP9sI8JsWff4vGEknW/hcs04nb9ijcQv+dODtdoZjStMv0PUwprDKLmMKANZov8E1+APhk7E31mr6ZguRmov76+8pmPQ+8cqnCmKFNJfncZOVokRnO+/qJTq/gh5m88l7y/q++dXqq56OzNXmuQ1UhiCfOESiNjNm8HoClAlYsIHgZXuwQpvI8AdJgNoInaVxp7NUii5MdfO0yoUQy+oedJSfI+Xir/NsudzKtKRjBa8CuVY9GG+P/F8fpEN3MBxQQ/xbEdOLcKK/Bp1X7MHfHH1wdVHt5WSKjzqumElp7RWFfsI/K8scBqWVu4qij3Z1yrfgBSV42bzDCJT379nWWvjepe4lsZgwKNuPoaQZ/gMFmpQw6umpK5tjYXg+VoCJWA5CBNTAui6KJtXpeBvvrA8BUtFeEXh0MfLcBi3WfDtDO+8cpOfstew5KGq9MFWVML47WLkCw0QK07dwmduBLYmS4EHWX4t1e44LC+XA0joT4G8ZPQKHs2sfl0oA9Dj/8oM078TSHB+bTkm5DZGrREdpx9rg5NteDCzKRtd7hkXnjDsd+h0PUtydTpFopOIU+PHWakokBOrRjxXemRmYb2ueFGP/Lx+59+kzKBwU4n9TRV/2WTzV54V+V0EdPy+VOWTrmS5B9vhd6BUmyFhBB683RPDcqDmP54yAJBQl9BPAhoaimCiX8RqZYKcT0O5HwGaxq1w/whJ+wrc7kuqxaBhcvR+UJ19XhUvMwuIpvzf21GEjS/sQuMa8lMeWzFY1QbHqFry3fhiyXpwtul/cMRSNCLnZzgbqt1G5DRn6Pe+Z05Zz8/CCRQbe1bmwX5IooK9yxxhGzr9PZRj8ba2EFFeiigxPSC1QixJlhmQpLp3AeBaqpHeKRd1lXhbmTVfmZVuLu/tNkp5VloOix1kMwc0tuh14PnR4qRP+6qnOzMmx6NqjJq2X5hgZa3CNs5/Ve5d/LUMSqykmuAHOTglNNxCmvX8V03Inau6ddHIp3jXixMoR5FN7Vn03QuH66mtBHkkajBn4zUX699E3W1itPo2J6dwqvIabZJn5DM3WGMaEknBP4bEXAOHREyrLlKoDpcaVexc2Km3UkpInYLK1vgKu38/a/L6zwwyS2g3TAeZ4lBMCsm6e9ORV/WBC9+we/I1MR2H2sTPGNPaSju85qJYgWXYmmKAgkAHI+UMbRNYVuzd7ZXlOkfLcmwar1NKnEMt/CBiSqBiwHBO3NWZgvOJJ5uixwehYsqgivpWSlrn890NMBwdbwIuqMAGqH6haVW7OBDWotk6LV7sefF+ynsRoxD2hG4nPwbb4tSCAjoD0WE4pyT5LyN56q5qZEpm+p3vmQ1lTeH5Wbxpo5A+qPpGrYsLuqRSbM88yvoA5vrgn0phhNjzQXqlVZBn3I82Vj9Ycgvh2qtl54aNn1VhsRGIt5y0OJRUaZ8zrPoAN0jjDldOhTo1Z0Xq3mhtg+NSQbnLDIg9g/d8DpmRf5AyO08jyXlAre/f4HxHgBu9No2sYlFguapVSGAayTPA2tUrEJo9N7j16gyhFaU2KZBeC9PCxUCg0w1spiMJwNeuWZXxnkMDwdCSgAnJw971MZ0/1aQC64ovpTOrasMiOf4PMPCCpTKKsGr339oRToFMir1C92BShQLBnRsCS+7fDa5QzE9zj6f1u+jxRNsqRwMwziZ1Ix/V8itPMJowW+d/Nrx2wTI39lfy9EoGrvayD38w0Kqm6gV4eSHTxjjyJTywj9kqlOay2Ej27tNiP5cV96imTX3yfj6+pGn1S2bPwtkMo/9JU+CMkq3mB8JZ/LWfJDtqF1JgXoVEROxXBk8B6llpa4Lp2/b3oDbjOSYMohKxjNI0XpSZBQsPDewjeCBwdo+edW6VRckr2NEphYIwY1r/tPsov3FkN+DTAWqr2nuv3GFUaA22a06VLYLZYBKwz9pIv5aSmu46sCBkK2eeHF0zzBwZHHztwDLK3Xk1H6BB1rVDGBRjVR7midS57s4EIfOCyTeI7XIaNyYNKy3enTJcQ9Ph84BeNcLadG4EGu5uXPhBLlppMnUeKJ7csIEGVxDo/uLjuPqEe4CeTVf62lpjHOtG/IBrmnxgG6MI0VwDfCj+qwWknJpywo6kBXDHyjrzVacwP/kzbSOX4qDYskbkoeFdBxTHi/dVWLLpvXWKPl+k7vMGgOA4Iq/Thjc3ZTGC/VF89VmsPzqalbcwJePKc0l9tqye43dhBIPLcovkfYjj/Eh9R+MdFK6Tq3IaV0enL8dJAwaGuBWCGm23kGt/s5tr5NLiNaKnRF0waYeAD2kVxXZkPgWSSGW3I3vFpMqA1BgEZKAzLjyV+DV6g9xdBgI1o/X0LpDVEUvCFAhMJmZLHfSN5v1PV5GmSa/X8IWTeJ3FACtiqiSdIl+avVX+rdqzEJvKhdBrYV5WRXPCfdWdoJtydsHrtYzPspnuZC9h7E8FbLvmUe+g2ljzdnthcMcaaES5WMtV0zg5aT5IVDppRejOZnbAQv7GxZZb/4vuKj8y/2O5IOhxJN7U1J2m6Oz+8J1ygaAWRHINok5433phkCw5wnT5gGlJlZpGEixUfgzvUAL4Um5eI2fokVVbPwwvvgvuB+FK+foLI0Litiml/HtkaaQ6bdKQ9zkNpg4XxtD31Ft7XX03GTcpw3HSVHuc2VoNqSw9DpVKnie8Ko+OgmzcjCOupuIwFCUpbb1ipst6wC1Z+2Bbu9roXeqGPNeAApPPOKcw489HkytrWo4Pru3qXVnbnLKjFAR4fCnrs4lEfhi4kVEHuSlflx2nx8cz0+XW8qyA/jsEmNczARCTp795FG9EMv4hdki8Pi7pOA4ENPu8P6MNo/9OjOLZ5LtU3Hjfl1xXISluBIZvo1NzuhEjP2SBBOO4Sezr0IxrFPbw0Dl2/ovNL+2JmRh48m8STQFx3t8qAm+2RSKhVmMpD6bjxRwz+yaVa+hhOmMKkjDcq1O/W5Yim2jXCOExEQOXiwhbvQV3qM+oC/CmS/yGFmZVTrVAhixYcnC0rgaA7eWt6uN79DAyr7H66x+74bOIdjQv/F+63omVezBlIKtakGQ2kGa9TYvBXHhniDpBgrrX+wOBvo3p/gI8A3hmWqeosuC1r1vvNbxAo6b9GmGjRWGvvCM+Q0+JA+Dr8ldPPk6m5OMW9dWWug4fbmk5O3AtGylh+osjVUgfgv0HK7/1EfSr87AtKIPanL1A51RT0fejkXvs2uRwhcLYRN2ba8hLBkTCj0CZGLQ/OacCcyqJG54MqpE68eTrp0FclU+tzPFqGmVQ3Yn4pvVfR4c5RoSOz7p6ZgZBnk3PjwBa8uXAoXdQX9trUpLKFQbm+9LlTKNwi7qtkEZ+Rfhq/ITxeRL4XYWLFKVyzjg7u77TffRo4Z5TjtCQm7eYe9OYhE7GHzM+86OW4P4YNrXfBvWkwpqOIDXn51gW5FwtkaKIn7X91vNTncNR7rlhlK3g7odjZqo6kRh0rdYCuWdAPCT+YWZcKPqWvsEJ/vnEQshvD5tAP2LSnWoUxqVs2SMIWtezzUYdfPmX5W3rlAMwnxsGbcIrbNpfEUHl4Z5waz2fWRyz8xz1u5aE9FTM5WY/IB7nW6Ej2pddwbDELj1+XUB1/MBWsXrfiPOJ2FyqBAJAzeckOltJbZcbFFCseNVzk7xR6Af1TpWrs+IyvLK4l7MYFu1Afl+DErTK+ScNwz339742Pi4D5adBWGQf5FBjW8LMwhhZPKBM5QY4XlrLTZE4vgCgpEpAYctGu9uCk9hRpdL3dR9kr2aDxCr8HnE6t9EbvNAJGjADdUM1XO5yGQ73fzcYEq8accmQ0+CqTPubbdDNCzI7W7K4sscKcp3hrrXm9Pxx4B6xSoCacxRFa5NWd3mGHXzCEoGWEg8HTuGqpjOKj57Ub3g0jbduef83t1DXZDS1eZnmvbtwphWkiAyihM0EQ1e2bkuHaeIFmYasy9n8nAoIX3Q0fGOxBRcyfqyfYuF87hODbxdKGzaofguLmS0e/+8TNZi+BrWmQuSmRtHoSCrIRuiihpVd1xmpieAh9+yBJjQOWafGc+ehqnduVN3cD5Uba+HNphaUXCOkA8+WBVH1rrG6unXfwcjNfZwMV0ZkHPiFy3SqKi/F5TnMdNLX19P9FSe5I1v444fZWu0jHgdHmAYfwXyDHd4zaOsuflnMCa9EgVs7QeJEFc11HdIX45ZrjLgAd/ohb6O97QSeZj/Ed/H59r06lEfwn4Op7Jz5RjtxCRHOX25arOD6S++9PKZ0+BYtkp5vuiXwl4RRgbD6Qc6XZZbI7GH6jaSKWXhip0WbopgicvAAooOZ2bYIgEpOqLCgejj2C7TvICsTsoB38kogeqLW7vEO664/ECTArZmcAvCHU3qB/fSjE29Rq9FPK70abCiP0S5aLdqAkMg9E0XX33VkObrFRTBRRURKJw6UOCmIQ3qzlJOo7t16vmYOJ1dQB7OyVBvrJMlQob9uvE4PsDoL+Ez9LfyFw4dNouc2nmZlwcH9s9aRyMVCGD99CHXfIFbPwdsv4EOln0DKyi4pQAS/w6M3bZGeJohdoK7dkfX6ab69rcsTeYXxKjgabuwIno5T/esIAUkgKIUv3LY/YrPn+BtHetdSVUUshQTMzLk5Y0UAxr1WaGBrlriyWMaqpA1Y8a1hDnam67Dytpg3bOOX1oss3bJIEoFTmh/PNb9sKeX3O+zltMuFm8NdYJW905rEV21AyQwFP78QS8EvTXClkTyBbzc1W2Qp+94VntwM3yhGPhDImpGVg95IdFrXNE9vqDlfld9ttzAxjyLqPIkXJMm9kH7ily3GHYQBqO04eihurpAWgz0k85J1bAE9gWoLqgjDnY9HR6R7tDmr86Xju9lJKox4boZ5lHvVUD4R9zMVxH5AV3mh1NfFDhJLVNGZsrI62xlks8zkr6zvnJeEB4Fp2RnLmUosNas5vs64BAAdulivzK5bM/5SoUoTAptbSPky+r0rfOCjwPbxn67flPoL3ctK4tfVzc6LnjzPYkbsHBI0r2USnTKWq1d/c6mJ4WsmKXgCPADBQy5KFsv95VfClC6yg1mqDiPCzZKMmmdOvk7H7IDNs1jeaeZjgRi2suPLaDTWhwX5XhRapKONRvEf8069DaxaQe1/RQ8PvdLA3HYCBBZWFqYwqDtPWb595FWnrubm3K9Lj9jI2ASO1JU87SoxfRT37ft1ayvZEaNaPD6icWfsagJRkFK/TeLtODJE4qJ2/krSF7UUGpPWnZ3/Jp/3AFLYnaAtkianBLNr4x+0WvdXtfXR/g6819/TtTE3yBhzq7kdsV+Tc8FoSZvo1Q/8PC/BZpXrvs6RLHuhCYDNHW03DxXqpD/ssAc5rLfajEQ8h/npZAea2v/3fv7/NHkOtIHCwFgdhaHopXESQGSASQ//PKCL3kJpzFycCC3eLOaNIIvSzYtAYueWgwVRgSmOk5yF8k9BcqjBSRwbHqRvnDJwsBU/27+WwM+56ciXLkJDe262esVB4vy8WNz2cK4hJ3dxsDzS0TPPJhqhYz0rLlTMoK61Otj5gvr498znLzuFg2dn/h+pk48TJyLzjyuUVGowbSrjkXtK11dvqdhppnIp9T/t7aBCwLYsVFhbjQPZTJoignRmgbeRQcb7S8g1W0XeL6pS1/wiP3YAfge/1/Wc6IfigC3cWuB7+O+HAWtJiKc7Z+mjpMvhndCQHB5j0Cntu7GoZKvvwX1DmRCsSlEE0Wq+4SMiYZ4CFliBJj4mZ/duAURK4UhD8WC1qacs4iusieL0PUJGXcLxaQ+rhnfCZgBTXHeVn51ruhgyFKpB1l7yIHzeFR+FKMD/0Ca14syqDX9O+eGBa/KalosyvhUHntlcZHuPQNXdpO7gZKA2Y2yPBNSaR/JecvD1rlgmpjhfWI+frUkAJv+Wgzg1l/hvjr8Uc7N+q63WoK9Pf2+v6xpNQwZl1HPU18eJ374cCKMDn0lNmGXnxpQcacUV3VFQCg7Ctsj7xE8DMg6lezYjnRTqh5rfGY3cEFLUSOlP45diRitni+Xyr+yClh/8vXvTiVWqJFA2iy5L89OmZ+4bn4mGeWUkso9Sp2Mgr3Xob7RYPH8vKCgr2WdnMEUwK1VQ0YXuf4mzE9PemPGd+V8tEMbcLKjXalSULPF/F/doHRJKaau0Rn4pqvw8YwT2wWICDB1hChcDdXzICnT1+WpVTCVmNKY1nqBnUv6ZpzjSIUnOVp8rsYrZyAWMZU1b4Q76gKNDWqBBdGYNXsS6WNSDHvcsZ1Y6vwPw3cdhRp3s7a7Gag9v13y/7ja+ynbzrThua8J1oSXEeciqvZ1YwTBBcr/DjgV8T6fqAlEhcPQvHoiePPvKDETXUOL9UCS+nXEgIxYWAniObTH6+VjyDOQeolV8zGCTqGvxjLFqVu1HVAx3MWN9JPyY9DKp72C1TYwq0RkYrKULaJD6IfHyUogYe6+Z5zagV7WbI3A+HfEB5sWMyE6nDbPodXIjblTBgVq1bmdiTy6+XCVkwCOfVpxihkwBWC8D9NbWil2fc2E5hrtTwYQUWRq4zcTUTr2zG3Ts2WmnJx60JORMLF1TQeisFVnH+nYQbtT/lKqVcIVCpK5ulIN44lMfatrFHvbsuTIEavVLS0gR/m4kA/xJDIHxz5id0LUbYZKLNtAOLcPPOiBkwhIQrXLSlAfLb2Ws7EdUmOsNDZacagaN6CfMBAvUlJTkMwgDjAty8HB7AveKry8gAPYIPTiinIyLVXc5VoaCxGEa+SgJdy6fAG+2RmhH4OUB8daBW+cpyxpyNG+ebUAF4FabG8rxMvkW8mBTbZeUxhvucXPH2WuY4nerrjJl3GCIHTULGnZhF/KIDzbVhfc9wwfPCMfQ9cId5CW5sZ8Awd9vSFtHton7B+tQ8CYOmVBRQJ1hie51lndvnvNs1d3w0uAwUvn0r+5KtiBq8wdURBf2NYXewQ8j5gVKuUdcvJyNbNNczErbqYkayTs5cVXY5W872IkXWwwmxEMBHiPwAaJ2M3QZFcUZYIrahHr6rBoRcpna9JIRpejAXAhZ/43ivXbu7Xd9Bm8rdRxfffSnZt4VadlJ7UIERbRB85M17aSFifC0u3josBBhRWXEDb2hzGYxaUaOec4QZ6UITXHi6i7K6jOKAW7uDx5Kvu9QiXN4LCUs4OIiq6nR7O4740zxerXNsVmcWg9Fuq/8y30Gw3jIM2AGHQTATeC0v9Y/mTykmaGKBPlX9GHAbJmkdyhoQg5XDXMuI5EbzGXsw1pm4qWygpSdAydcCvStbuAWh1b6LGbrVTVGtR4K+5prLLqLXORyel4ysgwVK5oVL4ZS/Pxu+6ARf+ApYtBNya04C6b1JQ2LVYBNCSeUB6LIqzzGMwUCl0COSWCn30jknIZG0Oy1HWWuEYTgl2bRMpl2wZIyY2s3UEJuGRHcWl8yed5PUd0l7bgLoc5Uzc5tcnK/JDBTv9mXGVrIYaNHbhorm5kctZBDvmvq1xcojtq84qjsF3Zl3hOAr639r7Gc5e6MrZDZH9Xnm2eS2Pyg5pht4W+Cz57VJYxT40/ZsK8sf9frezkUArwCVN+TDi1ViArSi484vevvdUEYGVUxCoh02dubpqMjMyo/TRsnjo15b3YVm+Y7A0UEr7bqehebBWQv57PpH0Vj/Rt0OjzSpf3SzsN0F0bZTgiAu5mu50tvAchaBnbw1V+5N11AmSI4rGmIKqhYK7TUA4Ep8JE4J0Tfr0MzQoxWqtvlLXU6hDGofPAobs7lIsvKIeRpfqtbkkqUgHBB4HDrFW4HPa7/TAORvj61mB7QNU/pAUh6TMKGrnhSLIRHRrPIUhubnS1lMWOjD3VabgeTPgGFXSAvhblgpVCbmpuTuZ0g+oJQr2kFiszOjYLXlzNm8tsajVRA5x/yZ6Qkwx7PH2o6SrmFYqIDP20MjRWrd2nz4zYAntLtVzsTfNdNR+lJztVFregnT1BFqoKyz97MtbSDmFZ6jEluVHWpvU8tHSuJGtQEpgXpALujm7CihOqtg6VRBBmd5dvwm4EEWi3Cd1v2xusbgWn3vNUe2hTmJ5TgCstq1/pPaWP0a+cotmyKdvc35q2Jstl5YWVIxnylmMg3Na+xhwz+88QmGlW/rlBeawIiCV0j+6fcmrFOSaoXMt74wAHPvf8oUSK4V4klmwfXqlQpxwAz69Bk4/5YbHIBDOTFKvE6WdFSi66xuOXEkxf4LBBADJG3kmXpIBJxd3Y/DXHQBVF+RTU2MjRjTdr6iX6+a7hoxmkEakouP5BhO2i9IajsyM6cDukrRM4DT3aB1AQT4WvUK2i3BZrebL0Mk9eupnVIvfIYighp0dOHjyCJL8oxaY+IjteaRmfGpqEJmdAhDPwb6pgdhvCQyPcL8pwmhz5m+EoScJCTj76fX3Asv7ZYjHZmnsPfufvBD5b6WMdxt2cW9frHd7ZDcN9gg3hhLvZJDlBAc4qwA7jU2dAXvkp9s8SeXYwNP2+CAsm4/6UYZ4hv5iKO4vrAGXOtKqpdygjh00ZMhq9zfZ49Yz9aUF+Y+zVrtOJGaqGD5wA0ocdoCba49AZoTOnqGKFB0mgRvqodDMQ9HSx/su23ZMZtDB+d3K0aJZq2C1p9lHewS+U/gSe3qJKsMz6uslqCjQClxZY7ce/1lgA5nkl1fEJs40RT5X8z/3u1k7g9mj1DqYUoxOOrTXZ8FiucrnVlwrjV5eayK5WIRo4HgzpcB2NsuvgNcRJd8WprYJLMgYUUcOFLfi/Va8wpQGaWDlkhs2D13WNI2H8JFvhyw1J6p2m/nEP2C9MCNi1RUnGTqQQ+Ggvw1IzbREtWPrgFbDM6M8mHvA1Pu+FARMeXRNfRh8asFddvv3afcVxUmNfvKw4GHUyrQFy0wrEEUwsxxy23dPQb7a+yNJrTA97KQ4tc1bEanzSTLewf9BDvwuNu5V9RjPjUk2NFOzArctHdSFNkiSWeKbFK6mqsUDRV+daqAElwFAuU2TwslTMoUrzcFILzon3u1JtCoirVWvJLRuY3bMwAnPVxJwuu2FaHuWVL+jCIcq+hqG/wFKYB1WkYqkoxtzHEw4pJGN9utvRS6zuyTSdV9EDzyXOJlsk7DjFxjx9kmXlR0LhPo9c0PD3oVdQIU68opLMgOjwP9VBNU7etl9DNE/kdlfcsSNdKxKaD9qOA4PmP3nGRBD5SJMOd2CJ87aXdaBGauVsTLLVaLw69M2QMh9vCTWWXYDe/fH5fKVO8Wo3XKWbs4z0+WxJQbqvJHtoE3y4IMQ7LmEmgL58VJiRBNfUiTyRZTrM+Nr6/FLusG6N2XdQhhNkqivN0MazgnJsFYwDGRrboiALr56p7nHciHIvn7MChqeNpa+fQtOEYLcvT4gX39sllsCgfq/U51ZWZHJZR0urhp2z0Ts9QbKFhNHy5DsuY0twNGVWDWGf8IbcAke5GkM5hN2se1oSAYsJ/NaRwdJweIh4BIZJe1n+h5Nwr3/FkxWQYZxGJgcptkyerFCTuH5IY6Xpmlt1EcVHY+/fq4Bq33EYenTBJvTP7XTJdNB0o8D8QenjCK2durBPrKwEr7OHF4uaD9bUk/26S0UMiF1+XFZV0mJIMaypD5EK7XEEOblXjF5stHGc7UBWbrASsEUGdTrYZjmgsjFnNVwem+jkI7Jj1hHroGcISNgD6Hi2C+hksyRpWk03PslQjznuv4qnp3nIL1o7wo+YkQnSbaL5G1hn1OqOxcgNGD3rZ3jY0W2V/eaevs4EZwKaLoIgb1a4Uq0Q10AOJLV79uk2/mUZnu9fr4C9urnmlbS0J/nck79nYVfQmK1oqGY0VpzHeq0pE8pmHxbzKnMFLsXvnretDmzNzTYntwELPAwZasoWyCZqo4SlfGoWJYexwkHY0vh7Sgos5AzBnu1giTsAlailcEGDlSfbDF2vy33xZddwfqek0cEpJDk2OtdUbTGhCoN3z+iAFCaC4nR0VcZMdQAvuqLpMlzPyXwuV0FFPucYQ+Cb91Col0nfOV7Ynjx0ZfePC5wDOOvxoPFX0dtJh+yrBcP6SoZkU7psXtpy8GbA8C6CNmmoPWjfWDFX9fwsix4Ez735a5G7q/RCgthhgPnQA7+Bhfl6r1QsVpO7wKFapWelRPx+EPwXQV5kSUwKbjnStJXZ8JIL8rnG2FFq8YqO0Wp93LoA01pOp1lt4fCrpSx5EGpgd14S49ftmDlbXVShoumTkMKlXP3Jy8ZRd/8zgL/YAxK5KayJu+K0rJHT5dQbDYKv7m0xtfVOQtzFqhDvd4lMXv9ic1wXx0ZRhqA7vUY6euo/hCPhkXdE//OLr7KvbaQT7yBCoW3uRbNMXmIdAl8OSSQDMN61osEUXON7ECPb/4sgcMbiLhoCMHF72wMSLC6ay8KYLo7Q54BSWoaut/4rVqsLYWMm1etE8TDrmZqAsvICp3DKvJCJsjsZvshxrzbVjvgX5QiQCIiGkCp6PuHHxO4dM0tflVxKZ8c7bfRvzl8EEUnyFjqiTsg7+4Xoh0CNSoaIAbxWp63cJAdSl8XfVEJyXIdRQK2CUESUap1oI6mtwq+3Ss8FApwh44+dweVhrN66IsrC4QucqjxJj0OvbpyYgdehdH0BlKDs4d6k+R+4SCL4dCBeJciYu/kl3lhN4J1d7ywodPwTK/3cCiBn7t8UCZUQ75trDkBTwhsT/PUgYHo2iee/9zufRnL5e/O6H8L37W0Qdzc7HWIpK0aqMbj6gCLRuQmfdtMhrERM3XmD3RMopdNLr9vlHwa+PXYqsRI06jfrC7BsJFW4yaNATSsiOZEuFnmG9JziL4aCeyAB+cDQq+HI4jpm6pGhb9PyLXef6QPkecmkDi4Pekd83VrPvd0nDjp4UI4vHR1Oks4qj+L9sYPLQvVXRLUVSQuJkxtO4qjLRzeKnV0NHBRXemxLyttZTdPZK1aiXnT0JmuRS9PVOyGFssVByE6vJQBnHXcFh2mJJkPAEdIUD8eGXTZ/UbeIgjZswFV0Ny0/5x+E3gZ70UwYMjMqMDxq1V8KatxG954h5RrxIqdA3w9iRniF2iv48YDFC5u+aT0ho04hiHeoPJz5rUs52t3aw1aQwFHEyqK5TQpRe0TCSxAszReLLXsbLRDzffMAT45CbIV5d1iDgz4QWhw7lg5iCXyS/0wjh9x0tL92Xt7r7G6Ic+mWS7V5uy5UP3fXs2bSbAlFahZSZeAbs7/M65RTUnuD+G4+iZtT0P5j/myL7rpJTVraywxAnOAWWEbMeh8Ie7+4KrJO1+IqEm/AOgo0sGfQza5IL8OxHj1NFRrSxM45z+AVPuPQx6e6PtDtMWH9gG0HAnUI/nxLOTVnqZnyuNtfLksLaCMHpRrEuzQbm/tq0n0TrSRE4BSdEt1Xu7ymaNFObOtRzNhWyhsyUzGs6xS/Z9LPYqrpOG1TSKS/C07fQLRDzNmr3gcnhCewad89i5cBpux44U9BUepJUO2gz5WgNwNZdWbvTpaaFQHSTvKDQ/0EznBeZlYaJznyIvyt3Y2xIO1InIPV92ULMB+lgUS4lkxFw+SXnKOUddL1jmMPAUgxKN7uiqHmz1/2HgWmLATLfxz6T0CedvUW/oIDHwXnY2OzpZcyrp5xhaHo+7XnLOcuPq21UUoyyL6llQlgvArHPt1sWaVLcbU6dIIUxFOp8EuQRrveETBFGBD8p8xx8XCnNiWMu4gqs9W5DIo8QLE5GwRPhx5dwjMt7pochAcL9/xRuOLtxssAKpAUR9D4JwMZzexDsuJGJledPhnGHoiXDh6b6fDyggiemcCg48TNT/IlUCadMDOoV7Al2+uwunNUapjm2naBgYBCZ9QnygZTsvB6l1Tu1hW1RAhEk5jxxlLcssyo5C0vzvUzIU4SIBRgraB3UXUPpemkjYWeaF9Se0ivaBG/uGDkukdQvyloUbYXjJwwKssn5w5sXOfznxv2LnENdspLlXMYJ5KG7A8daA4eqdkWkFyr8/erW/oWMZeKIadcjiho2o55IJWjaqgPN1YRf+MxG6RD1DJb3UgKl02K0gf9CuvvqYAJZ1r2tM9qsOW3RSjyTkrejFL6bX1iaUoK/ioHA6/ZLfykB889DsuEuxfHlYJfKTl5ze7TrwgVHTVM8HhIv/JVVEES5CmNSdkbK/qd7M4i5YMvawSBDLMotTLyrJODlNDp4S3zlMzhozypPcapPf52vEyAJB+tsUwoP9ItybIcARkU4QrNwQbPYIcz9X51nRRENcNOwSdHfD1qbcdF5aph4mUAREYZPbtWwPXfgDqsVww9LwjlUHm9JUQ3OXzyaAdcTh2LRqKH9VpQrjn0TLHUgX01/ty9AAINLWMJn5MXdK5xlKeNfUrZ+bON7n/aoEQY3EJaNtsZNtpT8/06E5OJiv2ef4ngGG5ADOFJwmJU3etdekvgpH8UOADZ6oRenZr0+VMpzR+FhIWUHuSZUflTwG/U+OC/nWpACBHKnQ+Cq3lW+06LQZ8TttAUoiREGwHkKhuu0I6Uu/AtCAm0qyLPHDGpICduL/b+fqVVfiR/zrb04LJk41R9Z3i81H6ayCaYPNy+Is7uhEtp2GFYE/leFXXiAHEltS0QpVbHxnUADLhfqnqEWx3PgLZCEkWBArjDvy9pgclUf4StwGYsiYUN3YhmVJexNcufhapjN3cIVaXUFPScFKmXTdn0nnZBm4+dS9fqzDwX9VjAluONsZz+RvYXhHdzQz6u7kEqVA2fKm96xVEuvqoetEGK5bo8MFagmv5nn0Jv8eZXGFkocDSGeAMvJuy8U77lEVsn/YsOiB+FpyYqLEgYRM/B7pxH4j5HYZQlr3lhsVxIGWXt6Xdvnd8ffPmIDZa/rE9wQ0xvAcoXhEtCWT52+ddPYsjKDgUDT7+DK5lhClxBWuZ8LdfFVxxiei0fJ4SwuHBFNmVpYTLkqK6iGpng5ACbcOwrHTb/Nc5F1jnpoR5A79NGPgA3L9XiZSQ7qizar0I+FbV1hacaxiYf61vxwNTpTjktB96yKg3weSEnNrrAmPxGRusQ6d2W5FRdqmGV285SzYiIRvXBWBZD4TWC0UToRtoSadH2wQDT2qgvQVGQSjw1n6tEE4EShS5T/9AzUTDaPJXsu/gjL4YAAAwftpPlwS9WkQpTqpJ698DxoAuQ+w0sa/7fcEzNPVmMICvjWccZUfsa6SS52GwBo0W25gr2V28Jz84nbVoIiNdTAnqseIX6/l4WxRHMsoRU8y+XVuEN+/o5Mv0cgfEEGPG66moV7MKER6rL+z3bqzdsU0Sh9UTrhQZdwX1IMKNgMmEmGQfIFbOcW8xG0e12QffTSjN22B2Io3HemFNz/TmdYe3lbcwHBGBJuONcw8EGu2jwRdELKWeKGx/akOyV9eBlkJ/txhZVyuHercydrajdYAE/J4kAURdYbKc9zxkenTp7ds2QZZis4Oo5bW7bgkfMJexQCbQ8+9Q3OTyufW+BVmKO83ipNpK4wN+grBBVaJ+LwHQk3m7OCJY0mjbdDP0kZ8qCVOHrumnU3b3RKtKXjVxVQ7pn/aiQUXKVmeBpkRqE0Xv8qxwMZeQE0ZcZUGGfq93VDyfHXYwUJahP8MU48O9D8qkk1BAsTaXBIra8APWMWcDDEdPtuKbw/8abVaArVt3VDzSaey9NKXg3bzKUaJd8HhQWKA9U8bCr0W4CqVhIt4UwAtF+EM0ej/wlaO1Xi/1+uHmWJ8qPCgHMCnwgRGwEUvfcDP4Q+5I9jcYiSaBvHeM7tSaLpdIyawN0lQIO4TpcLETKQgwc/msLK7dLXbSdTz8jGcRM013dZzKbCJJaiuGyqqhxpsCr3Knmvn0ZLntDHGmsHOedIj85bFcYCoUp+SheNWr7v3uywSDKgnUpvy4eOYme/1qn44wnyORmHGZRTX3GqAgaCT5INiL52U/5KxEK5WEZh+1ombRIbzwY4i8W//M1SBWHnsh0mZLI8Y7qz+NQUE+gYbRD6FaW9FslujWv86TU7FJggfI91YMm4bzle0TQmSxhsBXyd3znvZ9etPR2NNaO9VNJ18P5F+3ac1Cc2zmB5Rxh1NW704ZovR55h0MCHfCVqplqz5GRX3QeSV2TySTjhLKppkxy+sOFlE2vHAaB2BHSr2p2NnUZ9dyv2tlIsWVPBPCM5R0t1OZjkAXCcbRz/Txqyt+NPUxqqed/y1eDuHe8Ushs6raii7QW7b1i+W6e6aWK0SoKP68VR8+noq1A02eBEDOYeo2pEmVLA19fWz/tVB+bBtoLv8Rkg6fohM81kVVWHNepx5f1hFJbNBsA6Ht05E/mjIRVQiEPs9XWgFR4mbT+qU2x+RKRe25jDxd5FfVoH0MgHIO7ky9CG68i0XhBPHRHm6XUpJTgJj81U+8rid5F/BH2fvRqpNAqkijHZzWJzSdW4wbVC/yfP2YRKew0ewp3zxMRWtoqqsgARhUEctZTKj3PtWuzh8BZfB6fiA+xeyOMho47F08Mnx0g15jN1hR2LCha3sqlp491GOB4G74KbNMC+ttPFgcFH7XUNvw84OV9XBUu2qgFW+yOKeBs5fytCee+Op4hQu+jDinnYSIMgQ6ChMiBOv/8YLhaYcDSaAN+HftLNiVrr9A7hiYwxnrQxZG/EL/soH7NIV3O4w12vZVL1fgC/5G+jGCGYgy6g72FFlKJR1XqD0qs8N9PSKmYtfUS9Kv+H03CXSTleF58Ab2tsNZdaf+b7RedCriLTeflOUYmLf4PrxvelYl9sjaKq160VItQq9UaXCXzUdJdb71Rc2WFng/B6g9DxOzzJeVyqLdOPiCDfvJu0s4SsHLPo0ETS3AVDUm/qaEfBGF/bPp/oBT4Nu+yFwN0+ocdlCxGvN4jbiOSGU9FkyHO1+/93U2jP9cFrv4M1QbuYfsFH7tvE6DZXRT1As4GNXlgL1Twt1JclmfYluErV2yyiIxriZqsOvDU+K5U1/hWJSmk4BgrxE+boxKrZt8Fc4ecP8pXsLluFP2ngTYbdy+MPqRreeBIgi9GnZu2o3SixDd0nfENhT0pJhi2nr3yk8hVaGowKgKcw5y8xpR6sJYw5V2bCMAjtKzOaKQ4RFVBsBatlu44UiWHe0rQiBftjau0wu45mf68FbB1yF/v37b+aVKATz4VDOkvr1TtsR33p7zYUA8ffmfCyVZQtqnmYnyxfDoIQp+a+QjijwIx/gy9eq0TEJQ6Dy6QQpx/C3sgclv75VTUizDCeqasm7jzPWb78HZIjzEGtZmqnS3V3hwABTtT8PXdBqyIgjYQEhYVJOF2WwemdZnsm1UdYDJS3xJI7MIR5C2GWKpEioN3miAcny2bTCRMUZ6RSsyf5Z1zOdiUERRJo0ryPI4qoo6DMAjIJU1ndQltj0GXI3E8GDU5QnCzzT0fKklTIQMrLedanIQGNkR05vV+4kgTRrEyuOaYQ+PtrZUPrOkwjB5A1gpcMfPUY8hvWtHlpadmVoDSKFu1wuO5tzQpaUbEF2z3rQDiKx9xX9OgJvtvn3VdMl2H89sIa+r5qsnru2/ZRnSCltq46FBAOnexRzhMuwJrMI8RXGPkpABdp6OYKNzZwCcUB2pKQW9OSqlEBfjXQzTxRsTNrn5U/cr8/C+IyjRSRNKOwOWzkww+yK5Y5DsSEsz9ryJwrrvma4LO71ToZRfiAyeEVgrBlr+byInyuoJiFxpV6JU7/9/XueS+6FBtbB6m9cVqQamX10A6K/MV2uKxjMqSh11bQuw8TCY8OhbU5fwvTPlp+rUoJB8vuJVw+wEWEZGJPyPT4duBlL7UoXvEo/vgCbG6w0D+i751xgNPBi5v5gPw5fivH29qalwGsFkbKkYRJkdBVOBIWdENa5Jb8m8SHXsJ6XhiU/CZVtwvsUOOEQxERpjmKRFxg5re0VSr4tjFu/sbF8JtHoS/TZ944lcluOebXfJ6JsoG31f52uzgjhVIGMDpPutC7LGnHKL/WPG3Ppf/uRepkyFowPIZUQTcRa/CIScZ9zVymeGZhl/2xqRlzZ/M8GD1utkbwAPMWc+I33duWHBZ4Vreh1w90hrnuNvmJ0w8I2zlW2xnDx3Np7LG3udu6wEYxpNvlsUZC5nnvlEC0nsJZ44qtajfIBNS7IZmuoCzH4Hh1lrqsJYCApuLU7+ELkXJ3LoT/dfn7ciiWJPmb9c8DGPod8a3JFda24nWt4hDj1YEIbUPGYGX8UBqn7ozIYMdInTEB2lAYkLaMClgZHYR4L/Fv8KQ/E8WKtz7dAkvxZGRVg+IXHFH2g8rYVFEjR3nOeMiQ2v+JVJzc6zIlaPo9ABNXHT/chKoxRp4ZzNRCUK/Dqym434k/GNvxKtXcfIBNoGgXVzvMf5DL93ypYvW8uzJRzS2jrW25yDBEgk/m4ss1W20Vdqn/x7C1DPUzlDE/8t9I0bP/lY12+ni34mFNjo9pQlXbc0ZL5kxTMqYzd5F33t81CcTZFKRDFgXK4vBQh4kxzFtj9QJqYV25SPTR2bnNghPJ4og80c6Abdx991NVFUNW0U0I+5T9oktNmwjgowGxA5ImlOec76UQZShF2uvlVhbzp1EdgOh2h5vimzAwTPYPVn+8jEUZYGss0SywEkUHc7+crJQ3ETC+/Q9G8qc92sZ9mXASpJe92GTOhGeCvIVMCtQ1V6g/UG3yfdTzzieG+K3KtibPoKgKMZoEROLlONzq9pE4UVgNYF1wLNzr0MySfYD6bCdX4yK49uduNOZKsSlz1KH1OKZQiPda6hpTk=
`pragma protect end_data_block
`pragma protect digest_block
91b4fbaa21ed02f11cf2acfc0e4c3abfd28e49390bc87c67b10084f14df599e4
`pragma protect end_digest_block
`pragma protect end_protected
