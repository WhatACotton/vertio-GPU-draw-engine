`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
6IIjE8JUtiHj9m9KYSLirP7Vl1+59X2JhYWlC+BVdT8ykypH+Inf2XXSzcNXaaBgzcos+/9w2Ud9xClIuCJyVwwVsydgjD+pqq5QT+gyrU6EDCMwdbHfo3vMf83KpSfOsjgmclEAX2pwkeCgNSiP2sdLeU5vYRC01zvEKxFexvwh9bl/F8uc/cYBfaZYdPScjtglIQ77Mev1ntkGaYs6QKf3G4TsMzaT6tu7Ypugog99tBO8LdgxDUWIG4ob0oAEqYGytT9yWF+IuBqV5cjs4qJ+BR2p1xGyBBu/kc6wmRewR/TUE2XEIz7Bl2fw6XunQqJzFMEgx7O42M3PoZtp4wDMmVkwZhdcU9whVVwPUeF32DQEPuhYsA7620s/oS+KLAOGqejklgHV0Jxqsu4evIWYTDwvEohXze0k11it2hrYGSkJ2FjTEvfCl7eOWw8nLhL2wFxBE+dDk6qrX6TD8Ua8SO12z7AzvQTrOXHNbh7yVqVZK2Iee5vp17eeeAU4jL7/U2cHP7cv6MOOpRXvfbuVVRx0VBCc4MG8veNHQUB+TwXLd8oNrza0fFffJ5DA953bZSMUieY5he2VAjetE+D+Z7xRbMVmSXHDE98Q7eTbN18/I+cRYf0fL3Th6PmDCXeJwp8+Nj5GO2Jki+Ih7ixea10azVGG7Oikg64QJXUDa43xkI8gIwU57jTyGPItip9D4vIiATiy+Jr7+xlO3iShyac5kXUtg2GePHnU8fRYKIEwVKL940XPDxM00vX1FQC6yWuOepgmcA6QAJ4jxLR16OBtwV4IsyDqIP6zjG2AfgnUdr8fovOiOkR33QbIrQV9h+WiyrczJC9ixoXCvuYxFhPZG85r00LcpO8ZqatI4RU31re4CPBiA9lP3OS3w+mGdZtjd1+GmlTGM1llUU/yn/rllD25h+kq1cDyPL2+5CaUkteQnwa21+RAHEtH8nwN+91r+kLYscwxr4jZsBGQLUKSmQiCHvDXCPw1VF2JoidFcHPvB9mnXKwy9czv2H/DHItWECrte8Q/zdZk80JYnqlSjnbpIM1nuk2sAlInOdyiG/0Ok2CmwIn2bHnBSGvgqa20yLLTnD+phTQrIdnWN2MZ6bb0czGXRwDVbOmdA0cD4mQliYRCRc0VpGfHdWhY6aodtSemlo5qkI4OigNl1IjTmTSfFuhV4+UfObcXEKNySq0Lxb2GR0cIX+0sEfSOe6IqBBOAXSX17C+yA9rDUSsIjqYse+ZqE1PY+uM553N9/Cb8CFISWAPL79QcFlFx94wA68FXg0cVraZepIBreLDk8DrqmN8EHZjs2f+b+GJ5IErb/tYqu/znNAVR+5fqSKE54VFMOQnbkwidslHT3LyjmHjxxe3nwwIN8tgWjoJAFnJMD8pV6aUF5APk6lauIQAU4ReUgUmGAyszoDrBY3TjZ13RfdoDrifEv6QwbsxlM+gDf7Px+R4K67Ly/Sc6CfFGpmNAH3wkogd2l/RV7OjpKbUcQLEgDa87YSyWntRuK9AmWluh3sbux1EDWIrksq7C9udGYGLpvDhjY5vac56j0//vU1mh3Re+gn1R3wKk2q4rH6jMN0+A4LdMCiYLSv+j0t7dE0lVIGSzfkynJi1B7dZb00f4EqPQJHVARyUEwqu5qiQZAVHQNE31PkZqBB10aDvJ6af35VVoY9iPf4FYMmTRtxCw5V+ZjDo46Eh37HeRApVMrsslLrDtU1zJVlzzoFrhdue8U7dnyN+W9xP0/sOMOR/VJjRiEmk4SD4m5TjSB4EoCwDTXHBKSOB1sBifO6yTlcbGbTfXRN+YT3JqfCrOgXHUZZytgfwZIo1R+Ro0xwWnZkJKqkbCC5Ym9zfmMxZ/Q89Afrl2ACYabhctqwAovVY8AY6iXcz46YGjET6xAaHAt1Xu4GNzL0OnAngSLvGVFvwGwtjkOQ5vDU3TSo6c96rg9jSIY0hNS8jmdELod5p7UgPdovPyyILCL8LVj5l5e44dw32cJq5ZL5AdX8d+3B9e0Vk2ZxhAyq66HO8bG0byxQkbqtMJSOPyecv25WPyikJF10wpZbnm+QSWF7/BXBfvCMnPSPLwRVxX/6y2q+6ZuWM4H1cEJeUhBI0OacttmCwwY8e4SwKs4LgAbR0GMFNeSplwy7ThHyYNctSRgj1lbQNOqFJrf53jTguQe9VCzD7Tx8x/nWix0waFBPLXGBVf3WYjuVTUwDUKukpL/dIGqiZsGlTCTtu+TsaBPQxLdQAHBl3aAKhfDq72w8OSUcU1TYbSq5Ztv5Kksv/4rJgBaV9Dk3hLfe+psCttcKqe8LygbeBM2kXz8LAGphlJU8B4S95xxI7tdpY9F2EKIde4N0m72VeoGx89lSO6OpgKWGvPWqN52Yi6PioVWMjj0W1umJEpu0na3HXjUZ1SeI+wK2Cq+E9vrihtSWY3ExPAJbCvjrhF5LoI9CZmNnCTOagNP/N4WVq84H0gW4qG+P1u+MiGYca+bBojowFfiCxD1UafQJd4uDk8IMN2TtXkGWLO0CwOlUErR8Yv2SCNw2dwS2hGas5J7CyfoETNQ28o9ZeLzpRJvnFPzkKNEWAplJ0dqbKqsYh8lfWQ9mOdmAX03sPcYWQnGJp3qegG2h263r+z8ll5ghZa9jWE3lCTS+mlg/WYRwSyjplUjCnroPT3q7P/UHxZi+/Y8zqHpTbirns/RVw0MGc3hLGwzvL0MDETNyXXR7Z7J5wkDpPJNIRRUzFlU+nHbvKYumfCKv/dCbiSBgFqwuzmm7/7SmUm2Sgg7FC4KZxBk9B8g68ZFFtJtj4r+Yt5tGM1+sxPqM0+g8r9QjM6itreDNVlMbyUFYf+23VK4BdyV1rEVjZDq83zlKwqx8CVF4QJECSZviw/3e871HgAwbX2wedXD7scfcQKF2/LRoS+rlevsPwg7pQT7iNbNz59ppaPrkr3+/5tesiJAAtDWgGg8Qcsl0KTCol6F3n1p9Bv80bxGmhx0C+SdxkZCLFcTUJlh/iyOCLCKlWk9kF25qeEwPqtmqycU5W/DAJcbp6AE362C8RHdbcuXISD3j/DyJj21bTGVQ1DWkO/3mChWFz/LycU09Yn/M5fXvgOTpJUN1vIZ9FeuZiLoqcFwL6H6W7Ki5raB9ixKEw+AX4xCJSdRhKSPM5ZINrSRvJ2ZorqpqziEHVjSir2qC/80aQ/YuCjAwdBQeYUUH0uyaO1qgeYlWgNW8yX3Cg5rbAF/G+oPzd1JGZKguLEI0p8YWQwQFu0Zpn3RyuwJPTZAPIuhRI44KLCOLHlp3gZV/KOfX+fdvCzpZFE+KXUYV6QgECa9vXe3pWoN1WJkR3SYDecGZRfO+aqIuFIwe+fnoLKT9CezqN3EEsRS9CxqpzgrwnjihCj1mPRnkXFgr2g9DVcKT1DSXljOZle3Hp+POMvrLz06V+qHu9l9tTqWNKJbQuDBGfcVXWGqjE3O0NLyUczghSuhnFprjlemJZFa9PA2Cez35Au+gblMk2vLNDrYNfIMc3PMfMJU13BMHHpYvFKGQ7s3akpnkhi8jKLsGLM4gaF57DyqKHW3wmwp6z+aT3x76PBFjnAw/wnI0NZ6+nvHhGruK3dxs7Jw8Sgq0aLl1EmhracfdbMUiGeafBGUFEKvCP2/O8IPXDPkwbdi6OJoMibE3Mdy8ddoAXWOHKFbQkbkk6lll5WtitMFENQHJAMQcq/XpmYjIEBs3a2+xWvTWybUb1iP+suLoXTTWECOIDVvWy8kYjAXgGohd6egn96eFXwTautkemPZRyrQstbK2HUATvf4q0e7w9SUPVEjCaUaEtO9hdpz2Z0hbxxkpynGu4pBqVWW30waUsl/Ofj8NpA8TMvf430V0k8m3I5X6vXjsBWdOk/orKW1Zq2C4yR2BG3guZYlN3oM82oY0JcdDiVTYM6QTJiS9A29cgu8U/pPjIXkbSx2ucffnpqHmMDtOLCakXK9O8BqulxkDnR7+rjowOFpyE2Oqx6O4DFLF35ghEk/+fOtjIAySkqWjWlKhRXmdWQfWDUXnYs5wLhDLteoPuG4FMMYlUK6DWhemjCcdqu0hWmyT2yBmKFYqn97g0xJ31h13kwUk8OLaJt8iPbBtqellYF+ESYzjff49YZDhzp9NpoZvtXrEETX95gUpl5B3Z29weA4CJ8/jbcPChYTjIPsvCbSzY6vvtGuT7rMd4m3x0C78ReccVqk+IlsmWPkjqVTP9iojnG07+LifP6LnU+ggXdjum/+aHMoEHBuQsLAkWw+WsIAyGJB6QeBlrhdZjerZ5VkdkzFXCISMpD1xrqiC+1mfc++5QL+ekRBnEoDPefU2yN76a5CEbC/bSeoZ35q3JVd1kT++Sut1UkLttPNsWTQfj4jF4JZcRftoatiV8OyU9n5/EjnlDE+D++qGVRKrGYFoz38DKnR9rXuE+9ZX/8uDsYPIVL3p4R04mBfnR8pX2VhM6Ori/9TBPGndW35Bv+FMJ1gwF05aHb4HEynrvJcVg1oXTRy3I3k9SQIp15pbaPEJRWV/moo5vVm0YgWCYHuAAAqaGlbhk5U85xxyzyk9lKKQHq+7w1r2LWMtQpWAfh/RZup93g2r3yViBHJP4OfRPTuZd9vy5qzguZjtqtHvXjxY8dJwt+codWlq29YpXr0D7MUC5yUBApyNScfdDkav4KlOOI1++mvukdFrSyIiYdcA2oV24ErFfrXcs52s3wrrzyEW3xLdINaqEzyP+dEC3SELKEUelOLpDVhfJDhQmhYTKwOVTfvlBJwjikpXte78JAhnJzIEzyQNTSz+AwXou1BbsiVRxLuGuGX6qNka3DdBsEnI8zSGnEddvp6NaJHqE72KmUiRgex9YCIr7r/3Jpx6p4lDVQ5Se/5RNLLtkWYrqGayapS7eC79+VaYjinc9bOdvj/NCjkpY9Acgm2+5SkxyFHuhlnwdH1tPq3kY6b1mSDv3ovCMT1djeb/P7CAoSYxndquK4mf1wjpJ2Qq9EATrDtEU0cx/d+5//ZoCsLIRI2h/CqcqAMOjZvqa9hUCjUqq4g7SHbZfUFkBljsoavcDxv9sLOazJOin/dkTdnY1U6gXpebRaNPLsAwyBzVxXNypb5t+VvvjCeOiDVJOtjKY/QYVHgjb9LmyIxI43b9fIFrRkI5TooLHga0jYgxJs6Hki6pG+zfAClGB8HvQ2OvIweC49UQvO2LKe0X0UpA9Trd2/sW+g94FB7rU4z7NRydT0LnsF5H965W5jmsmZaFmxTiKh2uE7X0np0qCfCISeQiNPsq47tk6eAtntGmQ4of4IIf7KZHSYnJazbnVDwJqEl6+7lYKVBZT604DdeZB5MZp3kSvYQqdJQq/22UfR8Ruo/NFdJEefa8Br3b7huuRzWI6FvnJ/vYg6FMAXbPYqewaixxM3/7QEkPa5tZ5tV0v+Ao+17N1WyV4fci0c8dxy8ZvFdJOg22KIR+GOa2P+B4v8reZOT1EF9lYHyJJmFVERH0mzgGPk3lZMzBJBxV8G3o0Vl0cbrQfaz0V01tSUem89t1UcEBL+MEfTtne87SBmRW73+Od4jM0Xen9Apnx7djzh3Zh1caRbBPMB3PnH8RSgqxZrTaHucxzKkk7Oi/dczoKypgPAJYAaCnB7902gCmS6h7LB0yqh4Tq5GSOUQFIMdiZH4EKIshTVbVuRMKO4BuUtOL5Nxdq5+Eu6w17QThwaTfl+VhK3cDW2i8q1fyr+s2A7doqNKYAspRA465Cs9dmg1BFMorE1b9ZtaklZ7lnfA1bNSvdl+a2ipxpAGUCFyYaVQNfa9S6iLaNoHh+E3/XpnzmvfZpcnpabLA+4k+HdqWE4oFarmP7pbuVxAqdHWHUvCpQ2ArDpohEXmHlJTa3k6qFXC9dWyV3uOWZyQ18TqydxDAryCM0LkhuR8gOp2F/wiMoGdKTqya580ISY2Ieas4qbGyrdqDLGxEHaP2O7PcNV6MoEpsURF456tt3hWIBmvLxJHfCP5ePt8Wu7f++Zux/m88VtPDyeKbkdvfWYTojppkuOIfstOk3AZ5Dv3Z9fBrgy9waAv/YpGdrAywGerOKhdbtx1XfUIKKeGCpmX4ZVtAb1poFN/XriGaIotThHOskyecyJutBqQOpBtceGySxFH4C8obWgFQt3BTuC8++vk0KpnO0HG7E6CILE/GEFMY2OnTtdbSmkRP3h+0oxFo1sBBg+FluPLYwqeA9XeYDiAD0OssIwycU8vu4rBVTcVWwttJVuC6wILW0/HiUoDlizw1S41O+AI5s+qeEjs7pI1AeU9h0DqS04eFemeYDKJm95jD1m58tMRsXoZG821huzJge+SAf+Wp8JpzA/xhqMquQJ5/gZW8ocLkPU86gJ3nEcifet7xiyyc/M6tuuUkHWTMcbxmQCv9gm8bADwUy2HbcdHwYV/YdvTjf555h0Wlddy6oG+tMes615jiHRYzWc3KY3yeC2tVlyDB9ltAmYfxm/GM5lGbZ2OeQzg4hbsvgu0X8D/VU/nPgYj6Pg/PXJI9J/X41FtqL1pBn9hys+tu/bqcEXfKRdu8FzfUhq4Kb2aP99we1JMw00EYZPDw37D+ZEYViaL/XF5lDmNEX0VSzL6sX8ZvFt8BK+n8mhZrO0ucE9RYr1umkdQqo8rDfHtRM0pFqNNdWiuWCXwnTvIlAenbiQsBIKaJ8WabnftLqy5bRskAYlYbS9S7o/2rmYQrrEL8PgZXZUrIWgRz12gD4VQzsj9Wxug2IFYpR3JYUOkY1JQTdQTMBP73lBUV9i/p7H5tgBYcl6NEumGUGiB7AMnjwtDP5JxuqIx/tbs5ALv6jrjsGjvUarlJ5hCMT7tpLyl0WRZKJiQrAPZLzEaQj7GBL5FXmJh/wo8zlajYRUi4v7xxCH9e6p9AwIhRpxNpv5m2ZhmrREpoh62jQVAM/Kwo2JK3AyT+cvsnVQ8lph3bIQRgJKfcCDps0p583CpxlHW2XZjrcwji2wRuT7olK+Buk//T2AVEuftNCZOJGEVdPN5wdeqeGQ1WDVIJibITFi2/MSSmhwcHxq2jx+re3ostlXVqMhypuVyqSx7yt3jEzswmOq28FDnfMQytzjC29EQqenGI40x+FTmQq0t3/sn2WeekkqjIlWBLqpudzqtNxZOZli7EZfTZQQAr+QeW1qWEgH3c3qzXofdsXcg9wJ0puMc7f5N9J74t5GY7PhTjku05NYeDtDBwghvYLWPyfbDqC9ACxSKT1/2l7ljlLpkHZlT903Dbe6D5VygKOAwWvYqE70rVJMwtzvWrVuLzGP5l7EjhEkfmmePjF2NIGa5bLZtTDJ1HSnHoyR7eccRSpbvYulJVbvzygsuTxDhbLxtg9cdBmOhxOeTpg6natrkchg1km4xsRJB6T7ded+FvthCfI8dK+6RgwQc36L9Ny6db0sF73YsFO6/zTLhT8MXO4xifcaYFWiSxYaTRGhdMNcSHPu4/Almx9ofjCLVwoOObaxjr2WvkGoFh9anGWi96o+2zTeh0g8DCKGT6EMZ6XyUGMEnxVZNxROxl+vji1xihE+012Ifst4w1kZY/GCKOc9fsZVut0nWicFbOPdWC1p15OjmB+3XcaxJ2Kmwo22ZxM/10r1rDC0fv54+2RmhLmWQvHebUm5czjVI4K3YfnKyQNMMOe0ezd4PZlaH0F0d8WEsE4hfroLvKZgGl66cCttqsxggW6w/SmAfWJVwbgoRgEjL5uNm4NM9LaBaFn/63etdR0jSQgxwkDcG7eakq3MLiLtmPgFzbth5KEGHSWPETr+5LMCVbrECT0oHIu5IIAY535xelLm1J89iPiWxQB5fxX7Ad9Ysm2VQSR9aPVEZh2shoUcOEb5Op/tEa4bI1wSUhG90u9uuoLdROxzUjvF+IgzZhIrocng1GnxHi9bvcXgmGt1MbJLtHnMKB0dgEpFG0r73VTEn7kRPcKJQUuU+4h3LjICO9G4lV8nQ+GZ4va3/kfU8oU15SecA2v9GJWX7ouHzbvZGKxfrnZwavYjHWt4aHsZnbHlhR2MhRGj8ppA1lHDfkYkModoEZ1TO0StV+wEwzTCqsbFTaszXJi+fCXFjVz5MefujSAZjhtnlRzq+tx/m20+ak9pfcbMetsTSse1IeAesMKtCTsIT6IKiHBhhDtZM7FVSpD8esUrtyv2gVD3eo/4XXlyiWh1BzIFD3wFFPDBUPCxD42JK9tY/HUnLFdFxuNFS5V0xFngVwLanHGveNsqxBJO3jBoUmRxCjISA6fph20TKuX5xNqxjXTG4HCA29yHkvMjiCmoX/RSlKTgS+nkiSx7LBnkeL4uDqsxnoXJQmj0FG/rT0z66c0SCVUxPkSUDYhZ0I3PlOt5WhP52srxtxM/U82m8V8rW/baTVCdNxFemAgBkkuuRJGjP0Is8EY4kopN8xKmH4ctsrgWdOfCeGn06eWYKVNdxA74GY9m2nr/Bs1W7hfmEMbhb+A3Uir3Sz/6x+ixparLTFFbu8DdqGShm50CxyOBRQvEDm5U25oVOT1sHeHtVMsAmu5id71J5OGGvLqAcbRCKxCc0XE89A1B9vpIgDtqvZxUrcKdkzeHfx3v1ePkrkE8s1Pg3/SGAhu1ezkkQlYFOgG13fIvZRMYeW0VdoT4d0U4TwAmfjYgYxLwCFkZF00DoXHY2KRkc8n2w6ESWk5KptrVMQYB/1YIIJPJGLZRH7Ta1Ahc1jSKbMpgbgTUS69Y/rnOOQ6TSUNuFh3RCgcdJ7NzPaSTliNd1MXTKvaGgI3IQV2B5iEDCej93nRmpDWZYhuHGcS3wqiY4XVYss9xLuScWpAa6TsT64+0Q7EJ7+Iss/E7rf94OD7JeZWUIGEeWnDqp6PsaCjOxbl3Wk4rqQVYfCWl75CQOBarvnxChqFjFuXWPUeL7+Eo6qrI0EPl1Nj0C65OqgK10r/6yWARmdR71ZcrLQbM1I75KdcRYNxmQdSU47uLl6ZGYG0LeXXOl9yNuYB7tvifmOiPpn6rBVLXItAop7fqcusTBvigcDfMrlnxpoZE3xCH23rcGEQRMr248ZEmksQbfKoH9mNQUA7uZDOzPoXbwtQpazpUtns+Cep3+uAsdEn3cN5GHNpT4WGF87eZ2Td3YJ3GUwZ3bp19DKzkJHnUdk0c08H5eZd7I8zY/M55Du/onHfH6QRAK2E2xNHIOT3ovJeYMSSP/E+x5llHIqgtRQAv7nrp8YseoJ57JMh8M0lrWA4OXv5QnZZCQ4jrT3DZlFOmKDnxCppMnUW9HHE6hZoWgX68HSZ6YNUpWCd/Le2ZjFoIQZRe10qkK8A33kbaNV9/UlCAQjv31A83KApUVfyikWAhpg2Sm2Uzsk0cbpMlVjJAEmo24bnBaKauyfknaFGUc1GHS5oYI1miF3YUc0GDC/aUXBcudfF5cDYoy4MjC3QhbjbiYvxRZI0hmbONvPho9sc8XBhqcxehNNSnVUNBCuqrOwlYqpToN9UiUm+4Qo/bzOXFuZH2i0rgM5hUGXEtDwn04ph09ETazF2o8kLMqw3VE4UiuCWAYBHVs6qIG2EwR0gTxAG5Us4ZHDqco88OJWG4i/RlfkUVLacF9uof7GepkpZkdIeLQt/+dalROt3CEpnxceZaD4/kzvM0DsBGrWR40edRak6MlPhnH5TuvRfNDJLyFK1xhFLtf8L5kaJQGA+hc17fOTfIrdw6R5VwzhX6vlKPFRB8t22KJGcmcNm4FNTtGz8o6HeA6jE6DQ92AGAINkaMKHCkKSnjT8NAP8Y+1rIxFNFZSmkynvfaeNWhShpCRriAthLZy1vk+xHDhIThan0SuXBU1rylaGTO/QAeJ0txrOOvH+rbxbv2Y/1DnpCGiqHbIGE5cttMmKoUnsHFUR1XGeMtCVSfmg5txrvGSA9aIt4hlL0qz+pNQxt1IpzIr6bVqYO26TtLAtZQs7Qo7mfnb+h3Xwesnm4bZpBbY3UzUogP9jZVQrOs6ZcowMRgS6eNjgIcI/fMH+SJR/ZcjVqn1FHK1NuHCZRdN0vsZ3UIo/bGST6ee4YBL1NVQK77IuSmksUtVSVhYl5ERR0dTuR4wWfLGPANlbGUMOv9z1Zmj3OGzMTlJinrSLs4T78c60ieFd82UkY1wCMadX004Z8schD/NPut5tZC3IaHh/m2UbrLa6bMhtMy+UKedp3TqazQL9/SqKbaPX5Zat1AybA18CgtJajD3cMIMjfnh+sYodQ9YmEWqspVI+FBsVr0dpS7PZX/cvvyl28veejF2tw5ATs8Falkvi1Hhd+JURPiAWxMxWCIK9BpqxcrSQYm69TWhkxhwWkfi6XyeAFZMxaCl0h4V6gsW+s9i63YlzK2KPa+I+hisUMDEaVTqZi1QOGf6bB3S2jqIo6QTD0QdiFx87I1uISOLHT7Z0ddo5HzDUnYWMAfzlQfpkmdQFpCMiryayPY36PXmSFdazYLPmxeyl7jYB+hzz0bVwkaJmMUkatnKT4CfNzCzm8j56t6meUCmkP35cykrhDRsbl0VJTQjJqRpvvV4aIAtGT0wLBkMBAA/OQEJeKGBnjsSmRk1dIisp2S19ruCMK+fXnXKV5duNikWgaVd7qRrl1xOT+HkSe2egwARGjhsiQNgtXS5EqJK6jXeoeBTZpC9Ah6IxF5EUw0pDlyCIkr8UAR5YP8LQVS8B7jZ4/FgsPtXOa5DgpsvCLPYDyL4V1y/evhg+ZSJPr+EFmWnK2dmj2PLBqcmvRmaoNY2S4hLzV2pgSIQMEqWs3Ww8NtCBkUgsRs1NUjKfWgQYTdDsKT0DcbQL0iLNWHJ50lt3wKO8IcA4qKIfwxplLqSdb4FJEh0CPlRLw6gcCxQm5PN4LwggGnStLqfG3N4FgyJ7eXZHMYOiZVCpo6nmIC6vpsRRowL8JgZWvsQUYtWiIMl6WVuvztL4P8PADvcRjanm3S5SwCC2JQZADhFw/cJw96SRaMB9HkxpyQLV1aRVMlhI8Vpsubc7mPWZ0GoU/D53MMFQ8hegVJTY8/bdanpHyCvRqLZRpBSatmrJjdVu3fsLyK/BExsjgJ9ySQLszAJdsQ7axysQMUQa67ZixVnwpjiyPuy8E5ckCbLseqBnnSbX0qYtz1PwJsFa9kNzlkadbozgzPGwDf/jIkiYKa72squvdczn3XP5jab3bLi4egVk+rGRZ7C38CD2TRAEmXEjAaxKjxbdPbqCtIWhAru/pLijkCXtWIJiQVcoaFxJU4PsM6huuco/4jdjMjsqU04QtQIaR47stvI/dczS+GiulNNBUCXvac/qWSU0ZahzA10+RE88sgCn7lDXurkWfsyM+9KaXwTgfAS8SHGRcKa/0jhuG70Y9RswOl/Ll1UmCaYVqS+oS1Vji4haHlG8T9W12yzs4WqizunVD3KXXTrFPP2qz+BeY3frB7o5LHt5fV0gXPqQU4v2xsKNcXGcgTzpMioIocrOzCEFrUbSxj31EBZUt6TJXn202GzBcWFgXMv1oBHZJGVkXwsAeOmfnAxrFlK5VetbcDgbuUwYPMAY3+Ioi795poD+OiNFHq8nZdgYdJInD23LYWmMuv2vhR64uMDGx18GzKnzMrCbuUTROZNdU1ZEGpGH5INFMOeBmvFVGZo6LJSjBE/ZPWcr8LbYAr68PVy/dXoNF5NexLjHHlrBBZpeam9CoV1DU89CuEHbYiBsq8V064cfWG6Hp/t4NshlFG2c+SQUDpKXE+beuuBch66poFUdjvwCMpngbC2/9Cq+8eRcWGknPmbgobOb0iyABPWwpuZS/vSkyrvQ/0vKeZ9CGypHIScHrrgEd20bwzNim+Vi/P72BD338uQVtCymOhL7hm/9+6pCYIdYnqWmUEJ5lWGcoY3gx4DxQ7FoywXpzyOJCz53RpaSN5d7cOAFc2SKedk9zGzACGCerIDb/CgOVvnLo22mPpUFzBFSjpm7y2lcROSIYS12U98TPOJIGAoHhaxKwyISL4bQXv72mbC/f660cFAPXAsrGIkKC/yTKP1Q8tS6RODbI6BFR3CdKVpnnDxd71YIuZzLF2+tP54bezbTmyj+HU4IXtSMLqs4zqHNTDq+NTzVXclxnN1lMWklzuQZVaFg4vu93JLZZqW39gZto/tM+dNy4wEcSSJOsdkV8Ma5u+DHwgGS291bNdaHWcUFGumPlHDxNmoRyVpBSVeuqHwqgs2Lq2xrK9Dk6kvUSe1jmcsNaaSrf0F+PfHJ3qWc+SIv2z1nhgyN7+7yi86I0TWlxgEMPfoIQX0HMYZtrOgBeLDeNni9sDLbBsWIHuyRGhGZaNsdp4K+m5ta6xrr9qzoBt25bk+pBUO2CjJ2ypDSjWz4KfHe96vR61XL6o22BgIhyH8EJut+GCtpJHGAuTQ+nGPgfusWl0ledJlnG64tRtrcnD36eaEu/Ewkg81MW5h9K6cfg9UOVBT8G127y1ZWIGE2Ya0Fq82R4a2mN/HvTX3ChIPtepL6O1eBEfgOG1FpdrhR1V6c/vdpmn40yB/9Dav1gFl8thTHMJQeSy24yJN4zqnCy1nZpR29B1Y9rbaVff/2McIMarsrGf1NUfBQF1DsDvwFHdzSYn2r2J62qmHBkkTEP6Yoauhfajmd9TOwGKRfTCytOKu4IJrxNGlAkRfi1JDvjRg+nQeHjTdGcbieCh0me81NDNaJ6bR3mu3NJmE1Elu40Ol59BnKLUd9GNfyYqK+tcF26chAEhuJKw/JIXJZNJB9ZTECeQTIknrMIgCoFfKOL7apEGmnb9z3zo3dA+WLElDIRUe5pBZ8TKh4OkdV8JjMpDDyJGnfTS6bNNkfp/pHuXiWbNXYy0f3tRatq1dpgSmIXy3EEhDJcBcjo7vQeLoulyIrwpHyYpw0mcRJZePiwvHKLVWq8KL2lb8hKr74neUL5OTAIOHZ5rMa/cjQiDMMjxKJ6+xngMNNa4QFP/BenyhAK2gr98r67dIVbKBSmrPqMpoNjL3FUA3xvjtBZuMBFPwLLYuSj3nk97EAQ61+UkmrBMSQOWCwKQy7wsszdEtgkP2DQ16kCDJIpwGr4fbA8/23o+KBblskAd+FFbh+zVPt2ve4zJsEGkTwbwUSV/ySVqlEIf9z8s3HZyDVsSDSgo35JppebyGSzIPlFckn/DX6boJJpoDCQOHFJOjigMFeB9eFAHcO8ncRIXFSVpaaBpD8ouf1XYTGrsCSK6huxOTHIcfMMB8iYn3SmRCRjzS7tsBPCYKz6bn3+IFUwpvcOd9Jfbapg3VkaO33LqexnbLvfpB0dw2ow30C/eEl8NORBFYUYL4DNy72ZJPLHWFegUw4366xdvtGj6e5rKXySA2TLhAFP5pswG9C8WYNK/Bso0jTx1rUCuCdYh+fFshZExWoRAO4lCbgcd5NgfvB4A3qrQi5DisrLOETNG3q6c3MY+t+jA148FzRC6IAdsPKxA9jxLwIav6USG10o7xsAjYJuUXIgAQnY6ak1dUSJiogecdnjke0y/5sFbQC76n8GAR1Bo3TFPEVTKgHdft9uqXCX8fq2MpyoVvfsq/8NtfGf6xyaR8aRKMXPZXUE97cdauJF555eXJGw/fYdW4oXx1OA/5jfonZ5dAxB+xw/8inPUqG2vvj+AXCIyOFp8xnPkaUD2ue5gKASFSo5Vaz4+hIlDRdJQuQ8DJw3Y5oQdl12wjHNOdSh88n85JU+bUeiE4rgvyczKlulbUfHIbQhihgH5+CkS88V5lpk5LW6BWOuul2VoLh3f4MAluVRAIU6Gh2wLzEZsHoO+fcXK7JaUjfwaicili+e2kij4jfxis5JZqVb8R0GLlBVOXZOHqJdsQAbrMnVNQevpr7agSHTmerPAK8kSttaN67bUyCoa97aVyQAVY4xM51TELtuKL03qJCiVqI3R2EUzu9lpXU1aLSKrwXAawmlUkiOc58onKFMvYRxuDRiccKAq/A4FAQ843EXaGTqNb+7pd+0vHQEEtJEKy7TPkeMNB1I9AJsVIPYdFJKOB6ukY+lYR0E6ZJX42Tg8kyalJPLOogzufqmkey3KOZVmIGI4KNtb82jNwnr3wzCKNVq0d9znJi4sDeqMQWG1cQKjLe4p7UjIfuiGV3tJynRbEKtVwQbJF95xOvuil0BXWMXwx45lNaiw7mbJF8wgUVOC+qdm4kecQ0R9njPWw4mR/EkbyVAi12WDZZltJhK6Uq/7Sg+O5qPVqmIUffM9H05ODE0kIjAB3iAGII3/mLH22qCeXBm9FQlIRm1Yx6CNl1Fqm54WCn4yn+8Ff/PBeIK/U+pQhZt7EoQn5SuoePAyYWUkhFV07yYvXVuWt+O97eUyeTpo3NUx0OCdG77KqNVan9IoFscmyqK3TL+NdfXpAxg+k6u9I6vLKDGMUoA/V0GZROhuR6Mu2Jds/KYcx8W3uFLCrOZa6p+JSHHwAi2swrV39jZepYPWK3xinNqeKMvk9KGQ7NQdkWoKAekU7xbls/Xal3CJU91i/0OvljRg762j0F3c7V1dOhcmOamMFxqiQEJGu2tTGPMZ8VTjHi7mtCVf2HYIHId3t+CvexZpISsDX5aijZ3W6pW1Gt9U7a2bYLeBe8a+Q13CSV894EObA/PFTdJeCqoKyqYcwWnpbbVuFjRLBUo+mmodZnwM6XvUHO0EVwTm7yGTQJzRNckoUUfGNmxHtHzU3Ha3XPY+8TXDwMC2QuvnlvL/BS5NPvohW6piaC8rtZTbbdLWH2WGZI7WwDrW1VPfwfEiBfv/Pjk4SsTmh5uza4VgXPnE3gGU7HXKk0vs2VOgvzfVR34vG0U8KDu44DoF+hqJRgv1m5SSXhLwSpdvhop7s6qygPqJRc6Ik/7f2Q7QecppJF7OPJnjcDSrhNwlfhVddM342j/v4yGmOrwr7CmQPT8jY4+tjxwjb8LJi2c7lvw90Cz1t6ln/5N0GnSjTR4NBLgkqadGpNOTid7EpBj0cgQYXI1PPENDssDlMJUPhU3IJnagcYUWRULToexKfeUNcJT6x7srxK48Ar5y2GCdgCJtf70QIO6Vx3QIIIvbCziSBRHkzhUEFCPSbfs96hK1D4IHAQUqCyhwmc5LojV2xDztR4piD+pFR7giUtQhryXVmSm0n6PFM3IXPrNXy2amm7drRY6LkwkHo1utkoi/1XBdYFvEmXU5p6Ky/zmNmGidpayU6PrfZI/KC5o0JYw1JvuAl7Cz8/ChfOrbUXI6X6v9LFqdZ2t1a493T97xXm+2tQYAXOMbwrJDbMVmg1kXZB0P7fo9WMc3mWwcmN+862ztRtXBHb39BEfBZZCefnAjcTMjef84Go6o8SZ290g6d75Ao1TXcbwLjx0pTcPp7EBejdT5tsxVklpyVPxUkUKg/LDh+HoviqHhYOKGaEMEOeNfTLhZHLW0WIzXI6C0om777wrWnPN3Gfk33vBh5J52WOO84VaDWmfv1L2f7cxgf1t3bTbUjuCzb84Qpsjd/BE+G/lr1HQFPmHWjlRpJxgQ1pRUCdHiSVX7qDdt4zvPFCTkgg92qeVBvmY2EEnSeO3qDFXw15Z3YJnCHSoQJ8owa6XaA2cX9ZgA3MHnG5/vc0fhHf02rOzDlJc7nV94c6DlSjppPE8uUx8ck8wkVF/Ev78jLzat28uh9g32i7/pyLEPrNKcOle0SuDEt2lO/dqK4XsgsAt8W4ZgSG3nz0JsVJqW0WIfukUKlMfey1fVa09OUzGTZIrgiRXlQqWwkjC+pgxLdst05OmbQucHyq2cVfKl2tK6/WgIN7vPo0QSYogsfmDG2TZa2WWw2L0tzLGXoaNWuOx3cAdmV0Xmi8BWrCk+rV2a6+k2ECdUE/eCNRq7xyLQaXSDEOoVmcCxBbICxMqWgbVyXWcpC7qlFE6cBUGiBGYqrJs5l8o1LhTBvj4=
`pragma protect end_data_block
`pragma protect digest_block
4cb08317897fdc35eb72a0fbd2993c9c753bf4f15c73348dd35ef206e9eabeb6
`pragma protect end_digest_block
`pragma protect end_protected
