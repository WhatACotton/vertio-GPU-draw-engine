`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
wFzxnnY+zpJUH9SPojvYOi1qbi/3frB3DxO2KoowpbDBkWdkUxqsBmqXU6nKODsy9X84uW2uVlwJu3YZBBP6UfD3g1z1HwoRIL34EFJISt6VVUxk9YSWIJzJwRLDS86wrUf7WROHquNzVw9SIvGzB1dXspOoBofXWD/H9YtRICvaIrZeK/PHngfOJ1JGdRv5ep6/g1kU5kMbiUZ6jSPAbulCN/4dc1v2QHDykpWzbHLYrdhQAys57DR7rc5BkKlEdU8UYOfktKJ6glUbG03NNKeQCn5BnOtuJaYEEFqKbsxURNvLO8kPAF5LwFHBOaRXYxA8pM/1EBPIpcD0ghxwFvzc8zN8aVtM4UbMY4P6qr3mdvthHQQyI3cmt4pSYaDsV9d92R9ec8i7IrZhNGhBuj3mf/xt/F7lmNZBWfoTIentMQFZQva/7oolWBexqZAUqrBbejzz2S08PUo68B+h0qzi2/InXuVKWo9M+n6RuRqO+KH/nDf4eUdCjdjDSUC9q62QlEN0tnOw5h6Xo2zF6wgxW2O2BlXCgzzJ3Gz/Ndw540keKHrKY1xiewZWSZuNQ4jtV4eV2zkUjbjv+tJ7yBpjcKbdSBWcOiR4zMRnz6WqOADCMNKkakviacatjTIq3mNfrDUqmWmklrws3P+hPC6n/eFhJK64HI3fgXmpGqD93ZwaNyE4QECrwRnDfvBzRDYpsmCtdJ/qHH9YKkcz9hwI0XAuiH+3Z9iOWvOnLNe3Xs/dNsIEtDiTjOmhYHHJkVXge4DsTqHV3dfk4PsAbrrzfUgOeRHYlqpaTpNQIg1IUt+j5iAnqLRyAFIK5qz+zQefELxCin6EwEddlOLuA9zYkyC4OegmLsy3SDW+BtAQJGvHhkx2M/ChlOOvbssp8C4c7RQcMr958457uIeloKJMydJ322lsCi3Y5NlIFvFWcJUr3v9hl1zAQtCnHbxgw11Pg+SA+BEGzYBQgbxpBXwZuLKlXhPoB3EeFGAdLqrauIalIdlDi4frVtOip5Cn6e8PbPy2tk233osHfLrVVfFSB/ebqEPytkfsP8goWJQ5TaEpHXuLY9dv9qBr25yr9EbzzhbIg8tDw825VJWfLKCsAiJQWtMGM3DrKiC2+473Yw1wyaWUGwM4ptehmewXoRa6xdgLtowv07+XKngNjATZb6Lx9EtxtPMisNpzkhZxlfDiSv5Jn6kZ6ZSkq85tPBizSlB4z2sTmRMqczakl3z1e13vNds4Tjzmi42UyJA5l0v18Eedg/X4SpbhU1aEOJMl0S+kX3EIIviyuoPuzwrSXtYr2bMbOZ/CXmWkmyjrBtRAuMtHmD19ohvZxn4jC9cC4+OLQ4tNg/6yWcLYnuq0TdA60e6fokGGw1L4JEn1pQreLKUzPmkmbZJ51Gq6FFdEZyYLN/ZZUKQgym65O1gX8QiyGAQld4U72g2pBQVwj2qzpxH4AvHtGmKM7qBTALa95q5NMtwuviL0XUVot90QUfLctq43QC12jyX8dUvC752ZcxJ0PFE1ROdwj4ci5csHdGB3xO13nu372awNehe3jOkznkmGCjLecyx3dhtKzG6LYYSu9F+2mMchH06HqnsbYcSrtlKwnAwNCsaCA/UVkhUW8lapQyrl+d720X+M+vHE+kA0+LGjruVpYXm6bxb6wFENDpn7NWcdEIYHaapKosBGKOJwQRZG1Q6vCto8aCR53BO2CaOPsazjrsHNCqLcbi6rsh9OXtP0+64fA/1r/rldT4ly4tOaKTVibiqMtNRHpIYoGGo2ixqgSpuB+76YgyW7RMBb3soqCDzoJXNwfVwhs7bINRmoOMwmfVSdhg01DGfChrm9rtI+l1fjsdrSwDor1GCLp82GgGvTyCWx5sY4L9cnT8XRX3SjyJezsTz1s5BJUhNYw7wg2/xpMGAXCE3W9BHgmbGRBGNfNHGGV0INZHFCt9vfSAYQ8EK/shzj31cKObGUS1YpzK+Z3CPbfneM4u3Jp57h++KJkswAzyYnVcmi/Ohs+uMTJGNzAQK2hC3t4utTiCPIcv5lnSrqV073j0tfFVLpQuzHu2nQHY+jlatmgCB2xeELcxyOqIW7bCN3kbfAWlGs661wRqH3DK//2crfbQLrnnKiRe1XVIvKaw8NsppajHXAiQbkM1vJcvH39GV2huvsXpgXfw6Vr+wweuT1QKehD30Oei7mdZHj43AqaVCQtbouqzIkzkWkez8C8cnVreqmtA5Unssw2gY2WEQRTV1pP/OEROS+yvRxtBAwZz3gsPcnZtRwySyFZxJ/HjCuN2ylgH8N25mKqTkku5kqLoy4FdwGi3eu41jNhY42kgvYodVN+foKVOxGBDuJnddzF3tDzTl32ORLSupGdT77eXBXRik+zC0wlvfDdnsoJcBrrN6NhACVF8REGzeIbN/WbjUJbihM2emYHFVFyHHfQTPFyxBOL573p+7UI6ZETUXVahR67zRkcFuFgGOow8kqSU5CwVAoDBGZeW3EJHHQ3gvVmmSPQoAyGdMt9uxsXhGGjF+IsZTvh18oZREj+hG5DBM2rguCdzfdVogi0JZqIoDwvfgwO6jRDG+bfiD3xdBhNk7rWhqgmZqcW0VIBi/dMafuyyftr711OSHxX6CsLqHvjdiu3/+QegeB5Xg1lXD6MpCI/G2fK+Ta3ku71fNnn8qFp2D9xcnIclHCafBAC0xcHjGpeePjZ81DNSainJqL+gAN4CUCDojnXO8lPAovaUi7jnWkGMjkph9u1o+1sZYzf1SlEJezbeAZ7cSCpzLfvnxRdnMZON8YsYOhw+CJoqMobYuvIEMteDTS2wrSM9BV2NlkWHyznrOkC3YmYeeOTE99T69gDRWzwOYUXKMonRHfJAHEEolzY2PJ+Bl92yC74pDZ0T9Am9X+Cab7CHwOTXE9yU97CzO4YpoGIahH36tjURk7A7OFWGHq9HICHl3ddrvBbLKzdtRnWIQSaFtrM2idONdYxS8u8UzP/9w52X7kbEWnRhFbwtF8rDlvKX3ZNAKTV4FO0z07yvYvr+nR1APbyl77C/ylT2GAOrVQpb55dHJPe6d9kd0y3kXbJWjOcUG2CXfCftonrQzSj0lMsJUclxMJGuEAsebOl6JHLBXKAWMaGsz2OxSh/DkE0QxnO9YseSUDzxU+BypZsiL+Y48hpegs9IQJ++aBwukZP3ruWA9PNAXPpM6FfPHlh7TIZcibOLYQVxIEY/om9IHl7Z/jY6rdzJDPllqiciS5YUjGfIP4CcWuqtpkhUv4pLjQuPOg6zGngKvg9PacAgltN7e3TK7sC3Vh4LlV5PtcLgiDlqVXxNeBBnn7QWCFka8X30iRkAmyT5Lp7TrSvrpFClmmd4vW7AZ1R2uJQVxB+yP/QDv3ltFIXzCp/wZJRq3G1lxZ5EGstt3vJ66zgdWbR7Br9a2NkJeRbsrkSRyTvRoItzcnqA4NrREps1g0WFt/xkkY6ZtMaQrAxRkGVt+tY6f4ajZ3n3TrV0wRR5aaimah4JUttQc5q1ZBAcy+hzPmg5psfenpCRhMIlb8+ASvuOEo72vFL3cClexQvuE/nZQy646sx3EetEJP0zIsf2NFMFNTtFlG2AlIy3HWfRd5BhCHEqR6lqEqMdPv/unbVpv9XetIk0AlohpNb9ZKr8j4SZivM8Or6VzUWXedphasDjs4G7gkplwUOJc0FQK1KY+MZptOxsLTmh9ReonX6uue+EP81eFLrZLkknbG3ENaRsXLyw8IQVNSFfWCQRIqIfHTdFnuyjRavgs3vwlk0EqLBqfxEPnwRjqVlSegUHOOsb4OGNys8NhAHRzqYqBAJvFErstHJU1JSgYJ01+tJFggp/n5nFQPYztjIKFf4hn+2+AZOZdRQ1IX99k7e7AeB60UZfzrfzNPhJbQDZ+5J+WXDkzeQxy6GxV/kWdg0ix7JkdVEn3mQ3xoC4G96Otcm4uig8ue0ZND3Vp/ik7riVyYgmb2XZzJUja78Bcfzsk6YZHyt4+kcp/tFP6y4ez1gqmFd3WCtZZIKoXE0yGFYl+bzR4bjlWZqIQloKqaaZeBPJRsbcwHQnEiVzDXOywAuWo7PvfAO3i/TaV222yyDMHL0sTJL9J5dSVN/9Cqbk94zfoIjGqC7X9DjzEUqPDOywF22XUKKZFItKEueWOU3p7l6+v8DyWyb/2q72adeuXrLL+gvq9nc67iftpUxAAdN7fvtLoHhmW/HZs6V0zGURxUoIje9YPmYf4MzMi0QaYkRHSRDMUcB9W6nrVpTI10YJw+GNvjmmrFJuiVZs17NzOPSvRjWf2w5BWYscs+ICy3pfQfPfy79yYFim5SUdki+0zuwYfyt33SWdMdabKL/HUokwUbWecmME3tiyw7vrhQ8sra92/Lyc8zlVAijxyW4jWRqqXXefsdtfRqvtlJ4zuMr+82anzlll+jX5VItGy8RdWmL1bdoAkodRxKZxYOt3Ym/1MQPzXyw1C2zl0qr845t9VvOaCcR1IRkBUPJVdxVuoUCZDEXTr9I1MJJcEuxx2qkWMCqpVbg6Pvnd2Q4AvgJ5SRDcYd+P+snG52UPHye3SQJqq5S6ae8X6qT8nn1xyQ+sskrGLOEDXi4LywgeTbH8GO16bGbzQmMFoWkM+PTvTvVleyG+0RZlUUFmr3sMqisLlF9AKuYCdOMgN3htyKQh0GqrZryuj91LjLHBr9Ns/3jiJFojC9pQN8r0CLR5UmnTyQzTSOtv+Xk/StAHdppwSaazq1/j2U79H6dVKkrdD7Y5hpu7R6mWjgj+euARuPVOIZLVrA7rnBbaYNd/UjwKqXdcjx6rOarCtpkHiamU0/6ILIPBj207VO0VZJXZ8kwnCsmb3nREf8k1fPR9jr9+jVQCkSfY76gjjyQ3YQBWN4iuH1s3pmcHN310K1UpOeuCHAk0Q20op5nIhHRIFMmkDvYfwCmG18IQHPx7NEnwVLwMiCRcdjJIpeewiv0zH/nI3hY9jv4fssmmPFjRWolxUMZFZmtDClWfs8UdR4vWKozO5Xg3LmnMTp74L96/FUf5mIzPohxrLdV+ZwCb0y21qJ8D+z508BZyUn3iumdBMXmQGxCcTk6izpDdZJmXi4/hNVy7ZO57FNyXMoD+Xf2VxwP1P53subUYIpiGTqPrCg1hSncIywJaYQ6aHY2K/dK94jw3yuH72LzZeQcbM/6sCP8MQFaieiL9mnCmJzyo2F2cFWEvOEp9cZh16wNwHh/j3dK+OpHSMNiNGFlU5JssaZBY2HPz+bcPZQ0Z8d1N8zycyXPkgLSeCRD1j4IElx0eVlcWhrZkkmbxHQHNLBYJJH63IAC6/KuLc0i0/IZeDFFzkXh83FdoN9OyxuwIlFdm3JNa4csZkYSGmAk4vqJCt1vEq+KQUTx7r5ag2ur9dwZLhray7T2z1Nf1VNlCLb/EvZVAigCLeyhGwDBjLCdwtC3zUX4bf/dHGuI4orHpUffjzQF2zPYHRviMjezmoJjRtck8TVeefNCzcpplW1IqQhRRZVuIvCCEriOioaXalUmv5mIoVAUvGU+N8Xp8mbl6w2hn2AlkY4Tohes5Z2PhPLDNon/HzAQQW7MlouwgiD5+/4Ty9fnulxm6fJnhJ01Qb4guBFc8kbKZZl8E9V9ZXLGmiL8KWslQakGArmJJa/F3ZuoGFOMZMxjNdfsodmZ6dM4ALtQ7Kqc863up14xqQRsQS2HDBxZ5eTsXvXFv7KuEaxMXa/aKP6Jf7Jx5Qgn/6AAEApii2Uh022TWNoXLo/ygdG3GKBHAvatuim7dTlkfPAmqmtYzYAV1bvwJLx5pFSRfWc/XBxCEpN6meo7mf6u6yGpsDkoWYATGPud5P5F7/GrtMD+fdTbOocw9C50axEWLMFj5QWHikw9WZA1sk1RD9M7XYQ06wQIVJOV5BqPgyeTEPHF4gFNS64VAnf4JPQxVz8vhLu6csbxf/cL672oPUVNAjyXrqYzsmCUdpmO71jhVQ4TY+W1N5ybw+F6QiiLv6abA616jRU5cFo2Gf6eQFdxIjYRPTM9WgT0/s8wawXqJGs3hDeVidUQVBdT5Rw/y0CUU0t3BFfu5D/d7hEUCZe/S2gK3cIdFzSUuR367NR41eNpeW/CThcSkcg+ztx8+oRxNIHMzFBWZjJZYcTnqV10AQQYkN9JNSa7kFImGsGlB+UW/4D+RAIeS1MoP+WmS07AitimkvDwOSzUQxHdYOU9WXP/jsKOzWca0UM+40SrhUncv0nMy+fwYerr+JtL3PY5+xqlIGumWkLWfgx1zXeK0ILZfqAc2oHK7DxxCVv4qAoOGndhMWUMp6ge9nkeEdZ05FJa7Z1BFizJoDVAp+UK6ZTal1sdPV9GMLj0xaO2O7ZGl9YESJ+UzGG9d35PgdUEENpriMP+Vq7/RtlpNklRHdHXm/LTmRCKlbeOrO5PZj3+Y6mbNCPWOf3/SdAo1ieoEDeP66smuSf1P64ypfmq5OuuH9kGKSmm/BKyIX4Gn618hhaPTofXyWMQiVCIk6qB/I3JrBnJt0pEFS+Eu3VXnL0S6EIqHVnaQMrsbK4TUM61CnXSRzEg5TPl1VGw+eUXxw5Xgx3PQW+znk26ht5WOciiCoZJanXXM4xtVRj4o7Rgg3MnYxZYpeMeomxQC11IOyOt8TJVIQ2bZXdB4eylAcdk4zDjmQmmGTHf47U3BwoSTF4U+HWUE8e3J2hGqqbz/FsGtxXz0ksKIebpu3y7j0AHkK0NMwZWWq4SNx2DrpUyoY98ZLDAnGg7H7q+4UPbQnBNLIFNvv9CQPl/4LR1QVa6AR4+yO6jevymlZJRWUjgxv3B3EPDkLmqNxB6jREUjc+9kNa3Bl0VuWJetL1aH8ntrZ4uHNwOoEhDTYtFOkrgSI5qlVZG30J1d5wyHjPKd1Uz5O2iyfQXcie58tbBdI/EmsyGfllWftqRiXWugIAW3ihJH9nmOGaMxO222rbnBgc+jnFFAtffvTcWqlI6XmxyAcXBtUjX5IBN/qKE1z1DRGRGBcbxPMJk+Bz6vJ96kM1AWEHUrpeg8pMY0CzOQmbA5gqrhQD6QllohFrDiUUmLZXrOV82v8agH9ee+U9fxA87PcL8HgyWkjbyFLxhFrJ8Ssc9Tv1OF5mVOqpVayqJTPJcZhZIYsYNOBE/QNgixKHRWespvcHLpszBT+VafiSRbRj6++6IlVj1ng/7e+I/lZaBWX33ie/lDiYh56Hcer3ENoopbycEP/i8CgvOjywzn+vAjVToK4rtp9vm1SLloImBUK+dkxA/dMzxxZilJ0SJIerfznztz2kgmZCFCh1jM4i0XTCXzS/qXf6Ps+XLCvC3pPsAbwretwedseJlsvYdPRBMUmHEKRmuMI0V9qu/mK9pqV/8cVvSIP0JLmiDTf/TUZQHg+A4o/yEXXKNcpeQ2DrUOeZQjR/8a9DajWbfG+5WjHrR6R5fPLc11g+PfVP4ugqsp8SaY82DxwaoAUJqxABsClMntfhuZ4sMeFVIZC+lPqcYneXbB3vNPeJTz3VJsK9XPbf6CvVCed3TTOzrZTgnzU7Za58E9EZ4Jdj6YRGT+x5KWpv5oBQay7oUIR5mIap23+PjPPe/QnaKLEBGbWVSt3OZ71VUMCetz2dyVrc2Nhv5E8zkHzihPUzBjN5W5upU3paQoUNLX6HR6ypTXsKwnDCmv0uGg1ZyfDIVkC/KpanxGBSkTr91ssFLeW7/hBdI2DnwBbb3CkNUhYOOm3EifQ7VtR+YnBEh0drc80JM+QRdwnejbNPumpUMI6WC+ayaLcdr1agykjBBAhVQjCwuEHQM/1oJBLftFKsNHbKifaAQ1g/v3BYmO/ww8fxAgJeRCs7b2N3ldfrLz4DqHJ+Pke6OwpnLyN0vqyVZFT1ej3koKSRaDusgXAith2RoCdYWc8o5Wz8Eq84DX82vfrbxZhKoWr06rxtiMzVqt11ol7ZpdhZcaR6l4e7qKQjlJQ8+DplGz9a8sf+zkqp0oQGJmHNDFSXibiSe8DSq+bRhdNiT+IlWBHt+GpI/yX7jDXaxk+vjLfEUyGqrbHnKhCUuQwwKn+25HJtMU4grYKAc2j1/rg1k0ka/7Y9nniiCeIEeNfkvopOi/H9afIgK0IIbLjquiec1+MdqburUz4YFqA6rvQsEaTujlxe9IO81ES1OdTZMmUJVx/VMIXVzADFbACUkqAQV3kx4sThEJ1p7BasZgFLUd0asuUEVmW+2aMve4mvtJ/xxGVanwaQDqM8TIENrLNukGQZx1tgpEoGubUHzh6MDU4XSBoGCN8JmFra1edeLztOnZ06/hD2quZCLFWu4u/zCGHhyMdLmPjJuTnPyNiW7UgQskbp4s1yPZ0Gw/hesHY/X0HjKXCSOF4aJivgwhswEG6lhtJ1bEVgh2qHdehLUNO/FaQhi2Jq3n6NpZwlSfVTSxhx0FVCqR0nh142ExyZu29X+/NySvdjcqeaDuVb3jtJyzCz3dF2yapvuA043/Eop0mhl9u9hb04aDBdxaAm0/cF184FuqxT71zZEJrAFyhdyCQYl4O/S5dtk7BTpRWtGUxxrnpNGHYXVVklBRLUTneKLAIgpNkMYPV0G5RJNQxCaKIAg4fZ2QH43Ic6ZZ6TK6KTctAHFEdG/W9g5FjdKWNp0JO5JzYtj63E01+ACQoUiosWsIXFVa4pr8Ok++6coG/Sb3HMSjwlnw2dvFt9RiMsQa9teFxY77CRlNT02cWxD/Oy8gzxumwxJtcZ54ML/ZqkLVgHAYFkobLBPQ67I3gwIA0rez8mqdWYbeLzBg+jKsBAMnBGw1Mz5Lbaw5wvKV8KmfcqYuxGQotqvOIvUcpc4mGUaF5OLE5Tu3ryQraFwShL4VoPVWF+NbdjumveuUCGJwbgRWzeY2o2AMOa3VC61vUt9DQb9Knx1KEOJn18bEvYojwTc20P9drZAXuQwbRXXyHZo8dlL9xdi64Qi7SmGPPKTMc+EjoXXNC9bzrl2+CULruG+PmnDYzRBdaBYNzq34dV+qxMcR+wMP35eLTeWAoWMdC2yXObYep/sqtUu8TWzEMB+ASw6HPKXKQ+RX9EHfPvIKZtpvZv7ZQ5pSlYiUpAO5b02LZXmu4pDXF/P5z6nYoWQFMT9xcwvpWoNFI64ktkvfr9hLMkG0bXU857GqLB42bzDl9TAHtE5UAAdHjJrm/vTFKN6JseHyoyvB0H0+T8dJ2Z/TdQ8S/j07qmrlmQ28aKk637AFQ6q2QR9eluaKK/eLKW+hY1I9lqpHA7P6sK/MZPpj6n0EiNmx/alLpm6enDw3rAcJtnutkHv1TfQRxwaSpqKFP1IDsswj5c8q4o1gHF3QiLdPICxTXw1Ao4S97m9MRWLUTVf6qs5agp/A3nM3pPLrAupIBLQehPUwKn2lyeXeCqDY1KUZk4ZVsr+kl9VHjJoukaOhPdVxxVDtoQ9t/xMNm6fMfONOgrro1lpWhqN9W23cT5k1fxvSEnTckbmnUfg2crXtKNEAF+nsY+6pUA9yvgTKqW8nrjbqZEPBQRdpZI8omVxeL/nzUr4pZ9lwPUy4UDN0Xa02wUVwppbvB8C3rNGArrNFgxVgTU8ogbQlzpgdfI9Vk5OXll8l31T0558A+S2s9aX31bzn0+zQ7/hnaMESN9yMhV9D/KiProzbgNjTL9v7rC7tWfKeCBmujEZJroP1qeQLFmW3C8n2SqtfuOto1V8k5wVuyGCGGjYsG9OCFVFphJSG1hU6zFHwoMdNJq46TpsxqNm12eO27a2nupdCGFj+mwIIx0NuhqOTbgZ7B5Ze1v7Z04bW9EOZePIB7PcJMg3E2Q98/RBxOVj9/Q4hwXfbNNnfqt8qZfQe3BCIBUZ0g9g6sJ7fxgHO1D2+ivQiQ+bhRF7QM6a9qWrnb80a9Gd01lJ+0E6OOJXerMFBuexVXXK8zj5uIMwhZAMJbyKHWPHBuJn7nYf2N1eDWQYTvFBZHEaUFXFBnHWQsWOgpfekn2O+mTJ7KDUPSU2neVdGUYhwrDXq5IYM07Nr1dJMBFT/uiHw0v2RfV5VhWajluBlky7Nx61yjPXuGKy3Jcc3sEWGvWbhQ4YLi4a/S5awJ27jxC+lDnBI1ntyc7aqPHjw4jNtQsT0EsP0bAMFft40EM5QRv/zRkOjzbV2UQCDnW9NYujGRN2sSrl5W4gd79YYm4eV/9KtdM5ZCZF/KXmda6nMpTCEguAw70+0u49aQPsgRyYYp1A4F7S5b/+Nwg4JY0W09oI6Qagz5Lk04qLsPB4tJKa9OMHSArlXhGpKuvUkFT8bSTGQAbYRyenfsPU1hLYa3VmcbwekzcUoMTbxi44eBocB8v62au0KGLH26iWpufXxP8MLrK0y+vhDY5ivyZFT76Y8fUcJOIeIHlC1EDc7bsVRP73O+8fokdS5M79/cltziVaFWPGMTAWjUdEFXJoyMVF5nA0F4MRNFJAP5+bsL2CJ1pwpLWPieUiervVY2Cz4Qu3cMMqngkBYgrwE8B0Tg7vLb2+owI3p4b2IzFSLctYGFF7Fn18B2BOeq/8WbB68vMKKJNUE/bzU+pMAT3yElm27+SoMz4j+z6a8PFx1IgZTzvMSpZC/f88r6PNSg/UPagsobwR0NJgEegzcv+R2b4H54Ozb9DVbEUzwZrdzNcJjxSDeVt9/lduU0oBrBD2Yayd0wsjvUIwZoEVFTEKQb8uPutSDxxOaPYPHWvOEsjkshloz0UvmZ4vSmZgPmN9ft74DEYHvCgKLsKidhJeJcZ/40NpS6OJgetJv06RSNa47wd9nclVH0Sp8Ji8riWkhRofaBz2FfglU6U1gXnz+rwZBQZFUMLIs93HqBrUzI2WqLO77AdPIpjV5KXJnHxklbR/ow75PwEMEzWxKmaz6/sF40dRGAjC/jjtwWZe90GhxXX5jQocf5z8cuksEJepHhHQKDCoqYeYWI4FHeFPZpZ+hP+SXXakc/kAo4EMIPqEPz+e8io9amfzyFR54vzd/TAmEHje1MT85sx+cFD/aMZQx2Y30+GCIehSfg856cyWeOyGEdV9inP5GgDCYPIjcuov27WvHl44Ew53sEipe4yf7DxREhof6lFDEVi3gcBanZL6XMImu1lFe5+gGtI6O1HgV/0fqLJL35PUbWQV0YGYAr61EVau7n8PPHEFF614pULz1rO3U0J6qVQ4MBchmA5TGsncuWdrY5fZcBD/5+iPUMyLDmC3yvvycvKjD67n/YO09L2Y4cx4JPTzHOh7X1i/w9H09iERQqETH24/HgaTQOud8boPc9olwFO8Gs8Lh58pK2PbKY0pb214XXJI4M54vzkWcwZsQnUvDVorF109kfWH8ZSl0rMwrhDczxumk42Kvf5oaEnvaW6RdWGGVvoVONkU8rWcPmOlQqS1jv35Fma8u3PAa7S+xcSyhr83srktl/MAcrooTkXvJhn8jc8iCDy5PjarCfg1VePA1cMXcKsKQCeQPiJQswV9nd7d3/lShZPca+wCyYRpNSZr4rPAZ72coZ6+jcCZ8FK6c0d0kyMeEa4ebEKDa8/1xAcU2bZWtfoRSpvotwrO7z4LmwgtOGBxFAh/nZRDX4F3+HObKF6ATARhSJfHJAwU35Xfx7crG74dBz7DjgNHN3Zz9E1wqLG+UkWxz69Xzt1yxDAX+f28IONpQ/uL3FzBK3WjX5nkMEz/ZUAKT3L+Zzvui+OwLd8AHtjGESFO2O8IofVu1zJFdoG+gkaAOK2UpQD/Ga3ZNHjiGjTkQGEoNhsN93XS4cbF5Pe5LYBFHIiXRkGlW1BFqdvizwEDBJE9YtrBAKR9BrxWJ2ceITWchSiKg41B50jIimueL/bXUo95uvKMM3wJr3Q6+vri8oGtaJ7Ucn5LH1tgSkevl11CfcEXO5+aw9Z6W8lHZSxbMRTliLT+BGzWV8OIpvmwlucXvkdNBWJ49IU/QnJ5U3jIeFt610DoAttWdyVjEjO3A48dBKfVutHH8oouk3DlmfSRGqzycf0ve/+tkqrA0U/G0/Cda9GxpkzLH4X/gKcAB/9UBWHko5o3urYjA2hZRIGQxnhC5kUNkOw4KvFpJqGQlLBiIi0AMdKTTDxCD3iJ8so5Ca6KkmP4j34UyP0AhzcmmFcaAmxVa1THwWd928kgrPutzP86K26kuflwThzb4MKSSTAo3YlLBKlacUB7t4gdkOmAKyeW4bZC3sz1o/piDYtqQ683iDBAOfYHTJoXt+rlKU8c3t2waqy75NwpqqvRis4ZaY29/PoGFAEgNvEXqKbU0vracci5Mv66FFrvgAxWYnztmPDf3S9v7WrA1Upd8kdWNkZF0c/5l/OXnl/LiDoHf2CF6tMr0RJRQA2RbyIpKSFoNmDX6yYBu8/q9e6NTTF8wyZQvlWyTv9gfyaP6qmdpI0uljx8N/DLZ9aveXBLjb2KEKaJ4htFxz7wOvgin86rRqzIi/koOivwdylJFilrUKlzZT3Sg0Iqetz4L22sjFm9FU4aE2iPEjXQBUkh2oNmX7p+GBzBCPoZVJqfegG6X1k3Ii+HnG9HFMjt8xmtosP3BVlmNI1Mv6TZOtCbbXSuk1wD2/tfoPNvU25u3u2a9fSTLepJlVDzhb/7PfHCfhV8B6bMWR5GM4SM8jxpffVcifztt+M7TlhdeET8ml3jPDPJWN0A9OnM0PMI4vgqrk4br1b+Cv56deThuaq5Wq2tsxQ91FI0JB7BWwrRk1DOKk8mRQY44ZudSysAWRhqxChsYb/5gNiJTT8Zq+EeZ2eZN3N7F0QmCbIquEa4ixRh9PI7B1HWqiWIE2UHrlpP8dHGJ1ywzjHbF+boPvJVSgxHK7QD+4XDBxHNrRWt9jZFLyUWZTZshd0Owa/E3tHKu0+pmXYDnp+f56xS/KCJNmm2U7e5i5w4ewAiqZsL5tEFayzE642AxoKCvyyGFXmAVCQg5n9HNKqU/vDYEx8W5X5rF5/fG6mnv3fBZt3/p6PsAiK92bVs2imxkbYA3A+AVJzsCoYzwkSg1hJNhjh3AAIZmI9oQfVNwn3lJ8JZl5tEiXqI+Y9eXBdKHYFj5OzGf92Q1fUMU3HaKgbUWMhOVtAPO9bZwIPFPHkSk3uM/CDMVg5X1v24cRL2DGGcpzL1qMera/KEJdb0T/uR1qqoL6z/ILcswfXo1fc4x9ZcdOuwGQUUnWxeHZ0KHoBkonAIH3miJdbMOXSDyWDGTedWrEY1igWovaJADppsfyWf0OV4PCWhlxKubCiZ1EoXVESWW/wQ85LMiTY259lFS5/RBE3nQkHEoe98dBE7fLBLgh5Q6+gesVni435otdNeRTT8LWpockXevLu+Sz10dTM9cab0B79o26XBewc8kufWQfawmXnn7Exyc/BuSB888I0fnKaulGZK9yICLyTPIog/CvdjX0cgOSlc1SqN8oymwNiwrO3K6yfLF5PIC2aupTkIsD1Oo2E8pt/itD8WMRyubQt4exZ4rKnyDgB5BmgccKBvq0AzqM8DITUiESO2u4BcIpp0zMOPCH1+tFYHC4qhZcMsjsKwaC0GIzkkw4WdjMajgBRq6YCffLlnzEIB/W8pYC6WE4wXyMAobgJZJxQ7jdO99zvgifJEufm9nOVf1xTyqqTyEU8jpFI7qFVckLXmhkuEpoPjkrMbeiOfVh0UMF/GJ57fNIFAr+PyQUlMm3eLpn4mDOgeiwF2PWL43wbgqK9VqTkGYNXf3CupCOsDIyqQRsMG59bR2BK2d6aFR4f8MqaKzLVoVdDu5YGGPkRdwvnzdu87YxRZAOQtUrNe45WYroXtu3r4ma5NglMIwo04HWttw2tN+FELx8hhSRae9OI/08HTEBD3eV9XeK2lb1pvb4xi+26OreOk4gbz3eLZNbGYf0LB9vUjiRMa4EdtFUMwVHQcRdTJQ5rgs/eKtE/aHDbcD8SGq5egufLfEF2Q9lgPyGTBw92y2Ki8TAN6yLKYXBciw5YnxsDSCfu/UCdy1cwDojc8Q1BgrEmfzOEdz2k6woai48aFUIsA/m5cbeBIZy2g9uL7Dzf4zvSrakBqX+HqBQd4cQfw++K/Q+oxJzaHG9gg1Fc0jtkT9LBdd+m+LeGrSuhtV2v+pcXtLfyDoDAM7Ml55i2074q27Vdti5sSPxjNGX9Zbr/UjH9BTvNDLrJokR7UJkjM0R/OO4zfX9mM59pELkpYee68dnoSNto5t7r0GxhLNTsL6y2AptSjsZDv0cS46svCtt1qbE0MWxJDMnf29NAbFnrXLhAMX2QYVQcN8CmVJrg/RLLXpgqjflIwX3AlmAzuqWvvcr0fo1NYc55guVhQ0JmlHDt4gk68eaSnVtsm6yFsCO4sfj7bVuwYGWwzEkmrUFfdK33VRVMqy+eGIhVCyv13fcZNgJbvkNKS/hizOrLpBAjNbNWdxPonraNGymwvU2OwEcEm87O5Oge1uoMSDm00yQptjTGDnXoX1PxVUUDW8p/MSw083T8MkEb6D+w727vYTWcG7GLFiCq/os81Apd1R5ttOHSmJCt0ST1nRhVF3rg15oe6PpGcoivajQ79cK5uhXRZEBbT3XSRtVL4ndRhOiGxZzGlzMn0Jv3g6LxFrcOHhhskS+VcZe77OXRCLfw+LO8ehJx1tEiwuIJxF8Lrqo+FYv/LOKc90iWhr1JWKwxzs120t3cM0Jqzdbj68vIWMP+EAEg+vd2cm0geO9Sl77R0tMIJZtOTSV4BJtnJrPY1cJfof/E253yYoiCSHshtoQ/BwpyP9mvkXp1XwwJr7cVdcCjyjcn3EbJxKnVLi9z/mHwpA1jjjqLwK9G5STRFGA3bj46Ww1D4rt+W5+C5lfbhUUgreejtiKM5QsZxBH1nmxgniGX+xp+W7gBmCTHMlg8xaGcmaTjNkzML/VmydwUwIA01lZyx/wyXveidS8JHzTrsstk/b2dEvxYOxe3cFvmst2FSSHTQ5qHOUs9mAAsovGvyGIVA4O0gvZT5pX/UK1vpwlVQy/WkHGqDAts9BQ7fyapHF7ig20DmodhkZhMRHPEWhVyaw1Z4PxWsZPOQ/hniNhxV8KlB1QgYRAKfBdp6cV4jXoX747XsFCQJzl5rApXGCtXEB100rdWPkcHl52UX2snTG4Q8LYaDo7AaD1035q2+sgDo909fWVvonQd2x7rxlqbw67Ok124jWktm9ZM46UdEQDtkAl5tb0iN+MIRj/5weJY5RSe6KJRd4dH4z2lfaDM2m5jERofM2Km8JV/P4SXzDS4liKOWjC8J+bQEocTlr7FhojLARSceTp0/dExTf0A9OIoXaEo50ilF/HvdnyY6b3K26ePJ7ZZ1IRzszgverGe0wxBGSJSp4J5Zb3CorkgRQa3MuEP8o5xJ4DBKl9Zvv35PwZ0eDIE6zM0Zw3I77aSAhLaXCqS+SJ7t2IzC59jP15wtsp62CVTaWlu4FluPq6eP9dZ7bDUB9dkyHd5M360Rm1FCi6jhkb8/YRAxt86wDVv00THVAtl010A32DQIP1SRVYqCmUiKpryX346dWsyWWTNPX7bmlW+JPkjB+xkcnSYhO0ZIwQPYa/lte2rwhNfBo775L1sPjpEzY/sxxqNR9w6JafsOEgiNL8ELMWf4TGiTtwGgLeEroMdU1vQnNcIWlYDRcWJw32IYRppLqPBS3qFpZGaHaYdAwoEhR2Nj31xVWpJGAUXKMN5aqptb5qyQe+pllwGMWHhykwbt7byL+0wXgQKgy2G/BL2sttRcnsvg9cuZ56x1Lj84ZWfa9vc3Ye9aAokYz+hdTXj/dYKZ1a6NqJ3iPDgJS4f5xHgF/P9r5Cl7NHiAGxKSwzgF1hC5rnxJ+N20JtnOUfFUzLDAYtbOfn72ZUwMyNQAn2KA7QtLUTC1nSjI6k97PL5S6CyXXkWTK3Dyuj9InlxrqoYQjt9+wr35BYqDOh8w2y9mCY1VVPQxT30GRPzO/EgZpwy9TxHswtoDxHgFeITqmeyjVTi0adUhjZvSMq/uG3el9zPGT9TKw0m9sdaOOXrrYnjFyqd0pMtkZZOpZ4vBFFL7LpUY1YzOO6waA7vPdBmwygwQ/HuqHHPf4DFgrBMwjXoCcLNRFkJ2JbpfiOQfpXR+51XwO3TSaEsJHFqWpoLzLy7ddugouPkj9xLNQD3IaGFsbWf74HsGVkPgSmd65TJ4R4Vo/0wZ/M4SbBLpT0toI0lVE6hdcyGDQu2/Ht+cWdAmcdk48SrzQkSi9umu1ZsGIJCZ+YgB1e4C+olObhYaB77aGWXronBTWTulyET2DksXnbtmp0BqYYq1+DLJQOZI98YYLFaIcQpJzAqxz8yKNQHeZCqcbH8YPeTnXRT88hLwLBBSYDgRkavWdHvv//Uxjt+Asf9T4IAJKEwuJV46VWs1ZrUOx+A0eGwbwUnyRLvkF/yU4e50UyovnON/n39Ovhw+2X+A9CuRgELbKTMpPDQ93YbpMWYWzOgeVrz1wcGKssP+McFBoAguYX+NvqKO08v4tdiDrVy9SjgKT2It90HB1XLeMqw8HQdHmf8eSmVFrm/Dk0il/T47C+4Yn4eprET02i1DqzDCYLWoauvFVHflrfgnAPBeMhixLRG7i7bqSQeAOYhzEzaV+UMHL20eF20iHQt8ibUGzVqSQWWqwHRAd1Eyhu9l0isGl+v8GWCJkpFN4RNzeR2KF8Koprrv94OpC2qNezEga7uh7dWe+PtS31/GbMxOMXHvRbV7YfgccKgTiLgj2LcJAa3D6naiJGYpeN6CqB0/+XRYkly1+MksdJYco2Oz9+2i9LUkRc5/JEdKiyKgJXJOz3AUdvc/+uj+dWFtzKXJ6LnJcISkE54/QXRnd6ENIFjbamLzeasFyhcAiiEoVS/9rN+kWRTQfRLszpv8fxWg+sESLqzDqiMKYXOXxLIDwUx3pLSht0xtFfaD6QQ2ttKdZWZ4XBxIDdS+FgA1dKN7xZFROL3m76iY0WsvaD+u/I2P3kpM3SiR7bH9oXzgKTO1PWhuz4iE0XJ8/Up1oqel2gTcVAwI/DnKEH2fyQ1HNuT8Z61bkYc279l2HAy8Ih62i4R2fZ8J30BeoWd1516eERrz9xauQdtJ9YsNF7QA+5/3fisHIBY3iLchsLkzvhBBqaTbuuuWVLzYpbqOnVdGKsjYvTOh9h+jiY7iS966n7GxByNAZyyA90AccNIgLlmV3jR0qNxSGARCSPZYGGTCKmMTBcAu0775cbkhn+Q3GGFclpw87LEwzVP+/NJlZSLlq5vKKyIHPEWgBYQSL/YeRA0l24WCC67haYoMzRmqAtQ61p/rojhebjlBYczji7pDxwpm2SoDvGocbvA6qQ1ax6Tu4VKBTumj/zf6aGqyJ+UjdaFuL1S2eSUVG2/rJdziZLDRtMUmN7G6yVT8DEZnjtVhmGrFc5yCuZSUox37FRXN69MHNzyC7qzPeCdeGey+mq+qYS5o39WyAeDtYgdckuymXuULlAHQMhTu6QpEZSbIinJUbkaVT0oAxuLGLZn+VS9DT4EacGOH5A6kEjqRYhkVhS7UI49pQgaa9k5brIGRHB3N/V5lUIbsH97a+19dybJDHNcSRzCW4ek0X4dKeusweSaj2FJMiiFBZBtIYWh6nPUQyiKG6vQEL6lywLWqpCx4pHQX7ffDkRMlFRPwjyjGipA655c0RJ+Wv65FKEEF5IErAi/ak3bA3Pq+9Z6XnAjesgfvQkj89xFpPfbeBNFtkZhMzp9J0z5i/GqJRdA/yiir+gLOGlQrKppaNJXvifLqZkQD4cqyIFm1GIDS+LwQAw9mDhhob3AA2qIrqjAjtE1PyXBTRMoDPDfCFGWlfGY/MjhKdIvcmRXdWvFsLmcOOQK9KS1Mu47Uf9JtJzeMay9cJUelPLiZ7jRKjLNQsoZ+/Mi5TnGhlw97L8fBrTLm8jWoHih5j1SN+usMv+QcyjF0wL4hp6ko+P1PWDsVlPjZNZyiU+QSRq2QwAqeu+UeGXgCNmxn0OQZKmx213Xjr5PYDb7kwBGPgbSRD6y6xobnDGcbVcYr7UR6CD2GByymQJGfF6Im7u4KS0de8tccIc0kjytDwxISdeC7rME9gtdeQZYK9oA3Qi4iViwc1+x0UMWgdQ3NxFXeRxLzJmiLl4aNGfTndBEBlvz1RDXt6zobnsNHnpRg3zuPjVLL7UcUygkTm7JT8u9I4UNGSOKo8we9z/qUNGD1nb1uXCsj8bs2LV43Yprr2Pp8UxSYTcadbi0K+BUv8/m+jDoXhOeoKic/xDosqL7e1mazFIxsGzjmZN+5gDUtil5W5kNOfsh7glVX3Ea7ktuSKx/yOV1eR0Zm+2GnP5ubwbmD0e8GUktB5wfIvWY83fN6szWl2/7RVHEmtywpQX9t0jsstxvFfJywIujjx/s9h5jUQ3Fj3/k+h4LYc/FQSLyZm4IMOq8VQPGHnxDfYxEXW+MQdxQj4ZQqme1AjVD4ss52HOTZU1fKdN+vdTqdDYktaPL6zSI7GSju0JaUGiOw1gHakCQy30gnujJgtNstscgu4BmoJUCXgUPc9Wbjn6wrlnLzkBGeayw8lA5hAPmIEcyp5TbEZsLAFFs7tsgurfb0X5E2r4ac0/diCXSQ17yOzpEXtKmnNHBlEgoe9j9bD8311YXscXJceIF9Qqwk56q1Ue7RvCAymEPT8+XroS9KKA1ZS3RT2okex86XGYwxGw/gcuVG48XdnR4Zb0VsnJNfklz7kzT6gh4SsT0ozwsi8LwRbp78jowUNZfr1dRt97GO2vYAMe3AmGKXFOo7/k7nHEeC7qVC5FloCUHsDXLlI82KNtTMQhFGdLhYA6zhj5JPjJwNnUjTNomAM/vlnpY6MbwKmtxmigqrCWI0ostcvntxfzRLNqQzYgJHP8scpV9RE9yEfXfPk+zoO4DVzhZHF5w0MajWa+9ATXM2GV4r5UG5nvg5bSRAAHMOPU6k85aoSIwNoeQO7g6DuzqijO0yRQj9VAoOOxJ0bRZUWu9EnbSn0PByCBl9sR8gK0DTCunetWNr8bfjE1yH85/qS7yS2Z84iSy/b+InnaRlrCpoI6Zy+bYfRt20MEjAhZFfUyxGqxkRci4JRDeWjEg507MZLWQhO7pBk7IbZcScG9kqvXm/YC6aHHtQNs9NeF4Do6Gdpk4yHhzZTFRusBzHXt2NFZPENGe7b0zMuDq6vGym6C8Zb/772Vbx3tBoHQgOFh8Ji03qeFK2abMM1FFFnDMy13rSlDRKVD6QoxS8Gv6/4UVwzAiRqobfV60g/gVk9ggpJG7Gs2mFZAWitdQN8lAeHKfMmQGOfbz2b50UjuaouMOhVy3/aGl/+TOsvCkG7ZCUWmSCyWvIkfJNGHniVGKieUK62D52VyuK5PsqsEqtgWs9cPHBxWypoqPTnEfD/DszmI3xqzVEuk0TXMBdjyaa68iWNotiZvfQxCndpnHBkn13cgPcEQiYUe2xT9HA7W4NbD+Jsm2rFzgJR++g3ODgheBr7yqNETPg8NxWUUNCfBmRcYJNwuH0wZy1RPf3iyKE1emzQR+dqTa1fGH7VDHKvM3rVq0tmGwlraSCap6ByAIDw3UEBLQi29BIWLI2ckUJMcatxSMWR2C6eBSBgpOsDyamdWONKDsSCPMHUAGmSULnNuN84fWphzjhveBQLg15M76OugnJJopkiV1XrUwslga3CYhJVkY/Y/v0648aAg9LCQHGaOED0RHlodjxTl0m6z+LgTJX+J4GjPypJGasFOYPrhwiuQa21aAK85LhhYLlm5x+FjuCtSLWasMjoIgs1/EcXj2DWdQcK7GkYjHjQnkJw0GE89kFjDfWdyghG1g7R4ioKsQQDgo8lTipGzfZrIDtyPneiqjb5Zs167y/C9KW8Xw18Zi/Uz4LPn1x1B5ImiyLpzD5iGXlJDheiEYCeHkf9jmftLd7xrX3PUtfsTFqctMCeJUrxaJawlAFTDzZwvHo783zV1mKACxCSAl+eIjYoonzkImSzktGEK0zsT2j+F0PMrTWSJtFMOtAzcV0j/bQC0c3H20sKzCXHmqHPBAnajdL5Cg0Hgk+DiXuEJtZL9sXJRnmZV4AAEYhWWmojspMBVhgvCRWEhjiuxe4BXUIeuad6NznXNQp8au7cb9X3teLK9ftgB/TYHzNKH1LtXobitBh50c3XELxk9i3wPprKegmY+Jgr3ez6ZdTnhZWiDvBPeAj6HtL6+mWjV5iqaQzEbmXT3rIL8U6UPN06ClQ3VthSxeLz5r1C+oC2tmN04+WbWE4EX893AJhVNikGJ7d77IJfSdr1Fc89Zm5Sop1oJdtmdvBwnwUeUc0b5WPnL8By0CaSMoZOJeZ7SqNj9JQmE+c/XaeHYek6WWs6EoEl8Ph3aOHPH6O7YfSG/9YHszOZPLyeyjdSgGG2qR33F/Xh00qzEmWIUqXtKZhi/M99ffS3JWidybDrsB/yHTd2mXk+t7fXia31T/YJiRaP+ZtmJcVqqW2XWnbvr7h7SaZn2kPNA67gmR65KzMDjKTxZXLsRVfPGUb1RNX5Zx6FEXgeQBTQBqmfuDNViy2nDwxeccyjoTlbRbw2iRVlxKEgh9lTBVVGYIZ7Wf6o2Y+FQcJgbxltPkBK4J6admOCqzWWVP39Y2loMGcpumNHTG+r2LzLjb8iiQGdrup5qJQTmXODP3/oOlJMIJos+qiyQgYCx3C4Y3yYyVUZH8WiNO9oms7yKzF6WVfgtazByixc/R7UkqvtS8SIKiq8MOu0FcpNEVZUpAk9ZR+yJU+S3SREFPHriGQBo2pShnZlGbn0mD+n902JeKQ6HeeNa5h6+NkzLym7EiwJEMY1xJaqA7piUgTRPJMtk7ELanOB3AhxEFJcT/tq1aAmloJXBx70e4V2Eoeuuhv1y63NJYy3CASzX/ZSaCM+N4YAD54Q0y0wZi3MchV64fCyGhZIps7S7+9cSvoqTQZKYqWGpl1TZB1yXvx/iR5h97Lb/xu33m9pVLV92IEfMSLbOgC5v/qam3exVLP5zuJeYZMN7qDzNhdvFiAIpxL94f00ER4FEprdnARvGpyMB7hqSrsCR+8kb+qmfPL5dJ2XvjpS0FJwoL3v7XTMqHawtiSARihW6Mn4BAAGYUFljJn1r+H/XU2UybAfHtuvWAXa1/e2sBAHgiVn09a6fK9xIQNs58IqY9gsQjDodgRW8LPL42Z9Vx5Z/VUEdVROimxu6KfPJI14VNv/6pzosTqeyjx0HU8r0suivIN5hmoL2NLhiWrO21sxbCmQtXTAHK5TJtS5C3oS8NT+TgeM2r8a0vLQTHkOA/fiM9RyyJxTQmA46oY78P/F/WFvGboL8uS830/dsjgTLOcQPkdbsypF/KqliKnJLhqkgaxIQkakJLCq9QdwV5KdOpV/uxDq2TqTBiV3Cs7YE0ImhkPNmIMTXF8CxQ2K77o76Dxo1tL+825GtCJ8fg64lR6b6uRm8YrKhvd8EWh2AMTkbcEDnicBTR0x/k8w4HJi9lRc4QG3Ved0ERu+41qZL6v+jX3MgCVG7LScoLBQ0dyv+qQPGbV26SpAwj3JlAlyuwub3J+xkBhzthPaS2wKweiSiYDc3elywiX99nON0t7hdmZyAd7RcRw5DhsDVQqksITH1dmXao9rfiCdVYz1qcNAyhVoXHbISGJhZgZQCsi5HmzzzI903emjAAmbaViiWP39277d4U2MJbrL+hH6XtdaYsCqeE+G0MpOqsDvnqseIXIeblGyKii8FzSShwKLq3758VeSc893lud536iMxqVzsQ63T+bZzreyvi3yd3nBvgrVi3sxNGSBxLiynffPTGL5B9cEh88LlQX1/qql2Tv4oWIdF/LqbAXyEu/lll9IzO9uh/1tkCyMvArVK0PoI6atwKh+u1wsIYxcb7N/dYYkOzPP64o//uaKfz8Lvf+SghKju0qgAUS6v454OrjpWFa5RxAiqPig09mzzkFTFh45zQ7Sf9LA9q65bqLJ8gT37lNIzQDX4OCx3dAv/+ZHw5EDtsLYAhl/K3ZUY584fYYOULAgVHGGu8yloRojcvWHKIDCbYWzyawKmxnY/tN7KtWYH05WF4lop0LTaKlJj72fmoR4miuDPtG6h+7DPp+EiRxEy8oc9Jk3yUcS9amAVIo3UuffGplD8JSh8odGWM6ShgHyPhKLau9QgFnJ3sQI0sWw+rH0lOV5n3BT0273BtbBUaYM+QkBYfYngZMNtCHBA0mZzgf0lMsMrk3HAibAH9NVT7lbnrdpF2bFyCQfSkKCUYgURzuR5ZbB/w5bAQO0mMaMZU/wlXz+7T3D2ov7P5gLF3ZDmIknCf6TGHL+ywUPXEItcNUI89HMzkPONZn8R2MedvLeARjETFBahHfKnvAQHrAdUFkixOCuvg2yueWI8iND2GIfwdA9dBoXFuX9+RZqHIESmTqHRbn+pK2PYvaIu5rmdIjstRyjsZ7BzrSrJMmT+PI4rQG8sQT7SASGQ8fZRcooUKYP/xfQmQ4X0yD3uzdEwi/GRxv3+QooVLbu7iRLQpev544EKUJr8vFXcz4nP3V8AQHfBw3Be5JYz6LsP5cCG1JKjQPThKh0KjDAxRyoE+UfStRiT1km2NK9d/gG4WX26CdCE1BeH+KgL8SZrxHo4CiaSzEWIb6oNNxxeWNl9afV1QPgP2mAVDzg/M/zhKxgsBS1QYsPq+SRdIjs7wSLKmWeVbC5HUDgxIyVLJXljeBLLcM9xCilno2TC540dYlM+2kd6cr3jfmjYgPyfJUBa9rzb4PZMuqgbAdbJ/5crN2XqOscH2yEkx/UTtam0+bUbetV8e5YPzMvSLHlAnWeYnULcAQ2b6lPfJDh7SLrBs7fNbQkQshzJJ8iV8lougwediH+RRwetpcoHrqoNLVhZZLrwiEXs22fClDrjRN3zSbAseC6tqUjExmTPKuihPIR5kWKF0ge3REiHrjliVMfgSstY28M4/p+pIF4WY0qW1YrbqGu0960vYo9W+b6uLwhlyk5nrtJfgXFfVny6P7ZwVzrHM08fdihYfacOlYOZtAlytwO/avHgmys63sneVJEoz5vyeUJYLNRsxdpMpt0k63dZda9idmIx3oqiBWzyZPp7zq+xbit/lDtb32PKnFghebTu3DGA7jktc+753O77Qh0i0aQ4A7CHc+8Kvo/3ttM/f7P1PsY4q7+gYLFZ4MVbtBplD4GOEXeLe175EU+liP9gOdOZX4XwjOhIXO+DeozYqh3a9McY3PpzrDbFP/MWWpWR64Lap5nos74XR/i//5dA7aD0/FgtgNv/21cDpEFoIPGpUJ6TsIXmgBNpQ2U9gSzdLx+TVKadxNLNgXtqjLQ4UMY5SfQy0tBf/oS0KcxbnGERf02o/KQQ3lKYiTCF6vRKRDaHqBOVNO5rttv0jds8thM/UdjA50uB1nt7u68F3mW8FujgcXro/aS+FCpZ1YhDST8fwf7QPeLqWsyp+rRsdKd/grEqqmozeV/C5d9zE/cnQWQxCnU8IfxOi6tGH0DjzAVewg6zSpiA+/HqaDTULG+IkANVoUVz+88/Um8p6fO36tr/O4FaEKjvAV9d34SLo//C+Ftdo+PzCBEQUVwAONtQAw8daxZQ+UvtrCh0mU5ENwM9W9kxMtmEgIUAPwf3LU56BYe4rVculwFg/cCNxZpCDcglpK0LwwvZ7O7jAw5WWjpgph6HiZbf3eij+G0gEZbKi7oSVf70swf9xnOSAU8eaIRJuj0vFBFXuKOxRY3GU4JmpSAHb93BI1lWnBx/tjtWLhLnE4nDbG0o9AA9jjcnxde9XvP9jvVshV3m7KGVt8XmigOrvuVLjZmjVSQ8Dp+N/iU/NS/tCLji9B7Ne7TpO7Y5ZX1iXnaolC6FRuJzzMsV2MicJxvAay6zRRDb4wuUJPMqAOdCcTt8g01YxHpUqh/hJATFRKkqG50TKRjPMi2zFCRfM5g/bjejcPFU4uomEwz50ARxZr/op7yELV+S/kdR240L3dyVKPAYYyqotzhHvcVztMU/qACItLdccjBzxxKDQGFyTAoCW+IQh8kun5AfDYVHgQRFpSzhaAyy6J1HfnXg5fXPW0DhAkpFgJR28PQLkfowmsjsS4tRcVWbaGYLET0gAcZ7JGpKmqMs74AJIAW+ZDmLtwaWzUKnkFroT2WWN85OXBOwlT8JZBFMdo1ivzjkSdiZPdnwFMAbqEUO1VKbqzSRFHN4On/KPGyEXHctXuPEpc1UTwXbj9Uj/rVlyooDmNSnvMfNJGgLSp2puvK6TsDcPS2dnIZUbhPZ/I7b51GFZOYfGoWIote5QHfwDLkNADr0p0dIjwrd9JqQT5tXQzTjGQw0+wz1C61UMOVb/Avifl+czD6zVO89PESLKXy84JC0uqwdlLbBHn0FojNP2fpCCng73Gs9FdF+OUNanVW29PNl1zyrysIk2dNLlXt8IoJTuwfNU4gSsZB14N2nQyUE5hMwiLZM/GxfJyTilHN2wfIuOvdarvS+4PR2fTgOi9AAcFkB54JQMgTdiSxIGk7n96Q2S+CVUfWrIWiSY9GK/KyHq5oxpH7/e8SwySSRM/2fHgJCkdIl3xf/GZcX2WNmSBNuBsaG268vQ0Ws/9FwcgwVwl1UNKChBpME+tawsyqMCGBAmzOdgS+rsPLI55k6hZaiGiPTJBaXrfxzQCFsRWwKd2OdSP7xQiAaeeMhEfaJGyN9Uo7mTsmgsGO5FG4XWBd27JIT36AsXLcA3hz9hRQuB6uKbdxI9gnTJc/5ETpv7iqTpOb3OEw2NTGuB5C2qJjjJ7DoIJcyjgW7YZHfo8/OPk+CjTl8QiRRqmj0vJ7e/6y0cz0sBPZqD2n4gp2d5IzuyBP6IAU1HT3NnN5nwQBw0h7w7gxDdEywcGl6/Jh8ZRgaUE8uRhtQrfzomZ57cBgzeV3U+NGe7G2mLr5/sHbamUDIkf0pUUdhtAYkeD9Y+0fSgeA7c5iMQvUIaaQdyv2LcbQasgzB7mFBC7b/Xv6fSX0lLxDBWPp3zcQ/tDTC5kzVEoFkI7II5VWwD+OH4McecsQrCm5Rg7zGs9VQBwYvLAZrnXVG+W9clTv2DwPyuTgXIMOmHQVPUbTOTE54z2EQ+fFiv9I7J82XLErx3ZlthSbMjZhGx9rhKPTyrsD0/coqLB0DQnC3U5IC+b4K4iEnYl7fOGkB4fz+7l4Aqn4yMZdVU0K/eye0wkVFyhFN8jo1ROoenOOpkl/Z4sTyYh/CRHz7cZSTWMIwDE1PvFuPyutjvEVgyTdpwKJZh0Z2MVI0oMDplTov1ecifaceUFOblupUaigi1cIVnCPnea6sFDh58LC4SwEWVQaS5KHC7++l3MAFddMY+59vYhfC/zMdUAkLWr3E6edwm1GtBxLIiTM3mSywz6KctbcM9c56vX3Ge8cBRQvU+3fWTRk5LvG8ArE/AQGlN9r9Ll8f9YnI5w6tfBqPLuajoGm0OA+2LsziJJDfSRwWXUwgQsg3x8Kg0KnppI9Mzen/m0W2F/ODydDYQoZqVG8v5gPH3RkGBTAAxhPc1LCScjzfONDq+gYmShzKAoetSvfGTB7hfCGulXXa99XYBoZjK4OWkOYRKXb4M+O1O0m4n9tSlZOMMa2ZJOuvwXW7zpjVtfxuMK3t8Cc9OxzRufTLs9rymdwtVS0+msq043PXfqMa5dmi3q04aP5BhTkjnuwaRq1ijd5OBibwQp0VZ3LI4IcntIA6yrkqx36HhiOwZ7vgvEddAzuKapr6JY2cAt6eTLOXfjzNtDrJH6JB8PcV+dt+a7s5Q/8UaVV2O/yD1IYeF3RsDGzLoeuHlkHrLGAoCb5pBENADBE4Ibus6gYfMS0jWnYg/yes9zYMAiQl5C1+Jx224beTXdTV0k/dUsx8HEg0TkFsoHXxWJh/RK+tSCmpSZMb1Pq7BIiHRoEJMvPpxQ/wR7H6PvEhgmSzz0CHCfMK66Lp6ANXe5sKovIg66m4zXHeJkAvdMYfYWSmYebCQnJzL4LuW4yWbjhNVv+8LWmwjUWO1XwtSaStb4hGA1g3qbC0TSvSaOXdQ8ztINnsZQJ6tiKHcmmxZUzubeVuGU/sZaeKPdrAbCeV/DZmf7nGT4q58YlXhXShoArOGBJ/lclr+M+8uAGVtSaTw0x1t7Oe45upjxxar8en0E2+2Ml32W5SsZkrSsxcNukeeuQPfNQLrSE2fTyhDiXieNtBqRobxAg1z7kVdkfWCAh8hoH/S2Ekajvv7wh0xLh4Q8ij3KuH+fqufLRpt/lmjUxD0o9dRVlLT+A6yoXwc9pJSOUxw1XfGypxWJ8uIB2q1OvZ9ou17aTbYBfCJ6hb3+wdWWKCYDuq4yX+Ji4CjZYwpeWa70iOw9OaV5zBDYNoENS8GEr49Hs+w7SF4Cj5zZQdoQT60sXSZ8n9pjCWj1DKCY8GvFjzCwknzoxSNoYoN/aIXjFPw9QU1y8W9bJhaqYDQl4kucD0JGJIz7wjiDvVnjuFyO29mjKLFW9sPDUs/dSuIrmLQH/3IF6exlong2Qu3ckBCMi3yyr2pMvjbTq4RsRCHTjFDuYH6qga2E4edZIId8Djght8snonx9L8uT2dfkWaRDUIBnZ0m6Tcf8NCXuBiKr3YrJRdQxFyJ5qxzTDZ1whi+ocXucwNA0s0QBFaRePbVGEfGf2GNteZUaTnHkKEgM2UhqJbaJftz4ORQfk/4dO1tSpffWM767brUyAVXKpN+kYb+nmxwtN+6/AE9USWGtlXuRyGWbo8y5UFyOr8e+qv+DkIMmVsGVXN5j4wNghjvZklVrdc4F4m7AshlwI3v56nObvzqhG5K3QmycrukfmFeIyReJKcDuNyzkaGXI6iSV8rlHA+nLRQbJixcn2vMf5JsDrr1r4JiWz4soHE15XzAcRoNHeckYr6/8uXwlXD+rA4uvKNoS1YO3BWOc5Trp+oNAn5gOkYlXQVKToqwQXC/fkBe2Dmf6m/zzWgCEvwqBPaBVwFO1dkDMDX7zWYbYt0lYoPjwsn81QGvPE15+J9M6qhBOQwexP8ldS8Jw2fxAYRNoarm5uyyVfIp5o6Awmg5tezfL+3xTVnY+ez28mRmzyn7jMq0a24zVqCo+tpvvr2Z0yJ/8FjzzURUzzzeObWhJdv57m/W6XYlJCigLmi4tsXltvMVBUwcKDRZ+KKA4MI4CX+6YOSskwkfHLdrtySTTTPs42PJbFkVNqxSIJSLuZNVwAuRiKacZ7c3bbYr5A2H+t7TZhk4DmiIoEJhyPCvt/WiqcDTir9Pb/8shZAk3bVTAqSPqmQf4CRAqCBp59GV5mZ/tOBqotKTHvstpEbkW4zJbQbeC9nQ/LWHFW4ANr969yd7g8InxRbuzRfSCGkoH3myJQUeTBel3tRx/qrdFSRUcz2xtmAnja5FO7k6MMzYuXvcOFRcJJkNBMAgewxFi1+kuTNn0xdaI3Rrzij4Y+6adqv1l+Pu0IKSu3UF5Z8foxB1w1adbVT4/iglWXpYMc3RpS+amDEjTEtFEt28y7cHKWJ1q1Pp3mtORTHkwxlQTHWXyziWGtrIkavArhwe0eaUCaKn7cPE5TmcxfkOx5LLypcTKKfKIAhbHk1NuFcPOP2cMg0GooEX7iikASZSU7Kqt5W/H+qAzy5qYUU4VVvVbaFwdMseWiiwdawAVzxuPwfLkEvTRktwqams6nYMLofGDdVJy+gbepRqz98SgGLr2ookCofRjDp+eMFxdlFRQwloHT/3GjAtKLGq0Lg+x4paTTKCDu+8SKT/Jlda2KIxhfubO8KlnDNQNmcH1NyOrUG5NYL+fGgx6Gs5aDSOw6/8yKhnEAe3gUlOhG2/sKvoeljxQR49psO8LSMW0Vpwtpe0GrD4x0UCz18IzPMG/84tQv5aoi4nCmBFsklIaxcVpXWQgMcBqn7o1i4zkkKJANY5OprsuBQwKcg1REYbbUroIp32LGpjNHGm9Fuv93CumMqxKogufkb4FvnWagAgiJ0GO38K1DTE5l0ZACdFrfP9H0xHpwAhDs7QJbGQdo3ElqGfRfw0tPWy9ydadLu57SYxrnEo1553/HkBdvCthdo3MtY4sooiiluh/e3Kv2swxLLX4rEZqJBJ88195l6sdCDENlQYE61KjsF59l3jMVhI8OtvGRZDIwerEqLptEPpyUX2RyhMCYPuSZAx0rqlf7uTOEW5Ook+lH7yIc8Nnx1NrSvlepLoNujytLyUIBgSjCaC6jbbB4im6TGFuL+y7crVIUIASYcdppw8xJjZ/SpGHdkKlxFJiOU0e1DG/jO0FdgWBKVixRaKZyDqgAXY97XuINi4BocuyXmKRWU3MH33vFvxnBS7f3x6fMzkC8UX+E7DgZU46TvVDDDE5Tj8+PLt3fIqPvhcO/RlMcR8ow6WtQAAcUmErYhICIb+VtnzLl1PKI4KnLPvSc5N+hUQLrD7L8RvkSaZBWrgNpHupQfGx1xtbxBmvcc/RQCECqaV6B2sfUenbYUqs6d/PfCIsUNJV92obX+DBpcarPIwMsbfgP+ubAqq3vNY851NEoueQxXIeGsUkcnqb2VSJB0s4BdxCZJnPV9EtVwmcuKogmNX3gGoEMsBMVc/i0TCzdpPbjAdtGIzReQI9uLXOB195usezwJr2MofvOuanxoiZANs9i/e/hQdBAaKy3NtIEqvt+PWqqC+nE9tk+hUNg4oitmKXVqbelhYJy0x3x6AmFjczjnhhabECns+cDAvF4uVtzDhXECBwo74M5QV6tS7md54ftDG+6En3TBCACxY/URFUYLHbPS+F9VRUyMYkvmWCl7Xrl+oy1/+jB4WZIGoixS3o61rw5XDJwDw1wqElMzf7TwAqOpYs111k0MnckBmcCC9gkQdhSDSEo6z0/9RqNqy/GOPabq21y6n9aQVPA+Xn0N+Emf2D5OAtMxQCDx7Z6h9x9eDNjdzhgoBfOcNWoRZSUw+z03uMe+GBHXoVvKrhy1BWbIEADIoywMfoUudKyPxeDN/gm5wvfPNuoVJlK3hnAWR72leD4VaqqSvv16TwHoYOvrnDLUKD2+37lO1Hoessolij3onxC9aloFOsL1CHCSxoq4SrSzYYhsolAQDNTsh1P+Py80OGWmu7gtZPrdZn8hWvvAG3wX0LYfzZ5bGXj6D0LLlyAWyhV5A4d4du0Wf1KBrURFeIjQMeFbg1iy6GK6skD081chAUjCKW9RSDFTd5QpfWrZBYeTb3Wtjji4JYhpQQssn48V2dm32DmVpBMtN3DIRfoRsGHABw8j/YXNH1KnUOjByxPpkiK+OTtSYIay+eeDasqSjPvclUu6anvxN1MGDcYLASluw+0kpVg906f/J66c3QihMLpgRT3IBN4pF28r7UnIslw4cjdzr9M/2fvRKlpsHOLoF+hET4JaYUfzGYucQVpv7jfHs7nrYwrxpE5x0fO12nGk9KWshORLNJ4qR8Le6anwqQ2RTrFQIE9Syf50lle3XVdzypFawGNatf+YweKQO2d0dTgU1zuOD/AlFyeZMTt/Ys7Hbcd04eggmEPKBfjuuYv6+nVmDRUIsqrzCj319yDLpP5AlYRgGcVzXiJxmegrbVpf43DqA3OEi5WX/vkIGCXwRScDl2Mfv+JslmnXZOxqLBfVG2jcgK/L6ZKM9QfNPspT29nv1Rne0JcnS52+OE9atloY8t/f8PK+9BX1WlBI6HF4C09v3x67mFVzou8R3DcuVn8ut30IYB1feG63V12DyesA35ERg7obcgQD4uFnZ0/UCcgw8jCfNmAN8c155NBSCvNQKoU3YN39wD2A7DT4UIbKZ7LoRWFp6X+xS7VcnNdJS9eKwHFUt9ddW2um0S50NZS4D8RaIZwdc2pnE9d6JzOoCVIN+P9P56ToyaABAikNT1QB0p2+NHOZReQLqLK0L1vaGPbDGzrChFnpUb4XZkXMr3Ga/p1N+uCIeiCYcTpxw9uux/l5DT1SiQ+aRauLimtE78Z0EWILyyZHD5JL7frfCEnh33NOyUJXwr98HhjBdgFtxG8TcJt58vZdDk0DAHhIadTwTawsx5VqZUfQjLs6E+LZfwUC2kWnOU8uLG/YgreTIEENthG55PFlghob0H2vjbvjBVphtCUVFVgdHelASzYgE1Yi63iy4UUoRpG/Nm+BTuVq0YrZJuH10ZXdM37F4GYOcbD/U5WwAPfffXxJbxB3mJLlGZ2sjplePfCzuaOSILA4i2EcB/RiIAzshCpYbg9uwtF+u9wqNgBqOSB5hydeKbAQSZ7A+IdEg/RbRqG5aeXvvwi7bz0lX0RBIvC2MS4c3TvKrrtTYJLWld/fUt2YrIgLXUxRhtq/AmfdEzlQ5R3GHBHWYIBRjbsxLmV9qly2JDtxCj4S6FOCI51rr/IaU1hQC+oaR5RHZfwFIzceEAWRNhTK8dtLjA0j6u4DBKpIb1CRs2hspewiS3JWwAIyqerUESa4VeUOvXsEaRps3k/QG7MGyh13QPufVmT9U2Tf82hrWUP6w7hf6FOkVv7wys7v9vYBphL8/e0DWUQvV1dKeKpdSUo/jWoxhe1/00Ors8xmHzELxFITaipSKOa/iU6Krl0fmzQ+xWSi6LmKsxlEqFsnk1SheyRFKBqriMc93JNzzgQ0kZu0jIH4mexaUQ16taiywGA5ErOn19RrMFerXiECcXzNrK126nqWAuc9gK01gpaMAvfSSWru5PyAnIFb/reZMDFnngGAmAs1/3Fc52BhQZO1jwu/bnFeogIIYgfoKG1YxjAr4MG9vOYksiOjcL92dZv/AMFkTDfOwCEal2i2ik7YGxTTb6oT+fglrhpLARhJGvtLXRyYUJvysypUSoyTddt5R+NCdHq6hGc/5gMOjuoS6CkTTaizXt38F87ocHQCFcWjkPq3ouPG3MInJ3G9Tlt5zMEpjLWXyIsG8cc8gbOTDXiayhCNL69U/Q36Zsv5kJRbocjqV+EYO7wBUK/BMpSIj+V9mZu1sDnGkQ6n5sR4Cula43DPj7+3mUBNLh5GVLtJZ+YHUEJmdHE5tKA0lcZNSidp3hAR3yIhQetBfc1/frNcUXmOodBR9pUVMmZhBH1lCCbfja5yc4IamhpdnsY4opcwEU9BXAOx7IS2DfTfw01AyD8t7y90mB6iDM040wX2y/fnEFnVvsEC3TxN+AFeP0PmeowH4ANggrem68Vy6ejlXny5gxn3kYHfM7L7VjpNe+vi6PFJmV0lEtazDHsE+9buViI/KQSdDOLzUpPSAHH5mWwYE1OSrPL0kPUdV3VCKqlmhyGLZCWTodUq1wYHdBDxr71l1BUc14N87hfi9Sjoijq6/B2bN5Pm734kjWCBqRyk9mOh8YLRkm1V5lrvCPxTY8Om01ct/xZGoh5kJ+rgR73p5xTB4OU1AB4IaZ7uSlsScJu3+AG20lVev5WTosyGOlb06I0c/dBOZuq3KXcSvjlM6OtN6squOrBL2ysA7Xgc3ijugTf9uvXGMz/nVZJR6f8oSWKxTGSp6weSNWXIms4KPjnY4rE3QFAvvW9283HKoc1+GSWlk5b8Y02zcANGT6Bp0B1gKRkgZISNa+nJidwWflAl18eN+Bi0JYlk6ls2LbH8PV4ZHgwH3/nWo+ORJyjHR9busi4In1H9TRlGupoYanxBPKu12fWi3Llu7pgwdN6GeflFGJtbC0kdMxCrYIVXiSzlTqYb7dj6GYQHLdgM9KQqlCjjBRErIhjmUL9gg8Y1dyc2aLTMNcuiBkbScRJQvkZFePRt7mDM1oaP912YRiTbfuQDrJk4pNx5yGTaRi7aYwuJ66Lh9Jlcpy0bJzovvWeyB1Zc1PkYZ0LzdY3TD+0oNz6PoR5qBgFdDJTFeGBj99KqgTytCcagKIS6+PbR/WMkEzYZMibIhkpSL/D3FuGA46FOqJKh41JeqFc641fl6AaImJh3cE4nViKm+9NgO1+6bg1Tyg3oWEPzpOSZNlcKNaWYE72dhCrnA8dhvhjBUJPgQPeqSz6hc2sYCbSYK/Gr9P8RpSOmV/nrqhefZrKXOzuYDqkFfeTzl9nSiCkIydboU7jN+3ULLvXGAr63gwvi2w4WwvcuDcb53CgzrjRb6ZsHgLCFKm5JrPzivcHRq9KsgjFXXLOEG8PATQP0tMOgeIvGjQdgYuO82emzVBWfjzZTk/mI0xYiJigBBFSHGYzU9UIgQh8e3mWzxu78spR86LTKlmUdMPGcq6tAVdeCOhNOQpk35dKSLjpeXDF2jdJMHLq5w389LG4ptG7uUBzRnTRb9D9Or8Bj86/jzcgNqyWsV/Pmw2KO2ZaDM5kX+Lfj43dsN3KWZukc7bRf3V6u7hMSanFbWtEXxC5mHiSxCIZj6ZFAG9myxU+XK+6n21lp6GehBL71IvI0Ijd/vT/bu/It+ufyojK0Ya0EWO8dIlXBzz2tUZmu7xVrYeDFmz9M4bRWW8PpBZSoAgApxtyjBgg3sdcDat9GUwiu0gjeAgzxqE+x0qcyL7KDf6MnHxOgZTH2qjrb4TP3PBLDNdEnm0vmW8N8ubcT99sPU4RCybGuRfSbDLnm/WakfMAdlbQADon65j0UTD3aEjPVvtU/Z82yu1vFX3ClwV+k6LOePiK4+nLJUo2LV4lqVyAVCLcUnKqLC8OTyRfRb3ChIjezyWc9FeN+L+rxSivxsnt/nF/0en7qWOInWeNQTz5PNPIpfQPDNameXEs/xOPxdOzJkLJuiG3G+XXvlPPTjyNF1EGtAAddyH3UxcF9UAjG9a3d7jIzSa4tcJ1evPyJWlSX8DRxU3PXYYMphJWFSS9+xXDE9QHOADBAMwZFO1/WzvccMCDDLPpam5t3YDhc6qTzRTBQ86LMulHZ4M0e453ca2EACgP2xPeoNS+HSEDqo2w3EgtzcUkgpeOwuh8dDVzQXrzpd3PuSNWPEWwryFTAcR1v3e6NUghvzl95g9yQZUhHSm4jub/Tp38M2wqJDH4fSlaUti4niRUaBejQ/aatNCGqcplRusvp6B1DCJiEWVylKjPMX070/xufr+EKMM5p1FLirty6PPdIE0GfVR7tOjoj8sWVwgCqfbuQ0lzFnaqv5qGgFvBQEuL7PPx1cUxtVBxRBJ5VAu0eP5F646FnL09BGFK6KKiDIhhZAy7iLO5ee3NzcxoTLRC/goOVMOQAelJ7L45oemEjQyihDAQxpvq8eNCPfDCZTCezYQ1xQkerdFDOqSx75R/nS8jJaU0Mzcp0O5IwX6g1UzmcPV1XrNnsmXSj3CBhVEdByXX86FhMwYbtMjGmPIa0Bq73KWpkfljJM5uxRv9PF21F7ZjABgsdp3sSlA/ltulxEAJYM67cs5ZuJ1osNXNoqUbY0zTcQxPKHJZMrA6BSXNzGgfrO0OTUCG2FeccO2I4ydu6rBLEKVA2aZB/ClGNIs0dro+xyINFXMeQ1LdqFQmhjqOGI4rZyVsedIXtv2VcnyKewelH8+a74gjC+xx/HAC+u038LUPN6Qufh7GV8MYTY5y5IrhT91jtm0vdYxO4q/X1mqU/IaakSk68tVDWWA4XKxfwkL+3YKBNMBHZ+MPu91TNPXu4niue60O0FzyjbMGLZyeEHznalp5fSM6vBJFz2XvBKHng90a4EoHv+6/atFCQw3QJI+5sbeRBp8O/sUWZ02sioiZdR6bleyKaoag0cwQUvWP88g10HJoDlYybyEXMmKsYI1m+GSv17SbqhLCRmrP4JOShE/KFNKDkisNtGfzKCYKsj8DaCdpVOgyaEtlOMrmBoK/gC4Dzm9pW51AFJRUF06Tj2Uz06r7urYNPvVM2QfDqqptYBTvNFGkaJvbl3Q+IKbY8na2jc1bag2mkVbzZd4C0z7DVRTdxEGxNbvt5VWQGTEnIiIFrTRhFmD2HrYp1Fjw90epM5y7PgulSUznwHRP1U7q3w9KF8OlGcAiDdO2r7CZBVOKr+8VSON5Mzb2DwgLTdCSuPrl5Tvhx3foY2AaRToq2K7TZiW0Pidg4fd7ZHdGekX+9SW1l9s9g5CyvVas3G4PeIga0p9+3+2J3L4Z7yNhUjEUx9thDIOrKc5XNzefpUJ8qasyQ4o1r/ZaFpQ4HhcIuvUOUdLjM+7xzE+hvd+6Sk7QM7aRMWEZH3Sj3CLRuTNX0UcHovw0/BFTo8kdWGGgF/H1UWGxuuOw5FUXnLIKcKhP2mvtY5gm8Fi2zxzvjzCmfC3g1Vg/qU6A2+NmgO2z7Di0cG5rTDYLO6JHZThpby5FM84ZFpkEmxJNoEvkKiMEumSHSikC6vyu/NnV+CkQ42CBIasrivM269s7wCGwAISOimTawU6/ceMOe8LjAJdAovZnDSSKlNd0QxmQQfpYM2ogtQ6kWq1gPG1SBcwLpNFhNirEH8aF9j7BhHeK3fYbXl4kPORt2neshAP7obpHRIWYEja63O9ivOOdi765/Uz59njFlgaOFHK4nncsZR3gd4i0rj1LV/Mxgn/m9I1m04A+F8FrduP62a7DlFhsyYRouVe4/nXMVoniwI8yMGu21IN70xvwMMcPAkRcWVqkhCR6s1ErA079KW+U6vw2HbXxanhg4EkdXn7rmRxW3XWPm7exiMZMMA0XBUKCHt6I83IG55w/ua+vZei/9lqqOHZ4tpZobpfaA/mbkuCgt1dgFNDaqclRbpiiOAdmMgaCtIpo0Twf6o7+YIVV3XN2jZWd2qohCLAscZeQwsgPuoqOM80b6UbWY89JdHudVzZ2fyfm6hz7bUyBX/KOEsKOQ9+YViZHM6grc74yKmyEF3Zmz0bweKmrfpuctGszORlLfNkk+0BK/ChHoEcBpLucpIkRfqzzKYOQWTfOR+ttUPkkWjl4dmJikqYR19yw7y78crZD5iE66W43gxxXZPu27GrRRMP8tI/XDLfJ0kHGTEGG/NUfWwbHzXDz8GkPVm7PKfQexghwwSPq/hcbipG41pNqA5YKJPNs92WPHCRuRDAmRAB05zwxQf3Km8bqFRWDYpQQBqR42oMHUpKQ8FBJ3lO8SL8A64j96RH74RK2g4bcf4o/D1b6AYCk+lkJ/kFv1R5ePXZa5tuCi5ca1feXTunWxd3vuxSWfZVbUvSRwIwX93Eo3b4LrJszxYerQiSRyqE6n0RBCaIKo5PGmtp1KCb+ZLtwnK9k7oAalqB4EHCrw/VG4EMDZmBurXpH5qhhB9dmMsGVt+5XX3celUc5HSIxfHQeE9dboGAbKYLHyr1ptqBGt1EndAFtGF50mESOLf+7K8wO1tlIo3w0OlaTvbmWlEbFmFt87GguD7e73vsU5/aaZ0LDvRayColyCWmUL5OZwjlJ4sUofJ5ExTe/PKnnGuH4TwiwCrmrORzzCRx7OopM2R1Wh736xnr1Bbdf6yGETVuvG2u2Biw3kND1yqDg8lc5CnDbF/zWfGkX2NNzudgFr3Zd+Gu9kba4ihQUur7i4BTNT+UtVizzvVE8UDK8h8YXtTp/9wrKHABMjW8f5uExoPBERBLw77Ijh4ALcafnS06tT7u7lbD70gIb37sd0FG6HzmHv5zZIAK15DX0Nx5WqYmL0aStzfFIt16odlV8XSCRyRPx4z70umi/vQNt++iIanXOKeEd/O2n5e7oGNTa4/hlgol47y2G9sivU2XLGNyGTBlIejV7hbC01bGxJCFADr+eSZUODD2w7wlMoszsMsyAU4vE+M7M5u+Kyd5UlJxi6dP5CyhcX/MA8Jqo0K8fbbgGirYLnazzkZvKXoHhyVVXdwMtuUbE50aos4Vl/PzAwjaAbAbXKCc0Tx5zz2cWwPYz4Ad5uU1weIckMds/tVS0olCyBA5G+N6Z9WZljkn8qK+iFFkbvMh17g6tjgF0EKP+WgFLY17A7ac1wqIEfb49udyWpD33IWsPzpuc/VF2bPO4gXQ58EubSas14Y9b/AGbzmue+4nvM1PgaOO28H9lUHuSGLlLhn4xUDmOLg9hIe/9t0p/RmdyyzsWNchktw9+3c5OEQ3qGYR9SzukNcJvRIDX6htTPWncF7JlwUiydqXxd4bSxcUc+foV2icGcklBo4RBBeYv0fFt6PLOJY+NNETNSoPcB+u9/YXc4tMHFH0IaQNOWS6P27rHPT82lPUNKjoX/6lw1FpYFOjnC7zvztWU+YIMb2ppi3aDuUwKTn+exubb0dsdggTMCRoPWyXPAYg8V7CmiecS5n++dIB9qpjIVcjKFrt8QSWrTS6C/m6vWQCn6jQ68IpZs8YwPzsHIlVpbkgHPwiBa0/itWqcrM25Ra2HbBLI0Uk7Fo0y3dGO8RkyHDQca/paMGbu7iFGydsWk+fnUJxrY7zjPr6q5IKt+hniUzIS2fyh6II0i+DWkMZTRsRQVmosS4YoPbSvw29nGKm4Fd031nkzOyaWuN0wWXHtjnJO3yHrYdlakMNGP6BJxc1lAQO2zLraahwZOh8VYkn2HjfdK1XjxNNBPHO+6uE7YN+XmyWlXYzk4hXgtvBOkOtNV46H8ZJZjb4ipq0GhYFg/oNdq6SBACVsi2CMOWwlmrD66aXW65Rq+7i5sVAi5uloUknYFwKulizldlm+gAIGFvGTZZke4F5a1T9si7NuL9Rmm7x0t/UItfJHWBwoBXx7L+RSWuRaOf5wrBDRs6ICi/zDu5Mj7LM0PrCDDnLx1Q7568bkkvHvkEh1NTIAqbgx4z8t/b+lRFXMNIaWl1UVgjt5RgU0DBsJVnYeSsFrhz6VWbeSnH4OitPPxnGDoncWySsSPMDPpGV51t4NfZOGG0HqYwwmQV0vinExcbZG2qbUEilNvTdz4HliaOC1hn6Ggx83qauCf00bnuhgcsC8U3+3b/E3BDlz+21EnKe5IEC/vCDssFp4xon6z+XiUTuoudaZCdRYCZhNZY6zp8rU6fh0uUoFLXtST0nfqnYNKwPHiDhdNrr6rOnbjRGf4JzgyjBd0jtLux36FqogQDcYMgxQ2ePwMZ7WHVPPtpnmp2liRR9RD93poX61GUzL2zIGny4HaKj9vSdiZ0iLMfffw9QX2RiggfKYM3GR1OLAo31axeIbXsn9tDz2wMUbp7+pC+tRDFAXlcWbCnye0XxddgJEwJqW0lgRddczJoBXrG9HbuLJLkHkJEELWS0MFNsVx7ZkMMo9pkuIcK7bnq9MvEwqqksvys5N1GRtMwVpbA4NrLWR2zSWIQcCfWP2t4/zYBPwlYAUmf1hFJz/8jZW+yOJPvt+mu1fwi04imtNV6SU/n7beiMTeig290CHmo1YJQciHdrFlvs69R75MgoI3uHQ+BhXyR1en8Czgjjk5k2mhEvi3lsZaD4ZFPHxdkCttLh4FI1kL9ieHirESpDNPETT4xPaCglvwhO4z+e+l6FIi6Pz5bRiZt+zgdViyYpqh2U3DWFqkKx326kBUzGRakPh+IUPlhMWIweHHU6oaYfyt/HqXeKZToiYppKSMpTdQX0uEy9McGjNs8nrPgAXvG3uAdbQXNGwXmg3F9VAfIDJ4zZVaMI2/Tw2Xq8waY2V5p//R8p3a869abNEBvge0BZYNfDEBI5g6zHoAdfptG6NTxCzOk8zLRIZovAcubU1ej9VqAQRcpdzVtr2B2nVsRxJWgfW+dOorA7GZvWiQILCDqsNvo5tFv8PSUl/mZC93aP9tlz5BrTuFfURMBYNFODpmusIkGP7083wtFqerRhKdVWzm6jxKyzoY4Ry2uGwjuHkrE0/4mSNzXkCol1HwlJ3aBfdgm4fZ67wlhFSIII9j99KFvGJYFA7mlaWpTNMdlDVaxEgBIfh6v2F979Fr8Ma130liryRw18p8mU31zjy1sZXo5m1YLDo43WqFUHvQy8tzwiHTtmPMMAL9AQbQvUnFwcvX4ZYNdUT7DAkYfF1dVgQGMfC+Y+qHAgKxLqsSvur4m9q0IaNiSRWUOMzkmRBOnxftTg6vPbfa8dPZWN4jB8CQE6gADUFNWvxNrieZw0IN0jzcWtkVezoTS55imCj+9I7I/6h7nN03OmRS1BdsBCNE3tscGznC3lB79mKQy1Mvd/DsHYOSZRPv6h6o9tpJI89UiHsTz4gh6IbvRSt2RfuqWfQoUlBrwufVWS+zpIz+xHOkbNcdj9WTPMacKlSL7EbaWOhZhxRCEi9JJczsKGySLYfAhqTG8FiG4nvXhhWuLksD/EUTAn4jwDwo06l6zsQDLhX4fmELiTJX684mCwhImkO5sSGFpLxAV9c08n8XR8AKTP51DeKOqeC99mIqWc+HYKQsez2dzMI9T4myVv/1bKgPbRxD/wPYpWMNu/OayGgKMkQBiHUBLBtHW9KgVAnXQoS7CpSKZl9cMbJg/qKy4GLNVsX19NG1YUOIeWfPNeFuV2xvL3PICXvp2ht0mxme7nH5gaQ2i2VjmlV4HABZJeCwg9vUOcSngIldfYu8m/VjisXqvXSGTGw7mLil6EOCEeGnOjTwGLRef3wWioHAo6KNeiwIjR99AT8JdZj2E6ai9RjvC1PI9Qa5pqr/1goAThdQ+I6q4pitL3VlRdlC1+dNl/ypKDIV7iMMu2AKGROesASKezVxFy01cfzaA1puh9XMDq0xruKNjcuSgK0O+dRmFaQ14KY1W/6HM3fs5E7Um7OAdYW7UCzOUBWpsHt1BdEi14W5iVXKdqSmaIj1WThqdpXWzPmTW2mvSIozAPjN62EmqoYFl7Ck6iPe6bGOtvIep6HeVKfvVLCcft3NmAwqlT/bcXZR0ZGELHyDnDHxZ6807lg26O6SVAvq4fdczYblARaTBie6+HTTfn+o6rgx80EuhxZ6a+Q2nGS7iLLJeulXVQZjU4Z6UwwkUulCwY/I2O+uAP6CYuTVLswgLouaoBVksqR09BJGRwDmNn2+bfNzT4vwijKRTpvWZrRC94RwxrIDmqyiFCCJahcrxKg4/31FxJJDnaNbG3Al4joxbpWg6daI5yrmkCD3f3OKbPylbpj5dtQBJCSX/cAipThf++cah/R/n9ol4Bz38TrVX25eP8PEzt88dk4vTs66i7RZT9CB+Q92iZ+TFcRLi3gjeX95JVw2PqtSjNbJLwIgzFA0wMZyzGuFE2knSr3Q+fl3QoUgOPpkiDcVEsrg2yDV3OFa/1aT69EZMRANA3cfb+jde1scaOUdCJvSD5dKxyumxFEBAlarQJ85lGX3pYXSqAq6Pszg3dFFAG9SnLLubbL7oeLOemW95Nx4oxcgJnrEagoBYjC8B+8sx6ex83coULzOtu+WN0x2nsUEhRhERK+H4CUuSpItL+t91fPthTLlzNk10FDeOO/qbZW9VLwcxRiK+DVBPGrX4awpPwyyAjAElHVmVkn1AMkRLlf8K+YHXN6tiN6/uuPL0wp8DqVr/7+oIkMtBVIIGG6PsIQQoUwA8cW5HUxrddUaXG6IIfCpY2VpIc6sZBj0cPjbwFz0iVMJ4YUPZghxoDvD34EcJNB3pFloU2nKEGtoO1rmSQ51Y4mBT1jJp3XFRFqZAGhZhWJlWZDUmYpT6NRl5xu0SgVJPT332jlIkXptNwz+h+rJjLSEkTHTrDzfO9zKFd/cruXNpd7xvobxazTiS75Y3idFuRecGUEEeR7m9kEgMcM0ZjfP6JazBgAPxEu/P5A5Ik7m3AKFGF3n3OoKvzzGvN+Yy8lPzExizEOKjYlsqJefVEKj7yWFNSrWRRc/pEKV+F3dta1w/h1HU7dvV89DHfMLP2kVI7rtS1u0/kM8DGVVqlDJYEgq+orAK3dTc2a3Vu9c+PO5bEYHbMGpmOzG88+GHaGqC1muoXGNNjAtxycm69NuglN8d2JNYseZcaiU+EGKSkFmL5pYt4UaW5OURV2myO8zmJOvQyBL3xh5J+aRx6tRfNthEHrlRYt1TabErTHrrjw9GzB+uXnnxIWrf+ln1kxtkyZCCVhGxa6WG2cY2lXb1O0CCUReCrOz/UNAVdvp9jh+1sOutjE/dHvW+jzOrMM6tBl+yqvpjnI37yG31bI88xMB4sJyE06hY2a51YWfxePZ5kvgevtxLelR48ttxVBcAReJRlSh3sFOfgj97aaxVYSBiDq+YHPDAKaMEEgVsd1psoI2p6cBGTTiStmiWTYWVmqTUwq+RH/ihKCQHZlkuH0Fduux88RPNxHJClMCYTmQnJGCYWzON94UoL5jRWH1WKYcKjvAhyBm9j4WbV1N/OpDKNDywYvK4fwTT4eEpApWB9a745goQRku7Q6kyxFPu05Ym20EMmrr8bpxMaKj4xQwXPAvk2zRWavcgtxVLImBp+J3Vy81lebx1RSeiZ1VINP5y6k354c+k9wKTpuD2cZF6ogu0rBJH4fYTCzvUWB5y+mkfvJAKgfipIA8xCkD0WXHRm4CnpaHVCy/TNTMkvP5EFsyNVfNHiZfPSr7FEK6sqC8c5dOKXiRBcNfgr72eWIYxRKOE01GkSJDaVcPvAeCYPVtTSX5AmWOAJ0BXZmsay2an+wc3HlSObn+GvL+FGB5ETIw7SDJtRkuQcwrIsQ1lTVPwqqjLjgqs9vliRRyp/kMngwlHV3mWwmelHJ6yGhWttNB9VxjLNKl8t2gQEvcdPkMj6RV69g1d/+Oz+h4Zysgx83vJr+y1aLEtkR6Y9ppHrOVpa9LUn7mBmZ9OEQuDFv0JPIHYLRtteOD98wSoQC9FrjJeWPK6QC3PHLLLBmyvgSdjYjy4m5Cd45BVDqIrw/3/3lZ95EifKvSx6YwYy+Sm2KHrkq1QTftMZvn6IRTEQbjVga0alL/tE8gRGUorrbVkfL3sluowIXxeE/cBMcEsy7N+woNcNAGAN4zAYQHO1eTgrcY3GRD32etxNEAPqSt6Oz0xQY3z4GZaRKi7M27bI/65oQEavHIIkUJelZfqNrcQRLGOkuajNHc+QH2SIXzjBvMQyzTG1Hfc6UlblkBiytOo3qnzhym6woiSkDNzqtXp/9N7rKicM8icQOQygDYm9IsBzW3L8u6424uirCuYy4CjB2x1Q0KCCjdvZpq+m1HG7oLXOzUDuqmaJEar3vimvs6xQHoOb/Cnf7pjWhl3ffYye8LeUuPtovDBgYA8RDmGzhy5KiNpdcislZufDrnLJ1gkAOUF2GxE4CHWQa3zuNC+KVTgrrj59O74qixT/afRIGvKjNJtEiskiMMgWmh0tDcApUfbER+7V9MIShOxz7thiqn8Gld+MYgPLybvPrDN9SwE4kadGmlXI0Egr/A5HiL7mxGBxTnptBSHY7VyvPyFCuvMggVugR+K32MTVzERQF6aQtbUNovRK0/LcTFbsvyKzqX0ihzBmgvprqZD5wdQtMROTHCJcowVYu9400N21pxqjQb0SarHVpBZb8V3xcrulMcIitkEdJJG2A2D3blR6l1229laoTb390GHk0Bbppo4IOxO5+ibbR3HjdVgv/HgDpZWaNTt+lW/dQzp6YtETkJQpSVwZ420WuKKuHO+aaCzFeLdA8J/4+eX0kATdhpmy87K/V8PLZ8SqYWA9UXZz7jK71YWE7s92E5ogDhC3VnY4JlgKybeuMHPQRESMnPA1CDgBmv6M9D5cfy68FvC4QWCl2gj57zv6oGHQZ9+uSARZISNdqU99+NxA0+B05H7TAvGFEFHOBp+QCiG3KpYJuFaqDS685CGua2j29ZUFl6a3eZanhCEb87gljk5EJfdgLz3nArLPMswkr1u1nQMYF38PNnIQNtKdr6aNWJmeTwtOKuPMLzUQzdpy4+1REXAOrr0talVZLmG8PR3+xSpLFuV8/mREGy7fGRPT8YpBLtcwwmdT8dUwpCGc6fqnTJiSp/XKTvvM9+tmXShRYgjZm/ZqBi+nK7pX9JN8P+POR4WQFZjKUeCOt7F69OFw2c/icrPKTgulUA1oZaPm+CpCcRma1TbbcFXIK2xhgQyN1LvTRwah3YXAinxtX5GcGXN5sHXtx/iqjohUnOEBJCsSieJxvRP+1jMURE6HmmfES6ZpcN/BkPdpyRPdUEv9DqknYxyklfHROXaJn7AYK/XORDPCAP+q6NwLvgQwGXqkBFtC1eMbj4GSfsoa/OINEDP6A2gKHKcluuAfyNBZrVSW1TVOG3+1bWoh3hksjtSzxQ7nKTL0ofbkSg5K8lHBDrGT2YGqws/FOfAjg5BMnXJ1jsLsQ3UyhE+X8T5JMsdfcx2ZasPHWxOtkw/zO/2M2g/Em+3M5VTb6uJIqX5htPt1Ya7OPDLYqPBjFzc2V9319fNZeEz1iKIyiVqpE4AzjL+NT9pH/bMJfLT4WOk6FS9cj2Ib3eCpVsMyJ+0Or/lwiHXdSgLlqw9UaBKzkQeccbV+M5yTfP+CgSHHiNz+JVg1HeURicEqJOxQPPPc03u78n4M8FYSTotnake8J+X/weDwSUZ/c1KUJO53yEIjMIntzeYTHnZ7s64TtHh5+kiyZCQmyPU6Yb2XBJsg+K956+XV1IxfvGCIUHd5gcrTEW4m8yd807lNyI0pqv916diTuDCNPu0+dD1LsTwMMKK66xockppCpn6Gc/zhgKJ/ykrusT0WuDhDPc+j0xWAYeL3FERoOfiUFx+wo/p4D1lHPYjT1594rMvHLFNtA9uQrOV5oar5bz32UqHlZEBABoV5lJD70kleKUq57kYC1DVMB1X20ZQm9uzIkECPTOzUYj6nIncRewBo5el4td1Vi+MzUhjvKtTdA+x7OlqmegnLbw5xjRQ2N6v0/Qj60SJhC0uPPWcKpWraFJKQfCPAfLw1e3t9lCfmwoTfVu+jo/oANGnbUiH6Eo73+Jva9sEadZ7zmNUzcJJ7jpV1p8Qav+x4e40bvmWhUboxeE//qjSWCYp4Y/L83UijicjyjQcd1a3tnoaNr8o6Mfd0f6RhjofEA+Ox0Z26D417P6yuq7QVUqiYDEdS3d/RbLCfvsDaU4pPNcwPc7gFKa+/Inie8YpU61eqB6yUoxXarr0ynXkdSuNns6BuLgTQQCqUtoxPk90bj/KJ/MlLGSOJDYIaUnHq6ZDK9W/2Xl9sH5BmMefQlY7MbsRfbWWAUojmtc2EVIRBOx2ZQbfL9VC8PyUGiFK4h/fO6BuY/X9eaIFdHk5bUqTxrVLvhZ0Ggi6norZlt7l1z/KnKYbPGZJhcEqeQAAr9J1ku1bqaUYsk74WsnByuzfIY1HXQfaj5r0C6nQQ2cLLPqve3OqKzoLucrIzzlKYFqCK1q4lgGoaDcvIYCrZ+ffrsw1HL1bkoP2yvAN/HzB+wH6SN0SZtsTriOxMO0fZ97z75l+IfxH4kLCq15b2l3zj58N/oLQ4kUG40VbdhcUYMw5MMibdy1EJ01TQRbZvqhQCh+teMda6N/YrJzQYIxAqsUiv6cSeQyH+Ow5D+78+ATzGQBR1ZIMPQR+cIXrO85hmwYgJmIvdqUEg+IfJ+Ox1Iwp+HWSwBBFoqSBHpHIbX9lVlru6c6IktAGBo7+7X6pQLD8JMR/lD3uLFBX5fAdj6U+cOsZSKkjdnQ2YBACseboL1mdqP4WzvHOxcKeSGLWUeTr3/LIA7624oMv0RaAEQ+PZUMI9h+MTeAEep0F4aJgQPhgnAA/Sbq0lizUrYS3bqV8Z1aH5DkYSlqR41NODhtUJHOJPEq36FnWoxjDgA1wfJ0lTYrivab7pYkQFn4Vc8ZwdRb4KjNwD+bga3lPca3eALLyWW1nW0W/pfZ4qBPVI3K0tbcxi5yy9QWHXS60/A2BgMOgu+xIfs0UrgZSOx3vaoiZc8yqKtDgBgy1p90RyY34CzalNXjmsuaPn1173z/dIvJpymysnrDwqcNPf/LDRSYbe5xeFIRW602Esz7neGWQnQgNJ8oKW34ORP43exHLJkYkPSdVf05egJ6iBue/0k1LiwlZSaItuDymMps8Wkky09co0kghP1tIFuruOHKq1/zPlvs8pb9AJLmdtCrQPLx5bfaOeI9KbRFYY35eTri1s0i/rClVEvA8K1tNRyIVgIP0gfk8Sj2tUB5lbFY25s3OY9XzxNRBb6TnK4IeSjkxAjtDVieyhU2CTQjtvUYgYPCr71puFSbne0J22x5JLawjPzo8oE3GugkZl8jD9s12ixHo7eKDayRgh0BgI6jSyqJfi3vBHlo8DHMGrMiPGmjKIErz2tWLLWnmYYqJhXIftH5jX7eb4w7eDRV56qrbcxSftxs0mvM2LZ4SSwZawE/gsCmnHGPjxARxbBvSjeVfvf1c7wz2pNiRObVzHnFpHqOOvansArTNC4fD1EF1aFoq+DmSRGv8OcExlME39APhH7p0ECIE+6FnSkF2R63QSAsD8oboTIIhWf6XoR2qvNMzbZIVfA2PGP71boNY30iavPwiOgaz9Q0DeRCgLQdtam1tRXoRNXcOZu7mtISY1P/OghjnqMFgfJnzpF9eG/IOPYfj8DUoPQ+awxZ0P9+CVbqY2l8QeEbpLUpvjQ5IAmPQySfKT/G63SFxg9kWfW71vfy4QnVjIGby5Q8t+SuObgqS8gHZ1NhRXvXXctwyLJlHA4Hj11B8UmLNCUHaAY7Bw/wRQ+NVYIO2dYGrZWBb9cP+Fab5IiMUTUAiH2GD4GkcTnTBWNC3/2ay44o0jWDM9w8oTZdkm0TtuAK3lPwyAYWWAGXSivG9cYRCnMvvEYZcL4b9F6dBVccBp7Ziq/E6sgXz0crNGGhTRU+kDEbv1du0P/jBlXJbYeDSKoyXyTKIpxyUd73SzuknAPPif3r7glLxYjs/UdVBl/4v49Cf72OvUuyF2RkCMBo/5C/JXfQuqROzKDOqQUYeqJS5RsPe5nQr6arULn1XOaYwz8M4+HlHbf6++zXGrTsUU11nEYhV2+GKnmGZy2CkJkM9caoQ79U+6JPpp+achwYoKfH1icWosR4L+AL0ucuNlARtdLnR2tJDaPxIOlGwzKWWoIUXPMR9bkFejIhT5dO89z4lpSQAPK/+r0WqETTYShGVOtDBxk14pAEFskCaKX9NJNe5wKFTBHONshd0ZlmrK/ojFzkh/zAER7J7y0BF64TgSDBBoyL7fR7VNIkEEeg1OI0UP/Jh8ulI32L//V9RbhLbB/IEH/np7MYamJ3dUMKZFTZu1mR3ECeXuvf70Qfg/whld9F6b3KEfo2V4Vdmslspfq1lyOYC1JfEZuFqzjRDXEUOMSGWSR+vhjOtDCGEw6WG6ju8g/dXqmLIoAtROlsYJ1CPFml3AQQDwewzqFpExdNJDNnffr6GVEbEoL/LFOTeLLXbkNmcpiTpg9o68rO2VQoqr2y1QiWDc24WLp2E8KXkooLkAoYpUYFTAXfICmpUnDefnyOrjPUZcfB/OiuTGhIeGC1YsqfcKEni2oBvFtUWl+JtgSx4/1HgmI5OL2C0Gtx2oSubl3QYbsYIcj2bH9AFkQPd/entaeOAf9Na1ZLrauv7FQrf+m5y5NHXMUj66hr1a6MBquxKYxMeftmojbfOIDiPscJ1U2tGSSFPcf+wmMMBhER6XnYBNp0ekQOtZpcqZ2lPC1zvf79CrSExHxwGw3avItvYpVKT1IivYB14yEvR+GVoB00FPLD4vDRnlWxRNW1+N6MTxmy75CbbDHJNVOpd/bP3ye+Dcl/ahOZAv1czL5+0lAzQS+/2EGrg+wO/eD5u85N9NgGCmILDtPUoBFOQZnr6qhpME7ld7Mx5HOtwC4HC9GCC8FwHXs5Dv6wRmU4kcLrGjUL6DUS7XFc7tSTbV58nCKjWoz18saYnBo37RR3Bl2UwMQCK9uxCuyYx5m32xvQXAiLvc2ggenE4SUlSS4mf20mh7YXF9Tt/ym8uWzqApJRqIf2/+00c3KGag6ff0S5zagsBtsiQwtfFAMXytNO+gg9hPy2UPYtnHsDqBS6/F6MJR43Gff3AuSeY/2P3woRD2r8HGeuUjU2g5q2yMuk6Uv2EZdDYypLJQ5uGuL+fjYutzlbZe1Hbgj1vbVZlhM6FzPjFAhWyVAFItC5byeRlt8kfG8diTMZCK6lqBJhftaXfC+6oIbYZcG4Vy5kwQptPkaExkDvePl0uYX61c7VVVqOBoqp4eX9Un7UhNCwKfBjT9UCInz6699+piAxOkwNimwPL+7Cv3ur5duEQOHdlj1RwgXWQeHppkzk9X73QLr3Vpu6FFPwUh96vmY9htrYJx+YAqkPYhX0i61mxV6zQAnE1f5Ui1o0FTbRL9uHs1B9QNJ2v3oTzNQHRS3m6qpDnmecvUS6sR+Zc75b0R2mFEnAtvP2dhZZ0+0ct6wyRAjCfNwRHhGkNk+Sa+Ynv1NlBUL0HEjnAE5v8aH9EfT9ulUQnOtDnRbUd84tBQbfAaCY1UYTZO0wwnnaBqRNq6kZBdqK2I/Yqh2iKdhbhJ0kCDQEUCeUR3vAh4aGpgW1Z45UjyWCS0jQ3GPzR9PyT8Rlhg1wWj9NDzx21JJ4VnVsn9/2ELz/3ljd8bJpG4EOOP0wW7Hl0OBV6zdrtuClrNQBczEv6tXiIoSsUmt7pkA7EcWGdFmx6Y968l/CXP8R1jTYEJ34hkHzyNh5aNAPNqt9qAVNr4IDNyMmNK3ZMGb6rmy09nYmHppXE/KRK2xdFd+DHXY4nwA4tum6ZjeKlI2t3ZcLNAu6AicZdeL8QF1oTQuyWZNVSffQW/5WaW/KEqUXXmiI8GFRbRPIaAcy6cc3PkSuJpeUzlSCe/7z1Vol1ZjQjmsQsadqVkdrL3SC95wGyamyZDruUt0yhtja0A80kn/UuKH8yk7UujgC7XQY4x8W0ka/KonBWUxg10svrSw0UaN1RaX1nabUpMAHGRU23dAxZa9g5Ts+l8QtoOAGZCwktFJgB9WErF5djWQ7bRv0WYURY0VyIep/8eBHHKoHeQO6eiLsjK4DD5WoJfvMOn3X3OQxAa9vM9Fk5otoksCahww7+O3JYkV5EHIDm5q4uxC2KrPbmrsGkwu4alMRjofhST3jWL+YcXMW0VauvLr5pMLeggBX9Ez3JNgY03Pq3vkW8XWcOQWcjsUIP+ZdTZnHa1cP8PNnRyWg+p2LK0ZUbTgolWJuPqLUhl4EdWRkSx1n5ZvRDPzpFBnk2+lGakornlgLp3nCsmfXUVMQ5L6aichWSIqelDRVx94RD+e25RRYYI6WTbUCHZVWAl3DU7y0LomR8M+Ves20ziglqEu29EdZ3mLzSUmjWw5ceD5MyUfNGAkeDaP6F/n+SNInZr85KSB9gIshaUzqMmiDppA0xWKGtfSlYKGYXF4uY3h7IWNEtodLdCqwcQK4ZbMYaQ4cL7TuOyONi4dKnQAphHHCwAeONNYQhBNluaZxpEHD3yMkgG7rqXkuDGPv93V2Hk4MWMCcKWq2a24XpswepFwDkDUDt/djKCcoKRo0zJgR/EOrWH+mR8RgFxtCxwwKTi9pYQri46H50mW5bIlymu+tukogHt/e8YLhr11MhbPM8xYbDE1VIPSiSTIvzH1p2r38MFxZODJ93LDjkVrVa22dMjPs5/nbQpDDOynKCBQn9P+Phs9KtqPFsktj0H5hHPIeiQeiPoguQP3uJCiDPg814V70nWlMF5le/pnd1D8qkC5n8M7ViEvM8l+tsEez+VxdZwaKGO5zrNTXLrCc/tFW7ROgvJs3wtNv6M0qAPHPo9+Y2YsTxj6X4DpF5VcwDqghlSUEgtVVGJXPrjhBmbZ47MKTjuQ3voZjFQNinZpwjDcdp3fwPVMLbIGAoWuF0rFHkhuSKzebgiUS3n6R7slUdGaP0GFrv7dArmvR23CIrYvwi6UunQUUFhBMpkVeWJk5oPcxOSsMpdyml8VrQOxJPM0dUS44KlUBL4NeVsltZTjb8YWyTazp9cG/CjJbbh95nJLYWJ5sgUdHVV4x6dsF270ZJIVqCHDlLRx54gcEc+UMgf8zSIjkVbYFJZHH6H6PzNyGj0LK8c8QMZskgW+FwCj9BwD4v1i7D2EJGIa8X+1FGtLqQ/rqZCer1NTAgZ45pF9CAH9qUmOi4GUB1MvYV/Sric3UTV2l1RbFKbld9SEEyTQyaFZt9BpqfZlmis3teNlCrENskrDJ0q4ABepqlnf0nLUuvoWna2FBsUbN4FXU7jwP99pGW0t5EEYy+jgq+Roq9ZzYPaJUnQAcbTdXVqAd43xuoSm6saaRbDmoRpMlDWH+8xou9K6y21zVYbjSOnes5wnEFFKab0E67WeV4YWjF1jpI3eUUUwjDz9IxMWDMVVlb+6/GwaaP4t3M40qAX0Oqbq8kFmg+KAB8xjmDr46QJ9GfuQsxHwOsY5YAf8WEMTfsTq4Ms+6QTfpE2iRgtqoWG8laxe73SzJHHaSm3fGr7v2RqFMcqU8ay3yMBDYITHV7LpditEA+Bxw/8yI4bI/kdeV2Qy+DRDE2ySfN9VXg4tkDAc1dTzLAPYyDE3kIXgPf+fuJQ5G05JOK4RZvsq9nJ0gj/7E8QOPz6Hb5TTGyh+Wf498Yx4lepXdFtTSvSc0q8nhL9pidC/v7BFHlHOZv4ixfuuL3tWs8LQc7+BPxUzFCXy9dgVT23B62Y/g1loxjEVZvoWE6W8tgSnr+IP+zOm7Kzw27dx1H6UvPdBvAG+la7bUf9VBQiPg/ipEkvn9XJbUPvZyFFkjjgYkaTohBADtZk+IQEvmK2CbUiYBxizK7UmIl1NLOcH54BxkNU+mUmGFzhy481UNA+F8moE+39/5JWIrZCJFFB5LZkwGIVImW/EQ1rB9LjfK68I9EtsMOYiL1GFEJkkKF0YY3457GpKw95a5oLs9yxyRirvbJE1zUL/0jRvwZHHVgcn3dCTtvr4W5CiGHkxeNBO8R8Ok2DMB7NmCPglsqAx73FqAuq3cIT0UnvIPr5x6plaSi3hWqkLhq0I5CgkGQ3bIk8rXvEOPQSGOu9lyj0PLpRFHWFGwfeSfBLil5F+D+c/PlwRYOv7ZkG4kdx2VnWv8FvPDiTojA3rhfL7puSDAoR43+c44OQnMdTssOxaMTFBfJ6ldARXwAipT6cLV87SfrfXAHHzy0/EjRA6wCjp1DTZc237rVFiby9d9NP4fJDksjT0CoxqJ8mVhpCXOCElJzbrfFjC+vUDr9EoujqQfD4jmQ0TQusPYYebTJ9H/l+dPk2Wtiqg5nupEf+qKrMpeX7zW7nF5AjlGqwi4rKqPwSCkzFLvy/cawJx1RVwHoB6K0XqJiAJRuOSWoqxMHcXywlLYwejuacPssZiFMASBzYwKyg9Hex3guFr558MdVhVOp4Pt65fCim1dJpwAyYvuUMXSXHy4KQn6+G2Q/ns/CFi6CqHPP9VsmuTe2ukm3jpI/rTUy39GH049voG2V2nRR9SluYffjWWDbdJdwHSB45eccuoPT4e3tQDg+RPufEnCdkH8o8rn+lfi4moJaB4YftTNEWKuFt2ZL4dEyCT4hqz9Pxr1l0Mtd1+aq4KhhZQr821B/uHwmLwJBoBRDOumdiaxnN3f98hMHlkVFnkS2c0YTrTGhapYIGl2jbyHrcTnNPxaza+0I8ww9BchqHV0DW8jOHed7WM9hV12t4I8baRMrhtVTOlOt8VlCwrKb6Ny9QoGQ5tOkNsVsOu5hm/A/00GQFef0dM+p7ieCHmFf4bqK4mt8OHKokkuvcpjhvC/N45GLfAkf6bAfo5a3Ni0EjGnLokjFCL3vatkE8DdEAgM73l8552Fb734/PjYYI9dkzVZbc3EE6Sq2uz9flIR3J9kBnI8MDRCtlLLP08h7Goe80wDUtUniG8I4c7bauPPqPKIkRqQ5LQOc/Kwt/VWG2g3PKDPZiUZ3gTsTltDeEw0Gzxcm4pxLt7E6UQhNkHssM/DI91b41YQRYERl3qjFAMA9dhalKXFXtF5C/lUkFtNj5m/p2+G7gRjMhYKPifwyMwfesYYHURpZtd/96301FF2VEFyid5yVlam3ir4ltd88y+oIVdM70hXiOuTthaDm9x+mKcV6CeuHw7NY0A1zyhSwRkNLjOvskxcWk+FmAxXoZU6df1Yj7djkBUjzgvlBevBPGh4gUj9sQp83TAZbIhvERARp23ll9pkCauguK4c1bnR0EK/sQ3ipkSBN2l2NlUrOGWGZ+Vd4cBB4bqG37o/ZCucMO6SZBKLUl/vMZUQCAKm4KSj39bMETAiZJ88hZEk1SzxVOEE0D5m3yyMMVc1L971SWdW7Q3jOzKBIdbqrL47WMu50stwR8ptV7DUg/1S89i1D3YSwkQibqXdBxzGsZNSrFSS2WzcgkapBQEhoL63Ip4C48TxJqNchU8HS7EoAfM46iwCQQCcyzjUTTom7mscYRcVr7MDge/36wl0r/N7Yz2a6/JoPakBDaEFa45VFG8gZ5nwUH0gvz4ET+ywTznITD5GXnIFfVB7IQ3QV2WOJ0C6Ia46qrDv2ohD5tJU5ZfbjkqfqIqLocvJeSrUzr6cZA95f7ghTRdHBgWhO8S65s0HSnfXkQsjtNQk0hCgVPtUvOG7v6dS9lChbYjBzO08QDIkZ3YJE4/hdA1xPJ5lH9Toe8o3ALQHCdptMsOSHlhS9YTuAT3Wow+ICZ9j+LFMOBb6poA/P4Rniyeiz15gh2tTBEEM36NoV38qEl6IcvNdA8IyzkWxceuhQ324U0E2fNyvUUHTDF1/8rjXHHrC8PPWVbqPdrz/fWT3P7rNMH6dwX47aIkwFjZuY0+6v5lNxGHUlHklHSVxo5U3nAprdJQ9RRADmoL98PgjHAaF6ADaqRcfZPBsETdsDSmjbHQXNQvEaYw+y6FH8BeMhEypnvX6nJw6dmAuCrMYHOlQrcUbv1fV4ZYss4r4QmwsD6bYnLa002Z+KFfiJBZ1LyFP54yXQMA6qgLMO71Rsg5SShwLoaitBogioj2yV0fGamfTYEedXgfSvYv33YnsmDt1xUD7/eqhp/K+Wtu7jfmzIB2Tmfv/85APTz6OMiHE5NuvSMMGzEmHHhDYHfAXHoGp0RMzZyih6Xm5ITBq+5hpwGIK2MvNyzNU5nBBz2ryhVExcEe8PkieEvi+xTh3gLTTJYTvtoYllq5DoAXdTlo7jwv6K6iPGmdTGC8lF+FgHhz56yksLN4mb7hN6wKg4vPW54bGDVmU+xTq3+AdRk5oG6on0yIoVUldFoeJawQ6OeDfLZ+5L2UFRKZBgxElD5t2dC3lCX2bcwlUKt/G8wNNqvWEB4IHO2YReXDvNtM0NW+Cy3jdS51JPfcp3Tzr/o6AUDrDjMEmvpEwcmEbg5o9xHAepC6OueRLif7qsl9AcgemUw9rDiZM6MDQj1fdCaLfFbG27L70Ft5Zsx9X3YsT3Rs7wsVwIJMGPxULoF2o1JbgSny3IRVBHBQ1bOAqRAUKBLhdwSSty2WSxgMVlmKxsYqZQuvP7YUd19q6j6SEsKpnwyElqRc+8gpCB3x3NCUrSeenh1ZzRjMPe524n/KANzZ3xcU2/jP6Emsjrem7e+FQ1LXnNijSOAwzCYRoZNwOtKSooko1C0tzqhf84RSvCrUoH/6ORut4wv8k/h7jsR8Wj7/joiIE5AaPmlSunNGuy4+Gph6jqHmgchvHODaCRTRrdB8d/6vdHL/7loBGQNlN8qwPz9w02hXKRWNlRCRFbFbWzYY1zhmWu9icgiLs2cg+43v5GOBYKmPqoNXGsf8owUIQe17K+Tet8MM9wG6PRwyjJxWzF4cP/rSdiB0v//8DamtGyxiu//NVeBzSOXY0XU5vdwVj/VTV+Tut4c2qiG2dbIHUbrta9Gm+HXWpoGXq4W7XTL9NoE7oKUaQsOaFwnjkXdSFW+LnCRUMLCten6pgd2aubnooFnz+djpKTnJ0bw4NQTR/GxzngWghMeot5WP2ZXSw3WTt3/cwUykzr4JlsKOrGp6MWuSok9ifNgSXABmJ+AB32M0mU3VaPElgSXTCY8eNgwtlj9qfjpQvRnJ6ywlzuyapxbwvBwXPUx+qQ61lJTOdyy1D8w3+V8PcJ6KV6PvFS6O2QB7sUM5SczR/xl4BdxGJTcIR57i0FcyoTcBErfqooGVoLn8YkYZ1yhTZ0/qKRTdu4t8sdBST0Oc0jssB0c18gCX+UFIj8phOHo1qLV01pNZVyNIaklBabwaKMxYLiNY+KiVkgJi4nTfr8btjV/qpCpdBVMww1iK9Ec9oDonGS4971Ek1C2ID1UkCi6qGNvM6cb7QPyOqmP9ODpmTnAakPzCxB9GGNK7/qD4cE3HxD5lnCozsNb/JbuQsJW9PFT4XKp5g0it3P8X5B64VmC+5cleGd78ybpymLb4vxuhSPjV1dgqhi2nH53I7EYspPrjYNhQzzomg3br69599cGopUNxgFO6MKXPlg1mjoZX9T/mHxPH1Ve8iyuemh1Yf5mV/DvCsfJMUK8/EDNDiOkLpvQpYuqNqM+Dfbnhw6KW5wq8rDiOcyhC950DrFOhK6ZeM/ZuZT8Ofe2rcQOoXbBOM+n8+5RztGdJLNCTwVIotCKaA5/bI1tpldcaoShRlzBvYcAEK025SH+FgW6nFR60GRYGBYljw/Q2qsF6cQbGrX1A7GPHBKPdkl9l7yL8gqzu/Vd9Zh7EaUx1Ol6Vjmfn1DRHyY34b/5wjVIDhEaOcsq4GKXKbY+TLl5pFxtkzJ3MntVZQkG2WOYYXy8jFbfyiTimI6o1JKN5BXQFs27tbiB1CnHESv6RwGWFeLuVyRWEOclAh3aKhpNA7Htqi1HXvq+67H+8jxGQvlv8YedkJFiSxycNXG7EbC+nQ/9njLmvmdwn7qgHxql3dvbtFqdZxNbF6mukrnUDl4PMiOke00k8VsZjMTHaKGATbHwXDsg4Z7Yg/xTtQRl2aIQYaNFpU8oxwdeY8lCRJJ5693WGeAChvNxUTVHBqOfPYmwBbfy+vouPCwSy8uRsfJqR8YxAIXZlkpNYbe6yZ0Y/FW+A6dMDx4AACWuhNktq7xAkBWT/ZMFK+84Ps5g9cWJ+oiqM77JNmJddP1sTLDKkp6W4sJTdJmeAqzNvSIKUd9/GCnrqESqDsOJjeUsTnzhSTIWha1rPToFbFQlZi3A/L+H8j/455Bt4nZ8uhe8Iz85LhYmpDfCkEpEojRah96vM2bzrrZOH0dP6EHShBw81FfUkBgXSVrHc5RubzwnPSRHCAfzajSYJSW/Hc2DuQDeq51bW4pU8BbvMc1ph4ahINntuRwRNR3ZPEuaI8Oap0IY92XV6mJoNjvH+sSsyV44wZ6GmbDrM0pdC0OgpTKoP09wl9OWKnE3aFm8SrCKWmGAbK3YLyHStkzQZRb03YV6le+m7MwO5tzVEpjYmtvmmqfufAtlq5nxxsFykMNGGelGhjtqYwgfljIW20zTyUp+ZPGXq4LKlvPYETL1YA/sURU6dnym+dDYVjQnWhphObhgkuYQlyWQrEZaJHrv4MsMiqD4XOnaFhgHKqo3ny/6cB87TGMdupTdwBiA/OjyiKlFDSk2m8Rib5dw94Ib/fXQWSuzqxrZr947E33HtNYBanP4HTziD8T6i3Vo68YhH3PYfEGZPzMpk7TPxqISGxXghIN+pTMmZlUJ8M40K4V3yS3sGjL7QNzl0SxgECs3MrVegnWliMCtVqR6QTM9vITYqRPavDPUaMUMRyl/fCV03JqKfqorTjaUdRhJWFHZuDOyf0Czb8QNVTBC+dYnFFkLGMC6Z9h5XFSKtBtW4dpCNqNz/sqXneTdQ7YWjJb1lm+S6UueGKYh8W0vQx8yU3ZDDYXreS/tRv1uw0zIU6KsA5Xk36nhXJoJv+YnuxjXe4a4J2d4ss+AhL371MgcTvwFsE1+N+9tsZmjgc7DIjQsQ1+J9VqipRABe5wec5pwgr++FPOnUSj5aAk2CqsNZxUF4ZvdbmgZfr8mf+RYG6RSnW3Yh1Ig20wowf3mxJKhBZn3c8yVD/fQcoKcuN9JZaitH/sPplqE6ff/JvT9amTTAIxPzpdBLlCkbaXa5O3s/PySXohBrZ7ExqIgLY+PsP0Ln9GdSr6/vTVq4CZrqDjJrSJau+NROqdIehoV99A3sCzC48O/ItseRKEBPPfTj2PAFyrExyNRlGvRU1h3CWt4yjnBroIMRt/ZOHG5aWzZLXip8pJ/JmC7Y5OOhU3JKr8lvGCTTkfKHxIc8+a1DoAvo8zKRgmx2WnxSpCtmtEkkRws2mS8y1VsBn95rPQAqgKcLwx3tFvtbGr2G1g3yMw3lEHYm5z7HBGVskfWtguR1GcJDVkx0t/Z8AZYNHVBPecWhxqiEq//bJ62tano2NFtGVb9taLDpeHl+ekaFRmte4Z/LiVzedodV3VEGNaJgn2Aq2g62k=
`pragma protect end_data_block
`pragma protect digest_block
f3d8b127ce6c4ab48ba8f82487683ac66dd4753e3cee25c24444611fb8f47af8
`pragma protect end_digest_block
`pragma protect end_protected
