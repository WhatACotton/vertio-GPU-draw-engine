`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
Z+Ql5iraidj0dxOhwU8pYKYeCeQY3q1l63xBprk0pOea4ccH+73vEupsfVd/JB5fTmS67lgDSIUv8XQ7x6ZYfO/lHW4G9rWZOTypyUJ/LYLNihrTL56wkDJx144PDyDQoohYWHupfjmKMVKmWu2K3ZQNINfqzAvbZbgGvi7ssdcBwILsK38rQccbSB7Md7+noE5nyPG7Q+FMTmRQ2N6BKWzPdR/X1ZUvNSAZY88wKdGZ3sykOY8ahb+jMOEkoKjzT2I98oIo7YJtr5u65aqzU0G9E5NeANMbByd06yjCIgE3VmijU/crnH5NA7/8FWv0s60YD3P1jVH1dn59Zpu6upNXWBGYweKL9YImER7xN0rf/hOlzIlKZsUpmsgN93yd8kEiDZxhn30EwOCbLp7Z0RirsADPEleR+8CwPh//7gkQGnWJh+EZCx2ybiuuPri15SzvdmE/8xDkgeMZJbEY6KpNXCfHBdoA5hUOMH9/lzUTK7xO8t7dA0yhOz5s6S2lD2ZtBapdbYtrMLH5JKEHt0CgqHpSZK/bUCkONY1bGMvq+UcrPnFYe4dO58iYWbyg3t2WmZ89/WZhvkB1xabK+chUfBpnNXsXpe0pn7fAsOBa4gOquXmDXRVwjbXVyPFsaesTX4VU5x9CXdkStB9YB6M8CS5KG2WgWDbKGdY7dOlLSePqOD7SudxTN9PuyPI2hi8fxuqmttIKi5FhUSKSQZ2MmhqUPkgldo3S2Nft2OtLBd16YFLH1k/rfsIKZye8fncC/ltRpvvS6Oouttq2eTv2u4YVKqFTcDD2b57Nw29uuCWEzTNhIiAI8WmuMNEJWeYENVL2pLXntwE9X3U7/6lOmvXH5KmeWfsrWKQSIzgi55BsSwyiEul/b8Ym2RmKDEP4AfKEtcopYJ4SSRA5Ap/H3AdUKOkZdYexajDh3r6OtXOu5GueY3Kc4VbWUmaygRmY0qaLp0gv7Ch6Bh7OzZcNtbrbp0ohrpkIN2M/5Vl43XQedKvq7AnPiJ4jZxn1l8Q5O34XXyWX5CqUBSH2emxFJabCXgqDGEHlTLokpHxspkDAZc9JVbeYUZM6R9TVspTFzkYruP59c3i9fdsW/7NZ8M5yCw8BcRBFVTVFuUwYhu9oYYOXAB9zv+r2DNromJOAlEnqp4a/0CyoROM6HXJSr0S1rt1Kd0toqa0y7uAsYpfTo8lxLADcYPjtMBJI3cVQPBvNMpxP1yxk05Nzmrff0tsgDwF+wb9qYWtqLrhb1EpOS7ZlgTl7+JZ6XHtxrYLShRmJ60NmvYABn5PTZDpojO1TX5IJ4oxmOF220dhpfxMY8v89BWIl0d7SrBnglD0MLg5mAnF7JRtsQUQcQ1ID6SzdTmDHghggGco2G/pV7frS3OBdshv+hvqSb70GP0CpHrAYeJ8rt8k2861MefJWdlHpyc/+HEDUZ5z84PdElENcFd6tAzCUKLt/SOiCmnQng1vDV43GpO6XUM72xSRqNy4jD85pRP4RJ8L7ESYU6WJAIBVKOnjMLalLcYKvUHsusSt2oZOC1y1hrhGq7++uGNC/0wD8197y+wAwZ7FO63QNDJ91N9yUTQj18xwEfiREw5ff20FASQSZ7c3RQjSlusNCWhywCC20pBjXsKseAS6Ivw2tEQhHD3gR4wpGwdPLa7lIA/N4MU1VL0Z9AD0xbRXpOoEU0ZEA8ptMTRPFnBrqeaf8EqGcNOFXpLxZ9IzPrw2CE4pRh9CV9E330he3Uf3GotGWrsh0cqJ5rm2x4ulgTP6gsWicqdSXiFjyZEeqjDW9ASRb07eoeJ0KKPBnCSt0KTCX7wvBUkeux2v9AwEmz1/OLv96BPC4KJvk90Hlz/+m9VbbXMN8dkLa6agCPUxHoak9QV051c1lbwEBJI3LmSP85ghM7i1YoSmuCCCr/FicTWT9/i1E8qC26AHvsWh0nHzyCdY/7VeSVrZmV6WdXcaSBQ946qicgFIELgcDtVmCkjM7147gqk6T6cnsrLoLWH9JKyyRlfko7v3ib6/2kDXJsnujKU5hztH8mn9RgptOToY8QXkrmo3LislfmNh5prcqp5sYuJWZWIoSGFd1FN65slVLMnEn6apZ96Ua3hCaA75DGohQvDc4gCsz6vCjcgN/wZ1s5Ag/a8NgYAI/gtyM36eZbeAogG03mXC9AYAhs7Xj4tBG+vvUHZ/0r4IrJSflCBvbEu27LG0klRmpsN1pndCrBRrRK/+NmCNynunMgu5xkzJsYmMOTQbnxPkGlIKG4sACRYOZWVijOcsmNCdGoftThFWgLP/8p6C3X+SoakmRWCa8HPrixrfg6BTt0P1HFTQNQU3HJ/zmI+rGRMeKDdJd4kLG8uN90IjKmLgkJiwJNhvD8PemQZshKW3CSCua58Vghp/DHiKjAnTQVQkMYZUY713HO4YRKoEoqYtV3Ee6x8Vmrult7ZFBXo99qUylkpG0+CI+/LehDvdCgtLdQ2KFxgM5QuNcK6qtb1uJWthDEfytKv+WohEXsntipxttk7+lAIyi3KGyE3tPreivlxr0NFyADj8JvbdUg9ZDdWHB2OQ+gOu+tbLFxV70+dYu5SacqWiA44qJff4LgpXsqJBpGmsVl3P/OFAOn5FpjZq2p4G0P34fMrdFLaPaz0PVZHsWOckRZrIRaTsM0SgTJeSzehITg0bB+kFczwbMSQdmnA997N4k8uB36XixotEd1XJuNH5/YC/daOkNXu9r3nlwNIOKbs0aPrmd2/hRUB5cOMvsl+HQnnz1aoxV5Eu+w+cm3tO6ZeLElVwnZR8Qr2vy9TGtOpq8OLhRFxbYe65XjDfO7eHlXyqAX0aCBp5ZDc4PtydDrC9lOeCIuoGl5YlQDToCmspEAZ+mwM0wThsRXPdJTOFh14Qa6qfhR8C3bfoZOoojF56cvZC6k+y4i+RRWR7hWclM07P2UU66ZEjMCXmuEKNhiZS5USM6YGU5pPlA9w9jmClN55J9GuzDYCleaipXT7UVmVg+C2rOlvPH4hFni/in2HhKUuR1UY9eewvHmZb+cxHh/A0RXMK9JWXeREFkayuRYarwRTSPzPqUdXXN2bPNl5PdW+b+AXgK5G8e2goOKP49w+/OPKsUrid/3hc+Gkrzo3XDDRx3agMtfmVXbidITbc3ag0iEJ2rdy5dEKKzeyXK5o1TkFkxa4yw/knlxSe4cR2fdpH+IJ0rRFO6Q16hBnDZ1LQuvXVQ5TwhqOpwR1AHOABb9mo/sRwjJP1V0jYQtHsbVmOExPxKiFsRlryOS0uT+FpoBZnAFsVUFNpYIIVfMc98QTjcINWXSiSrZLwpH+UOIQ4qkyCWYXIYU1Yaeoim80gxKzCdYTx2Qmj8y48mIXrsHWjpmkakokWSlczAOeY+zvHuKcobb3BTsYfoixUokZN4aIAtuM3YtIrJZvDa32RcY7rzL4UKZ2NwRW60uLRwTMrbagzJXxgKqJP3IRXmOjPkjrT5Rrg7vnli45L2fudKDr18k0ptMyWtz5BSWQwNMVwyumS7Chl436v2jdA6fuxOj2zkOVb6rEFj5fdr/q+4UkqnAF7mLONMMT5L/TUeVy+QIPC5Di6FA9ciP3c2LfKVwm5HtEU/Fme0lqw8Kaaa1c4rkIsZrdVCUUqdsNhR57SVjgWezXxvXLTCgB//KGL2Q1YzQUjMNOhnEaiKZIKXQ/g/NCMgJPLuNIFMX8lGTz/vCkeIgRZc1O0ztl6aoKT19ZtnwAhjW+szSTm45b5F8qz2cRRk7alQhwYg4SUiPda8XSRNgQHCV4g9WM4frnXsYJ/C+o9hstxuxQ8Zpg4u8Bho3Tl+8acp9ZXG4QGBl0dOU+TjXyJTByAo7wmb4vwS61ugh+LUdM6bk/QLXrnjuc8SgmCx3gQNiujcIgon2xDvzieO/ldq3Yv7epEAjxfdrb5DKRHsvtVCfVqCxaNYTHibnaLjoQwQnnWTEg9V1SmIlXcwvkOslQp8B1YmdGMQhqQAScFLYDGch/FfH42tVgONZxg78seYhM22C2FuLuQb169K6W90ThC16kM2V3Qjw3LJAwrNdJHnscUMC+gStFDmKtqLtNOqQYkEPDZ3uv6FyTWTm1buBuk4Ihxn5WdXh1nrGK0/gq2ytNHU1bB3bU5oXcxFIJB6z9XvV36KksSHnAHSgWUAfNWR7Cad/SUse1APxfZ0X1PWZA+vSaVvekQS3GYGthjbCDNcXEx2I1oJpCisyiu56v1fhAhWIgumUqmVhoJkVTMcWKdo9rKAdxIREoHJFpZUZtckJy9AyKPHyl0Oc4cGFoJWGiay0gB+igRdGitTZhGATt9lp39uOpgZs5HEeat1fklzZSMrnVP/lIrnrrEVb3IOxGuiNZl7ebY5xOKjRIlUxg1mp3nHWMZJ5dWLvr1tWDS1GTv/m+NaSlaD3vMQrk5YPjXfnNiiJwNFVmb8jPyJg4EBTWYl330OGvxxxTCviEgJrrEGsFWfFV5silx9buWwOEEW6DlWvFkjZidRNjPbLITQWl68MGncU43jSixyve8Nh87BaYVuPoyXi6zm7irW+OTqdQPQp0ytGrWfgzaPRIqGfb4121zXUNEp9M+yByIHAcU4Ai9s+9mS7+nSDqHxSye+V52UaoQEXBQ+TWx4nRKsEYxXlRQ+G+uabRz2AGirwc2tfIfPWm2BvfG6AYI/6ZDleH/gxb4Zzf1THhj2QhUd2v71UIBqMwjZA4Ig+HsHkftyMg8xoNKB37PzKD86jyO0XLnF9KJydNFvLQBbXXXr4PkQ/I+ZPzA4s2z4c4RKNyTR8AlO2Q1z11Htx4LaMCPP/hKvHAPSxJCdJSbMZKVzSD4bhdR7iD4Tf4YQur3wUF3y23xVwm+GegSnWYPfyFq6zMsK/6c9R4vMJI2bMUnKLtU6Lu0PHNPqeSM2IMF/gceqzS9Lv/oeUgEcvz0Tf9tXnjVaLXkjYlWO0iXBCEvO50KVuWqKO5CCwGvviPJXbxthPm9a9dV+4kn9mF2alBcZ5q2n1ATZS8r4+/jnmiaXpOzHalnSJJqiSl7aKg8NBlpuCIDMyPUbKKKOneFw3FRV2vsuOMY7ujhKFmsZH5uKh5/OQGVTN9q76NxS8xNaAzzw3dWRQMEsHg31OHEqLJJg0h4X6jWnqQjxH2rEGq4YD0gfa0r75hIdUvYIAyeRpKj00eCuZdTvGsnViPU9NDeDlBsOKpgd0u/xQvh5LdvM2eUASUqe80uRaZzSdELcTHqPiMfgxWqCLa3XjwcV89J/a7rIZLiFpxhvllyRGky6j4ClJwZRz87L63ctya++lUdYro6uUC4tpRwV8FzERF0GY8OJBhwvk8GGKl2v1vaib3CcqMZG8kVmTcLOHw1SnYAsTohHSbUtY5O3+xL8DReIPjo0NqRrwYZaqICsYfP0+/r5ag2Kdg61dYF8nKO/6muO6MAz55CVrj9GwPqPQJXOm1xgvhLlqSbRaY5kFB7LFnoXLdhwN7IfHVBuReE5/h4wQhM1ITcE6/LexczI7kCGk7IFCfBYaeUV/fW4/LXTtdSLk/cRuP5LMFymqzGUYXk56Ul3EhTz+kfo2Xnaud5e6CpaSmS5MpIrFkTNl7DTCH/Sxi5i5D6P9IEzRpSg/rSYUcMkMHPIr+3Vgjg2xWVW6krJCEsZHuCmJVcLlXNcpLgxZv+W/JrUYPNzY8jHluiOWx1C9Vzc+4TEAEZ7HM6FszIpvT1U/7sKjNHBGKYPYUjzKZ2FCuHaDiu3KRRy399Sbb0CHNiVGERWH1DeVQ03EssWA8uZdy4TU8FATg9+pvMW9mgWNd01bSzyUg3zQai8hC91SChelacQaIfYueVT+yzzT3WeZzKnW80nK6z4YktftonUnIoQHwrCNcvWoGvdOE3GSp260fsofby402lRlOOmQlaa79ZZ5GOdJuE0hRjS+DUxgvisDGufQxaj8qCmYtGFKvIOo/boIgqN9h8cTpYTd9wOrqMaZvflYyDDx0yaEF3dlWZcaiS7tpgN7xx6bIMQW307Z4bUOWwkXIR+I+nKDOfGtbeZMY7Vn4LEc3eKjYea7q5ysb97qMw10VQ1JJO4E6PTw2+ZjJ0nTC1WG/GF+xgM6Gt+oyCmw3qmbp6FsyTDMRJscyKJjixEz98rJv9PxLRkArTSgSm1IIZI7Tbe7C1tII46Ov16Jvl0QVua1yOPrnMBUdObEn9wdzAYz+2yTLcw3zDzvhym0zrwH4e6MYUPfmn/mq5903gcX34Df30CoBczGZb2RHHpWAUwSEnjgaYsMZOcmmjXrWzluVLpqGW8cBWzseAIMk6SKebEV/+ItKSAiU3PXlAcuT+gG4QskVB5THEiMkZ8At8sw33usGY7NMyPsD2DW8FogynaXcF9JhxV4zu23kzIIbFfwN6iosjI3QxAnEEpD5fbn6x16P/A9VKTM023yCBJ6KEVk26p9DWcFJGbWpWVdNjjGRbdnBSU0pgz3JkqIg0GL10WRkVfQvJfrAwexZE8UXO4sda1X25ZnYXwvLBTRjGKMDl86CLrsge3V0jk1RJjTgq3wqDo28hNMTeK+my+nssvEtexsOOBPNN64wvM+k/tI7+rxzXPZtPj98i+zqrIfCiQzCd/z9GbsToW9RsOG3tqwOAjM1S5RvVOtCO5mB+2eH8ksU4vVKqH5fgY+wIZ94ipt38fhr6BEuQAaZQjgNT+X3ib8rLpWOJRSgEUswV2cZW2OEX02VTSbG9kUkvvREOLFvRYwnFFZUs3m3ywfF8XAOVEkDzFWQiKistFAH1HpYzcemmptkTDSIt3j9O9HDTlkG5SGAc997RWoynk4iFbVdKA7dF6A+s7wkuexPTwD2+K46+WSk9dhQK/TFed/zVPtda67mCub2/ktZ8QdNam9aJlq1sH4V7XCRyv7eocIqbknwyUuDsf04N8glNkXrTKsIPV6HxTLviJlui1E55dzKLkZTyXKpVpF+rDALlEbD12vsfb2wV+Td9rbvFNZFNq9McbIgV6Obij7UxkyUELcmg5npmnqXmbHP7SJS9MFFVurPCfYiJxO/SViDCQU7xpMz6gJnU4UsUNeX9bP2mzNr+isfBxieRU9KqqZVb8PIAIj5q11FRTkoe72z4U1nGZhXivrSdQvvPROlm9ztT+/3UyDQylFLbXcNnMSIEXO+nfAT7kjkAZSMHX938mCm64XLGqDA64tBWspHMmDUqmb+Jk21IyEVOAnkw7xXeFVfIFk4uUUNXV4IReCi77W+5dgjDurldcKQ4N+Ufbq2lFsA6YD5zB4WIvg7DRg2r67bf2tkoGNSvFFHnXv15QIG/A9w1vYl4PiQJ4tHac4un9fMr2EyumjzYm31p2mzZEOp4gmU+nMBUsJ78POWk0Vin37Fjea93soTUliXJjPEVGX1DBZIMMysX34BcRiGGJqccqFcYtNWiiOY/a+iXzaW8TWMwIC8mfLT1aBClmobfgtkyFhz/4TQ5PdAIg+FpYB+J6DT58L2oxAwrjlczAu9sWp++X0zECD+8Y+f5Q/42z7vk2e8MPlxC+OhYX5/88nEt4Reegsv5R3tZhgjA9LY/wlslS7MiW73GYTwA2IoNx1iXn3Eds5uSgwRBUd7L29vo7qlZsc/OlzGhl6AEg32eAwnB0k6ohtSKvG9kEI8eriTABmGI9s/uNYR/AV72BvBcFpzajE4jDhz7crCOP9WoQvpAAr3pQ5+QyIFHEQZ6sTCCgcuXBlv78tsRRBigNJjjlzroewGycYOd2gX9VQY1WeJqc3toQvgqEZM7kJVRWgGvnv1rkMclpWnSGP3qZy2EwqOrgiEw6DYxyZZJ6eD8GGs9U5CCDD4j8GUfuTwvU+FAc3NRhW+Nrhn1vHObXbDQeqRlScb6fqa1noNf8b33ynaOdp0Udbauv6bsfcJGdiqJTib620648ZMarq7fCJnJfIbiZyPbJQpQP7irz1Jivxw1GK73xhmfu+Y6wKyWWsivaaKCs7l7Z+0zCk94lj2EdAiAQb7AW7/Ql279LpIPkD6hyee2HP9vn4L5Tqgd6Do9wUVm/thc6ZusMi674aL5SSwKBe3aU69TJj1ZPgwyzupQdejCxgZ9V3tik3I02FwG9oj1/y4KhlfjL5SWfZ1mNGURjTJNCr9FsNrLRbBlZnuLgyEoo6b/1P+TESN3y0nPP6415VmDLhXtgHNwPNy/LljSm3X3KoD88WoocEdk8D7GNl1QWykHSzJVoQ5y8qbclSv8NQPG3ApjIAAE8kNcF+Qaud4E0M5XcjIscMWprmKyLWdqhayWGnU/GkF2b8IIsPa5JPsJFqSfOxcyhod2EW7QVhE6ZBzXc0hpT48jnvT6crEfkC+BIKjhBTFUE3FHm4vpe+WIhIRe6nbVjxRhYGK2ezCE9NhIgsqLLv3rvf1SZSJl2w+zm4dXZbshfLiR6DMGV4I2vIFLBKPYK7vG79T5JtEpknFjAm7OZyPhyeaQ8hM3LzmtvRmdRj0ootgayObpamtHsunrdqcbp5rj9M8qz6ecaqYhrSxEWzHO/Wi7LyiCMLuYGgEkWNsVMssRT0N60aEqrZXGl3WaE8jVKE0VHMLxF24/eGiaMik68EMzpKveEMYdZ/kJqWjqOsL6I3O2As0QzJ6ufMYoQ9AgYEkKe4Ax5r59CBpGQorZTcI+Ri/uY4HCKSibKDsDLA91fzzkk+QJiEuYobI8kNfppAkIpl1Iju1zdxGzqqZyW/EGJquX0O0v9TCZDEM7RO0yPuV1wzqNzVtTrq8iNy6xma8PU5+Iwi7Vc1OYKbFE9UDSFjcqwLCT4h50+FQhZP7AY8UWpTjPA98ryEJwetQY9XtEsSZx8F+PElu9HNd0yJzN+99wdNiC+bhc7j650c85JV6vM/EJ8j/kwe9vz6HGTytHq/0LUPZOUoUn3o09gtBIyLztEijGrR/Vxi+j2FaaLu3KV9fj01+iLZAhS1xy1eUvHS57xAW+LlqEAw68sQXNhLjf1cnyVwk99Ev695137Z/fqGIxfoqKEKt3WhEyRvM1gbZ10Y2698mSeTM4zBxdB1cEyhEY/hm8vhx3MxLswgYqcCXDjNeFbd6FUvPtNZCroCAh6k9ntf/g8hh7cd1Fh13F7xrj+Co+hEMxWvMwwr4uZMH92N2iFxeDiyxO6UenXebNcVxF7LEbnnPtyILiRLDEt+LCC0NO+O41ZSNB3YIvSsmkgCIA0b8njhzl2kOz85NR/WwZBkW0Z/Qk8lswtxKGECh5U8oDLmz5npVDQfeIaGvVSUWilAaFtqFwGe29+DxTf3vbYld9NfSZ4Ru2GRJo2U1bnN4fOXJTs6te1kVMCEcQ8UAV0y84xEkYC0ZaucoShb4Bs3el3Ey3rXAeAznMNepnas4ciK6UgssqHqpOitLtT/wnaTfMuAg/1KSyWI2uPguBjFi656K42pzOy+UUhNqfFuHppqZPsSHuIcD5Zt/udvS3sQEMIQWneQbMnatdInyVEEuYbCmgEjRd1B2QSBhI0lOFVprtZZMpFIXD8uHWxq/5MukzCYoBOuPioOW7xhmIeki+ng5ffd9sOJKK4H8J0jMUa3qPSqug6L7zyE9EzWRZUxNx9pq5Qo0d8ZPgNgobeKcvGkaAKe+H8sUGqmKtVlYkUU+Xdz+33GuQ5rtJEvboLGVQLRoF9ZaA8x9HM9WC9EIACwOFzO47p+DV0Dkim4Pc0JjDLevpyxg8Xda8dv5h6WnOkaCiqB0fjhSmMIEKYrS8ryNX4WArAfg4wqwhEjJCQ/foWF0UqZBjnUDuULnID3Vj+o3hXdzJS9Sqii0oDoP+cAZoNQjk61Jdyx9D4/Q6SadepDmQgh2kCwjDjx4cI18v3Gv4keOvHfzsZRK/rD4AjS6lOtXTiyr4mYO51vhnvZNa3yv1drX1vAtc3JtL7yIdY8OZvA1Db5WOvqMwmUaLf5QBNN6iZyOytzX0aLx0=
`pragma protect end_data_block
`pragma protect digest_block
f56ba48c7eedb112f71389ed689608fac5622a62a8af5848743ff34d0f96b8dc
`pragma protect end_digest_block
`pragma protect end_protected
