`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
u7FUUfnn7QoaHuxB3QvbUciwu97LBfXoj4051FZbfobQaxvEGoc0ykdebfSnxPqRLYx7TF3JY3fvU0GjSq8qDfzD44fvixbHaVlde1b6mPiimAr0V+dWgDuIN370cLWSN5sUIcsKO119ireVQcM5wHgv62qbLXyV5jctumh6bk9KylGEsuDofPb1eeu6i8s+qJFO7yegO1/a7YJeMisXr1zee0blvLfkfdO6KKkBVeEInN1MxCLrwkYpm+XmXhOfs+XSLIFdjtnACMwhyBuVyhU4uQTsG/Qic5HLhRa0K1K3kytNG//Kux/0q9M+EkaEkULhs4E4LfGK406vkrwtIRgnndUxiUagFITUJQpWoHAJ0uTr8ZmrqjEJ+HGnJ0miUGjGs2b9Qb1gEQD/N50JoqXKg7T6PvWBJnKFTqz6WbRc3EWiKUWoRXhQhvNtiWmnJ7sGboQz8aOLT9Vriu+KchiaFHD0/aD0VfBcLQtxhYpGDjx+8FBDCXDzvF2aOqenXInGUzr+zpZUQpaUYgWOvsV0EjQOiaWGtQSB/uB5H0dbRNSw0K9SORsuz25M1NXKufUPRUYrLEWPTRxVkH18U6QuWv6Q3eb5jLQtca8KGwUWGp6A4wJlfwPTo4xUpn2QSFwFhoFTdzLevCLZFmK7c4S3U1G0XEP1HGKXel/IkFEW6sk5iVHeSJyMTZM9o2GXJcClJpeV+Uq5//WHZzcH8uc3t+QhpY2nYXPcfKUoItBXO3f9NueIIjRSuQYpnMp871WKL9m8Pf6g3vNW7jPeEDmVN031g6VHSjyz35LpRZ6ZtVHKZb4Bhf8oHHvPbDlxgIcXHzaweEHyXjLfQIJfH5pXVTl13i8nkbL06wZc22ALLy422ZqWwK6FBcOias1N5alWHjMxH7dLGmHE+ahgoQrFHtmY0I0ZtbDwA/0eSIOCmYwXQpaRSv+skXqz08p2BA5mHAeYlzWRVVNxNDJsGoR2Z2HAxn9Ft4iXawFt6xUzwKpiTPILGwKBXSNJWNFyLy75xGTJm8u4qywuM87FycI0RMWuCJTbiKvMK60yLF0lHwy6wa9NIG7yG/efKQjg2OVcNNWi9SeEW1CT7NcqJj2nqZVIz+u1C0CjSNILfdEWsbczvDXB9N5zYsGaGjH9wpnjQMojxJO9IC4ZhqzhM02ufp6wFrN2dpPLBuwZ1vNhEEuFoW0HxTGXG2OuyrjTZNvs0oiaWkyNCRj4O0vD8y3HcHYozwezqKo+xBLInaVBllkwSJBuKNOPfCD20+HxVgiCVZFqaEn07AgIBtb+cM7ZRhhJdYJ7+vwJY0Spia2PBcRIIF41Biwbnu+fDQcgIJWdCvd6cd63+4UQPcn2NuLntva8fghnuFEsLpEFp++HfKzMMh83FLOixZrndPITNj83y4G/cC3aaNc/Yloexp6tTeEnxRVwx6EyPjIZi9o8BMgg9NN1BWt4IpjJ+VLsOACgI9B0He3OVSYWZJw4u15Iazm7HljrKaNEELT54YKHWSVykPAfyCVlm1OjnMoIhK/Xz3llRgeQSFNTJWzkCIX/GQFFjqhKnZTlaVkbcbEviG1flOLiuAz1qmPtCzOPEpdS9HqtLFijC3cVP6PTT8RY3dMIBx2WHlGbB8upWBAb9esL4ll1P2w1wMHW8NUOe9thiPh+HELxmyyJR+5c8N9DWCb1nIeIsMPGH0s5H58d8HhQpGIiaMrV4tuQBBoh0b35rA/JgpOXPiJ0uYsfF2YuyCHTqQ9LmRDoQljmc6Xd8VxJkq6wNRRS52uR2+01EjnnS6mrlP/lHe1fCEGKIq57UdmfDbI7kOjeHPCEnRHqFr483/6h2xsrjahUfkJSzu+/LBkyqNeVOxlhw7WtQcXyVxEyMse9MO37Kv4zjwR20rpj64xrdEABdzcC2Hljc+owBvuTjbv+kWQEmMKjWB5KbQoCoShBw5m7W82pOx7sjTJSabGN2IQG1VvQ/A9kD3KY5LYebQhhla2k8sI8DVqoGAmTfxqPNVNp5jOQSyYnYV66GmuEHbnOit4J4gEh/d83hK2hAdCPJozm8bd50dd3Ye3sbNZ/lyoKdrF9hTQNI1lPNHDPgGUbDhD8xK3ZgrrtBJiDf/vsU4gFEmoh38hsvBNGJ2McSRk3Ei4O06iqqA3H42yUIXZ606rzE+oqpXtRz6G3/xWYrPQRYET0arlPIkHgY7cHWdxiVVXZK/VU2BYYGWjhbAjusxzO7vW9SICNDGpYMB1urAD8JAskkqtRiklFcuRHMx1I3w/vl7kD7uyH1Xv5v6m/kr5tQ1euGeTaOAKtYDV4Obdgq9D2q39ca6wp/Vce3Bj20aE8MEZ/nV4g4yQWLrnUef03Nuw6YPrPZAFlowQ0xV8v0kpHDPD8jUWhbeP0FlUbvaU/jKG4/FqxHthjhHs0srqfKk9f08vwH6XSWaUBPA2eBU7s7RhsBhkVv4U0szoCwYO8xgJIFBdViFJbsS/5bgsKQ79QShWVbSHwHzxklghHPUh/8Fp7r4C4+5yeZDVU8jsi1HvTvs+ndkUwDthuaLPT3LfjrsPm4hCJgrpJog9kHmbpbhwHFiwlTR/TWz1H6vHEot08+0KwHX3box2HPIwvJ54hFMuTCmraHYFhxhTR1iL8sS7Y1QawSHkedO7x/5huJDzoI9goqEt2XMUxlVxJcaGAu2alL9zxw4nTRdzhYENERQGdXqztTSmnGgdWOKatgg+2T9zwfaQx2kr9t88p4KHqPDr8K+b6MTC3wxEpd4HQhuxAkq/igsrWBDb+RcHaLb6DDcq73utMzxjI89OaF6TUUC4Qecl66xWJPr94svV65kRb3Glo5eXnpuwsH0mig/Vl7fEM+8UYIf0c2hOCH43mlAv+XkASuoG6W8TmrUGP6wBXN6RNf/FfctuKipeMwfG+LZ6NILrxZ6EhgQ8g23wv3XSFN86qcHSeFBAIescuz7zgCzOKhh2npQLr2J05JK7JYtON0Epm2+xAbcInRe+gPjqY40jTZ1+r1qDqqQzmKb4I7QLhzzcmqqX77kI0vlKwhgygnn0VX63RpTg+pxybG/o9tmrquDPGeq0BiEo8giXTgusvUZUSfPONryjSgFaOvDXCARtxypFACWpbpziZTMq/5necUZnE/j8UN3D0j7ALxF2aWgSqvfMTQCXrPHPB0FptXgAr6L1NxioQBf1cGWzEfOpsJy6IaGmSapQgENUJPkp5RGuXOvK3qexDn+Vy0z66oHzfusieciTEaIvgP9vPWiielyJvYyuiRS3et7AfzmHt9u4ZO2TYjT6Qei99EuQvj5z74ebgAt5VA4yBNFrNj2pQwz25rjRVqj/+leuMl2JLxoaHVNm6FmJ9uN2S1fKDTcicRppSb82x+tVIM685isQiCMQvNLo+ksbzaBG43GGdYE+qGjlZ+ab7S00+HDaLVWmaru0grnvUi7u/H/qKc4HpRwXD7To+dDob+ilaqZwi9isU80sBU6i2olSAtva7zY5zww46lRAoGb88NrChZu3TUvf8uZCwTki57xdp2epIsa4rfwzT/QveWSGmJvNr2KSbrkcYMFTJg2xYS5Y5KhQmQ3c+wM5BSFWFpG757BllV3Nolu2GunN/f4Z+2eUd2VMVguSNUQdzmjvb5J7zU42xI+UT3V4tnrpi8LTcLA+sk6K9rSjughuPt8E15Ca6btQU9dC6Qo3Ph1hGZHpp+uAdc7L9xg4QWeXWyiHELR3ChDrABOylZRXg6PIB22nPJRNPH75ey6UCM7eCO5fx0MkIrGbyPl2y4aLP9Yo9vc2Wl36emyPzUkrO7Mdi0vqrTW1P1983pCCgtQE7+5PUIzAQRHBkDxCeB8jJ8p8RVjc9Hk293yGy/ceYDTH8i28yurW6IrrbUJvxG9s5aAKvfiy8OlQXaatp7eHXMFtqAOrX9om29d5+69/SNRTlO99BkMgsvTYvLuRboPDAigpD6l3x4P//WkW6UCckyzmosj92vD1pVUNiKjtVXK4NDeLNB2gxalySRliV5UGpZ2MVL5oVL/+bu9h42FY9qt8MI82BF3UHf7va5/bi20Q+KY8xGmdORIg/MQ8kV27sTpoBCCCbbA6hijCo3wdIBzX74VGIDolMubH/mzs72U3eUUd6TQaLvwRxjp5iTlgFZbMNHyUvbuplx6YJOlaB6sK6LTVtx28CBmV8Kx7zGOgCwgTRnni2plY3mUX8z88Adf/4k/qyQpJhdSD2/ahgXU5wd9Ky/0yHHIE7YiBihkWaRv2v9nmd+auZItlFmjW9k+0lbJpCQDqiEPYvhd49Y/Y5k4/vNyOVyaSE8t4W12XkABUT3ruFvZCq4acYXxs+OSJZCJM9+N121FslfC+xKMsI9eWAP6nFEp/3j/YzdYetb5ECx1k4ZLylODQ1WtfZgVfqTrFWlpMlCkWkGHtYC+ZBQIDIvm6vzIpEfUsh64Ec4sIpW1TtbWh8oYQRFMEZkVi8ve741QP5LEGEl0Jxw7aSrFGvemI0hBFXTNhSHIcDVs+/+SCleDXX2TBWvJyF7Inx9/qvsPTRPX8vmSAGpVTsuZBC+W1w1Xxx4VedHJ9q983HGt4z+DlzgRanq5xluafJhb4WTTN6jffeLLe3K9M3CkFVqaSxbP5l1wQazy6qq9E2KgwaaO0FVk8ETyW+xMb57gzKXXhHGIg2aMMlrErCWDcYnYgTG8brFPm1p5D4uh3D57eBvwshG907u9yZTz2PC5APby9NLu/LMallT6U/0VzFr10HiXqez2RfKSQhgymozWfbTc1RwjegwscOzKtMokvg7M4Z37EtwW7U0luPCNMlYclH6gMvRAZTmMT+7rJyCgnAaZwIPWY1wVdombZj7G9PNVQpWC3DAZ1j+s6QQ+6Zrulq+F9ldqPQ+3nlGZizkiIhbQnhYMZZ3SoU/3eLupifzR+kYmciiPQZ/TOyB5EG1KEZfKaBKaC4iCjhOkjuhvlmN5nOeutBfE+aKL3/kXzkzhyN6thIEh0lP3dN0CZ0Js/qkFbfsOX5u9kaejg8nC5XvPrl/UJGEu7Pl/yXJmVZED6qOkxPnpixoJkrBaKLllkm8A6+awL88aMgdqR938w9iVCYB7tKQzsTSaBpa1tT0r7pw2sawSiVlgSW4Y59FFwERnM0pIpZtuNbeWRxN71MWQfl16/8e6rLYFkAccp9avGxW0b1iEaM+VphTASrIB3DtaGF1xZtmlzDuQjm4EaTy3ryBX7gbRwqoggKl6BAjUlEZbSQiVJNftPcLa3o+zSZi72MzFU+SIcP9Wd3Vpwz169upAknlnUviAsSu20RKRU3dDHJxgpi3OS/+LrEYv1CR+Pkayxo7F3J8FXNon2yFJAXb+f4ts0xCm9OOVVBMQdFQsjuSvGj0kHkkUGOeTR/k9eaWgZuZxuHRlM0Xv7onKJgAWlAeUWf1asKBuYHI7bBVN7QNdExUf9fakzO7o+C+5vsVVM0mjgPptEDRG1CryoL3GzqAjaXvLVggup0rcSRZVDoiTTX8U2Z16Tq3rST6W3EAkW+sv3Q7LbYfnNV1yY8sf7MM2Ey0tivTVYxGO1UCvMuaWRzu3Xjlu8dV9MZdl9Tg08VEvtGQNQawryhqYBV63WY80HFWr+e5vGVwbB3NwVQYIPXNQuob4b1AYeOwpr4CY/GIjf0lif8yyABENRHrGqFz5SmYZ4jw4+wREtgI3J1p3MKHdlInq3cWzshXP/jMuJNlbkUitaqb4sNI1uZY8pTjhuk6kIT3Dfqxqejfq0deuCmwU74KUA0drZAZ9OHdXO7a6PEUg+D3jFZiUuEVss7yd8eZKnAZY269eTtL64KGsVW7MHFDAHTV8jalyz3A/QTbFIhzC/nQiSj00oPSEFbXjUQYiO2uPCD1m79em85B0/Ti2rxsNH1EyhhR7LbXNxN02R9+e1j3U0y+BAvg6xkvYELg9+MFQYCfxDW25Ov3hAB9x4KSCZadLZrtXJxrDvOQFzmliTx757kUoEBx0c+t+Yp2pcXL9Ml8nebQkuS4vV5TxLBognC07ENmVyt8WQ4l3jg4YbnqOtXmLUugx+bbKKqoIlZRUdWniGOnB1YAL9z+6JfUU3iLRmm9DYkZQwx/wGwb5X0ORwOa1TRG2Hx+n6PVKSvCvbxuSPEoIDytzxlel+SXPgH3qd2xlgM5CnbEEjy3uIg9uLJ65IWnqLT+R56K2Fkilx4BfSSBY6rKbTB1fkQGpOanrlvzvKgKsRTffaVhowEm6XS50FAX0ecY0cXw4VdpDFSRXo7hwnG9zDLwivHgxWyhnD7An+Rx1C5RzrYIbcKYev5vODhwsirwvawH0GrTDf89QFCjThmuvQNkkb9lZ7t1bz0pmGCrVLgEXsOT/cn44TBTbyimvFCSLlglnq5tJ6BuWFescreK1A9l1JzVbNf04h88v5yQwHmPjg5XTXwcmvWMfWE/uUthFgbdCZuby3TtutuFtQp7I4uBEBweiF7VWSSXmLLJ/6VjKTccH1djBMUznObzWiDSY3+HR9k1g+rGbuMmWACvP6mbRYiooZbgGJ7jHNrYQdPRpBJriH+MY9jAb3QfupHjFG0oxt88g8zK25uMl9Uxv8iK+KPvf4jp1VVvf+SuKmTv5kdnEHDFNB0yM7KxC/EUjOJdqEmI4cDymuDRQvGNkK2xBf6tZes07Sy9lQSOEkGZSRcL1ZjnzTsrUc/Esk10oObAqGx4IDHyQdQyYEMEjV7NBYE+g6BI6iS76ZMyeV5cMVI84JHE6dT1cppOBhYzIJUJz1G/N/LZJpd9dnQe02XhpqD883Knb42ChIj9fh6flHZ2Ah78zJPO5NxX46aNfxsxNmSkgKu6ci2dQT1NavX1VGL761pt+03Nd9YbP2xBYmlwcGuwnti2XygryK1QAoLl7Z0uVO09o0XImTt5j0mr0f2eeEL/rGkOZ5HM0uGb0I/HTuDsZbnQqNvUwwI6HAGfg679giSGe2TpYzul2X0YBkA0QZ5l2g81puMLgsbYdiz0uX94Ft2M3uzQImgVLymInxujUnHSIawbiHHGJb97Yb4UQpZT5e4oT7wpAfDuZWScf7TYVWWkA9NQ1sJlfyoGnGaB5fWVAoKnei8i3Vq0ZFI+B6UGlz2ktHN8yFnYi11CAyxrko4MPGIhwb+VUy0mEvjDMXYnib+8dh9CGXVpNBKf+KdtAbK/+W0qEiWB2Ou5I5TQjqqkH13UoU2xmeInNfcSSfePs5BZEcxGpPfiuG0MEh8s5XuSezimp3zGldZMJczihRcV+I6e/D+JTl9dpr9KrfKUjW6NEzw2hlAiHvVZs46p6vk5lH7YPpJtcBoH00fDzZeaWemz2td7Cz2zWhMRNBpq8sV8dOQTQxK7ND8drYLeWvteiBw+WeoY17UweZvG5FaeyasJ/ov5NyrZOVioyr0zpFjUy0WthgNzxURVfKXwhN+0ZH/NpmN2CRdHtcqOhd2VByXLjHvNOX9Ubh3CZMGQvMBDsWo6EBJdeekRbWkoTgqN4iK3zSjU+zhQJXLGPvmugZ8XoRz/d99M0pTjb0IzzGI9jJ1Ggvy/2p7AfhMdoj08dHcrbcHUWPvyJZuazbcSIJPbh75mA1UDCGInL0EDHXPRIyPwIfKl2jJLohdIRRdqr6w2QZ6SfZ6A8SE90xcuuQFfVAiEZLazNJeQbBlB/lDAN/pc6Rfbw5xsqVmMJ9152+2LUCVPIVsgZsoecMz28bjqHYemQR9cvI73Mq08P2D/xmQtGtoKxKLQjkbcKeNAviqCuMLpwwjXBy26sliHqV2ApraalVVlbbaV133LYO52ia3xBpqMnGXmlo0aAS4alF0Inbw1tzGc47TQ7MwluvgWkGv7NzsaIMEp1/hMzZ2vyDJJ5pYsvYOnmxplQ44BxJ3oX96CYatfx8vqMTwE0DHdFX28nP8PFcuS1dY6HAlRZCrHteveprbvVOJ/6PSY6RKQxMVoIwWgeVPh8+f8TbJ/ZTGjIxTkBQbD41krhCBqrCPhez1QHVwAMUG+j+oXZ9HpcpEs11iH2TtOBlOuuYsCN+Ps4eKe0+yQYoDuN2ZDxPAfYRfVw/xP+QjkXTF2nq1VggyHQY1C4Z1lbBNdspe3eFXAaVolJOANkWusoB9oy1dbU70mcHw5qgpWxP4MT0wG+WEVg0vZDJ1+jLiZrMJSYSQNt/T3hHk/zs5KNB0h7eNs7gNjjk1K/OmlZqogBO6TqX4QxeDi24hgiKT32daZRUch6Ep3q1vO+ou+XO2X2yOw7nvixsJqF6dpRRAa6clCHk0toHpOviWr1UrfCdrWlE+6gk3Zvc7tLp5f2+3MP/fARY+I+Jyx7OS2x3UL8fwt+Is3IM4sIroSOIpxzvU6DEcj0xtp85xbPqFqMaLoPmRqRd1xrtFUQX/qgbz5E12hjgQAM2Po1XcFAWs8YCkOryAuzvDfUfKaKj+8j9B0gbwP/NsGBzp7pLbuwftAqSHJlADvhFHFMp6QxhWjMlIoSHdpKkf8i0wBZEBLQCIhWlExEvJF97jNNtqxGJ98ufYo7M5QjUyd+CORl8+03Jn5QD1jiUkOcVP45SvNn2J1pTFFCG7+TRC18nY2J8c82peOyYMnF0eKmMlBTDmbvjGeDnAakduWyvFvQd02pf7g29HKI6ZoGjqvs1hwF8JJMhYDsIY4cMb9FrENx+cOUWppLlttgwtE/u9PrvuPWDah290gHfCkdZE///pXkrNV5mr5KBxm0W3vP639+Paij2+MPhBr8+WDHU2N4qClcVMWA2LnOAM6ubgsRx9fgU0+gVYfvfEcoc5SFUCVG52YPV/74v+PmS6ts3+PBI/uo45ZDZm9N9SPBwxfPTt8+WuePidy1eBE+CADjM6NvvDpmXQjAvqHChRvg9SO56ZN0N1fkXDFd/MKcQJWc0kfV6HtiAXfZ+Ib9Ks82nowbWlHLvKDK0a90GpBQIx44hwL6VDLmQYVK5jJP2xMe0/rqOWn5gBdbyybLD5kAqduYIabvYGlWYYHLhig7QfQ82TWOTcEjCQ8NoZc0vwPt/gk+qWJOnaW6S/b6NbXJejOyzHMbvA4+KNrDdjjTPInzdhfbF5hM3AWIXM/j1HL0STEI89eP+y8e9AMvtpMQcPUe5ZHRqf548gqs2ji+3VCQWhbrgJUujoFnxteVRie3uG0wx8AuJSORSOP1JSTS+HylOYrcdnPCnPViMwQ9DTkfhdVDuP0jxkoUe9H2EdtZ8W35RALCrk+BkWDO+b839U+ASYJtUgcS33Nk/Dy6BD7xUUxPRuE5JTnLoQroOQMwOSljtJme2eouq2FLQbWy/NCTUov99gfrXUd55Aba3lX1SM88LNhvpV6OvGGiQOYZSn395+5fMYggLSzU9Xn+NilX9z3pl8D4QKLnWjOyyJjbT35Thngh+QMZLvhVIc1U25w/GSW2JCNmuTi7ZWMPKeyUnofWGMlypwbcaPRhypZEYDImEpEep0rcaWPm1YqFuHN6n3gmIAezBrCYqMcs4FdxNPw9I2cCtSvUworXiLmLYvvHi+6+/5aig8glN0DSf/4tgdyGY6RLDzwlCcawYfn7P+DRBV19vnZV8i8PUS4QP7io6AXrKAARYH96FfItnLAZlgX5j6GRfa3wVc20REM/+t9dcqLtyi4XVzS4IJfSpuwi00Lszw6zMb+hdShvxl3Tor3eIBvoYKBaOFVKfmi0tAXoTZGrtqB1J65cn0sZQlbTgjyg302mtlSWqB9D8W/SWNmiZ+dzOJTcZqNzcLNlJ5kyrxfYKgTMQuRSsPrkf/g6j7iM0pgrYqVZeT9ngM6jBkiYXtUYYBQCZwgxwAiXrV4cA8y0bkE53tBYOsueSi6UswdPq2hkcFiEqXUBd3he19zFWpEZwRiPtT6/N/tSOQh0W3Jaz5cBqv2c5Ud76wCRYJyjx5fG6d3MRRasUYUv6DWAVxXrPC/bSFLFSk1wNKZj5HLtS95V9PED3nRpGOiGxApcOXF9bR7QsBaRsE2CkcoOoQyxDD/MUTSfMPsyBjHDJgQ3aALlQGXt4ybMzgKgTgyRD14SaZjl8AAh37d9dzQvyRPm2qMJKjtJD5Q6bnxRNsTHEWtjWG5WQe3bENNvIfOlXwa5RV3YtqhZX2zFiYeDNAQXWuge6LarTD9fdQN/5M+VLb8WMxTdpCHYtvlW3ttLgNcS2zXxIrp9Nv6HPWXg2BzCXgZL5gMkutsBNZsmxFLv01LjQh5dIRKnr1ZOlrQLVwf5YV5+ctEcJO7lg78RqbMRxBFNjYuN5yt0OvDmbKbJIAKFCMoO/WSouT/ej9ipqlCPOvKjHvPKbsZcScKGpyk9AsRc0Hmx9GL5RWkFQTkb1bDsZX1AlsjSVzY6MXDT/d6dMF1ymqf+f9/pC2+FpJLLqgosKYa7w6wn1JFfrXP+9ntH9BjL67oNKLo30fdFWdoIYBpom9GmSO2tfrrecnB7VVZYx1to0xFpnvuoflC1WZcuURyRENesFkIc86U+0wHDLTKXuhmhOoNZ+JKQrKnqAJpAxw+/wCeyyT5UPyESlaPXV3qOYFpEVxOsEP3fhFMFjcCxvEqr/fgy0kg5gqalBqk1yyOpFUA6ClLq6a6siMfOwt31oq8DbjvW+W3yAFqkEnWXQOKwkpcOoqSQO3EGRqjyZrWvM9XnYlYK6z5FVZ+rWKX9RivK5MgM59ufwFswMHio0/n0Dmd1GsjWuhhM5v86WILzHue3VuuC3bg9y7vCpyMuDZZn7GCFJMwKKjB7Xx+NiX6LmRHNNC57o0lgrH5I5bbfMDpfri4+0B8dzAMEWcu6uA9zMWAZjD1dXe42/JBD4Oh+hhz0s5JA1qYYAf/ikywhex5iETs/qXMcftRrujj2xyL+IujSGLbWH5ET0Uaukzdj1E+nSg0qGussct3jq5hKFBAT6FzkUUcI4EOhlD0262GRd0LqP/czEEN6gjkwXE+DYXYqMC+ZpItzfMVgACPezlX71Ha9hauMrQQmbI5BBv5U8Ds4FLa/vRieg/QMEC6rLo+gW7FFo2DHzPDhKb3K/6cuvl8CEZ2f9QmSFBpce+p2sfHNaneAJHtcWKRf9sfuJtOePhuGccESbcZZ5dK1IW0v7MHXtUQPP1WjCx8qW6aOWBYGMAm3R5f9sS9knS7NmlmEm3AbNQykHm7CHCdeHFg1r3UvF2bQzyDo/xOKeL0TAYxNov2GIH+k0anHzMx6giLPALjz1ac0Mw0J+knganKKYIIxHSxqtyipcY+hixuvUvOsYcE2oGsaxJt226HRA/wQY2pAESNZf88oXaQNYV6j5hscawTqClVG0qz9ZtYsPmfRFzjRK/l4nMxhYOHew7/cr/7lCh7Da0CJkclPP8390GB2H9Jk4x6jM/B/gDvqW5aSNoPxEqqm2tGEeM1fnSo1tj2T7Q9LZ+G2F5A/c5/wF9Ovxnfkufx4hr6qJeWiPnY4wMfv+ZDeWhKoP0M9HQw9SMUzJJtYcUnomq5hks+6fr0wbu+mP+vc/D3kZNi1kd4saQ8lmK8TYnorFFg60gkVaiKe8/bnW3nOoMdu9xI6gKtOCZe/sFkfIatsZtLotH163Mm+W343hh+E835jwtNTs5Y1lo0MtelR0bO2jhw8a7FAS9DVMj0V2flQl07QdM8U0xZWmXs1RIOEQTSlA+53HPgFCSxpPxblLXmn5E2Nt281Iptb8JaHHxR1hwIew8UlSplH4nw6LSO1PqfLgeJ2LHEQNqHSHAYIXs5EsT/LoDu4LHtPu7g02r3lvqFAr3FMRU/VpHvQGNTCAZFnCctOcT1cCnRVHDOHed2YJS3TV8fgvorKcE/1oRdUzqFxLFut7LjmPqU7znP2XhukcEiZjpJFw1WdKu702YKjZCpcXqFMy5hWomx1gxuZft7aIXZXr3OrkHLIdmH5dWL4H7eBUaLcbPvw7IYHdDSCSWEz5BkFB8N7GH393hhXPO1rNGkqBS+4rVzuxVXkhS2UDMfigXqXw+vcDtWWgaaVJYf1vsycOtCk19RipFYKhSxqbTzK1pY/04xthmzV2fnKyZXRKIcpz60zV0JUPwyz4/K9Y0TB8cJ043qNZ5tVFm15lOSKGb9ms4SGVQixNFTKFII0VXrJUKpH90iGy70JYNnT3gSwPluXD1yc06icBcLwel8ESDd9P+3mJmbkhSUlIO1+DDXvmw/PqZPMAR5sG+Z5p+ELP41OsUppbTELmoELS5bpWeeft7e8GbxFHjcNtlwQHRb13OeE1BmmkdUpZEMS1MfzqeO/5A4MvaVzAAbeCpW5b2x4i3p2kBTuwVR0zEAQmfWB/Vvq+YXD7v5b9ZptEvqduxIipKVAXE0FhUKHj974G+w850gGUc8MzBDAkJFdk2ktgqs3ocpu7csQiavRKlhs7uJrFpxDwS6oJRHmvO+jATwVMUAWpu5w3oI2O0Dp8zZYLQ1Pq2cxZqv1002G5OovwpHYAt/q3WittOL2KRlI83nnYCaV7ldgR8zcXLbJCaej5AQPuWRUb3TyQow0gAOpzAlgpAUlNkTsbLGX6CoT+QYtmXGC+or6S1LSwvNhKSO6y0BUztdIfdsG7YCJeZXUcnHl3NIlXBO3T53ztbtpZsYbDwQQV5bLGAV/bktZ9OiMmC1f8H4kSCCBb9zzxy4iOgXZSXsh8KFpVoFjsF8t+22jVwBxBgPDmGTE2jfQ99jdE0lPNwmaDH2weot79UkBfqU/j2O8BQMvqfJUbPqEg+zYFq/B9EY7+ojZzuFsU7T0lniJA1xhG7CKMBONpY3jUxyF9vGMeJcMhaZZSz8VlfnEBH3gLv1DuaMf5AbPK3vNq5XhdTKkKJ6ozS7qWnMQTTIEd5iW6LCqlDvB4Qj8AaxhDY00lO8CEAXyN+i+wuohMfasciEHv/ps7uUdya1tL97lSoqi3/SfqcSuSDOwcTn5lBR+C959kWzpEmU91C7OCoqO4cpEHvLZpCovvfH+QF34b7ltk2LURNAYMD1Fg/uaMWXs32jlQDu+ft/RhVHctoa8Msh4KvzsSTV0PY/0mplAnyJ5m4t24WwkR10vswQq3QfLolLrMjgl3hk6fP5CGpqj3RyfsnFDZBsKut6jiJz3/Kzy+AQ6ob33Gu3xu9hBpSqD+0QhDiwmhIEscVS1HAVRIKj9+ylpRVk0kgRG61iqfmmmOmIBjuZXaOiPV2Wx/kuJQ7+B0o0YU2fDt/P2Z5bG2hpzXfIDO5QSpNHRt/vcf047wKYzpIGU4PAtIC3o4TMq4aHD2I5vEaa2hPChLrerpRRqLfTwJKu7olJkmRcO0zTAczFzkwPlYggRoR8LXJT/HJc4l190NrYy27V4gqedXwiOG4G+b79N0nwQQ/OtEwmjerwuBM1GUobafurf8r8Hqx5CbRhzn+hTi/pwFOG3omcAFTTihtZwZjilbC+JqwjqKKmW1tWZFggMwlO8GZvFcB2Pz40mBBEAJYVDEtFnngRMXbf3BNyUSjcydzHDFIIsl1c4DKn2x8wYPLrvKecdys7chXX8ulGKkRXurdh88nNiNXsgRQV2+Y4Re7Z5VqQL7hRWVnk04nX9evKcOVKlzTnIsXIRudmhHytZEeL0mNqD9W584SZGSepyfBr7jG64j8YZ12BOBcU25w4r8qvFO3F/NgLEAX7Z2gknHpRUCdK7nQd8aV3tc2jqcGk5WLIM+3V+d7kH8dsAzM7e3zzsDhObJ5+aeFOj+es7Y2EUoVU9mOVixud9Zb+veNwz+ATj8/d9HbmY/AqMYQql4LDZ2Rv9DCMuLmWgR5OFsRDIJhvP0NOXNNOoaNFRGLKpkgHbtFi4W/aslCV8ideg5sD9Rxgp79G6RJf74ScRjqarZ1OktU45gYXyla+QU4lOR2T/PsMI25ddzSnQvtFnx487kSsYfY578/v0Zpw/axUW1XaNmb4iNnxkZYoqJZHO28BiKcF39PQ97N9pM2Y2Tf/gbyxoAtKTnkMXQHe6EffWidmqObTJZxHdvyTdI2uIELFUNvuy/Wu53Ew1TY8tThiMvLBr1Ha5s3Eqsq6DsjwpWRX1K0jEEuYkEUw15LFA6JjQgzGFRR+e1bzcj+0nMH9Sofi8NMgLg/CXuJ+DEmEXAVoAs11RYCGho2++6pPXq43YQY6G+JNt5uN1QDMxL6uqL3GCIRQrMBizkltpFZ/mQyAr9P9tdIWL6zXoMXes/hzpWTkh1mxM+aWFo4qM4e489ZJKyOzGtELyNrVJO5nCH86MCyX3UhSRRvyH8b71MvynRaqn5ZbLWM/t6Iy6oaLUhKR3ikPOgQ2hoy85msFRe01VlpelYujO9Su7EJ5mvBuoR1KATd6r2rMMb2C5EW5w+XJE3ogdzcVsqR8PepBsb6bmVwVKoYvACh6uiMPipOZ5Um1yu8IY9HBxYmyVNB16J00qMTWt0LCp1RWgyBbNzyA3mNCcQ5ehY8+KUmujwBSHpm05wEvUjsYW9LWRGqyKq7gqMr+K2gmtitjqXx3d6QcQn79kTCeb+gG7MRgvh811dOns5Jmkumxq0Y0MYmi80ZbBImo4MYCNDPt7CqAkgs9s2f4qG8MayOoUG2sXCIfTMMFlpsTmGJGOxOTZSOoq1iQR2ypI3qRYc17znJeIHZXLTUwgERdFmsgBhMSZG2GqLiSi6el87BkaxXtMQU0GSS2rvbqqm0RoOH3GhgbdQUXmVIl8JbOg6BSPlq0Rl+R+FqOHOVXYEAJY01q/fpHB4dPCboi69iSvli6BxYBb1N2t2gpx1HHQlhNAnwqhphIpj4xTLiIINmWhglFU4zcb91OgKCIR2BxPSZTdY9R3HspZLC8wXZzGl3eF89uSzz+ifH5lmpyMJ4++TEprn0kPvQVddOTzAEsksCJtmaaEsJ06Rp5W5nbYsAsujtyOWoymQ6yhFZp4R3j6QxXkcTUHnd6Xi5WNVFSExIw4YovJeAPX/eD3BZoSP7eRbv/7k4szVRh47T9YtVqFYzIMG4FKh9g3w1ngUHfgGxYT5tdMhyGwR8xM6i40ut5GRxPJIe1MFPvuUduMi4891LIRMMhwnV+vppqH44p+Qcv+L0JOsb2e1/4qlMXM4ecn74t4NyDKUcfZVlR41b181HP8EzVYOxJT9uMzXTbYVNP+GFeaqnB9roDOkMHGEISgVD8VnNmGw+lzH2IYJnKTHonkzfq9NzJx8JaM3/dKvF2HG/AJpN1YCgbkXUpJ3jqH2oH/Exd/of2TWDbR1ntbt4v6N6AMnI9UE8SI287myk963/WDMuiXAGlKC9rIhct10Zfd7Tn9Uob4kLLOH/kxRfkoMn0v7I3lCBEdZ5jyz3HdCYQuAeRhM2OGePhCn6duNVMe0Jb4t1JZPa2zVGj+1uW5JALKUdiCAvRSMc2xW2qLkv4JiP/hfVO8IsQlsWv9EsoUqBZ6gSCZmkqap+5DtMdKF9j2QzVYL3AmUfblDhwiTqYLZ92LyatOpaREzd0leq7tkCvs3LcZOvqlYRXzb5YH8B5csEGgReb41Ojwj6XLP6jzIq2BPQ1pEsivhMUbLQVdqFZNoUUebJ3vnPXeiFxxaHe0SC2GVTQ0dQ5Fb0trTYP9EZhx7LyBD6k4IOv9npoDfCZH/z720Grf5moNmZr7pAMFo63VUBqKBhNmjWS+sqiZTCroWUjTTEXTfOlHdRmij7tQysdI9+/hVZ45XbLPIcNl16EU9/AmVkzqfxca5BcnfYcqs0LUnWM5NM++LtGwpNNyqcvL2T6O8Sh/pGpBnXiMzBQg5cxRJP+ooioIl+x1nemalsZDUsnkl3nqkHf2H2wb55ha+YwYxBcEL6iJXJfGYkmcQDLwbLGS2vSdBjybQpMd5P7GBrfR0mLbSZWW9JN2uwCY5GR3thEoGOq7alBLCLmmpA15Kg5bDpFOn0cxfDim8=
`pragma protect end_data_block
`pragma protect digest_block
1a89046d0d87dc3e0dd905e5543b04dca677352b2c290214211f9bda3737fc42
`pragma protect end_digest_block
`pragma protect end_protected
