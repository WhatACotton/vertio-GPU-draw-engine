`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
ZSPBXaa9xP86yS5Jkw2v0hJVO8HTpjdfXXu4hOy5usGOT1h+GYZHfrCM0osYONdyB+KTrYQT7ZFjB8+pUGDFsm3oXo27ThFxDoFsgY/wqhvBNqaMoX5BMMjinHvO+zZbTKxmSYC4M9haW08gVasXSqiQVIEORV6cgNevS4z+XKMgyP+hFH7l2YhR5rj50VUs+BXYBu0laT88IPj21lROuHmgm9XzWifHcc/zpFENX4yhdb4IcYCOmgGaZgFcM3UJz5BrFQ83iB3n5BXEk28yWuXs13a7rai2K+noVIL2HhvRNvFiBY3k3QojvgoNPNLRi7XTj9k2E+fzmyldVTLm1zg4Zq809rYP/Iu7SWcNLsupZj0bPNcv+FJ1lZF17e6gVw39SocgYFzTSPCQZ1F4m6SIObjEpINhpzpgJgubpmt5Rhsf29c2i1psGX1J0sHw/5nx7EmUXZanXSR6L+GREscPO083sL37+tAJD0xbLpLvvl2Ybejq5/RG7wdUod54K8jn/PeyGsDV+OFyrEwBBwvI4XNwtjllR/i9zOsMeXLeaV8O6QEjRhfaX76XWDx9/3hlIT5qTspOwU03ltJ22+vsPh9WvqMy6wu73aYLAhP8MylI/bsaqx8z3XmqiAoyomNMjpkODWtiPLgjCTuH4Lv0uNDrIV7OjVsZv/4keSTr1TK44uu/0dK8UlBkkzCIEpR9j7+FVZHKzUQUBCUtpfZv2e/f7jVCSEE+wAsWdi6R1TQE13yz4ZCOvgbrN3/jMy5NeI5nXJ/ny6P9n39LdTiB3eB+9JdIjxfA7WhsjrHVncWW46hO8Z9ZY6a+1ONto8vihCv8AuEFCKTmJ6eb9VroQXXIXg4ShQlyy9hZvBjejKKw60aXZfKJK+vrrIgQDCdy/jBHQtR03IEF+Lhkl9ys4yvm7Dpw8GjBsmulcFka5aOU2UjgALiinHd92MaxcjMTxs/Ga/xL0anwdFxX4sq+fN46Y+Zi0SyKNXnv/dXNYcV2MEkBp5NO65UtRUhw3uB6usK3xHDF7Jeau+VMx3+XnLg6iAV+ElrtZru53AoqgA6kGqtvAVxi0KIfOd9PBLm1LPXWCPfoLLCEty3eIyGuR/e2bBljbjVen77cSnI6BWr2pQy/Dq6VotzBhGed3Ar2J4uLQXc/z89NTxF54/rMdORvf1ztIDN4MnJLRnJLw3XbqhKs1fSuKmS+5bQOPlm9LZOz1O1OwmA6cvWBfLmSQ6d+EtN6nRakRgTH0NsIvNYtfs4R2T6gg3BHOXz5bIgnWyHe2CZ/n0V0ZRkeWG9h1LvnLfrmPy3e5I6vXD5vac33ZVHC8X69P6JzB7A4pyiSyJ9FYdlXaVg9ePu2QziJEo5x3713CR0BGzGXoGRBEqCBXUq0oZfIwYatco+5NGbIcXHOtFLvfbCZZ6aWv4q2D1gcuVckhy5C2/vAjqlnrT+SmsZ3pEsnXPoJOldGc06r9/MAM/NpnHA9gIlEwk9YpVDUC7M9tnQA4IFcVCObe0ZJj7aSMX26+ZhPxDJBnf/PVQKTKcRIpPXE3ui4Wto72qEIwqyOsEDYZrTEqp+Qq9NzYjNGOvD19zHFa9eVjKQx6j49mDrMfz0AI6x7tj3moZDZgQzB8AzQdtli+U1sjasa6UFJFVtgVW4bXIkwgVvn4BN22SE35aNOaGUa5eErc9tU4ouTG6nods9tx5+AjgABJfv8Zj0KBC//HYpe+G2wJpgF01YfGspR5b6iH+f9V5nty6gbnSSWPDDaJD9xgQ8uxIuKq1uVaDKNu2gcXovyuRVI2F97A+aGYE656crE+rfEsib5Hcx2K0Dtlh0T7FMqSj9ll+9610bP29E2brhLeifbBjMzSy9cpZUow6Im27wF5RpszP0Ij8eN7hLgBjtoQ/Y1vhxwsn8A8B7WwODaRHrQ5GMr8C84hcCJKUIMK/Sa1Sc8hw8dZ7IvH4KCt38WzqzIKiat3kJBYADXuknZI4HbMFlMUygyVFZdMffNuFIa9viZk3EOsYjUdd9tFsu3wV5wws+ASiMJLQaycTBRDtK3L3MzG4NGYwtZOncKvcTGHJDWhFfP7ctGSDBNsiwwEBiTTRabYz409B850GYkN+VfKT+fIvH5S5UWS6FYLcaKUTHq2MkF/NatYYywKH/nuOLGc6PHNxXW/BQ4IcGaK6NXvNrpi3gOusZNcCHii/UlZtHvSiSEfhY1PxSYraSZItyFzJZNCw7DShB7Vzuy7x9H9/sErqqYe9e8gKNQmqFOO0uJZhybk3C7Ke/kz9LcxUn5UNEYKcaPoYnWv1sb5ytqJsBPDRjb1kXwThCp/4Oeo77K/CQH3O5tz84QfuxrS4sBQ0WSQ5Npw6o/xt0tVrdBJIzVzb25aN9YH1ytk6+kSb2co58PqF8EpEqGkmQ/SjMHjEgUcSC4YSq7IZc3OszizaGJmsoQg4qGQNz/YqKDnOLPCI8cZLsjP0RH+aEJZrVUDqs1RKEuMR19zv0b5Q2ueJOJqkxpkWUUa7JKlntpbFGXQc0pHBgHT/lQ8+PLGVpIDXvrAJiQjhzLlURsFoVfxPUb2l2fLP4uTbXssamSnPL4OsEJfgVrP/OsF4IceSqw29pBDQhlc2TJxNyEybQMRH17Nh6hdrrV2ueF6Tavv5PnrXMBeLNMhuxTr1th7ARjiUzCZfDj9b5PvByVVygzpUKC6JAOBIe/eFq5PPnxb8nmGpAqVLCvDPIaKJYzW7sq/6FOGfmMhyeHudz1j9wX4xM5rhb2Zj0lyG/nrqlVeEWsjCkMBv6ynzYhtdooKsy9J7Q8NxriuPR9aqASjd8ijf8bk5yggUtoWirVPx2B8v6WPqoyOMy/hcjsjS+QMCUfwlDs9P8LGR4pO7Ceyx77f5rKevem+Njsr/Cw6vbV+wig6qTJJ9xhhYH31BeQVc22IgTF/WaPlK7EOJbCEG/eGYublQrT70CWmRYxwnIoPzJxpHzbZhtWOiBsE12gtVP3nigkiu8RYJDdU8hoLq6R47cKKUwFJysfz/pSNOSvvsWyOx8kaMF83/VqQcq6mltVpk5a7fThTPD6S7agyjR7J+w6QUF1wvhXTd6k/j3AAOWjyVIy6Nhmm3VqAZVSK+/of3WCHy3XNTnUlUKXd4vbqCDCxA5FlBif8slD+fj3P81qs+JJt0ESSaYzQDcge8YnpI0zjm5xKHeqU/DCZc8ctwbFu/MOds37cjt8dUP4sgx3u2grkD+gTTDs12I8RWASUf7n57zdkhRnSHCm6fE+DOM0ZMoQ239tsibubw+Ctg5KiJwZMfT/BBnzkzHtFOK/VPrkUsxJMYgRt9k++pTLnFlWLGIaJDsUVLra1/dTlPAfdyYpOcsqp6yyBNvO1cjQnwfKlf7yWYlKVe0ncz3+AnZ0NApc9Lh/egP9Xj9Bv8d4onjrVUAH/Uq/NnB3f0F8No87AZ8KfI3twks2SZkS7hRtQB02rNC+aA/JKX7wgsycKJukOJSR8OYoZJbd92Nhg+sVxCwnrDDhNbEBa6Pq4Y0uzZZ8cIx5PZYLx2H+5IFp8UZtYVxktV25Azsb9KY/33qb7n/sckz1G6kU/4eOLLxwbnq+Sp2yYrmnNPudb9FfCr5KFQF7Jzf5xjEi1XoJgMo5+G054EBwKwjzJtMkVuC2TWuRY+EESo/5Br804q2jKA64YWaWNYDylLUf7E7HzIcsQo8H6ppaXUGynbsZkZQPSPLGL1QF2rR8pZOmWKF8kp2HcYKAzWpnunvaZxcwWda8viH7X4NkoRRR0Pw6CkwzHNnBpaVqNVAk4faIzE/Yk5hmyUmzg6egrD3gvk/fNu2OTbp2dtMDfH2I+VVgrl+NxKgnodxzi1fXgh9dSm9coAeDIqfXKPgwnMxAw/BM+5tPEuXs4KR4iXsF4kFpKNMx23nvGjQnzFgSDfszRfuPzV+IRAYMGat4ta4Nyomuq4okOp8SJH1Iv+U2AEaLNtSvlmXWynTx9Q9EaQA+SRPwxlnmyMVpFWE14NtOu1jk0xATyAl99ZLa181bvp4hpz4j8JPGkbM+DmC7qNNMVyvzVUnt1RiSf2+tEyFDpyPdf6PO2ik8XE7rd4L2es2dHRBbz0HTvPtxqtpxAino+Dwq/NLAmrflrVQrM/vmQ9Ma8jj0mfFGAR2LsUNJxYAx6qv8pCzrewQtXECZYZUZJkvLzYiHVnaGyWOZivsXb4cb9/5CXVbp7TwFy4CaTj5o2jWtFmf5hw2NkB7z3CRJxaFmHrffX0tr8zpDz41KU8iSiw1SXg4y7PBSPEmCqFOaYbhpoFGgZtO2rGmchvy7IgCxnzkXCU7u5h1MVygv0H66W6bOnl7HDWhVehGWXtnmC9ueCHQmrUTi0F0Flgo/1MqSuTDqDNKyIaKFp0r2jqeh1a8Z0ds0sRAgK5cd+/9BL3E8nl3Rz8lSkCiILckUEjk+UrK976iY00vN2WNNXwZpmEzSBdKtcLfuC6V67ckTLSD5yFvYmAHRQHv6OajHV80DCjjM3cldq+touJopfgpiibYXPYKdjmPr0ccBtSZ8eiS1f13WyabgiGwiRky00FgReIP6oTjCwL+aGOu/R0P0umG0jksKqZis5MSqx7zddlnLhMeGvHYXRGqbnav+BVHu5GJrXdn49nmCe3VfXLvhQaoUgVFC6vT0knJYy9LAPtPsH6K5CMf2W9JoUbhx1d+HUS0vEpu/1hxvZLvxX+hwnnn5hAbKFQrf3ly2XEq+/Y8q9ZxwCx15FMQhqFq4iNoF7siOJb272ZGtiy0/MHLMNKOGaWi+897vrdlt7B6Zte++3jFQKIcSxLWiKh/G9xCWctpjXB8g5XewukQ1ldidiVn/5YSJI1SBkQHKUF7nNmv3tXmxm8+CPFW3UVE5jb7HJrBNdqz8O2jtu6tetwx3HtVF1W0By3oe4KhcCfCvWdKx1xBh5hHhQJcLyGHsKEwEsCQqlMnhZ7zddCmGf40yLRyRKsM0cNzJB2/ssqKb51Zzv6sfhtbWAvsy5E506pJpV5V9IA/B2DbcTiQx2VpVOFhYgMrjXc1z3KLsVQoK79wiXbDPDVabfMmREukQGEWK+dB0IDEBOn8u0Ug4sB3ELv9iSSRDyOhqy0tbcqt47EoXi0pGwPVaGFQNEqZ3NLpyhvQUUSxxCV94Wsf/33R58x0RIPRjskcasqRAu2fnDiQwtvp1XtOPxJy+//n3qLUmu2sXEJhiJGpK0tDYFT6bPT/ca8zPeAU6G9d8tSbDZWf4sl4NDT00WJdC52qC0R5f5Pc1ujITxbPMo5J9AZr2kamnau9ceIAq3S3FExeAJsDcFd76hoDv4T0lLxJG2PqSlpMpRV5eR2GE8oKJDkrTmKrOJtLdBmZdFQFy2kGbhDZpMga+jpcsJbPGULrQIbUXaW6hcaM7OYcifMg3uot9ASO9eRSCXtst9Tji73h0Rbyv8AlrtqtLUbW5DH2arCyzkhT8GGdPje2E3fgK/jFfFY55jSOjlFVSsqA/YmmD00UjV99LIgb1xHZZ1vMVb+n4hnnII0sitv4dk+bEmYdNEpvSudIu+E4AhzkWvH0HcFgdoWgcvt2KmpL423HV59/CBuGC4bvBY3sAuu417VVeLzyZy9gYPQ8onJhg8jvv33/mvL4Xt+OreFmbnOJi0Njlc+vx5Rzrh4uy8IaLaJxgqPJhGSjpedGNFNXJYe4FFk75C3g3BXIFERQCKIPDcr/9tj+hxUFTJO4/q/8wuj7LHGWvnZ1Ty0NXhjqGZ2Dd0zshtETET7jrXuKd+GI8U+v18N20SNfLZVltej2m8UmN97+Y9kD7d7MCjV4EWSVKpgrysHUvKG2p8JIrJUId3pXLyBuDnsyo2LE1qpho07ClNdUClkWuQOT1h2FJc+XXZ5jjuCO5AdLuwVPgA5s9wMeITf66tMUp6+345u1Zr6bBWqD9vZRO9uFcfdz5jT6LeHjRNtbzviGLLj+GinUmg2aCnTZC5J8kYQ3+jGQv0kcomUx45Hjm6S1YRBRnjBlbZmxZwNdjvuOvdmSQXHogv3fcDk88+YR/+I20mpJteemiPPIrI5mP+NPMTc4gzhxVruRqeaDwKYzSH2WZKN0BSkg2rh1EBoNFaAKvwRtj8DIbwkX07ohbuie4++EHb1mcFuDHxO73rCvdimY9UCfIN/b2OqyuJcjVe7vETKnE4ic5VqTmhK3njWEoHXQwH/W/QNemliNgKh27CYT3MTtCQTb7I8vUvo2npILQvL8sBNrUOQM02lw9+t5NIcCEHobcKgswJ5yAADdUruWqkA6JvuLVjhhW+2i7M3k8gyV+aZ9ad+s0jyao9RAQVEapiYKLlYhMVVc6Q+crud3KvX4G9TjHhYa0la9tPYhNe8Y6PBkmyh2eXMw2CaPn4RogJeQVcJR57JaVsSxr7cWgmiMUuA/MH1623KwDSG0WdPEpxIK6NcZQtWkHKQuuArjF6c8ntIgPckgv/ouhgZp4y9eJaYY7HtXUxvicHbYcIM6HN4ZYpfBbUAx1VsvMAP9d4leuihLnS76AA/Z8ImkqJ8eScDY5Pk6Hzd8ZDE4lQ8kwMo2FTN/AXFm8zQVniAMc/pWpqmWVUv190EJ6QdEUgw4SEB/s4bLD61QTuTKRcYVgay16+aDYQYpKxmpjkOd+aqcLJUSDkAOZ8zLXQhTgQVfZ6WMHjDTganxH1IA9g6TQ8q+CXtxILr47JwmwaRPnMHzmI0MhZJou5D3U3DjAjaRsFBpMC1J556Nhtt57Qwp7eaHxmrGNBwJdb3zZfyBoO3mR8lcnm74XMTh2+JWQtsdBhF9QN/IXlD9vSImi2Z2/x9ObC1pMGwxuAW5PVGf5bGzDGB9fe/DtKaSuVraluoAw0CamqzuxD8q5+4vTrXX3kq2UeGDIu7gakKfcHTIzxbdtHGtJpbg8EkDVxcSUnI0hy7gwd+pY5O7ZOUTe5Oh79NPOdNorjW37do5eFkY9WFMtmiebMV8IX/cD2cOHZE1qSpJxJtino5pyZCuykvzaTw6CQ69i8Zh+GxyJiBdH8sGjzwMUB+CtOHsvKQYZWGBeoOHUkPBsp4DPBFT6gG7nwVjkneSPrhqSePxEXysAd76r6bg5253piyIkWdGqEAHq+bRONRyrgMUD6MO6QlnD93JOUIWbOqRtPyOcXUTIG9nn89pEF5LDG64ajwrdEz69mxMak8dkkEh7Fgv78wNIY218I5YoysXAYF3XMc78PEWTizsABdbQmSecynnU4pNsFgbxiP46GcUoQWEWvaawN+x9LKF5MdHTouRGhWeinrED+cz0jtfgAj9abFy/McBB5+H7txG9/ay/CYvMA9f1TUO+yvyw9PxeJGL2e7lm9327Dqyon8r0EcbxC0wtK83K6BkZvUgbUvaI0p1DTPXVnI7B/2TUwM6yA7tpADgEMqbNa5qf8h6sUXnEsq3zauM4HllUiTVE1bETFDPviZbfu/wUjUKmDZivlXOOhI062lE5vrMzhklrOHhaPD6A3y2g8dUCNuy5hZZj8yYIUOelH5073XXdA1Kp4P7FzoN1DLN5eNokcfZ8ZWFwTeWCCVEwaBxlD7BFUtA03xt5+UOow9kxL7sBH/R9qTtZ6hUqEDrxk3m3QvFCj04Bss0+KDUJsWd9v0hlYwNy2u6It4TpkfSnup+e9zO3xsf/0KiOfGs5yUaBByRphKyNlUZVLD8F+tKdjh68vU9ORJdTQ+FFPl9Ze5/zf9LKa0bKp0WUbwq4vjxEvRwrXbyxFqJkpZ2K80PcSb3yzYwk2BQ9NnlVM3cR4AZdj3QPSPkEIi2KI4GIycY4TWLqPrT9f3W495noalv+ZFnLXXIbatMm2+I0y2WLTuGIRQfwikMC9bAuSVh3NERVpwpB9KwMfMEg/873hrW0lC5tGDxT2F9/vCM28VlAURVlvBvZSw7OINT1m26ifavR6kUpoK3MQ8IYHGoO7Rg/tv4Rg78vdpEkilU3BWFawot7cMduZ2wQhP/NQ62WwiJ0ROocze4wec8M7O893MK22Hi4ipT57BffCDhp2H6lou7L2FqnkWpEEO9gHSdkGkkqyeD+SyvPRLrQZ0v4go/w9LxfW3VU+u9vgb4xDtBedz3ea28+M2trjIA14yb7Q9m7jfj7ptfHU2ZfCfRVLEi4djY+M4YXOekDpqPKIHKk390hong5LxZgnKPq+qUpGGLoaj8ZafZa8/wBhoFW9O9KUJTUHu07C6emWE0UfO3GLBnP8Tni7RL00+F/ulP3D8ar3NkrjpY4gDAiRS+I789RDy1Bfqn3Qkd5wZnbmY50zMMo+Q+tOk/hAmGhGF1T8jSMSe+DGxEHJ8zts/gCkrZTiXTvKwvcDidzbdEBX13ORXiQ5d136GnnHZtrbcqwCDKPX7l2uunhiXXjBZQsEAnTA/QJZRcP6st+BygZMFbExd09scNI/qkfxRmK6WGZqvou7L30RUeu8gzHPtOpq/DFuUqqsmD6DoncalUE7aRrMbCH6ZqQbmT5D23PysTMTMTplIHICM4Z6Jpm5ETiKTlodc6SUd0okLgefjlLEHpkbB0hTLKCKJKTLTq0dRGDdhhxwpQS/tpiF166FDgmPzWFGUtsBS03fdM9iL5MLHo3qxHWBFCWSkn+ybieOV5ORqtYgmBZPfcjWDlFN7yF6s1mDCsHGTDqF3ol3KX1ePDpX2X0BJguIvkdK3uXdyJ4FQ3eQDA0FH+GAqx/Z1ECQ31YNnfeahiZvtgKdbGWkBNGh54GnNIVbXfwk29XAnT4BYZZdj4lPPPgyepj84dp4dacKNnMozOfm3YGb3phF2OxZXAU8VAIFyPxojMewVN1RC4f35r2hyyGQk4WFICPL/kEnkmWrWqM44qUYNs38CEFK/gQLHwakDVEkJ+S6au1PMwz50UVT95sgQKSNiELl8IFoSNrbzMU30dLdCYWpfmGoNPxvzModSxTUqvRwk7uXtWeVFbFgUNYK0OrhuvRPuHS4Hj9ljrQ6RN+Q4vnQmc5fVhynnzs9QlRZ/ZOnjq14CcMrlT/Q60ql+UvJZER+Euj8fTvx6roprzMLozmmc79SqPwqW2DOIo8iQNQXKF7mxgUVYJagpxF/MZufB4uDJzPwG1K6FonxR/pP2Ru36XenqzVLEWfOQVhPZu4xj2Fa5ym2SxQtcfVamyOK7aYhgwpccKrwNRmSIYLEgWLKh44ceL56tTcrAbmtOb6yNjVBYROc8C9V9bhChCTPaXxSa4CESRJPDWx71lLLAMmTE6fruopf6XUOhxqiss6bgRajadvsSnAbnrOIc5rLw+A/Xw6/I8JN3ff8nwyeOw3LhVs4ii7k4qrO63miF5ZXI5D802TOAkdxJYSp3IwKpMdBvK/7qE0DiVipi5ogkgXGODSRQ0RHvUVKsqQQ2K3xGuut4CPtP0VqW4JyGmprgXogwBGZiLUfIGBzEi3Ds8eivqzvXZyhOYKx3UBs3qRxMXcVl6EwNygWvpIQNEre8iDAd5iRH7bGZ3w1PVLipkm+UZakU1Ww8mIBG3JSQpQQq2++eX2DaBsfCkt5hHmGJb8VA5VfuM/jNpZ/KVnFpdpchk0euJoqYciGR7wuIwoXsUHpd4U3jDMXJPOXe8+e8OR8698zu9mgLI/AFl09BvVhxp5msXjm7p/8/cbNhc5EB0I/rYvvcDoK4g8nXha6EDz8pcclgVXjfQRcHbd1hXhuAHE9flSIh5ufAdZGIUR+HYf9WeGyXYzFnMbKSac9mHZov8+n+LsiSTfnQ3stMu3G4z2RH3M7D66C2gv7fzY+CY6e7GRDff3Emnv1p2fGE/ezfMUj7PAKa2bE+MN/qnNv3/ZFR6BSZ90hRfJeeUjKSNOfEes0uyLA/s8T6CiX4Mx+hOB0sDG2uniOG71dt+Og8G4S6e4dBYJm48EEdsQ19q8PXYHl12Sp3ELzbvAxzQg9h1NpB1cC9pEut50HBMs74r1UdCzT4vtcvejAuarfI2tguZiz+7grHvkWD2uk+Zd+XKLUsoWQ+akaBsuxR1wf3E0108HEG6bGpoNPcYscmQUYSO89l79RGMN1JCwqiq3d+NCB7VEEg8FAZ9cXm4QoIWGckuL21X1GJ0fqIHl1cBs/WHnpepT845Zm24U13MBU7BHH8hzebDioR9hNCRkxBl+/vdCAbj/7kisirOW73KsR4/tCH+agB8ap1Pc4mcy+LR9ddBfJqU6S+TfEZttXVR7e8puakrwjPLOMe3Ky6PfpMSwRQhTOLxX9KsqAZzol66AaS/q55LLUpoTTGaKqGMfJRRh5fvQjiTz5NxzPG6jgpv7R6lWc0aNyI6zYUOyLjxbxD9bgk7Nzf5LmDXoq6SlUSv/bQaYaamwSuSDWpge7YInlW98tggznqufDNhA2qLe+iw1j1imP08qUMBN/ctC9/8I7c2/F9ZK5T+9yFpA8sVV8mhW1wPMJI4XEHr4pduLCH7EpU9AakzSNY/VgZ83ckri1LL+HiLhQUs11/W29SBw8ZFQEfyrnkNdsRK79uJb1I8g+Mq/nJ2INXBYBeMmc0eiMF24WMcZm9jDYaJZ4RxZ25Z5g6VD8UbiMzgj6jZtFMufGNxJlQ1GYw45BEkF4i4+Un2RH+8P53f8gZ7zr3VmuVs/vxuDdxLeaDcQ8uq/Yx23aog97mg5wcCQUGANSkca+CnxbFlmu/BY6a+TYY0zzoPB7P//+CYs8WOwU1O/GeLKpMOZ/7mPKukf6T7rqjCsIWAbR/U/MW83LQnafGyihqPJlHzD/Zd4LuVD+3W4+8XYv09h5Btys4CRgVOh6OJ0HGxap/ugtksgBG0IQ+ul2s9kKxtDBQGtJZ1fHm9xfNanpRy+j2epvwf9mZgv7LzKBvgcLz+JYbdQkVExqCziz5jFyW4IqI8U7PerZAtjodt+naN/4AqgKDPEdrAqRXHlXmsDh0UGseRAm5TA32lE+pfYdmQGqxiinSaDtVNaxNKIFN0EqelaZqMNOFtC7vvXY2QrPfG//hhrYlUpM9c7yvH+NKuLwJJ/MqmMCSNbHFP2AmPf14VWlYzLVjRAeD0DX4BF64ULeIaAn+Am4rHOSO4aMjEzShb6p8tZfHZkrrXSElc/ntLrXtCSNwkZwDjcYJDJaBH8OOF0iumnJv1ePCezbxRfc++GKU2x2hO8TMjpeKLl1qdpY7Ydp5hRW1lg+ZPVaYZbqKHJxNDNILkUOxYWNAjv4wQXQKPJxuCNCYpIO6CqaPhjzQzXGrVP7PpJaP7sHz4PAvuWqfftbyQzPIafo+NLUYJMefvcz6/x9qGbmposCvQ+tw2fDR1fQCmrIkm9LXeQAD8AkN6Qs1hA8Tk89ufY0AOG8jllT3wCpLUBDznDRHjFyTJS9nYAuTaoWXTNCd0MtdUqvH/KDYK9dw10GBQrO8xkVjWbGAod7ajGzbysdD0UDZUl5hcXcw+LWGyRseZZjBmpZe+VMASe+rhwD0V8fTP2KHWr5UrNtebJaGbCE+Y8qIsRIxZYqyAZFcw+7HV7aqPpkSARDW+mT9Q7Rk6CTo2HQEoDMcGJVQFNzu+ZybBDqaOToVcQ5cAfClFMSSo2gCiaUMtEaZxcdpHzp4fQpJ6Nbhx+Agz2WyDn/z+fYE/BljnugRbcGatWnDtG0tNHG7v8luzrJRjV+puktAHRqGoaj7vgKgc7kvpjy0Kr+cJ7jU/9uJB2FQbNjGYwaxPaanaU9xShq476FCSTvfoY7mZO9DNLlqWHcHiZZFCovg2P2yK7q/cXwv1/c4oZM43NCVA1Sk2mqpV5kX4+DXih8pvD/+QmUSRwhj83OPvFHl0G/30stfkKxU1rzTd6AQWzys20o2S5tM3JY/qUtB6hLACvy9Y1a9jN+ALYZC6KS6caFyuFZdgZWQr5OsTC1WPVkDVHxIcVZFcL+rXwYD9ILFhm//VkV1zMHD9MefxCozW/XKMsPpBPiQNhVSUfvsEa9TcicmF5Kl7Zlst+YLKRREUIhg2kLeKpv+zNYh6FKrR9zaGb4bBZNme0JQX+T24rqJgXOr+czn4h8JEIJO2VP1uJHtEKuKN4gITy0Gr/lyBFlwCNl0tpS7C9fKv3S2oCqd+aN0sqxPbi9XJ3RSOBYcnaRoRtQEXqHbLoop8zAdvBgavtVogOtid4jPztzyRsy6yDWJ7CfQW/2ey80WRaXNjsIKA+NI0a/SYwPM6zkDgpQYN4MIDOGnc9bA21EhanK77iaebhU7/9N0XSmTfvXkhCGpQbaAt2As17eIw3NtZscSLelmeM/MZqrhfwb9pZ+38i5Vpv1D74EBwJErg1cPoNO1I+gC87/sPIZbH64uUfbOXzuQ2fNW+SplhJ0z/uHb47WDeN3ZW/F8TeXWZjXhybXsohKbalQ4c9M1wzC6gurb1NPfwrWJAqqiSiIlvAPLSkYMxArfrHk56anJ6bxysVpnxrLPCI3+rSh40z77boA1v2/IDzt2Oz+V5WPN1BUEfMX9xKTcKDjz5fSS8TJ1H9rIodR9pkssvZ84F7+ABeEGem6Clq7n4fapgLRAICnbzBTLWdiaH0XhkLFqjZJNy363z8yzNt/+vFqvFMHj5unTmm0djF4U2sMaaBWq8KdWhCjiUnbjzGKeNMb1m37T1ng2NgIhFXU6qllGDmBEABfxExU3ZYIjPC38lgTF9E/yc//NgjWvTtyPCVygGv7mrbUk3aXtPXYDHh5WZDTzNDsijjIZmemWRBJD69Xg+o6Nqp7/ep7zbivPtVl9eithj+rnEN3JkprVzO1O8HtOVTtV30npbkiVDzw4wYSJdxVIPRgajrsNJjlC8Vb1i67ZoCOHiUuOhokyUpSCQVld8=
`pragma protect end_data_block
`pragma protect digest_block
492bea5d64e0cfb2ad809c430716c87efad1cc23ecc9c0e051237dd3e8dfad20
`pragma protect end_digest_block
`pragma protect end_protected
