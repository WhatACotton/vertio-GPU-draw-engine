`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
AOMYTQoYWbmfugaw5aizIUDIeLlhQ7UJ/A9YDIdRcHGiwkCknR9BFQHPmByyARS9vHuO+s2mqdc8FO73nW5Tu86/fPBThOEMe0eVqtDUPM2ePkV9AKPSs5on/7GSwuQrxgj/itVur1KGNS5SFslIjhrucMPBAXYnpC8CY4IcKVlXEq3eiVff5xvTiVR0+xwmwpsyFn+bKj+UIxmH8m+kPMM9yS682xPCjDewgXkvmsjJV75xHESvoH/f71Q68Jo7m6zXVf1wVoZLpdQiAujEi9lC5OB95iRaFcJ+mbQJqg8YDEp8qgAWTuarrAiJAmOfBmryA6HLeMr4YX5SfxOnoxv8iTzSiwVuHFCWWQtGl8sU/1GD2ezuConDL1VIVETNNCFNxPBNwu5SgGpvywKsHEZaKYYAppPHRxEf/mNUhB4Ku7JTQfopTKJ80FrzTddHgEnHP4tHxa+yiITblXy5D6Po8i0bBEqbtvdDZ6dFABs2xB1XCKPtlILTggu4SsQvQKhp8kw3fS/Dlz6KDOJsDAyhUF0KkcCk0klSZdPmuQ/Gh52CuxHBBFVAy8lqZZ2P0+HAqVhGfCV/bMDb0/pQRTJW9KJ0NsjIZijdGrmXIZb+zWvQRqoET3LJCcB7IRSBXmDdB+0SlU0vVQ/93MoVT0iXytod/V42Z+OMJr9Bc1qnqgsRvJh/c0v6hDFErRvlStlAK/G8mRzNrYDXmSTBpznn5h/2aeh1IQHuEksXVXvelVEIUAlTXpBVMeEN/y9s+9EY94Q1DiG1qN0J6ZTJ+qpfkrSYA3G7e3x3GiMp2q4Ot4WdpD8jCbFrpcMAJhTrd2RZTshOJ9jXJt+RB3Qdr4xAjQSH4ZCe8R55OlvhQWonR23kok7D8590RyqPZGPDwlfCYVs4qCT9a0dDAvn8TLoxyvfEdcwhwj2nVAVDAciY6FJU/uG5g7+9PKsw/JY8BRAqAq+F1bkwZLxGPW3slPgymwAB02lLfiLdl4W96VxVkJJ4nAn/kAG69liEpuovLZMiyN+yxwcdeodnY4KvK1OpDFXxuKBAPbaOXR338PPEGQFB1FDkLTh4pfNP+3ArzDoHP9tLwq+AmAjk+Uwl+HNo3u4NTxwX2XlsgtlHs6YZ3ygksZEqCaBu02WjaPkS1OuQCTzj8bb/Y7fUYFvEKDsi1xLwhc6jh8Zx/IwphZ0zD6hu4zByayHrT7yn61ZwiTcuA1RospL9Bpnwrz/gODwcS0a0bfor6gxDCLC+LHxn5XuZCL1IHdVZUInL2KoF4bT0H8WLq0mF6mWHFPVF+wsChIKgD/jOGgBg3Zm4hatU+0nTo2Ws22DgXYPI+o80cVx4sWGv0BtqCnTV14uTUruFk9a59Oj90IiL1YlvX//mQI8KdA/YP7s+1FsUOfBwe0pxECJD7NlFma6Af0d20bx10LSHVKFfCQ6Tm2mNtH55wRnJZkIX0ArQ6cLaDj8IvIRr5pkotNia3qxYs28wnivWiYpWBWD5H9957aXUw0SJTLFgjpnR8eFgmahAj0ubWqB89kLwnJsf2MSngvthzp4Mw9B9vPzMvODVQUgjlU7caCmVmYPM6Ys8WU6Oj+msMiD61WRjzxyK2Ck6Cwyjj7TDK4bzMk1RA5P1sGhFALJAAHuWOjQ0U5IA1O8R0mcVDVOPo5Uz6c3b4JCcVwc+oTiMJREy0Mxge0U0j29KV/guaOnJwd57s4JiWThvsPkmO52lBWHjVfZsybqCsS1wWyA/BRKqC+p1HUg0GFZy6SmBdEXougHvBHmHuUu0AmCEvFLlinQ5Socpgy3bCn/9vzSx61YJhrxx1EZ+JzrZbfxZfhuf+XmQaSI0BN8HHONaUXYrDMUG+P+NbZ9aeRadJ3vGrcb7jtY9Q4Fr7qgyX4Of/WXbwz5wIRRltap9omjfB8CGR9CHZALPgyLhCfAoBpP/TI0uHe/tZLotqXHLGKVw6S6N9wE1ueMdBo1cQFVftyO+yB/j/LBWv7Fw2JHzhTWtTGqmPtDZzvGryEHlh9UTtFlDAtrKGGFHFLBmVTMWhEccwvI/tjnT5KqR3S4CCHzTI4L2x5ZHT2foBbcyDQuF+ODnyLgAbM27I+N+PTEk7gGrIABWgcaN5Z+tp5pnIJC8NwgnDY4C5Skmflh02kVmnvc/nrjSLxl3/Hmtf7VB3aXlhH1kBIAlWd6lJ/8TTnlEoxk+WTL/3sjuzYqksYC1IWh7ljZ/ptZ/ysMOpftD/sQVQ21mq2xBnlk2sEk9i6Kz7vUpyHhkKEbMHpT+4hmwAJeUPZeS8GSxjEmOXwYYlGLCaIfUVV/HEqxhxkAhzdH3/kfUjc5h/BK2CMLhg9weC3INie41D6fn0pTBNakGRF2LhOsuOzOgSsjJfc4DNLGKTdAAh/ExSoqygCArsp7OlbvQ3fx9RGR0AfRjFU0Nfn0gt0NKm9mhvwykRqAEBxklYS0DOgjhJ7ztjq3drzPT453uwTQSOTWgPrOdBCEAso0qK4Q7qlYRZJym15qoAYCp155rHXBYXUMe29DhVlJM78sAomQ/U6Moyt3shNLHJO4AKdE7igP9aVfKn8AkpZAd0R0oymH5igu42ZjqUeGi00sTGwdEjmP0Nbrggw8yIPpQ6/B4xyEIzlFTbTvS/r5CtwJEnLsxnngvF66+n2OQbMNlsGkRGsK/lsRtmaO3DzqOgv6e67RF2UaxNID9UTIpxNMXD9emJTarhdmG9UHjgRKqEZvlcoOgkvsLiH/iiIeJoU7oiaOSch++ASQCH00ziaqQAtOt/07VrShfsrm20MKahWSLWj4sI+6fzkxsM4HHGmYa4BF21GxW81ZiNx0+bsXJiK7DM98GYy/Y7RTpFOQ1hzOdehO3Wl2hr9Xcij5iRtAgjR8QvnFbQcmrnBvGw1gaAauXVEKPrq/bX7ptaAt1i1ODu3nSjDo2TLK/YDNBQsDZbVONMX8Xihg+oyu0eUqN/048cAFFkUQ8aBc/Nl2tsYrpZaald54nCHzApUrP3Lws8AgUvKePwibp3wCkZGTnM0TRHHlPEowjAW92DCkYswPxE9w7YDt3NtUMIZl8KVrcsA3Y2LEn4zz5xbaqBt4ZWzTH/fRELE/GGUhlu+PmHPrszIHH6Ob15yxWZw22nAiUpbCfJFmJeW5jMRkbz1b6mU9Sv8/f/8pcLmFIhveCD5wsuibisS8eQ9I0GGx06k2Uz1exKaK50DeUxF9IgcxQPyNn6iJLkA1AtCsgoOTru8Qrn3e30clF/gJdizVBw4cLTyfxVqem6uR2Upb9aJeYNKGOh7q0d/emtpEH6buc8Fimx9UHOJhzOqEwykCTKvb2JVJVLUQfbWgbLdmjgpKho0/TPA2SSDMB2YrWkNWHWFuYtQrGjZzgCKV077Mtp4ysl7cRGCj0nKmHLThYriEXvSKe2Go5Nig0+rBB5rdWBHpmhL7rCrZHIVeFAIDxJqExLOoqODnX2wd1O0tkeO826XFuLDJFFpouv3JwsgrEdI4jYC+GHZTBmWga/mww1SfNprHVFuXSlCkW7xbR8D+dvOlINLk2YGCnkWaG8CanzcZq2GxQFgnIz6BroCywXEiKJxZTdI/UugHJ8Ow+EJLrSM2SQpKXV1V8uckRvxEvr72r75bSzFKe2iw3U+VdPjvfOufqgbS0aAUXeDZ3VsRBVXq/1MqcZDE4bzg4gpuk+aFcNlyuI/gK3HXmilU0vURJlB/++l1Ei2sf26nN+1f1T4ybxqXEfgkVwMRivYn9svmblRzvNjudx5xSYJr7eygqKA2V3Jmsagyh2/jtUPEmoPt5UggHqaaq12t0AaR4jyeSXvkY7tGRi7hYUFG2jcc2DjqlxkCOFYFA8vz1eoFMEeSATuAhcZEu1hJmFfb4WmLCSnSahYwKDIxQI0EkgrrWhgHKMtu8IHGECttm/0fMYYq+5YvaIE5Ni/aSalj1I3kyVcGVX1OsYPjBvCkv4Ua6w7d4ohUqAr2HE5y7lsHZGPjoLSELeBCnaSpbklL7supZ6kFsPteAIP7+8rnSh++0uueoWR0dQVXANTvRYFMlX1fb4zdnXPz7TXpfhWeNZSOohg432mCz/Z4neXV+cHFv0iTpKMnLIgDlRWHpPV5kcrTOXxn7ZtlpSVQ+kfL08wFrOrxNXXblXQnlaZsfWCK0eSz5tQseMTIY6LnzjHEHbQMSRtoSA00Bw32N0BBmpyzyYMwwC+wDiRXCNbA75GDmKZhDgcGRkcvO5zBI2fg8TvC7qpKqvIEyvgciO10BjjDnxy3vlqp1BryajQ+js7wJCdbfJAjlu87fLBpgM/7lA6lUrdPywaRxFlP0hTPPJ8+u3jPDvVSyDAT/c2NAWuuyXh4A1wlXnMvgG1NIb3u9V0Yc8HBDSNPQDJAAASb+zH6t7X7oBk64R8hrjWDtYhuzVD1daTVKn0HjmwR02GTU3ecaFrzhChgHmLdeXP2AhOGshi3hey/GWrCSa/91vxpEZx/+Gdtejyj0Cpd9YM5lJay9YY0LnmJTlyf1nUUZ5rjUJhOoOzpke4rrTya+2eVQTKoEPHrx3zSWCes2GtqkhRQT2Swqb4Ht4aadgmAy4m9pj4wy7IxKe9GkZSrvirCTelg+EMbkiJIH1zUlPjK4HCq780Oop1AoEIBX64+KN0LJilToxDYI/cirJe++ntFyzia0n+lqz3fuFPaYD/IZZn1wGhiuEtnJ4NNO27BO3Bsh64Wq9Lc0Wy1+qOq5VXmr9yM7UC1mq/RVJ13MTWEZhhdBL4IKvlZcoI9laMkTUdNakjsm0+VaPqA9YTvxWOLUG0xAcZ2NBnz9iLaMSsLeFd1kqV7lhzgShYmePZk9cko8amrLoYtetitOhi2jhauS1TZrFuYQghkPwqSEYnHYRaKOVvThnSujGmyQJc82s6SSqGU+0RNOa7kd1FWbTrLw5+OX5k4pqZB9HxYYTOm7Cs94OYlSTcQ0aWGWH+nrIz7tJrEYXcBJLmITZGwQnih+JkcEyHRD88qrucLEzIu8Df6Yvi6Rcqk+gd5HQvR8gLd7j+xWjZPtXxXY1/7fnEiB1VRzsrMsNyZemCqp1Xyp6b2f5KNkXT6AwM7JJ8hFxmu6I79i42bgCRKp+Npsyaff+oAMQdSUTKe4LQAsTatK31T0V2RNHqELfcHXowEauiH8CZKGTTkNU+PDvFKc4iFygbzbPrrYjF9DGDIUHdnpB3Zoq2v0oAhceDDDiSOftOeKwhkdhjTuWNF+jnVcVa3iJ+HjANchX8OfnzWECV7opiXxRg9Ek7bv3SyY+fwRjE/nbz9D9odjWu4GUh5Dfcj7Biqb9j8gB+KEjeT5XK74FJTTEm8dov847O7F1m5lHCYQ816/oG9OKIKz/ZN0CRjeDmNFQUx3JRZ8PxoSK3A/UgICtTYmCTswaYsiR5IGfGJ0oqtiZqivXV/ms152UPna/47QqdzP5162eBL+9iiduCS7kpc5lbCGBKh3It0ySWJ4c3A+KR9EoKNCysXZnrvzdicsg+LTnk2gV98+EhdGb+Xn32C/PsiyJNi3na9O61RnQyuuBC5EWo6LgKL0YgCdsL4WKoANNgl22EBfpFGXp/fTt84rG1T+wBwHPebV1IGQZEX1fJJt3tdpLYmwu31QLzYsp3/P4Lltlm8lzvbQ52KAW2cxuat5GDjVq+S68BMEbZdh+8iBnxqzAq8rwmJgcLMsOvagnFjB4Ur3NspljZpeRynSMAX3bRTZYGkvFwvr79VvCA3jwxX2T9JZ31wtmX2v1X6PepZjoQ84DgogzG2hIB2BPW2pimZ13zUA10s+VeLUMn9uYSLNVy2C3t9W6WIEVulHEzjIFkGUD62FV3XPpTYYSNCm7+UNjht/GcDRvefl14SDmv8Qiw8EQaBWg54vlO+SKGBKzxREKyWbQ1kXhn2fUKQGexMpfgBv7UXtBd3972J1bKorVL06zkQsinQq0lTI+oL1geAWT/cHqCEAGtW/XhhmA37qzlmdD0PxfjoQy5ZpatXoHJScABHDcjcpmPD9/gagD9RKeJ1ehVutujUbwgezKYjEL5sGyOXvmovq8xnLP5MGtj490QpAOIMHGE9twqr7Km6sL5bSCIiXPpf/6hMeea0EgfAdEBHOqNh7Q1e9azxVuakUHymo59hQHwZj+56Vzg7OV7DQsyzekSEjvA8uKrwSey54JL+Ig9HErRSN/84+d5Pz4gU6Vsw1wBBtwW4QhJHsS5nGWPyfDjCOrebPUoVVgG5Z281UR6U3xVx1SD2kri/6N+2CdkD2byIT0wkXhhd/5Pg2oUSUchhcXV3YqZzM+XdrSw2jsdgQXAbA0tGIE3s2tV3uKRbBBfDURca6fbCkWnYih6IJvXufowpo9fDsdmfPHI3aJg0WEKgikcXvNAg97zMNZGNHsmULwFaP27QTsnhv+N1aY3LvWDmsxUwr857SfL5PZP1t0r9PtCTnfY0F+hnxTgYj4KDcaV1iJ2DADGhU3G5pIbnu7QdrOMGzgD4BLiv1dEpFCJTFIpuAMlB88s8BL8vBX7gcmA8YntcpDonSp7/FaVrmXLvp6zfodhfAA9vC+ujoFGMwhPinGNRjGQwRmirn14htQbtZ5Xrz5EXp3yWCx5PS+ON5ok1NhVoQySa8vchbgiGhlsJeIVvQjj7gNinzOTixRXZVLYhFGQgwxJ8KYbm5zymJ98qgwRKT6UxdNf0o71hTJSwok4WW0BwbrNSXDbbVj/iXMzgNOb7FsDzOSO3LfoI/mOQo/6futcynoh3WP1oJaNqrxVgh0ZjemUxmIABSuM9QMg18vOuZ0Acp6E6bPbFRK8n2eitFwTLzEpByQIk1vDJP9ElnIO+bHHosBbXihDRTw4VzuaK3NxSbkLiJg1vmJj7br9Qc3ruyDGyFcq29R9cCwterKNY7DEAJPiFuhVD0lu2Yw67KPRZXsfX1Yp4CD3sf+0bXBpOwgM7qEq4DX0xYl9TIAB6MVbcCnHFQqjYAml3jjZYHQU4nyjZ0i4WqoSyAvq9Jwc7XnpE0XwrTiO3qu8Yr17UBD/RYIjajmsxCouDgBFX0V4mbpAmU9HenN5OrK7KIewYUMkr7jtJYSoC6JMmE2QKclcQGfZing9u+Ia9Y11IaS1KEvsw8RLlm6dIRaQvmYzcZM+jp3rJbn8TfLBQ+oK89NwQzDw4kR7rv1wANlxTQL2jH3ERjzAFl6kceztN+CflQVap+G/3SYO4Ylbr/u2xSJrQIWL2BkcYXtx3VA+oWYUSi36HjFKD8gcLjtsfyyyDT8EHrrz30RjSb4jokYhEWKnDnclKYQj2Wxv2Jd2nf2CM34BOhanjdz6DbO3iKd7IgbUQYepvqnMWXrA1soSP+xOwT06fmjMqvNwQW2FZf1kLq1i1lE4s8mvkesF3fUMBPUNKwJzNaziSQs26nEkZC2PNVo/mPPgtgG2MsMvVq5PHBk0Ejh/f044A6GpUjAaTCozrAfUEpSP7VYM0zKDuL5u0lbSe9S+CvJ2tTyxV11WO5KKk2xhDXOng0w64ePBpmVueXWA77jDvQWPVQyvthrZb0kjEVPp53aN4tTF6xJe5bnUTY7FCHqtC2Gy/nnUur+d+3YuiEFzZOVG7wJt34Ph71pPGeeeo9X+hIXlVKh0qZGrHnlels7i/TDa+LSK0JHdLud6oREVMgoXj8mAcuEaWjK8ou/k+ajfgwZ9toBhviV1ML7+3UG4ZZXERAztw68SkEuNKQzJnOQWheL7fNMF7powY3QwUvqhhNF5861LDrZj+4F1rc1P5yPuRWvVvCZgdJpchXa/L6Mxdg/G1JvPPW4eLQrO2ioTP1MZj5lwQzGcinf7o3vGBXUGHgJyW3izxfF9n0LDJLmTzOSySn/jUYzXucWzWNF03r/vsf/mDQ/gLXtgAMeLsaYDC84AU4YHFIj1dpJ1F50J4JyVTbhewpqiaVMlgGkbilj/R1jT5sYVcyUY/2NCbZGLEZbr+aePw9eF7WweTTqsjBTrKLPRxZ7KEU+TrWZqFaSdhb6Dfvj+FnFMj/Ukjmmt/YxesIB11BR+Qsid7m3k3HnKYZGx0m5u6GtPJ+NnfndoeBKoe8kxmIhWzMYtkQAGLQnsiP6QEQ9sbXi4wsY+MBV5JNwEGdgA7IpbxsYCFgcskjKSnwRuU85ZpFCPM2c+TodOHrxK5iKL4VWAv3Q1vIWijNJSYKs9oM4+MC5aH1QDaSDAtfXM8Wy8zKrCYq1CulLQgDius1Qb9LEMALZiv7k9nA8dO7zknAWQ6tcGdA1dqK++kpAhrWMp4Zum+AkupDbIMReS4T3F7HLO5CVHk3cU8FfZvMrAGvb8LcWg2Kc1YCeT1unz0MeJ4T+uZYcuO3AMJ5K5fR1c0Co1HIPaQ3kUaHGKuWTrS8oGy5if8Uc3s9aBWrDorvYZ2UrsM5yTJVZFFWG9bO0wwYH/Pa1jrLgw3LVqgGQfQNKmVXLE3a63pmW0yveT2naYV8Y1+TiUReb16Z8LacZ7sUknAX26rc4SpYFdsa3cHakyf8SH9zDJYQEzDh/XPZ/M4t2hmIprfryC82Pfe/Psqlfr2NWHvlmPh1ADa5EZ8pZYUo0yzLxKKlByfP7nBT4v/uQdZqSEU0wb1pIqbllsVKrVMpv/cSDgVFwBPQXfd7GUyOD3yGCSdfdBarDv1dKyS+I6QMnOfyG1xK757lSEAdy9SqHdt3Z9rc/nfnKtE4nysKvT4zdD177epMNtRYlMPtOtLjEt0ZLmqdSh3iQFGQe3gxEDA6R8sARsikZ32L1a1GrYYL6czhVG50sMteh3wZ6p+aERP1Uxv2w6vxLbqQghQuP+vEOzEG5xT33Qg0FRZIKee8wQtYQU1+ZU3RYjhdOtDTNJNnO5oX/MgW4KtGO2RCKAzPTmZEnZb+ZMZUibYDGwDzdCK+COyH247A7gEKcnp+f17JJ/BcIxPzVTSPejHK2kDByFoFbmVyVGzTBYnYrmHRT6Qx6lHxPYvLH0V/N9qvf10o4SWMy/m1EZESh0Xklxl5voER+k5xGKIN1NsM+k5JQvK52+f8dn9oxKawENDfhPqeuhn4s7flqepHbc0gX3SmOPrbIAAGreX6vjdggm5ow5Mqwutr3asZCJ2k77v0JmzvtA8m2CEffsxPGLI3mwHpcjHffcbDbEBlRGi/MWxO2NFbjxq6yYoHHFsYWL/8rZLl/A6eU1q6mmuN+Xpv4mUKig2QrXpU7yWnqlU55Y3ExL+MAaW5MvVup+xiJbM+gvyc07zqcpipRIKCnl6ckBPRinjfuWJJaTAW427+kIBYNoNSqoGT0jmpMSSGl17Zn9jGA475UVnCH2rSK4OnscCC2yJ8JaSwn8GP5Ejt+xnIY9obKkBk7mSUVdKZcooXNSRg3Qn5Pq2eXdXExtBxKKMAS+PNeGgTsLDKRZe3WNgqDOOuDJCETfL/hDL5dKVdt6cl3vDoDJusXa47zCWALpX+0mZXXIxh8SeisnzrojmM2FyLuJlts75CVWNPXZJyMcOPP2eisZJxhOZ5FF49wYZebNUnNAXlaGeHVa53QM/NnovgCy2nQQBybmfRllcVcACT3Ihkkk1p5WA5tMw9EbxaeWBcFGuANc8kLF4sey0+JXDPkvNlrQzVL2JpwuispiGju2e5Fg/sz8XlDLcdLWUP/eXofmsmzEyjys992EKymjRhUMPfflA7WxUy5RVKTngGV9NMwGdJO36tKucuU2iMebKWAsLbgVlH9yq5uq25Qbb1hfCWaogIX0aJVhsbvZHfVjD0uITCFvqAG+vKiwLnOXiRalZWcGPiKldrWOKbMBm/03rp726VM4QDcjTTjgxjYCvMBXuTFA0OG9EhNJIzyQp5Tmg5UJjc/SZ7jNsY3pSysenMS0Ed1eeCHYRJv+IuTrmVYjnexaof/Jrhgj9vZUzKlD/SrQ7fJ99KukkgD5kA5Mrea7C+XXllwj5EsKHC8XotXtlADldAm0yrUPUaQyI4fNv8VIHCMXMcYCkt1eqTvJk+BkxHrnqeEnlWAghulZBoxltIYS+05NvClAnvFfLSBmvJFa6CL009/JvgNtxDkNXwKRFj9ibI0mt193b4GuFLaRTYBuq/aC13YBn+OpMmCcGWkISRtrchAF0KG6UyA6hyDAUu4hpvNS7j8WN/LKZblaBh2lFARaNE5o2hTQAjM00dGJayQe3JU4CW9aasIvHcE5L+4tCGNyBDPUjwLlDxdl8n01cBaPsq7yhfeeMaFzgof5qMe/YcZ515ukmYGUBcWXemo7Flh/rFuM4/j1rw9hMnnFpSOT5ln5HFixd0h9w3SIswaPDWxwHvV3QLVMGQO+Bz9vpGiVt3BR3Vi/L1oTHbKwFwRjmbuhmFFA8UFNCf0+CH7d3MgqLPfcwrtZy2993EAfctxwh0BjdpQwRZ4Vb23PmVCOJIbtQtutCyEW9aW7DgToNRS5JjEPCEvLS08IbVej/l2aON/MiBUkdCbLDEVHrT9eMoMpkrZnuZK026mFY42wyRnUVTTAjgMtqm88YPdEdktx89OyHBzAw5V+d059aFONTldcu8H2aVZMufWY6suEcRlpwAdElh/wGjulL1t2MItTRXF5UXLVIzq4f0dRKPcYwXOGDWRFjSAH0NrT0wvk6Dm2/s5INujFWxLRLbRFHtcHtoD28JSoiiY6MyZjBee07dTCJKsHJQ0d9LuRi4kdlNU4hmySJJXHqj8BAthdjz0PIOE8AOef6GsI1hq7J6MMiJmSv+3GAahP/fYF+/BvVu+R7jV3mlWYzfh9fFEgHj/b+yx1i4BVSqb0gHD9Xeh1LF0WttBvCH5mXdRsXpxwxM9Q1a0qvC2SCTxtnhIodMXbr2zKNR179maQJmOqUoiNf2PaEzzf0kS4g6lOom46I+YNeE+ROeOvBF9850XOOF5LjMQ9LJHy9PFSw29onXcWR/3b1R8BSG8zc18Oisfv/q32lQmMlHsEWPdyVAJ7ObC39JYGkTalOUmd4DKif0ExkvccPjXHBBKbN7UfZmX2re7Tx3PCAUM89n4cBUqBFkOuoOGtdvwPXw++MYb+fcT0af4I9hdRDpAC5STdX9WP7+OLHTI37XzsyUX8KY2VzvtHDWHdaWgSYCx1CeM+E9TheR0L3WfAFlWm/x17jzO3c9U6fH/PFEFMu75JNvpdNlHJXPr21PkVqmPb12WFCnBAtoT4o/y7IwTAKYpUSW+4TXf3ex8HLzhlftDwX+lrKn550ewD1VqkU8oCE+vsXaK0JzH7wTrg1BGHs4f/S8fmwjJ1FK65lBTCgbhoEYoxfvG4yHB40IOEW7rEbKSsvXVrIdjL7ouOPYMnG9OFXBqXgQrC1ylph2zayklP4UmzPuUkoQxGEj4swcyCLXQY2kobXy0QqkTFAMcBzgLbbgW+yDzMez+qCvHmOi+4seGoN/168eE3rPCBj9wusRfNGxDriBPraWOw3Tbqugtho/n/7KkXzurMgbSBTPCGCVIvX6GhtVTB7hgCxsA+UKv/uMCPvFALc245+lp5MNm4lSXB2g/GVbjF0eR5LTSn2wh+N6lRF37naRn11C9f2Sgkawpu2HqM7wMG+/auCwkuqvXKMer/gsY2sY5x/7fGhkyWuk6mZ+/6+mxid1ifgsWknLPaKdXgwWtkdsjJyJzfbyKauZxds0g7nS6yuaxD2J/ia8Kmwg8g7D4YRmJtCeC5ySXMWVaChXdPZSgc4Q7hO0IIyPYCfY5w7BMIZWWrZ50qJe5DyzhipzOSDLpzM40RfbH0UgwcNafysWkRRLhyw+6yFedfFnpq7ZzDX6Zf2oaGBbN//yO92ejlHycHMukUDUyZowS0X87pqg67iQ2LNUh/TzjB8NwxupB5HeBWWTd6rLICwpocfTKoJeDZ+OnaytGjLdABDxiZ4pGuesTiAINOv+60ZFOVaGKuZ4YRn9Mn08pGTHL+2ZhBke51oTkWyKBDdDaRhe4wgcqBNC+1o0O3z6ONpGs27sK621/6ENqaDpZKMMTD5qVoB9j8LMJjYqWyFdEYfH16khTrSzYFQIZRbHOtNl+/boFy2KAonC2NdTHAiQk8L+/1NW26V768xcZc97DOSTCTSJIIM3wZjCTf7YvAQ8H62xNQvF3eLqXtMqC9SeJZ1rCC8rL8QX5USIR00ipYSqq6TYFdamxsGkrGvMHpkMo7rzZeFMxobckMW7vtvSWueQekyVqZg0XGf/BjDdrzdfi1Y1YmnbrF7iR6fSyvaFW80gygQJOXW+wNxRJQExgF0nMTRTgNm622QAzPQoFDYACvZMLCwoDEPACpI0MSCFX1/DbYBdYTnQ9kYXE4doQuXg+UFT0snRIJ9+8Iyn2f260FSH1WglYK9rDgfGwPQD2p3CRkGLUqaZ8dc0xm+9Eghg35ysDZkD29yStGBcLWkfTm8stTU2MVaDCy6eJ/X6x0LEKNEt8Fkd8PJR1OspbBJurYFuVduL7PJekcBan9mQUQ6Dr4U4qod9njiuuW9rlP4PXW+TxCv0Jhkbo0rZZGrmRzf3dJIpdd7F2p+2B9dpWXZhR7/hY/ST3E3XvVlG1dRkz96YXbJoFEL007G5CedcnvWeZmPTpBpBcqVWXUxYfFGCJrby1CBxX4Wo135SXZJTIsjQJJCZPu1cJ4sh7ZTfkhtaTpQ51q7Q2+WYudnC6s0ycl9BrN+v4caVim3ZTBSTyJ7hipQ5BQl/i9Kw5K+/z9JvsEV9rAA1jZkjJQ/kRs5o2QfZcGEEbD6Ns9/Qz0y+FudRD0SrrtuGTxUI9vBcjvQWK0o5cSf4LS+vqUgY7czc4feirF4zwEaQ6u/PN6SVt87O8VB+VsThbdwDfx92CgS+bvDHFPjUJ4McgzcD+O5JS5LItqHvV9mCQjsFIwpZXyFnCTsfeLOWaC6hO1ncGe/dtMPqQYC5Hwpzkve8K6fpIZsGUM++BS+EU+qZieD52mdEdcOfe6QuHdOkHNHgAqBBj4OVw9jD4Qm6yCOqfLj1IkC56RYQyS4PR9+MMi5VCUBwyYyvNm9JBXgJd+LmWpUAG4igwlycEr5LkBQxTFiXEqPGqj6KCh5dEnedhL9HA8aqMNY/qoglywZ0Wgs7dQ3F4OqaYctW/Oynlgl1fxdNU4/XM2nH+lJPc5g/p8UtQDr/p09di2Xw06fp9E9tdisN35ZXrLFMOAyntF88cyWM4wmmFmzEXlGcFZ/TZK0HwqRfANV5lx45C+sUEnVru9i6HR0xLtdVrLViq8KCWHMbE+p0o4baXGaRM1edlXxTnvz+uulr0fc1Q7oSsJFi6kvsylD2DQ8F8OCKF4GFmoFMnS7zvnW3Saz8IaiPIL0dXZBZFQROe9Hc8TbivcWuR8ACsd4qE25bsExJ2IHTXcKXh3Fk0mxePAm/AFKaMs3dI2gEj15DMSCmNbsjwx1ZRWz4XMyGna7NhL2PvPz/8l5F2xl2jJCVsBxYgukYGPbawayUG8c8kufxFL2L/KKJfKwNQhh4jX5yDFbiGZgEqvkoSwP0Ck0Hank3SRy/X65KrS6jeSFjmj8VEmPziZknc9zLyw+A1eitLOk/VhDdb+JB29XkGa1Z6JEpTZ+CTS9f4OKJkhv+droCP4XQw6CEWvHneiIBUm6k5XQvcsvIEKdAcpQr16EP2MAg/+OaQWeo46tDSFHa3OqYa8Z3X1sIVRDSnG3a6ZumUG4NfhiuAcDSubHLVARv2jxMDOOqJ3vzb4c1U96oM7smhV50jiH+RZyY6lIH5GAhBkhRRe0QLRzvuCBODptyUaNsof/jdbQ6Pw1EJ1rBPsuVQoDma+P1f3a+iGNhXPjzNSz84m6CaRN/pRhULaYYwjvk99dhPA3lxf6AgQ9DIDBONboRi0Rs70810cV4sLnBtnelh2LyHWev3a6Gt3bYDnFs4+5J25CytqDD7pbc4YJtR+aeVbWxpG24IizoC6jVjWjv6FnEjd8LMmKiK6GwhBUcfTFBO500SaE9KhFApAC81GVn8DAdi1jlr5bwaEf35LuNy0JABZ+QE5bzKyziYLp54mBh1gtpoz61W/OaTPWbOz1w0PGhFEoTjYPBaIVXk13ijEN3n5ovjf9pJW+10yZlnMgHEUvZ5sQWnsqecmrDwlnIPg/9XSav13gTR1V5+9WSoxy68/v63s2J4dvo5pQxp5GdRYiH/ckP/j81AIKcfBw/v4M4V8Ps7NixD0GZZda7nC/C5jN3Y0wheD1sAgwbp+BQjvg2UdT80OsHiKH80lOhW9OKugxkwebnKzyCTNGmQu11SGPXH8ce+iKAU5wS098L9QacsmlGgvuEq2PaRbQj3Mlc0RLZfCnWXt0oF/4peHgKhGbWwZY6RCLU+s9J1+PbYOq8hNf5LJd3QKxY/Tl+91MJkz2CNHEaHQse7V2YNAEkTWauTF2xXk+CAHj998uOEUTHAchN4iP/yeeVGyn9AYya3I0TZBPfzsx0/QXrVyofszpHOA7+cdjiAbinc1+v/r5FNFnz51dvbV1mlW1VB/eLqqW1f2+/uCOSWfoQb1IuwDKogWk4ebQGhzVlTs6mMvm+P0/5qKd11WhyQ8KF4xmgwVxbXGi7UxPxxMXpx86fJ8u4YRZ4gpFAgOi4azmSZbQemqqcCV9LSu5DydIyFJGc/WIvLtLvBTl8p8ejUPt72rEmSSxYno+WEDjs8P8s8l6ciGaHIsqgPr/99LdXOeFIJQJ5e0QsgCFXwE54O0u1A3p7qcgp8+CB2PD83GRVtR+KWccXnlI4RN6vGK918iTqbjucw64D0bhctyYSvPGruRRzyVHRcuBRw2fV0IYrv9K1KW7jkman0/eKJOx8/ARtegfsVjnYIpJ39uPQ8mpzDBjyDGGTydq5G+3ha2RDTOPsaY32QIpgH+Ri3ZyG1AxRqPITmijSEi9f/vtzIjeAh933FqXgSWnjzQLF+iO86QmdW3lfV5fq7NbNOjpLd8LCYSnNXDwLoGsOxc9u9kRYB/xZFdjPM17xPSVpSmO6pMn1Hhh66skRLeTw7+X3/MeU4rBuSCRgOTKw+wisggUu2mPAcLx8ZUmEPCdic9LyXpR4rRr80U1QRw7OxXMrREzXhTO/Oop28O6qBQ8vzAZ1IkE/9NDbtCb0NKULpT3NUMEAmwWAOcfe27JxAyqaEi7hBdxhYOeiFhMTpfZpOIDQ4kXDsuw9zWb3VWAABAbbk+LgXsGwvFhxgb4eRFn14QvqtbBMSFeS+XCPTc/ttua2V3aRHI/rlVm5vXtHBfpRrt0HqOvEjaSjoSzCDiK8OSadK+Abcpo1FTYq/qQHhvxpG5O8kIlm1EM6vDwKoTZ+yaeBw4yVbA67m8AEsOM+1NWsksxbwTmW12f9JtaR0OkanB0Tm3cTDZM9bGJZ8CpOpnoYLxn/m2SQQKd1J1OrRVqD0J8icZ6J+ilyyo4oNtErThz1rOvIe75QKCi99S/qORMZh1KYfZicw9cc40WB74qm0g0efNnxEGGBAD5iEo6oamqy0jmWHtFJENaKUOUFYMhydJwN7ZZwNFOG+hMUy+li42ZPkFZuh7HRlJxuN8iObo7orq8XeUg2oKhEnMGVf/q1+3KW49tDBr2e9nXo53L+y+yrj4KH8Sy/WP6whEqfjWQ+tKCEirC+MmMGx5RpOHAXdxt8Hpm3dW3OiwkMEvwPVucc7TZG3rI1jYJyyFyVzrncuWSsFO92lwNNNVmGmZ9d62Bgf652gv9znYnneLT/uBuv9XhqwMPiKGaZlUE7P+fYY0qO43WVNBdgVV74nxJivSCzUIzZGrlzFEWRnVzf3ey+ROyU+jcaGF6RHnrp5ZdOJ74ViqbGDe3WVLMmmJu4a29FsOQluEsdZbvpu3HR47ffIrHxwwxw1zKKhU2XAgYIX4Q/jHSpfUSqERnm0959iJKs6hFQGRaYu2Y=
`pragma protect end_data_block
`pragma protect digest_block
debb1dd2822a5706f11574fe52d962a2e62066f2562d1d76f6ff771bed28e13b
`pragma protect end_digest_block
`pragma protect end_protected
