`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
4gDj0bOzm8y+pve0Xdpmz8hOdZkoWLD0s8Wi1hQPsdaXA/2hh+NNDOKWDBG19riQGcuY8T2Rr5IPCKdnWE+zlCLdD5bNgnavjlil1P+0JVZFcgUmvA67Pvmo7R3LhcA+cVMCzjXd4ih+zo7zGQ6XIFEF1BrMXmtlNs1wUHrX3HKYQjnwaa3jNsL8HUNb51mj6rJBqTZFeQDBwT+MDIxY2EYdV7Gd8pbmsB5AFzBHUtkOCbDkg17oBooa/v/KsaqhYbm79xvob3xiaMn345oJ1J8y16FDJmtYI1JUi1awgvYOxEH23Fo0EIxOUdLWaf6l4I3oD18F/OW3a1Ty1M55hgsNf90aNhzFqmVv4lSMTJAWDqClQjJAOItNvDqZxoyB8HELUzLkmOdB5DQm58yEZetAzl18w64vNRQ9D1P2noqBbrM7bWaJsez25ZlaiGetggijBQ5yg41fKB0my7P2davKhRJ0Aid0Z04BEGAMFltYH1JJ+IZ5daWZ6jOvVPvjk+9eSW0otR6+YFCvKpuXLjgZMibt6iUYuDMDyPbqhv+u9h9R2uBebOoe7d96Y8YzW/FkW57bal4BxyCrQNCq60Ra7csFrQ40xLezxmnC2EuYorHWidUGl3un2B+XSxcaaaVGOPInqmno5JWrNIR+3JeHWxcSOvz6p3DdYUEzTjrbkYUg8D8vIcBvMjrwsMWvfDHo6NEGYVxU+/mBFxpARApsjhFpgiPPUDPBYmLcmkAlVOWuPNNoeJgE5elYLIwxHGTGngg6n4ppBgXf++fJwkG2fDvJ2B1JT71BtYVnkbXJ1kI7mxD3JTr8TQM84ilNKr7XjWpn+JG3OfTm/ArHzhjhooy0UNlMZpdUF2Iwyn9vmyLBS/uz1qo5r2NctCMSsJE4rRkOSwNfQjINGL1qkKQkNzUtk2cBWpp/9dKSX/iRGeSoRxwYzR1I80XS3IlKBYOYILVWpnDZX+p4gC1e5EUco8/QBWVFe8xgAbGFhEVUF9gIZS78Op66pK4eygKElzR0aRSu9r9i4S4+sWGAOCHGeiqyI9w/vTN4+z+2xD6NWarZRtetFpm3xWxti1m5y6mflx2x0/xxV+8c0FqikjCNwVsGxumM2fXWMzC0jHRCLplm9BKNsySBSr7rCawOFC+w5czcQJXGT5DYRT0w5wKmdp+M/LdKt0F1okNEC3bf4YBV13WueYyl6dYlXPHlKD5ReIIUlfh+fj6ATOgmTRwhQzRh0tEFWJPACf98DVDxVn4c7iyDCY3aEjoZD9IlSTHfo7SMa5Xe3YPxuAdaxMCpl7ZcY0d++EVdzKNbzwynLx4k/ZwxWZ9RgqHNXXw0OPMBu4FCpZLBYx/28ZDPkIwd6Xc4ZsW6j9TcNahrgxeppVM5Y+G+xO1B5+O7MXKrny2Agi/85vgnKCtrr9IyM0q1Vl1YLY5NSfZ1PuXCsMdLrYGitobUvDQISyJdVYT4ql8sUwNX2chkD7SsNPDLdY8YBAneIe/KA+Qq92qUO6+dolkd/6vQlhL9gzxVWP4igmHoHDfcnPOCGUn3iH/2kMvtG8NTW80KHKfOqyQZtA8aejT+4vUJsf/80dWmj/0FAdHtRuglSVGRdbHEC3ZBMeJDsfRO/cTMmffpqQS6k1JMZVsWjUs3h6rzo4sCGC7ffvpKH57I/9vUJFfjUjdEStifkejU7IyPS90E5YayfEvbIxsn1ayE2FSXmQYmwPrvEgIJBrRT9sFLUvWVZSJiq2JvubGSjGDBh/RLFSUOAYtsTGwEIKKxTJj0mfoKyM4LGYqh+Rp9Jk7dkevJmkTN5A==
`pragma protect end_data_block
`pragma protect digest_block
cf3f5494da8cbe6125c0cfd7e9ca0a70f9bb3dcd97329954dbc4f65745d1d8e3
`pragma protect end_digest_block
`pragma protect end_protected
