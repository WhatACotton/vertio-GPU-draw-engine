`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
TrIjNjG8Iil5GZriXPEfssWMRcdgIRm7XfHIKqqwJ0y1Svroz4ysj0lIdELe+f50yYQF4G93udgT73hXVgBShPXdO5E3n1KGg/pRO7GkijJf3ykI290ES+O1qFPH7OedefWqAKE7FAbUZ8PbakM0R+NUrSkb9HIOMYgVwMOO4ejzY5WX4g3+CNjOT27pvOtzdUsoDur2hZWfeOqdQN11wss8kz+3ipn0TLpEXMKMLjlMA4DXDjj0rGEFO8NgRubMNNbQ8jXA6HrUAXIPJmm7tGNxTUyfPGPNbISQsmzWqZFZzigBicbLA70uvNmQ0TXxsFO8+DFOmXDKgEgwrGqbFOdg567zKq68irhVDxLDd5sUB04wEiUD7iDan7Kg6Q7o3uF6eCmtQ+ZKt2AZPbaCwQhB4jyWcAdYUiLEFooDaThjY5/sIXi9swVV75v/d3CUb9IN6ApGyzukCdEfM7JT8t0r4POYmqiSHrkTkTRWHKBWGFqu++A7+FvgcpgbFu3zu6/5D2wY95onY/PhXNvs1XmPy0TfGoQuwwssqMSCHiNs9ZsVS6GrfBOIuSYGW9ysOfPZZTKTvD6yutlJpi6lHTHDJiuI8E1C/ASwZ+0jQdjrrDQV1PMhULCArKG2i3VuxONIexHMeOsAKrH82E6O8pnQe/5ORUoMdvhibin5tAyA8yOEZb3hu9f9pySHsvAUoXt6FNtuKOpjRBUkBGE2ou2XneFSGHOvM1IkrEEbMorY9xOAa2R7vjaXYExVplNXprSFS2CrSq68GnCtPsgEUsG/jSQJwdGGdzuari36JsjHFG56zMZ4chaFghuXDcEsNu3Q+Z9F+4lYaP6j7pgI+xf5RkRg0J/3YfsqUGywnQKDpMwX0kHKAwxVoIDD+8G8PhI6++jaUyLA7peX6c3VKhsgkTjwexTRp9ZhK4xzMYaIeAhpd2mPCU7fXHkRwsYlFsccVVoo3oCYYA+o1bDnMQyhLsCKaEmRQPWfILKmTR3T9EWi4Bah0tpdAVFRWdLa4gd9R7WITah9Rqazf1330bC5tLqDJfjl2jorVoDaD26o+XRU+6gKCcs9tKkuEwkgJO2mUUVPDINmi7eBIhMhwFi3PsGNrxl1gVmfmmRs/aY94jXhqndLD/VSOkOXtb7iCC3SdqvrY/wuhn0y1q5JtnwMbRVzVstoYFmTA0SeZXv4VNLGnIeduKTAqqLWyAU/u1aboh2yS/7M3Hnvs5S8igNP44sQ1l/dw/dSkHco48eQezqi9JI/YoCGME5+W1tz1XXZOsW2Y5jfx1Tx+ow8jd8UXhWkmdOOQawE+MLpzAr/qxXor75DOiyQEehB+WM6MvpC/jiCLt6j+XKpivHYVAOl6YPY4eYQcxzZiUVSLq2boKUbjwBXzaSdBsq2NJzEEaTkb+joe1CHXDIxYgx6265dpYsN0KuyYd3HrPChVU6Pe1v7ngGVIKDpJH6ctTIyw4vhXQPG7nTZAE+9G90Xf2OTd16K7wI55jz3jL9iw8127zpqiOABlClTIZH5w6RAvLVZA5uNhFHNgfP1oj+KZeBoQVdlrqQTT1jc718KWVz4lhM23IyeXAI6NRIwy4pdM9MG2atK6AgbAhQyBakc55fWUYb+Gqlelsn1jmsrG5xZkMmGUbRcYbzLC8FfkWTaHpWYDZ5zb1HcWjaAFISJb1YNQZHyVoUD57m/wyOfjMQOzEKM2vWVLJ1m0Jp5m4RtngDcWStFuJeh4ufQoS5/f9m1zHy7FFE6J+spjpxDGZ749o4kNkwfrJeEydi5jr5H1wXbED/huInsOjZOtpY5E2cit33lBOSeKl3IDR4zxORzOvALmsWnLFl7sUrcYTxB3/QtfYXAdikOfPXDPZtBixif4xPiutu7sswfhgjhvWoX/ZPYG1EBsuQd2RTlePwc+i4gt5R42Mj2waGtlZ7mjWRZznQfvkxhmCKAjs/Bc5gG7C/Mx3gLkT8riOWBChpzB0KzSRb/uv+M/HIdzq7F2Wi2M7CEBqlZLU0VMDhaw3DNrMBKtP6m0jwfsJTO8IVbTNwJpppcl+St3eCw/GVS9nqsGcfGA28pzM7its+MK7X4C9aK6g1oUWwWaaHmF4WlHMDrGOwkVtVe/qyj2emyjAh3FNRgdZQCrpDhRKJBId0/+egpgl05FSwUk1GAPUVvzbN5e1p66t/lQ2Kip3WR46s1oWCD8H7pIWLUe1OnNhhVfU8iTq0txy1ATwgaXRd9wsn1kHDGmtnP+CNu9mYn5st+9AUC1YHDBcoJu2QUKQ5s3fiaEm9NgCeVuOLB0zI983eiPr2wbHYkJiyao/yvJkUZ3QAIEE5h9+Qbq11jWSQzGMYF0G7ly3c/4WP9GwXKMx2iQVYqWqU0/k8qoLZfgBkTkJeLPATKvswZff6iUohrx3G198iuSQVW2O2BBsxqAa6oCSl7zzJ+A3WHmi07Peuz+xTLupJYsXQXZgrZtO7h+mI3rUP+BRpVIn/MIBB3edvCQjQIaj0UoLNDCyU8kkA+Gxc18YroXf/cruo6kH9+wfUBzWl+dxVx30fA+36ukbHZ+61sBH7VNkECAC/bcqzsFYygyoyTTzLWErCV5Kq7PpP8UuXE6eYCDIKgz7PHcbW+8kyFWDD0OCQQahejyLyLVgSuwVYzyMP3eve5i5ymMzCEas6TRUCv353d+p6w4jgQSXPmn/41t+Vx8V0e/Yiyppy+eE6Mpt8tMJspCDgxh4PN89iOfF/EDxd2OlwiRtFNZ6rZh20yx9khmPM4rsA/JM9gxKzOt7jUaF+T4PJg0SVmDenZMGVUkeePv+ntq9CEOHHJZkuwDrbUBqF9VwjTaN+71WkHLHTAV1MHsAS98nhTgn9KJpBfM88+NVcR/TL210Mhpn8SsQ4Rn6XlDF5qc7Urasiq/wnJosNm6210Cl1QiVcTWAnec8V4jV6c7LxdcGEVJSr2RszDZwSv/VKQyrGqxVQqP3XIo5i+AkU8Dywlxh5DsWP1M1XNzGsgb7qkBUMyLm8xWBfv5JoPKhMWS32lQkteD10rAzphLttzbYdcGk1DQVkf1No2qlpzAC8EmRe6vO3dHVgvkgPRk/sagrex/CcTVBGkgY54GX11sjK3z8hH5UT1JyMndznNtMSN6qPglsKUlWCRWMMyBefsiM/pElJonzIg7juaiueogmEY8h7aDaLp+PyQxUBhgKJxIu/xBwfTpKrXAuxrde7rczQg6yUbpYGO77SG+jLGR/5ZRMTJQjo75woqu/smXne9loNg2gkTp6LqY3OIBEQjDRQNZ4GqQrMuZmJXOCfFJb6TycmItmplidbEJxF647p2ZWyksIlvcXLWzZe5ABytcJzE5W6hP3hgFaOe6syeU778dqpp5rRa2tGX64Oi4rnNJIMJanHwFcp5SXOoJSYeIeL5FOkvbZq4RPvyrbZJHSwsDggnGVkCgr4X4+b7s2wMTcKpc1mA96tw/EUfjQL+fVhIxu+ZFxFMofGrXgyYY1yepRyC1almcesZ10yWj7U4rwDZAp52BnPSprA3n7mI5P8RPboZHMvVo5ZfePcEPMjy3SwRkO0lDwvPfIdki1LPXavV16vaAbiSRCj67gePZOq23+SNghE5HhV9MxtQpax5LXkkiVSPisR7PEAuaPPAAZlQ4/BKgvrvHOnliw4rMTDEOXwpTUH+i6niDtTP8UIkMrXElnPUgLANqhYyDpFVamWMXXi6nA/evkTTpc1Kjv/GndHSLHtDgjfcwsK7D4F7mb+qM4HYj72I4MngyVsVRJKuMVpyf1ux6rKoUcyu3xkayj0wiTTIm/UGIvJqtUlWTsiHkXWHGFDkhpk/Ba9jdhrcGSmawERhzo9YSopqhOB17axudds/BGglT1VCyA8yxSbIXf4L7n1tU508k08kFgtHOMTYdSBWsQaTp59A6yEKQ55G/R9+4ZKJWeMuSuHP9IcYffUXW7e/oUaFYlvnvmAuR4F4xGAULXwbvlBJijQilILYDPrgs4SjLjcpMk6X2HS0M8JNAIvRu10KSj6SIwE6g+PFAZd9OBwQQ+x43GMU8iMH3MVlkgLWBSfMUJHXQ/mXrQBk+4vSYI1id07fc+ITHfZvT/R7dP3ex8TlAlZGuzCfALkgKGQvr+1/6xl4MW4/jC1D8l4TqNfuc5H5F+bzIqSYARdFjioTS3V4RFmfhql4C3pwKmvhA5RTLWxv6v1WFiYzRDdgazt/NKlCrUXiPQrrotXZhgFR05AJXBIsFy101+NOUMfreNyfNzCUwaMVGurSXER3Kj+xR7wpk7ZWa2eXmbdx59X/dEFVTLtbLXwAR9hCK2rp7ly+51A51q+1TAGBMBvd4T5s/JsqIz1WpVky6tMWqv/QmMgZ/c5ObN8sVBXRqJTRqnLElzbUiMsu5YdmxMOhnr+828/I6HHFSx2rnrIIWBhyFPvD/mGDb50jNsRU3DI8rMowAXS8sfxNPbnoHNf9mzFRRnxdGQ7GkAWS1pY3dxFBNXJVlicxecuPFZ9J0f9qYnum2OtnFExa25RzCbYt2OWNC2nLe25ztXJ1goMQwFmb0hD0bYX/txVA2CykjFRNms5gHEbncIswJNvoSikGjUNrhvLcrmUV0aPgTUiskAwY9gxYGToVpgrkgDkqmqahrjf9/OB1P4KClUGNDg9Qw6xS1FPOnGOXDRO6Ct4tsbZ3RRL1zyVq7Z6ExrnbzcfRr8mR4R+7QiJXZ9FTxqE59ETq0PAScyB8eJjiG1E28VhOOdmRXkCDMB8Ve/qv81tyQtehMflZ5WmeKQcktapTGiztOs6eAx4fy3yj2tLjqdVSOYe0uLXi083G69YJCWCbFi84ee2FIiDr5oKCnBUnqn4D4PfyxeUzF6yqhiSkp4g+kRUXYdMoEKe1d42inTls0FpCQtAgEL0UIUZRGTftP5wLbd+GuMHI5319PFkyW+KMjjbvBXOa5fxWB4T1FbW8aH9gLT3UgOGf666CmT53hKnCAJTQigVG4ktTAukBc8KPsmsLLN5QM7EDDzsGpM2WavLnggVS72UOc3+K/7LDHWfBWoeAAugHrdwsm0cdYWn2JDOy4WsCCE3zf97z7xg356r0fQ3ydlCAszITBy4GctwB/l+X7aMLjhdbMqH7w5LS9aTC8/wM2QREQVRpn7WRAinR9TcTZnKDEfKxfkQaYUvKW0IbeyaZxfF9yX0vwpqF1P4ydh1/pfZbLG2q3Pstj7bGIvB9VzEMgGc1LkmygJgXhRpApkmdPrOzoIfTzACPMsxRC1KV2pGx9ZJc2D+0Woo3aX8cOAOOPo9P8cQlEEaHwtF8QYQ+SODRwiF0sBsma1IDd5Bh1hCNmQUB2utpLJkaAxs3s2GBtRBl5yxrpgytVCgUj1bpzlmcuVNWJB37uWclfKst+CMZsHchajM1DTxktnIh1kSqeQFOFnoxRhrUITUX4FyeNrhTws9AzndJ+FZRot4KFTBeH3+Gtkz7gSekgKB0+xtG7g4wnqoa7vf642c8MupnhJIFcPCzxQDdY46L3TGnvno2ndnPKP6vENRBbXKiSg/npgK5NvYNRPPfo0mfpU56PZGZseWFKtsQHRGJ3OdX7RJAwXMlIqfjwnYn7KH/ijNmPp7fW46WtZZGNnLoX5+Ngjj5jPdpqi4FqgjvmAIQ2zlk+eZX8hnCuCfRS0Hn0UJeQ4wZD9arFCoOFJBF6sY8iirnYKTfpqwBJ4yfsVoUurITIbNP8oDcQ/bsFvBihGleXjX238DvbHKCegpvWbhEtgjzw/XoIurRZlTepiEL8AEBc+O2FlO5S+jsKNP0X3QTszCLq6AG5x2cRClHsTRN7gBM3Q9HQ8tIi2V/crZQOdruAxPuFiXNycYDfbRDP2kszX3fcrOu0uzwLZpRC03aso6zSR63dMqCFBOYRgS5+9B3BVIXkAxc5XegcMLXkZiLMtfhh/N0trCU+dy7Zk0HSyK4+9enbFJ7ly6aa/P1LL3SNDoaibXC5BbQDMrW2laC1t1QoJvNg94wx9shq1sBncQYlZTbBkSXaM809tnnuoEY6C7rgi6dPbJ090duc67X8rj7oQ2IMHNvMb/yO7vjPLcS3qKnbzLa7zgzNom43RGfDmv6O6UaFtTWbNSj/JQRvvaAtVNlBcr30Sprxy7vDtW0CwEUC7b9Q7fTszRBK2MRSlrdZJYLskmvq55jbn6QFDQjyaA1LRpuL2jbKVEW42qhK+QoqnA/c33GvHs8bvdLTUeCEux+AKQWCaDUZcuaFvtjrZ1Rcm09s2OSEysaS0mhICkU1ZLUd9C0Xopv679ur7Vn90roVwUh1BCkeWE/++XulNP+Z4ejRMDczSfC6Og3TPe9+23gRSSZh+N0i3oLafDULhzW5pjqzX9JVakCyYSW8mMQOoz2VPK+a1OWj+ETkOfWXBNkxqDBHmnBTHv6hF0ZvlAvFf7iybd/F2HUfgAPmSInCD5iJHVx8oRy5c7FuQcnUq8/1LzBy7A/EtCBHaQFwbgzCY4a6eXQzq3WvXuR7xituIOWRLd8TiSCRH/OUKI6BmbXndkOAyI+QJ0tLisTm4vIYAVC+G9DP711SzhcU/lKt6DowrePvSqYeBc9S5aS1iPzZGZ3/gMWvEvB7BvZmPKErCybSrZGqOjZiR4tPvGFeoi8eetAMR7Cpp6MO57z5Ae0R8Woo/bofdNUsrtZ3cfowjVcbksAgQ6P0sOrzgbxboiIvkfYMjr+FFMsal85cddiED3rfZChK7nSU/7yddmhfep9yNW69vSO8lBj+mjSvdm26L1h7jupl38g39AQiCi/uvc8VjSvHigySynqYnH9HA6NEdiObxvCMkv2l7Hxdk3VDMJPkM3wF8zod2DENKsgh6I0h6GJSJ+/xfCG2JfHIdiA8eolKqpAg139jIXyUopihSrvEzf/RpPiybNa9xPTFjilT90gHf692gD7eGqzgIpjM37xiwtNko6N45Q5tzNI+6XclqZLdP+d/wNFXGD81HPAdu/nS2kpRiI4JKF/mRaQv9RThSL3PoBq2wD/GdTwfil+0nA86P/oRImFkBHiegOHVGol4zKcQNGbViGqP1Nu8/lg1NPXJz+58RlqIWypXLUJ+FXVnRRtyE/Ps9JX/3xiencCm8JxH2JuB2/u2ZzBT7tgS9mzrJTOAdETsjwyzRQ9HIOtVXI+WO5WvwgL2fdq9d/3IAV+FJUltVGKkSqvQx0rhcCgMohyO6WZdDPsjI9e3iGG9tlpeRwekux/LSaRuYnvJZlKtN+WZSONgvj2wDo+Jgi9IXpDaIG8CGV+He8yeIvReATsKpY3komab7DwYvDhCQbZLmlyUaR+/NE3mOQB4QfVP2cfRqoUqzT8VYfAtF6TYjFuKwaJeqGtT1OcixZsictcid8vykRJKbqxocd6PkJ6gYd3pqLkPymM3Iv/AFjuupKPlvocs24axo25reJIcRcNmyiHtSJfzuSD5FDgs9PUFl0rYGuyKT9tqbHMNGgTvIDIoHBCRRFfJaZAH1mgsw4zAGQVasuEUK7SX+bcLzaKdXIAPEXn6meSBX2sqO/Zv8Umm3MC+Yu5lm+5VANKfmI5XQZiEnZ6fDxKRHMw8/7hFezH7KCEG7hHnHudAcaIoMRffppCKz7FOyyvfLyTC4MoY4HLI2PAXtSzUBq39Zjqr1wmDUBX/4VlZAgebPebRCbj/bZniZ2tO3Y+j8ikLZ8Jc/phz8Sfhct4UEgtZjr1/vG4HI1BIaImlZbdVg/980oUeCO55nLVXS2AlopTyZoDCKtiKGw5j7dhwNq1+LYpB4OOYwOsH1Fo4OjEkIXCoGUQNiaTIZ0qsWG2pa9g/jG4EyTw/4gPIF/sfQuegaqE/J/AdiJuZO8raWsT2ZBMiakt8Mnr5ktt6gkvxM3+/CeqNI5GAwwJ5c9heohK2gGRl1KPnAE+ch1UrhYipSq6mdOV0yejSUj5Lsozc0sX+TVfOF7AX/mv7pqNDNnGJHVoQ1YfT/66fclmlIjrNHY+6Uy004fFbYxJvcB0Q7bfB+z6tU4e10b+zvGFZbnoip891aPFGy/fR5jX1yTOTyXp9FRqr5/pOrm55t/t4Jhee5ptK2Hz1rzSd3KPpyZ1OQJweaZh8AWzFfqwgiANkkUbsIrsEaoX0ThgEb4wBWAgmADZQ1o0dLT9oD+AOMn7tPmCFw4Hx2u6TY/HV3MpS9aBsYq4Pr/rs+tSz47+UUEMVncHYzJS0hBe3QOeti9ecmtaVW2hvSztnsJOHt2QmrTt3IAZGXbrT3MvG6jFPQC2Q6ma7HxlIaXAV8UAmFiS5ayLBjNLDFhY0Qr+b1cIerCimQ7FpiKTSba9XtIhRr6kHKuI5dbRY3W35YuGE+S/rmNst6w9WKAe66w+2LDNy6yGvEMjHMEGm59c27JlG3JEssya/pZklSKBuMzXo/yO84t5u/7KjUFMB0GMTHo5Ab09wzhdDexbOWUbQnvTRODORNkoueKmFXCtxlmvlsH0GTol9sr1VZaQbfdGqDlhr6QhoaaWxQBFSpWeQTtL+PZAgVnhSSkEqCb3OddNrtWARdNsB4vOZta9+CPeFon/Cl39uIm/B/rkoP2Ob7ihsKbO5q0ZbHn7llYoWx4slVUhNLj33EohYSzYKOwoV1UhUUzj1xQkC0q7NS2Qtab5V3COjmqwUeFgvAeulXwAJvK34y3H7weDPhIHx2I/oXAHcgdFybZWsFx5DAVtQvJLV+NjbZhBKLK3HMmL4ARy3u51Hh+iYGY19QNrIOW+Xk8d/Ou7Uinr/YZ7d6exNY9QpkUwjjMnJu4v5BH5owgRZG1TdLx7aTHAXI4ze+R6Zn8BWJZblce7zM81JINTWGt4XSQ0WXCj4o9O40HYqw7IxlQ3xqVQci1QchgEfNgyHCcwu0cyxkU6tAaQp0sYLJqXFhRfeQUI58AskXSvqTuR28c8SJayncgu9gAAHTFXhU8u9y2azpEInyXLsJdiR1V6hV67sAmFgmAXtMt8jlNggrRSZrbTB9MWRTD5X5vU9MszJnMYQuC1iNg1qNlzC/exlU2h/8t8RT3nUnmeCVuxZwOxTjwsUM7J7Rpg/ykh0OaWn9ezFkx6PXnILCBLG00jrM4tI6RNlZ9ZQLK5jEauNVlKT6+cQ8Msxe/QvmehSsKdD/pw4yPy4nhhN+lSIgbl/KkznoRT6Qm9SmBsMBoq1VlF6xNCidMIRGeb8OghxB8EOBrF8wVJ41xgAHA9eeD2q7bcXEJBNijNnWEo8B1IrwLisf71J/4EBdx91L6o6XDJ8x4kQww5tbVmvwTgXLs6vdBX0sCJTt/lk4ga1UbKLunoq9b/etyWIV255mYkYLa/lGsBL9xTBjd9P2g977OZrPPnNcMMoKnSWabmz4dedjpCHkDL3cuxjWc1FrTGzMsKI0+7kSS16RVaxQB1L1XCtQQnR0y5rHVo3qXQQzH/Ef3d/HiPNS5gDI66vA087YO1Y1oHqU8Giw/RpzYjaKOb0xHLne8gCQ3eJ/oTcd7BaWNiSmrxP9rI1tmC7poalOBK99ZjEt2VPewHwJK8v5p9LtY9fduEYF4NIzQIxtHq+uzPGdaYAiZKg1TMoRZSPs9yFo1fZ7wi4khr5T9WT8a9EDv7NKHi3vitFrtJfNqv/8PW1CVLKL4I8b2pPdOK8+t8uzIMl4NmsFDayRm3KFpbnEvKA/7XZ0OX0GJ3sjJuEtTd3DlBDJJn3IMWWk2DUNtt1Y0cJMP0a8qbTgoBBPfnUg/ZHHOpHLuNlcgRzL48zO5p/IYj2usao9f0ahy0EubHM8MVDRw8WPMrd/PgRLMOW9DLdziHcvPGUCTnbE68PDHn7WAAjjkIFDx5r21aDQIEhK6QymJZKbl8daLRIq6nnmZs/sJS7/2Ts17RU7+EmNGI3DIQL49XB/p8wL1LKXGJKNiIoE2Tr9x+dCaa0mAtt+PPmL9Ro1+NELwKq+EfEybtKUUbMFGcMjd1OOCv5Oh+XZFw/Z0CDvGlorew9OwtBMVoPAVlh1c4QUfiKwghNzZz2uLgkIM3wA2F87SiYq+Ki8A6FBQLXCASeocVMiIgPCxVfHzqVYDdGM3Uikv6HCYxUZxhUvEoOxjJABoH2qq7IOZMITrO1VXh2XbaFSJ5BZOVsD47L3RZiVf454UniOhds+Nq+mU3cmuvmcGvFTY8MsTT4ZmWfnRBLNhA8agnBbR0IlAvM3ifpncqj920t2PONL4R8aFVl1AjytOVGOCRxQypE/pMGpvpM7HL1+fmLu/Fs40/bHOtYxDpFA4/MEIOe20Tle/aK991DioKS/vZgtZBbjP7uaaOEbw5EosI8Od8OwUE/L50zEZzpZSUY0qN4k+ycEfa09WWurXKTmyRym9Is77srpqFN/RgIpegh+e/ZtwxtBa47m5zFgUuoW4QuZpobgX4NEQhGvlzf8ztew1Lmmn2hwJpwt/zuzvjLwlJiTtra61nv1eZbvWll4CfRLKfeBB5/riW8UrA7S5V1wq43e1jaBN2PJDrrfVbVKTBQ0hm97OHdbbQbcN1ujl//p5zMWtos54/qiw9cgKsR1ZUKEqp+kY7f2TgJIn3dy5rdvnO6vOCntcVHUcm6DeDem8OYrJoMlQCbTCPEwpZiafljYBbzl3KfCHT24wdRahqVR5DgiiISBh3udN5wvonqCFO29BRGQyi8Hz9BvKktuDc6dsX5P2cNQFRU+tBq6agrjOyXj3by/5oV2qxcJF8rU0YZL9uFK+ywLDS2owH6gjqLlWOgSvODD6Z4+pmZQBRUrcIDk7k5MXrfeme32YcIq0CgE9Fn5HhiYiy2jZTiQkmJ25xu/qlYHW8hGSe97YqGbykdUjr/iJMcD11w/oZ5rVLz/gd57/ZoWqLEgaQA/ePVBuhaIMwjRcc2N33RpA8kWnRHSpXFmmmb1FlCJIbcb+v8uKGPCiTLuOvrm5cIl29/zBR0qWkIFSjc5HCoK+yX+xXYWtsnyh3OhRIcHT2xOk5AkRGurwp5YR5ZvGpVSg/TYI9/QOsYAY95Y3fLPmY8Gyfm+UXuN9QwZQH5Aez2TAMBPit8n8KTFFt64JmNqT9VuE3JPGPmZTA+G+f/9IOkkdVcM3qkCmKZsreQnkTReciLaSjXKTPLyIKHoyEzkOzplf15fqaQ02JLb+M69PjxlE/de+o+B7TNWCx+zWfXxsikMDT3qC0/xQMhKML3lomDH9514ldI68oUgRGBaTFQHXiXd44Xw7D7s1v0eHUOQhh7VJTpGmp/cDg2MPr3vnZnOXCVt7VAKubJ3FH0uyGnPeLHlopaDTC0gSjtaA8VIUxBQDN+M7oaxDN/72NOCDqiChzhJ1hkSz1E41FlyXsccoKiGG2Gx4OXdVY+bww47PyU4265uFYi12FKj4x1FmBWiBTH7irT1H81jIQS7frED4RUMX59XehylOJ/7YjEvLQexmShAULQ4r1Iy3dtdDYvHvcEwjcFty+Wd8yoMqmVFP/Rwpg+0A06rJA+BjmVWjRKTzufnO3dJ6D4xS5kmkjqBF4Df3n//obAUL719S1GPODNuBrOxFqCkYmhpWoK2DhhpCLp7eRSvSpaWOldM8DmxtuYA9TtIkKAVlFZRUME3382HBfF6q/ds/hLMbXgAqGyC1GfGJyVfYXv4CFkrbqPLDaBCyG5NrsxKw/1W+REkG0t2qamq5XuxI8ijA3CZ+NYeP5bJIQB1hnQPQOJdCLUGjrXurAgzzSJxsSQ/EFG4WIXVPcXseZPjJrtImMqjlgY5Xj3o4LWw4f4NV/9ERGLkT5Dj3pmG9NiLBf5NScX+Mz453W++kFX/yRjRb5LloRnYXmDwDwFCLKV3DX5rbK3g4vO+r2xOoR7fj4sFeZ7SE8bjfwByupCRXFVx7lp5LrLL3arb2jw0IVAJ+HYVLuRjJPrxD81JoaHGiiiHmGX1TIDq0qNU6BoI51X/Uzl+q5PGNFQjfUPt7jjjycRkDf8IEYSU+Rtx1x91q7Oz2bwFt+zaHocDnk1B4ZGGuGSKiHh5r1u3ojNyM2ZNpXoGpHfbhx2n9XdERRmfIVn28IQDARTOg2PMY/ElWdsfG7F8jzpteiqE9aYrdvMGViRZuVvkJmypjt2rjpsr/M5S0bMm0KLVWqJjQucACHF1T+9xs8wNTRHVpV/qrvGqKXGQkwm7aeG5BxBOTv3z2hz4RAvmLdBXbMFwMs9l3zHCWDpgzsNzrWsWrLZOsorENmHJYUI02y4xbygvECEeAzdinOYbclAnMVoU/Q8BiKWszXtJodrhirPYLW/lZrOyCD8WfKRkfoTb515VhLKqWuR1IHgzsvzXOXNv7rz7IE+hmU1BpwrmkJTZuvjifMoQTvEy/hBWKdzKPG43CuVGzooHWkShVydEoqPpumEKdSP3wWIZOsVPnVPPZ/+yS6AEO41Snd5uiUrei1z8HkNpsyBtJFWmZc+ohf7hQ0VMQtoOV/0hl9sGYwIiup5l7IxRF5BzVXfi2zmYMlXq22L61+I+cXbYwQd+RLBr2Vg2dLpprotH9d/JEVm4673AbUb0aMjZLLK4aLqtVXEwlB9KgG1GX3A8zLKkjW/ZkxqcwTKlCv0d+7vUZbrZKgIG1KZOycHZy9yaOWsKo0q4J2W6BCHus81olutePJesumivhpMF4iiC/7I2XrSzULRJi3FTp8bmD7IxjoncIicxLUNpY2LEIECkgoLk5CY6sL97Ef3q0t8J97OtKvFvWXe1nbAEXw7jDJ/KQoI0Tp53ilsDBrHYCZ1hH/8ezDocP8Vms7BJbrfrd09dkuY12WOWTVGcEvIh7LvHsyt1SjBLUmHawbBF3FqxeWwAcviVpMs5Wz41tpeWwWAy1mpdLocMJY38LBdNe2irDjdsEOw1/LTQDdqqXeTyIbgHsMeLYY/wzl19vxmq93EIJEkZQ97MnPi821Frjb3ydI0kk+7eWdeKNA5dNW6Rj9Ovl6MoQFfZHQG1/z3XBki6m/HDR9cIhFA0YUWVe2QF9q/wNj/NMnyv/0By3HVYCi/UOtKseaM03NP2zNPF2fnDznT/Io+HJhEnpaybK5iM0BtEL75s6GqP0zW9E5mSXG4RPtf73kdCvwY8DizBgENWpqWUQM1UBZZ4/7UwLas6PMr0Smg2T4tChB8GX42972ZfcaqOmevTkKjeUaCqRJAl4VKS8J5d6whFEnMkkv98klsDQ3EMuAEhhhzz6Mv7CInw9btsT9UttJPnUactmeasQrFNy5aZarbp8jwM9iL5tGOyWM5sCNTfBRJ7L1Hu2SC4iruuDGu9PmNpipYOHppT8VUfXUWzDOwhVPRZMaB+TipjtpPyVUASIOs+MOWeTxPwX1SFkH56GtTjaPEUPDDdJVmNg+abWuPcBeG4iYOYi2BVGL5thtWyVV7hB8BfPZm1Xsavb3LCc7zq/PLKIuJ/1uBkL3iFRuDEt8Yqv04sPTNkndlaoH4DPpozVRGDo9lNcuQsC1WfHf4AHzoWSGClFdhZYo1tILBiCFn6wsM2zB12KCUjEuwKlWr4N0IdhdJM6oobCnD2fruhp7FIlqfLrzAz6hbYNivrm3oamhnqilvg+03aFLVqx5k0WyqioAmM+5sQ3GRJs0ayAGFMHsw8u/JjB5RmTTNfeo3tmt++8tTPjceq6BaQ4fE9ROv79STFqIUBNA6XMm9GJUcF4OMnflr9rbEMpWJbMJTj3UpbjlqYut+wB+DQzgIdRsjsdJ2urGjA2GbORcShSUVzJoOBOdw8IPKhs8x1gDFLYoXD05xrd+tT2/qA2g/0XRYwA0OR0hg5k9+dj42Nmx2YL59gH7o/2FsHn57+LSQMapSUTxIqxH4fOvuRAA9rxm9xFZkSQIMbU7iyqOEcPTjJWJ94+QEDI/8/YRNDKsUCTo1T2GYH2uEIHTvJCQFgFha1HrCBpoehsv7DDDAzgUbg/1HslAUik/oAdaieb6bJJohKMJXdQov4dLbdyv/fkc1RZJMY7l71yg4orCijpI2WPiR/MRD9Q7lLb8TDu8b8cxbDSW/+Y7/AtkhS42PQ376zBxRAQDhfmNHLlSlndSQxvF838+khcP1C9MUkDhNPW58fL1rPXYC9CnbAor+UGSm0NZ6ugXklxbR0ELzUmVcAh740KTyzp8ZMmukSvFKNS7szCa1tYN0dpM/PxiAzic8rdtxSEm3W7/7t3C0C5nXSiSBjy8VvJk5tXajL82T491vyNPw45W/+Q4vp6pOcW53sHQY4eB2YZUquo4vkobscvBd3NfzGJsDibryeVFwWuBMEH68JmjR8QFAy3+FarbbvCjJhIvuFPQ+QC3QzFpV/Zt1xMRV3Et27uRiBUkLMJgaZaOUdEmh4NEa/etPjakoprTZtsn0sMAa2PaX0EbLelkX5OSB8Wfjo4HEXWf3hbmWnHGnReVNXYYYKL/o+o3UgI7Bzc1C1YZb1s4Q7HbauAAgOEtL9+ahUEsMslNz1hU1+U3oqtPWHZqSW+rDUWaTefzBGVfoBTJSso596IW+XMv9eT2/6dHXIPUDFcfmDVvvy8jjiMPV8o/R3zzbJIKAtorxxGvDQffpss7Lt1geCqdtcnCMX/dwq1X+PF4ohT9/xgL2tMiWMmAu4GgUVxD43NAUpVOusBxhFx03ezZLUqDPugYfTqyGs79tftNwJ93o6Iy2N+OLTH2xPNjNzwDqaC0qxWkwq5EoB+zq+v8jRd1B6t1eVmECluXklsK0BvjT8j+MR+zvmMy+Waa2Vm56jyUoW8hhpMp5G372pzRrYQwby8yahUr0fd+9u4hgiqO1D7AQHLSbnerVsDRNkDkU1njHCwvFwk9MIchheWtMaZh8pAR6SkhqisCfWdVQGufTna6/b70aRwmdTwo0fYG6/2Uuz3HMZNvTNKng57nYxFbWBbzaiW03rZ0Njh7nWxJMLn972X03hCimxPg2yWtKRl6fKjRcQFFjpjb0gjJ1rl33AG8p7fRLEUMrKtV6407Ghao9MXlSUWDsrUE+hdgplbKO9WCQvLyWjLZn5Qe+6WpfpoPoImPVOGkYagjmfa9ySQUUNTdoLzzF7wbOeXnS1jiJL/jhlGijPoBMQ/ZeVo1oTm0WNN4bRR4KG4V5EjelUh0u5BdZTAhy1M3LE3R6VfwCQqhUAsBjtBGqvbbTmIlXYxNZfHLXK9VLPXFpyxXtxyutxr1NwKWm4EY3wN39nYWEDoXUM4rP1xbnGITjzWrrxmKIKTa8upid/XwEewPqm7yjxOnZL3Hn2P94UwGpC9DsGtsJjfIECoauZnInUEHsBeskNylrkVtYn9c0LzFnPMST+tD+2X1TGLXn92Z0MZskFl1/J5phmkAPrphmhUwiLI3THW3Hbk//QNd1z6gkxDcUZrjm1pyx6mj28QaCRn97fV8rOIEbSJJp0FIaMzX7hnQ2BMvemRYegzfuV3lP8PZif/sd6NGbViTyDK+22yReZCH6uCkKVhN2eSszXfbjLAa4EwzXdlUHnYUpAnQ1LvF9QSN5vZwt+2lUgBo3txncYJtqEoC+xj5CoAy5BXgNNj8FF9FlixYFQUBx/VSXPFzN8XoE3DquD+SDO449OZ9RgUHthoMhe+bYzYA0pyeQRKcWCpZvE3ivnCPN/5ipbWAuSLaERDltojdnADDPhc8pSKObsZ2E4JV6cos9vU/U+WcsynE+tc8vDmJkpkyc5nJ5KUN2D+EYrF8hBTAu++S0u8IJ9mgqftCfE6RKEglekVS8+nRQkjmCe1C7RF88p5/2UT/cxrN8xJ20A/unBaUdh6M4nB8qpowXUUUV8M0TF7U4QFjXjg0jp1M3FKz16L99iwaUeUkJlf5vJXCzjLmqLXN2TM//XH08KPfQSQOEP7ewn52yReHRMYbbzt3aXFYZyrljZvlKMFojzu/aLHQXpphGBnHGAVtvzCUMlrSy+GTQm7yZFjygUtcp51gt7FSGqmheS09SjSsk4MznWc3sFHcClbzvTIxe5Y7O0oMy1xTAREiqu0rLWb9n8/IhAjksMgEtfnN7cEBVwWY6/2pr/4VglCJJ/de/vGKnhAu5QC59y8hNKKhVMxCLQzQxTPY/yAob/D1OQZo3us6Cf/dNENI00FQm8UmL1Wnjzxk7FcqjGzNM2R/m/M9tyii2dr6YTxRZB0MjNm+r4+01ieJWRKNmwG+p2wwRrMYhgI8fJf3YZJzppJlbm5BOD7iCNTm/AbXjbpFaet6+MeLKZiVpiNtgE+Rtof5Coqg2KGmIc8VcJ3Mf960lYz93bfvUTCPGrpl+HRrHYKm8iq+5bb/vQ69cug4Bta+AC2CNt4xv/9vxl59gLW1NKUT1ErT3Mu9vOPJsqRZ3uRQwX/LC53G2HpLfGAfoFYEVD/eFBws0by8vDumF6qGHqxFvcNYBuXbYGK66opeyn4OgaQPWLXK0BkF+Cp7s0gVIFEh1YW027orH8yrd3bCwB4uWDkanfmq8dEirF9mXKUne5Obf2jjOW7wIBmzRW+wuabosr5Or+Q3Ib1adbargGeiwf0sTOICegIl2BQCQ5tc2xsr4OZJsJYS9sMIwNvT+Seub1fP7xoTi+wzo3DxMzREgm35Dgf1LjAlYlHF7H5Ckrk1b1+me0y1bUCyiPI7wguoijnvlSWammmiBXV0VUgXt0EgHI9v4VFhiapvx9gZis3WzXcEUfdNWjS4l09+K0C4AeFamOB9MxHNqhO7EDXdn4e2AP/cbkztzKUPGWa/vBd9dImwCqjvpf3qcyXMW1pV4pxppAzfEBx5OtnQWrg5o5FuaESsBLUzTNe6hbmsz5uCr69SyBMd+SC7u19fZB1/nXmINdQ2vYh/GuWZ7Sr4LiYfxerYmAUjZBuiFzAPeXBXcDbZpm/pXtx9n+bj3VH5g75yTbY6wBZ44BA02IL5FUky1AC15zZ4ufxu2K5YMJU8coCqvcbUgp3vVNxkPN+yj2XMdXqGDBAtCESDZNve2pTq4lHp/Vevw4gevl67BZCnP2jQgIFfdEeLgzLLHquKHWBzzpPJDLxNXIgjtMSDVOLoh4HMe2O9IahoYQ27L/6E/vrvjfZsrnypeqlBRK5UEJXniw28jeo2SEYJ/hwOYbljMFqKEErpP4cq5uX5gkpYWViHc7eR2iPJs6dHMsabRVhATLZY7vIqjDP6cGJ+8RBKpEIEAQNU/fkMPso/IEKBLZazdLhdQ7L0QR0RhvcSDp6i5AoaHqolrtBXjG2FENYNn4athl2e9nFkrSVwiLeq3r6/tisai4mjvtdtPbgyB86Z6lNArFU3EhmA1Mckpv+Utq5msjsKdZtV4VakfDqJEJyOjg2b1AY9Pp5J6hZXUAGPYIoEtk5jiO5du/m6BSTUkyC/14c2K2PwsSzfoKQwXemkZUjr95hDxwCzNi8DjhaYpynfox8AnLAvY++FwmotxeZIi5BF3oGi7Dvxd0dH/ZBfLKKl9BS4cysk9g277wswBYBC2LtTtS/JBmkqCgy5NHHTCa+jD27cNJhKYO2V/fUnwFpOAqvmMBh/Hpz18jVfqLhEno4z0lqed9EGVacNmk/aNXH+zxTkv30+JMJOlH/1PYR7UbpX9LjzmbmBpdGe2eSld5d/H7hQsHegRjImOOUEen4A0URyv8fHuCYY6QYONDpvoqaRqxDS2iXK/0+ZNKV4NoPF19pJTboDJjXINUbEzvXpH+XWePBPQwp2xrwF+QDGMiJT621pkU+EROwj161EpQEQzVRRxj8zg8I2eLk/mcyExFXSdTir63FPJxG/SqvmcBejudq78e3eb4em1uzlaIkRoSdUxSv1Pjuoq9mGBG3LDn9IsREy2GgzPcDITsMymNvuQ5CB3XEVsvUeDfo2I80Inhb+sU0DkEuaMIgVOGHvejuKt2xYbbsQ1WCn9t01SmGwroXoG+91SrpbMaFXIkf6vH32PaXoT+RMGVK5UkxUmrNir7k0IS5aGiediXkKlSjnnCu/VneCHEKPXCPBbHDvifqpWOB2J9CixoUyg7H17I3UU1+qUYMC+F0w6ziqxBu3XRW8LklQEaNWZTp+2fx9uYN9snp+sCM4hwQf3OZibx23EHIDqSWsOHBBU1+EfmUnvue1/XOrEnlJqDd8EvV3k152eWWJABKoKDzg2r2F53en5il4n1hKPxlF/jQiFiEOj6oxm0156O9jJSeWEANUNPwrL+dm5cDquTEt4eOguveTI6ZSY4FjC96q7geI3Wukr6y2FVLzlla2RI3qitnny7V2A06d/QcRZIvvW/pzS2eryghdGHUKRe7JyiPY8Yz2C1QFfUAM/HBUN67Nd/IYkce1su4g+4hWo/5ij2Bt/P+U9dl0hBh4sS9C+Og5cnTi0c/EYykOJSYlHKPGMtH2qCFtWNao/toPqWwoV4Fwn3erxS96s0ErJ7T9ohF6R7RNAKlbCGqiuZTZEaUzG6nFG/DcIuh7nUGAU05vdMPjIsmA29et568448AJgOwhqiFYa/KsxJyY8boWXjUhv5X/16ddZo0/hGrsRwUWAH+t0Ipe8CP0AD6guYMdhIGBuUe6p3twnQQ4SeTjkVGG909JDww8QTHQxlANYToveiirHhcQte79sTzHn4SVWee2JtEqg6dKLroPYi/1WgTBy3ronD53AX3I/0v1RaOOwC1YOjKS5YLl3smmPemZXYD0I294sUn0PE3QQ1QSsb8zRMA3I03d84AOHzR+iQ+QKxFnhSdcVy4YOmG2SY8a0oaN1Rxy4atuCGzF7YW4T5aHwPa/3bevDM5uzBOYnLgDPAmIA3UzAElHG+kSrgJm6G0NUy1pho+Dt9aZhoC2W7FR+6kGQbnyWP9HF7CtWRFALmODeS/E3/ZRkgB8mtcPsKNLmC5aWzqa3HV1wmhPPWA2Fvh10RvKzGB4AKH2rA1wzK83PKhvbWHsOzflouso2yJTwvRvn8djh60BN8vgPWR27ig4PpY/WpNAPEDfzbS9NqI0WrHFLb1Hh2qW1QOajq3v2yBe/XtP43ccTjgDCF/nVhhVYsrD5Q0InS8AgG7U9MI1rtN+roim1ffdSCD98UO0LBJ1SKpeMUL7MiraV6pJkOuq0TwKXnBJHw8Tgx/vLrnfVyKMDu1lkh0LC4TcP65RLaQnnTSBSN45CcRZv2dpXqkb+z5vN58S7ikaXGvhEy50bdO81zl6lQa13zRqOB4BQAsClHgSHvnqh4HUWIU0EiWI12gVwCwhbx56P8Lp1H1QFR6rip8FjThBZJZVI6F8qed8IV78jjF8Yl9WTudYezAh1oMKqcDceKEo/UP1o6FgGquI0ld+6IXBwOcZIKXVanuDoXRnwmRZeaZgu2PIhbh+z9PKRLY8XsG1a69p+yIBBUbH5UVoi41snFBp+EWFnO4NbHWS3Eo6Hsu8PrEmeJut0M9Qa/Se8EyQSdT6wHnREJS5fktMsN0hSE+A1biVtVirmQKT/71PnQCJVonr0IT8jQyU9clwcc2rNzP98NSwEGBB1z+Hz18sV7+0NWwJGjfMVFIExg28joJdUbpk8DpN0TasZMu+aFfYYMfF4qkZJchruEecgzDDuZZpsBUcv9p+VMDSW8jRO1nZGeRtcuVJgNSaIyFyh04OwfyMrLals1ZcL+ZFZGnE4HnTC7wdhL4cWShdWIy6si5TtTQ1lLYF621xDR7bhFdqlS/6cp+sWlrQNVjuJ+Vzw8jxkZB5UDA17szomuXXD2ERCtPXIrteEpFXwoxMr2+2SrmU/kzl/dF2lp3d0GLEBUO9MBtsIWIP7/YF56SwtR8TW8O7U9A0JDvzxbQcVb+i2yVORnP8htAV4Psw1I5Gk/20HGgYjYeypWYGE5fahHQlWK1WuLxCvUEDDTWyt1KjrVR3CBoEm1ATKSePZIEUKKSrUNWmaleUGTmnmLhrv7vRAi+1ZQ1Apx7tAQppHe1LPaQnzjuTE4wXhtvNG57DqLfijY0ipBbuIbu/nSYqEKdIdyeSGUcDLf/rrR1zGTULrpnyEb2dRFXHwAB/H74pEmFUrSJPva4WpBMrsC5seyvlKkOiPVXd1/VnNbrsiprcEWNG+RUEHu1eU1XcDN+XuQctfGjAqDzWZdcQTXDMD0PKqL01D28BpsT+M8UznXx2vS0fsrrpefZ0UYKiPk1r6qbKk+6OjnXiZhUzd3j5ku9L7U3Z7JL4C55Cr03hF283/0uy7iayixL1QgGLAGck/xpEVeKRaoyMYzYtcDcInxcusy0twld7EPk7W7bmYtznI/o5P+rwIjmSeU0vLgZcGS0xwDARZUvhqGy0iLV0ctjzCqleiMOYrPfsFdHNZt9N6BON8VJ/r0nm1ucHtPl63EBgjhylMkGCrTFrrjZ9CTpta9FaUJr5H790sIPVv05hFr9TablGTTPtSqmxnrHwUCT2rWjNNohSz4pxp1YEqNJ2quv5M8UWig+WSIuSerD6WQtQF//rGvneW2UzZ8twBBnEB88mx67BGBX6uRF04bOJGBy+wo38cxumMampPFeMCm2OCJHcYXQd2nm4VuKlarEUIvRl61F9+us/5DWXrZCdPn2l/Mwf0rFsQbV1+leTy96eqXwdSaUs5v0Um2tyWWdArNW0s0STWKZKnBGabiisjmbpRBxoR8Bq/eo7hmGcCyOFbdvBc2SHVSuf8Ed44B6CFrBGcUAG0pHil4LTaP8JFdFm6C28uF8IVI5LCw8c1BHxh3Lgqu2XjVUvvVEMH8w/U2P+YnLL/hHAZ+6iOCs1FAlRCIPhqSxCypp7ooTiIFqXb2NoJk18WHIEAudI/ily8z89Of5SYDtCOU377KzdFx0zkOFluowYiRtR6AaPY12o8bZShXyX9rqxq3rQ6q/nVp0GvzjgCNyDRCnZQ+4N5fOdAgRG2PFmiK6U6bQtKP0dD8uRlFqNs+8hCpyq5mx+cpgmOJ4w7S5bs/ZIhysKJBebtG/amHd+z2DB9dyGzl8O0tNcVxNTl98cXSkqV3XGij4xRb6BgkXBXZfVWPc+AhmIlxrw4pZdHrrfi09CpOkx3kpMsyoU+OocAuy43bGy9/jJHKn6ETNkEMYNxi+xGkb0VMPzHaZ0oHdvbvkJ0HMWyIywmhMLf4kT5OEGnw7iO6eKbeQgqXcYKj2QaqGRXq6OCqaxu+K316u4SyDLNicrjPhlQSi+NoeofCD6GMSH4ubL7NIoiWGJTtslrv/cMYD8X9R0OL0zplkWB3X84ZmM6R1+ISPVvhvGmh+O18BdPmZoSHKDgngZeNiPGNbx+nC5sAvaT1gohBCSHx+92E9twyQ+bRBU/KT7Fn6CuutKJjfYBuGAoBJkBJM6LcpIen9NTCg34sOlIm/cMA+0jVnpUvIZFN60e/sohRhcrEyHmneP16K+nt9+xWva68RmNDI0LuJw8dWykD9JKNDTrl/QNDcSt2+QMNS1wRO+GYC55AofKPd9Zr7/J7EuuT3KPPKf19nWtNQcw0GVjgiIpXhUh8/WAJL5R1F3XYxJ7unX1Hm4PGxg53UtUSG4wJXjR0+OEWAAO5EQHopQL/OpPfo2+Xp4InFtx8CD9PTccHX0hrsIhfh+I/V7gC+7Ws4qOHZ5NB467Oi0sJn7w4qRHKAKuv8C8BAiGpViqSsBc6E62sVRCiTwYrCiW6ctPcXW8XSJRjDCmOWJLu4spm1Nrzyr2u3JMY6Qzb2msC8/6mdgSyWzquv7NeExRQRiAo6tTTuRZeg+46yl2LoB1eXDAuPQBcx7DEixIW3YbMFFgRSfPyp8i6gjgN6aWcWx9YmPC89m44AWXiWz/M26j1wIqo0X/W0C/d2z9S6+2JfXQsFNfaI5/2ZKKc0mJoijVo/lmn6bL9/BfEL62fJT/qboA/EGcwKCvaScv7wWxUKIqzgn4GzWFB2q0m4Sg8ZbU7GWtcVnvfOOpBwu7NzLahlT5Sk7rxPwi3WxpTD9Z1aZOp10Qa6Bsc7yweHID3rOolEC/kjRKwMbCcXjl31k2/IaXnA0f3Wyl156YfZCRePPFCQ6WdbldQ1J+34Wt9/JN9oZRrbDhkTmsW71MuOw51m7INwuzbMrwes3rEFS2karv30YgdWiIw/z/eWOguazZ7LV3U28NatCDOeiYF9dkTD4exX5nf1QMLQMn2+kFYOnz5VvUoce3gQKL5RdnsqlG9G7InLqQVqDeSYTogQSXXb8gf3Eb3Xb7wiBwkcO7e9tzRCDSETbNwUxlCWWkMX+FN68JU9YI6dGjnSEVz1okyzHCGVKBxOh9hlW77KzlUMmyJOibrKdgq33XL3N/1IF41IFRWC1SmqA7kwQrVQ16uePD0H91WzNbzThZzE0Y4YghLbFCGTpsZJvB/KzCh4N11ZivHi+3mpAOL00ShfBmBsUorJN8hSQLYvP6iSFl6mGjhaFirj5yFX6N07e3MQxIS8/u3fAp8qkSz6Y+gwn7aOqjSJ0+Quri7/UK0p+7MXW3chVXnWMR+SvAvDbe3lg0MCE438ZnT0x2AjnjBVMOQxJp8F5p2PahV7ZkE0UEtgwcWIhtplJPT4u+RnBTnghGDU+bsQXtwWoQ+5A+J++us+ulfpilsiG1vcl1vnLBLWr5nXK7hdxuDTTL291k6kbTnp6OIMI3OmN5pOSqKp0Ki6dYsGqIOOTnBkbp+HeMXZPVCMmom/g5KczFcBAZ8+2pficC1uDcTbNSL58hzMzGqQZKiRsmodiXa9ocrQY/Pp9wa/+HuXG6tyu8PyknA7vROAVBwwICa+mEoltZqKlUOQ3zUopq6Guyy/DYiGxiEbzQA/3ylR6vUxWdP5xoVs28Vn5MLNQikyhq7UBJRRgVAIjjdyNuNois2QESFed/6ETaw5S+rcWupHZCfJ7Pwf+jTYalPeWLj8lfdxizuMUV5H8/WEnFfD4w1QbUW15ysByXoyp7S+pMf2hkh1OXdj2LWuQdVQkOhc6rO0jJetXWgNRZ+Wga0AqWRyCXqVvgVSYg8YeKRJde2j21HlOPacqmVSLQr/Tv6kahn6h5x/FHt+gzajNG7eSEWM5uTTLCIC39Q0U5n6mzlzSHxPbI3ka09mAhfOA6ik4hrmRW70LgNevp/FsoDKw307UN6JSpiqYjNU8lFKIKea4GJ8NyaCZbrm2q1i2TYXgh/tSVcPuZ9JQyUJRhDX+wkJIw0klg1WkQVOzv5QjmqZ6tBaN6XNBvDzxUmtn4Z+C2bPNezjFCoKjhehFc4oSWBUMOSRvwdyEi+PKTKVc0UI/59atF+HOZMBsYdjGy7GfXPC38Y6Zwa+Cb5v4pH+VTPhAiBWkf7X0G+quBho8SpwQ3Rpx4otbZaqsc6BQ5mg+2GoF/hPvHjH2YyGZ7z2J0BeIkRMMXhdUr9XGBFWHKyBDLkk1U6HoVZ59sB8sSRwb/ukc7AixPoAhueY/JFmkWe79ntOWfrwOYbYIA+R+BmqF9jHsTd0ObMt8Qoyt55pQEVETNdjX8WamqY0FEo3IEwpWx2avn0fIEYjfV5oj/t5NK5RuhdHUPsYawjt8fwjc4Vf8z5dfqNUxIrxPIV5hpFx02gMRF9Naeetfn4+rcKaevmc1XXvPYZkUXtUW2hQV22pmooBM2r50Ca8NkFVQfCAQDKlBzh/Dlzhe3ija9EMWymQWxp9h2ISZxLkhlP2x3DFP2p6Yw9IRDGEZnI5MM0iyELUI85Kk26z59SZB06+I9XNIF0TAtaCxGo7JkUABGLzC0HxRkpn2djBaA6IZKVKbVJTjmSfVufZHWyTQLjxnF4KL495W5iB1TWMSD/iD9TU2QXG8kTwThWWvhT0/psgD4rCw3nvcGV7r7v7W85DvN42gnNBdLR2OWQAX7z6ITTDfR3rlwS79wWrimyrATYTUd1yl0yAhgr6JpFN1epjsxXoBwfyZzYxbiSVpM5xF/FbXCD1MGzJKheIGTlX1V3uT/3OvNaj0pX0dr/7Uxzvpf5r21H11wBFKXijNgJY95UuwLLDodSLgiTNHxZXF29YRDojT7Y/cUAQs2avrdA7gvGAMSjNBskwuN67WzVc/sA/rDx9wrCmokbz77/iCNisPNHRDE9pYKo3gskpdR9s/w2d9J0QYxEgaonjQOJyyrDuuwwNEE4YftclK2n3EyTnQwdJpQ3fcpuK1r9mSCdOdWzqC3w8+BUC/cHSK4+IJ7ETeQalDN3tkxOLQqmyGF24jx/0uuXlb5z5H/QJVTWONWxfl2mW2uHuGjWNDCuXU5ONUsAQn5gn02JBamBLWqeaaxQAUIDSohBoHr5kOu/hjPhYNi4fZFm3wEJJY9behWzZhcZE+ft3SazHzXcN4xfW/doAy8k1RpDtkNBRxKVArnssDdciRyfkCTG04zixWjPa1d65G9Dj1aJE80MS3wpX7WR2Xz9U+M8uQqTIo3feCbU8i2LY8cwQwiQrRY3tjvZI+Dkh14yLfQ2Ci9qFv20gd0jfBO6O4CgpF4u4Hzmn3QORzNglUarxaneRXPBPix57FlNAwsisPlpNMzavqWiDKi/kTOMioVVmTRTm30ye8J6ktZyXaIiJTTRZeqQzpLcBArOP7HXDXxg+QEzhcH2ZiI2VT+SGOnnzmTkANBuiBr2d3d/ltgccrpDzsFQSKTgQGnqiGR3pwTOvQ1oHGC3TTR0s27edp0KQ2V9Xic8GEPEZ9FtBfqrLkaYQHa7AJqL80ugzovkKDxdNjH7GkqSywg49qwTJA9qR73rwblJDEvrT3iXpUiyY9UvfnVXg6Xbrt72zDD0rllw7cAu3NvuN4YVSF0PUJx98+DzJOEa6Ap/hGsF5CKwkWHIsk9EsYMtFOOFiVIVWK3QLweMy5hyWxrMlFHjXfmuHb/UfebOIVFkIxpmDJzO0jyIQ5yknmPthcMSwVoXBKRLGF0y/b8+WpL3sfYD2h51O9QwH83+bx923+zTkPrLzrmIU2WIu8rDFZuCy2AV528hvGiKPS5Cf5btUIw6/81rTDP1f9xWpACE6MNLnKcutMZmom6qdhk+lIozDgF5fF9lvEL0eEbEITXHRmohljNTS7uHpO3Fv36NgJMyYPXU29UIX8m14O5p6U+woMEMy+rp3oInOAOyoZNVYnCJWfBQb2ionzKx8oWaCTQSrryTAhVbxlwaKDSayvulTTjNfZeYU745dpzd9tsKsS/y3YoMVZUdJ8D/VKoyrsmXupQywegOBqBktYWpfu+Y3GNkPcqd0yOsxCMhZM1pTJyxDxjp3+hAAJYXYQ6igRIi0JSgJvSatFdVko5K1gB/q8MmgKaU2iaKZibuE8XoqPSRAhflgb26co30h8OOoQXOFtUuv9aRYMplYqsZwyie3Vb4vzPDpMdl8wH1ULd938A8L/OH5VIGuCj+bwpYg7Yy+e0iyvpga+j2eJt+z9FBZAhOQphuYoYqk6AaiplQk+Gpf9PHm9BToilf2YhhEOOC7ZUoIitV6Q0KsPM4phe9o1Gql3O7FRjyvJECNFiHS7UHZphodrBl6LgO8zvJM7OQ4GN0lz3naOXS4/jsoobizrZfLx+/VdHm70R4zO6gxwqAQjZRBpanTR4s7SEPxl42XfmggtQ6SM0O3DVrZSeJ/WC5seC95JLFND2F8JWQ6ufwmzLc/uMGnbCKxUQPZ0Q5NqzQJncaTT+1NK2LwRwGCNGzz/mxssA9KQszW7elVI5AfTcbh8fum2iUaUGbMRwzTqE4MJls5UVAlPn4KS1D/40XjTTO2vGdehUFedg4CI6DnHPdVUmXWERsuD6sikdS6Gi8wAVFQqqAh+yTje0K8LTNS7MFEESPwd5lcZgjXxaBfz/AYKUGPDzSQlWur+1pSoZlYxus+JVXEMoc+Myb7VIEdWfk75X9eJoFoOWeWYuuaXvuslctVsbTpPseiw+gF9SyEuxJS9a9NZ5DtsB9nvUsFl9698GsLoZWkGe0Q2xzrqZduq5mLKkk6/8nF8Ad88NVDOGJFjiPjr6ayoQ+xeXz9QTWskn7ne2c7v0Cq45Fj6o3BRKcP+mJjs76jkyOKcLQam1F1Dl9K+AYcdboD5ozY+Vyfk5YNfIj1yDWuO+rrHlJV4OeEFxOJNuvpbsnQuc8PwDOr9o2VYEmXrTQStWYr8I+NYQJoV/gopiqfmAFRXlyrPLlub9WPyEXU9P1RZSsPe1BAY/jQ24MUrWEOXrTOZ6lhqEqVpuoAa8rC5mmZFtF1kT1V3yRnH/LXdNZZ7YFSkXmblwbPopYFiKbiXU0zF/YQTGlYMRUMt74/L17TrP3MSSsh79qbp8KY0WIdGh5AcbNS5d59X1t2PNWxlb81qZ1Myvav7N1z+VQeFKK9gS0O7KzjiXR0qFuPNqWmGIxK6Y5gqwiUmCjA4F17iu8aa5dWyMrq6qh8ObSTqq4Jv8si1GpXB/435johWv/T8+ePz2UkxNNaqg2j8X3d0sr1JsBtiWIn0Z9t0f/JMHLyWn9Oo2E/Y0OJ+jweRFlwdEkHUkXm87ivgATz39flVxWFx8HtQKpn/bME52CTDLVRBufnUdPqo67+n4vhVWKO8RsceuoioohV/Ps2rHz6t/tWY+DEx/geNUnG3CpJMT7oWqbvmQXjOXvENNFKCRL26nEqn4H5Dg3CS38l8qx2WqU+eTT2HYYlNFbSr6Ph/LFELwIh4DTXpHJ2k+MBTQqfVp5ZLZAQMVMR+GNADrWpl4SILXvMxiPX0ITdKFlbFpCooefGyLlO4xXU0miywj1bGO7l7AtXF5oogHNpDpCEGhY7AnlgF5jPJD2/OOviBobH3JdocpcIy/cP3rIHwaamLTNhDDMQ582u9ohBmffDll3OBRX5R/WaXYbsi3tzqhBjztP9RLZ3iv3/vg58KDCpkYBiwCX5zNhA6tibpP9a0FzovJihWSYJ1PNGPrlSS/m1L+Z7xUglechx7EZrw19ow19j39NSrlg8jbJnFc0vjqqtF3r4nz/fRnxLS3beT1KegmsozzGqQE1vySu+y/IUgANs9pObvsd6Ee86+Vr8MvRpwVwy8g8hZi7XI+jgmgRjMVQKbbpRTc6CsQkk3o7C9dAk2nw2AWVhAcExsEZDn8nuRwvwIx5wA6zEyYQYNDJ5wW63OA8cSd14HTygGdCb6iK2B0DfNBSebR1a1PqsJy/yaqKWYIzYbSBam9TYBNmlqw6tXTpBVrAV+KmjsSJkmESicNeHkBdgID32X+6vi3NuTYn2W+ARi45tU07MJ3x9hKFcWX/NupPHNKmPROPkakJ9k2u7kdiRGrkv9928W4NqubCGfb6DUj1OJaUNUoC4vIlqJoFM+tTy0ZAZByMDkCXN4dKU4sx8STDo4+do6vwgF5cLFMYkjjMfL0PwsRehzSLxdiAuq2wLie86/8emlCSnBN9pg5hWSY3d5HRPht8zzkD/hgvcE/fPrlQavzdKWv0Z9tvIhLtcQP24sPcDxIFC7cT1SVUqBTwjFSbVYMoRqmhcBbsfcEDxivifUfyUgT0lDe6ECectcAX43vn3WlUXqUnqLoCYfN+MxiAnEEMrrzXfuIaXVm9yGd00suJKZvGnyy7/PkboaqOvjjzpSXLQvjkaaFgc1L9QUeLMnwUDntbPeVdj538ia52GeiC7dfZ0wg+J/+bp0p+gA2jvOKfVyhvangNUPgiKHIkNCUCUgOTI8IToLQHyeq/NNWxRVmGPHOm9TP1zU6ruPC0kOl8Inx26r/h9rP4MxPX+K4pkpGzFqWiAdeZIeXnW8LYx5xOnNPz1+E2iKfXRZknCs2Qs4PLoC3KaP8FT4NN0D6zKVMCG0537nuz82WSawehxbMLje8VelF8GECtl/yDOklXuGqr4Dy4fYVqoJRQEfVYr61GlcxBiYYuH6Dk//D4mQNUdpu/BFn7QfddvxVYuJC6h1bBcofyIZz/llR2qfYlhFpJxDgZOG8nBMQdzpOkPVtRtzV+4n1j1Lvf5uMaEuQs3z3W39NSlPzvsLtDjyrer6vver5AUMxzrtBMRlhVL1iN5t+pwdSRr4U+OKG8m8/jdCJ7L0Y7Z8nb7F4/EhXhYtp1w8WexhVP/vOpE6+6piKPd+GlwMla4UgWk+S6M+2xkfl1pwhKeOGk+cdw/CkhhdJpjaoPeD7q3hZE04zuU3j9BNwQF0+bIR6UaHTVnlhTuLX3cJtlcpWtKNIQuzp4eeVGOb+J1NOnBIaRPaZjJBDSLhEr1ThzHPfERZJszGmMmuSXIFcZYGucW8ck/WCjz4vgnBUHb0mqkTpV1HS5oNUh19aajGAVHeWbgiLDZ1C1fc8NSEIfJUhW1erFxjrs3TkKA9qM0nuodyBnRlbPX8tfE7lovRMrnRmv2FZMScmcxT+dtbmI0g1oc1T4NCFOT0x82LFu2l2kJ60g+mZlBfH1ns2K3nqof+vGFQXkAkgefY/hZ/yJmnPN1r7S6pcK7hp0PI3eSg0JP37RpiSKEYLY7CxGm2aSveJZrPzjU85hucuIdSNO/7QndTYJP2cENycmK2RJC84Ar5hxImYHgc3/AOwTaxCTBk7gczD5zJs+vac+OgnC/CJpo+CVfhQl2VdSqjB9ZPFWscP7I3iMnz5Znz1csOzwcW+Hh7RFymPkmJfABmmS/VGGbiPedKXKj6HBnpivIoQgJpW+qrqOZrompv4q37J4TDydhG212SKz5yfyO7E8Bg0+5j2ZDlIa5ljz3ullOIZteQV+CiqNwecIPeWuSKszqR6lQ6LD8xiEngTzcCMuGfnipu4wkDcaGPhHTmOhEvMk0dCoTfUQNkKJNOtT80Z9q3poiHPAe4Cskuq4SyPeVdVAijtm0XPNGFdlzyRZLtaFqiTg6bbgbhCPurxGTKo82VofDYfoU0b5eRkHUrFyhKo0KJfYQdY3EkkPF5YUpxcSw4GgKAktKMXdodvlFGZBBfoPf6flrrdDyL/37Ajq0KiSAm9U5FetuCPuzQL7A/EUfPy3B4BiDItNEt/x89vYYESczq4l4RwNXTx/A1o4u+MFuzMz5ASidLUqvcX88LyAUNcg80W62c2nZrRPrHcdEZy8vcKUkKNxBibF8QegSYJ050sUv1YSIMXWFpcizYyiJEU44AzFLuA0SH4eDCBuPUjvT64/N4wNOcAkrNZbHD5GS2/nZrx+/9XhUD2+15kItqydKDJ4dxmjll0eamAn6bwWzoEsNr6LAeDk9LXI4K8jBOoc1rW7jP35w+U+J8V8pfKJ1KK2Lp4sRE8wZ+XozZfLLKyOSEVH8wrkDRDTYrXg87TqaZM9BF1B49928fLUArmkZnfwUyoNsgHZ2VQoCyl4uqRtmrO+1nHLO0uujYfwtgizhCX3vgAa+/uL0KT7va959PdmTM83/dJkD0rlmHRQYBcVmY63aV2lKkVCbP6UdH7DQodKgujlk+5kb5ByU3gs6Bu0VicL6n2LO1zJR3+rWmzLaKjeD94sZ9QKw9z+CPlnKTYVvRk3U3YW3YQVIkZ91peM5pYqozsjF6Z7F2yth1s6/wKgS8t1q3dZxjMQJ1xxQirJKpQ6lfMQF9yySXDUs6X0XMRrER8WxK1QXEBqUlVLOEYUJSPmwqC0HXXvgG7e8QaxOKHQ8i+TLeaKiK4ta9SfLMLdVeIBQxeUTf56z2LdMF9r/mgLC69v2QUMN/zaWMGxndN5RV6Q0irCTRi/KF2auyshGRcta4gA15q6LLGYVdH46G+B4EgVDz4NGpaSruWvvXKHBY3DqXHvdxuQmK4ZA4ZoB0J7/9/S+k3Ojx3fn2asj75cZe7apd9G8FSnR6Th+bK+Lu/6cM80E3ixDVcZwBhCriE0XNXvEheYJMRz+qsVUqZl0a+7encS30RQv6yPuJ2lYBuLdOYT7RmsHd06XvcLreAT50rAjeOMVHQ3+RYVU4tFPgTOvB/vj340iJqcr2K6RmFF+YMjES6u5J+AyfnfHMoe110W+uL3ziyG5saLVIj1T/f74PpqUqKqFV/+EGugw7Wt2quREAuo1CMCOFmT7j7q6YqddLdfvU282tq7+TkZCis7dYrZcDIayQO8hD1mQXAwxwnahHIc+FLsQcURV2LfWAddkp67kpyqSX8P1Luj+1sEsrbE6IsS8mhdRU89evVlVJH0YNSXCsX4iUzakomKVmZqMaE1w4RTKcVS3rBpHYPKy9baIQwhUbcuVJUav9Q+rgyiGxIdUqBacd7JxkybdF01GcEQ1Kv4SvV2Z/H9DTI1GBwP3XTBXbc71EeD2XPvKnyS0LXOYXJfauqdkfWqxPXkOFSwV0WoiXgCSLFFHxCKEpXa/DUxaDEPjFAujqjOGzwhLEV+lHtlcTRgtqgEZ+hsYmQbYCorrlsChMKTbaTzT7Qnl02DWMPC+sBaVCDBygrGWAaUJ0caYMKWtBY4Liap2INk7ESV4n2ddTDgnK9mX366lB+OGkuLj8Vp5+NmwmB+BkPG2WRyFiFZMF26UxY3vS623QbJQEwzQtrUdjwpsZXUoziM3/CmtOLEjk1WCSLmLY/9J2dDwtO7smE8Wvcf704uzdTots8Cz3NXDgnE2qO4ybl44yU7Gmsz6mhJPGvO1xtQL0177o+HwNyTfl0HAY9517Xx0tBHbyEQvaxyQiipjpwUBKSb0vvVTmTXBx3nfzQ9Gkri6Z4bFo5G9RxVy/tb0flbJNO5CJqKnb3Kcqjdz7gyNDkfe641Xli4guhq82tCj2XfKwKQRUIz6QqN7pWWpwG9t9drNWnIoLV/fXGlYuwa17eXA959vLOxZ/M7FI9lsIXWmtEsHsaHWj9OCLqCGZ+MgpET7DwzI4/86soUQENmA0oDiwoojdP/pKcdwAoTB0R9nbxyjSqEoXAGwSJ6FB0SbuCbkMG24rBznGmpii9mBSJybZbgK92Sa6C11Lgy0TiMbLtpBYrvUE1niPBQVwD4xE+XzGalv+YV8SOdNZuJEKxcr98Kh8Db+IeABknkk0vCOI9RqyPlMKrKU+AiNrM7AvQ+fzZbW/nDXdaWxxL6V3Kz5ji6aznX4H3QmANaGkZ1ms+XMUsJxesDQ0x3C6WaFjcRsPKN91qkyNft3JmFjoMxmXPLFPkTT9heYO/EYALNGmBKao9N6Q5K6ghRG1aWTG+96djB8fE0/lQvq6Gl9NtGvG2wQkMFfLvH+T+SSX/Z/Zd/pMpKpCxW/tBhyiMNHXODSM6R9rhHpgmiIj9/H0ncOpZQLUHLZpClZ3OWA0IIdMqPSSVXchsyPiyhXVHPcEALfQrATXw/AFZknSM7711qXgpikEo5lVJ1DwI1JQDGDMLV3WB3ugBFWQMcByw3uInK7i7s/XUczylfdAvSVHey9Uw8cIuDc7o8AZT3gVSMMb0IqhzzQs27hu35OIrDDGIGlsm9GSG/oqONOnSEwAskj4dZ2w9jKHMcPZgX1vldhMFqq/xe69IPggxXNYvWiyE8y/OksmVG6gScRR+8BJusOSCt9Q+qWF45hruPj2ssRobIEa807q24JYN4act08Co1eq2CD7HvElbv6RscRM20d38susSbN44NSkMLnK1Zx/eoYo8khnCTBPpRdv6h4jnOtC1VbY9gMNjJwYq2CH5MtK5oLR3pK8JU98qj5dVUicat5Fed1p2MKmKM0Vgud6QmmVbmp7AlE8xto+rGztV1J3VLowy39Oerai7R9v4CugJdT8ZtPyazIxrxDIb7Ln+opjqaJSlPJXdxSMUCCh1+WaBE1OjV2pv3qBTn6+vk8w+PxzbrdatXw7TGic6kGP2MfeGwKjWZMx3LsNS6fQxty+FfwI0sKSw6jP3WZwdqD/MzWwYzq6xZu8XnhM8DTfGZvpIumZ/hzpU7fkdtMmsJAkdhe27I1U2/E9ZBZL9DTthrtl4Fl4AmkBRMuVI+fmxgxCRNlwS4vsKL4n7HtxPEopqctANXfAf28AcxhuJ9iGpgwimwYT93xihXKuCRnEqcJ4ZEBKHAsCd27kHeDfmcWB2IZLHeZ4AvRKDJuCj5DAZNyx2Qvva1jeLTkoHnBVar+3ESjQvhaPgfQfGED24dZayaPLUpt+Ksz9fdDj9EADRFuyZpkrvZFG4bBKtEzgVInZ5I8g5DGN3r+diiXryp7RjD1C/CVTPRWLmbdTP42V5n0I66WpxZsyPTkAX1QyQacGkBPfGWkwSdC9QjxDB5fyoVMRGoR1YoUxt05rE71FjquKsGLf8I/xqunFvtPIqpg2U8FBBJmZgDqauACuxe4aZmBKBhtqOj5K9bDWnWAxHI1JK4sbcW6ASTzRuGGSgy49z8RzATVu7DopfMKxPoJnp+ix5uXZdwXxSWbBmmltpdsORNqYWbIqs37JUPeOxJXDfcI9YIva+Lmde+7AHZsdNWiGXUWYBFS3EudxMIhMR9k5uaIg4iFgqQltFOD2H0ZNK7Ke4IH1Aet+leXXTkHAxRkQRhppp/Yo0+clPKyLNBhWlTkQqtEhyymTIETfQGSpY2VPK5KEaEXixXweuIH3bRKpJdXa9d+VPGw32GIki9D8hJ20ZcTErRj9thj/zzEK1m2gyc6y0ePH02Rvcti1ydEgqhJDttr6Uah31py7jDA+gJ3fh/sfoqOQrAPWRsQPa2VBFIPZG8mVufTj8u65fUsV+IXaB7acCJ83i7ZPYOjFG8rSwpnAW3x3/WnU9ZVd0MXJNfXxJiRupWnLA/SZ3P+6JMUGKYT6RaZQDRLiltJeOPk4kFc3TQa+ckFg4WneupLZzZEcMg4PN8Bv1NOlihoiQKtMjvkV3I9DSXj7Y++nz7ijz42BTOMDiJ3iHl+UolNK1JQIlVb8vCXVLOCHHYPqiG0O0gS7N3c23H3T9wkIHaljrNYiQJHu+SCKE/dGQ+LJws7DLR+9sHb9np1a3bAm+e1FFwxmsyIQOUr+P8S01oDkswzQN84tk9Hs70UqH0s1EFWOv4xjMnzOhb0xA9rOuvLUldkJVmG0U95UCgYt8UQQHAe86iIrCKXpJi7Lzw/LZTdl+g6nhwFPUfnDAiVLH2WI0cs/f2DE1v2/7NawrquPlVVPCUYjZuiNMBBGTQ1pSQzA5DBBRNPDZVOi/2Z4Ud1MW64nEzyZIYROkqUizFeSNyRbHrCVBn+9BcEPlgK2Ovw7cjLQPXL4TWGrHkO2+YeyPWGE59d8vAgM0ecEJldfC1g0DVM2R5KuPCFoTHfavmwJJZU0WDZxUMea/wLeuAUZx49aR7WZjihL88qa1MOzCqRK13SBGPnwbtmwl5zIORaN9pfH9P3y0miq5uefF25uQIz15rBKg3tKyw01IUj271MVkv0VYzGQ3TBRHt/fpcVPc4H8tahZHmu2UT4bTInrKQ6oeVHPMXxTh1DIAdGD/uwo6kkXnSPhaoCCZq+CnTb/NGeLDCtNvGntSkK00E+H+HCvpRrZvM+LKBJUkmpD4OxNjOVAyCK/c66YSQydwgj5qaSIfJ1HXyOhQmy7N8XoleW6rrF9dFqhs1mNGO/a9aJbP/SMl2I8lYG5Ut2xVa32AlrYZb5gEkpdJzB6T/SJu/sUzxL91S6ECX2a2+5eax6wdU9iDJMrkefOnNqy4KHOe5MyYHo8MO183GNFnOAOcL+W3QdEKuXsEoYqrJapZRQwPRa/kEEXXEAVbu7nILlTN6ssR6XjJ9zQrdDsRcgDJZP58jXl5gHLPXEZ8OgqLuE/f9LQ8urRqdH+cPh8cqC99CD8v4M32yc1qeuLIOQdADm2O7AKdbsLtzSKlMVKlPhiMxpu2e/E1OIVUKz6s9M8pVtRIF6zDLycXyubeNOCipA9rAYbcsgeR3WzRWKKNFA0Tj8Wpn8klTl4sZoFEA2vqkkSVyi1Yvy9ahokicWluGORQRu81ia5zMbKReFV9XvuEOAI1HJRIDHQ0s64DRkOmTWgF9MszPUX8/5h2QfR4hwD9MzBkEUoiB8ZswcnMmk+PrJXmLNM8kFsXyqpNSOMdLF1BY2y8qqK0TnzHGXZSW8q3el1Q2Fnrsx8NmNElqDdQVSu7XyBwoE778Ciyf3AUcENw/ld0sl9ajgXDAm5g77pVfK/ddxuhcfhFBX+ur2SrjlKvFw5GQDmic6CHHIn1AxSzHmLFMwkP8+csgv5sw3pGyxzHU8VZYGvs7R74lP3uC3dkQQR94/2COjiThcrmIwCEu8jMnxt1oXijTS3uY+GOF55LmG4+mKf7nW7RXYbvbRR5AxSgf0zxDwK3IHSm+uN0oQd0+lPMbPnh+lsVbqWHrE5YYw/pyRu9MoULbnlLizGEn9kAGyYCOL6KbTVRV2qepU8ppzP8bWpqXMvqWmdTh4/Dd/eC/uAjQHOd6fZlFZYHIzvK46cxRTo4OJ3Lrr0agKCN0+iyEu7LkqKJpPFwUQkG9GaJJwZtWTZu7lE7hZvh2HQV5a2cb+Ll8qOwqeSty/b+woBi4S3Lw1Eu6ix6ZjWYYwykf2jj3H2LCmo35dYjcXIAgWPXhHap+VzqZ1zIBmqyQEk370bGYXKLnabY3eRXdnRo3+XXe2OhxJZ4g+3iMAzclvPsV5CeR0gX/+fx5CQRxt/G6mqZyrGMeEpJnxj9ZsUOVuBUtGYWPjhGf9oe2YUMiOkE5+kK4U8TJXUqrcL0Q6CdOnjNRZ8zQbI2aNfM7dqXV5dEVgoTs34njIapF0YajtsIBuolb1i1iv7qze+G/FUggZIRBAyn41NXKXD02Uiu3sVOjalRaBDkLYtsHtPErWJ7T6W8UmWDC+15Ihr9pMPdDjgQPlUnKvI97LQ+vAPnUxMF1tL3EmLos2yIXdPZias6c6VgB/aucDVT08njJvO1P3kBqPldzi7tWjT/Dq6SFRmRwzZmi6T83hZBcHmsnRNM1ukU005fw7B+ur/04nxj+DIepsudmAmrET2u8MYo1u4zvNXC0ZU+r9PmilaE+D8vnMJkAw14TTFNI000RZj9NA90TORRwBwt+zOOxF6B1ugNPII1za/K6A2oxiVp/TJ/KlcJfVQ+oH2lE3JdeDX93nnmiOAWlbwQHBGSmoAwNkOS8FE8OGvZIP5Uf9InqgAno38ra6M06xWFD1u5cwLKFqk5s8z55b6vCm0HJT+F2f5sjLfaHuHtJQ/nE0o1UCyfUPN6/FqySKdhi226K0p0sBhX1FdeYVzZnX63xjylaw62amCz15fMK3RdKaPwDUmlsd/+eXnEQT3lP61NYdBBJY/ZLzfFxTOINFyiTje1DCf/GTlRLyUOl3QJZU3zeCszMrwC7VdzhNn0n4LqpV17N/m3DpXzTk8haZUKoP68PBwLAPxCQEx4wMsN9dJUy0+KuN9HQEuL+GEnR1PdE+KcNAqPCUwH4eP+YygPbljLLp/2pUyxovz59OqA1VucVuV8r+DP6fnjR3PtB1+bjeBlZDrQdUqvFjcC3RgidCHvI+Ba9R1eVl+EWAGcF2ajJbx08aOGA7ehHA/IFUcQFnG16hDcTYwxY1BAyhKLAbQh18UP2Tb6IdFQC1jDvCvgsNu1R2CBCp305DDeX24p87243lV5x0O/V0NpE5xWZG/FKjCTw2dmx1igBUWE9wCFzLzDVBBbAT9D6bQITbsyiP7O0VjhVMeTSHgKwhVVf21pUTebOtVPMGWJe4ki1QqRx3187YUovMMlReZ39/K7AYzLGbxsdZtyvubdpS5SjA9LL3LP7/wrjTXgx+7CcC1FPTScpIR+L96RIjnmMFnHax/MCtREm63sXVkDOy4MhY+/tLrBfqPew+Dm6oeoTq1iSV8re/hc0RsT4u1FM7IMdV9KGalt51Sv32yYuD+6C3skhWTmOcDfjvOWOVwpQoaEnlb2LAH35c5+gjVMcTcfZN2hqhaAupNLM3Lnm7VX8bh7sdVNNGUQG6yaPbOHku8sNA4Z2swxQuGZn+aOFaFGw6GV5AqPG8o5XGe39QkIvCr/GHP84hso06Si6eVgtIryvoKXIE2z4/45ABORw+bsHiiLN7AQF/SuqDuJLK0By5wjqLBPEISuHiDqaDV15K7n8Mtgx0PhB4lpzJxlm5hByqeQzUINWUfIMQUBys9cg9qZ26aD44lirOZ7fnRaXCVy2VH2qdvpiZY5ZDBsd20MGsUmTfjTlTt1yD4wRLUdj2P5N92b1Z9/QrB1O82PYiN5O1k9a9OItZx9BYnoNk8jEnNnkRCrNRLiF0uQ6qFA6rPZI7vX4WdOPIcIIqzauakSdGXRvlQmWtJRysV5zeUtYDAZmP/Qs27iPnIZP/vQaGxVvKojcY2T6BXjXjyRBYsT+OcIm/lyR225XwCZBrCqE4l8pO/+iwpsOYgEJLUvwjK1DDmDK7OUj7rLIsJlZWOytQuIVbpBTZtz9J7Y3boeVqwRctZPSMTQvw6evn7LdBo1cFmtgrmC3UFg1+57oH0udzdH+sVdniU4FaFDKcAozOeDOTmPVY81TC0NfQGBg4xmBAEfQW/fakWsdNWJ61b0vL41ywuiAdr/lOJgTc7WqIc9nkGUMeYkurwxqF+2RveOtcqh+fAn1C8Fe6gXaYfgqiSDlLilfEu3j7jRnnh6y/CkJPfLCS1KKUntl5ira/vXeY8NSCFrVMlmBbA+aF2TKjS8bJEhs7+zXoyqwYvfm+Dl8egOYu3cFpAErDD5iJBSGYQa1JU3YdNuwpYo/qVkmpQ+HRxJhwTWG60UByq8rod7OWGCtaJGQfXeHDZD+AYW2J6WM4UHAXpVP5ezsaAA0SpnHfOyyvHO0ZxlHs2SCNjxLLIs6MYonfTRuedHVjwP4MkHAe01q/153g/7tSnDlPMUoBP8KoYQJvwoT2wioA1QMbeVaGpHqaUvzIgIhRzA3krEorcsuPCrglE3Fav9hJLlE/6znM0iZ1xMtjgxDDIjEAHw5MT5IfTR06U1WoeUVLUzaV23J7XFpoJeDCRzpvpCPJfHgIgkoXZW8AzPS3pIkcskWGIeRMSJeAgPLPCIIUG6/xD4TFjgy1zzbLFny5+4D/Thre6ecytq+NXmd3i4roySH0V7roYxCu7P2elCUYX96B8Ol+ARYvZt0yuz/VzjbR1kF4XYkqoeYPr4RYnMKBWl0+JmKt/OsBYlFkvIngXzRQutzJub2NwPEZL/1VxJPMh6/ORqdkStXWeLx8myWHRfzCO9LctB5ASwkZOFb1L3hwRofeyh2aG1HC5HKBBAFvbDFvRMj4e6p6TalrFO7ypXEk6zklFCl5tq6Ggfk0vRDJh7nuDTWZUH+rbfDDD7u4qiA+Mw0FH4hLHDzD5h35s/OSP725DzJlPAyg1KYBWL9fQU/7USMji5tWMerSXaWrXBqVRsBHNZlJA5ZivCc//VbYYPqZ0aixX/BH+GC72u5gX5bJRQikCQOuRRggc64ESbIf/CbjYrcw+T3ZiYJyohOjrt/2V6dPvJrRYVHI2zz0hiKMA6uDAi+oXAQd+A1SSvtmecA578RSwIrFIABWPPa1FstAShWBOf1nhUDB3VPlVktbjThB4pU/1wB0uJw2J7K48Gos+ojbMSGkht3+bwAxHQ9rbsx/R0vEGV6mjHzimcXJikE90Ppan7RExyR+VdBZ3jfWsS5F0SjA0wNPE+N/4I593V3igg6QpN7Jh0qCU5TR2++YijVy2y+7UMqTvTj+Z60RkQ74VT7c90mnLJq5GVMgJgxvVa6jjEK2Hx2FzYvxp5fbREbZ5LFdlo9OOKg63sl61plB7f+2gc8mXhJ50ZEzGYk6tw9M25DKdsTic6eqoIIFnXJB52mURxpcSKQrT4hQXPFBBkhwLnj7/eGy6JdSD1xtNgO6DAs7cuesz4EZxrWNcNyc19vdE6rl7n1QDvdGGYusBKb4WJl1YECjw5Ggyrw3OQL6l1Nr8LTzMk6x21nri1ejyirzJSOY/KB8qRaxmn0SDg0QsLLj87xk2xA12ST4/Ieow+b14S8Ivkq7/ljs2w3O3uw+3GyxtjDfkqtUPnqYCuKKob1/zNVUVO4p13Ek6Tq++riLmEu/M2ick+TYSWAeTZjCnDwEA46SfqL1m5jq9xaRGLrzAyv/Gn5y2WnpRNU75uZv26EXfZndQ8zm8e9rC1y4dqBepW4MNDeIjVaqf/nxl0TgOUb0/As3mhJu6YFqxoPCPARQ/liM9JPA6wOqzCCh6nZWIq/pg5OykJW8DC51k+bHadBfKKikRtpg+tFEEMjIVrwanX3kCepwd3pHvzWMJSleUPjSqK06k7oEuvzzSnO0aGw4FoJto9RTdFCD8rTXN4gxZ1e5gPfvB1o2P8iD+KCEdDoswFWvtQEfacsVJAXapszFhPs+aIxGJhdyn5Dj8YAgfJM96GUN4juPA0eV+CGPAhzNPe4uPJZXWEcZOLpF8IDh4FkopIOl11cfsjgp4qqwSVI3Z2LEycRljgqSsszztYvXEJhgnhOlyH4W/1UjXC8MPuiqfI/53w2npQMrnDDxlV9kN0Qbi9xmHTFbBVGk7YiHJwCRRvhKaD1OafOrQqbeQXRUk6X7woIitlkcYfYsHzccTuSXcWTlKKhf1JTxN/COQcPu8DKMrsfxvee0fYeowSQbRNKCmIm8Kg6paQ3isKgR9JL5EAeXDQL+Aml3Bqo545IpuBAS4lXLYO69SVdOm7kzhxKr3xp8OlgwzgWOOP2MHn8tZCao41Qwr8Sl40EI4jSIgkVzjQMNDSo9305jRsXERcuuNulVAVPMoqhy9kpRrTVYQ5fRoWvGJV0t/GZZU56xsREJgx3sc5gEY3XX3JANODASs0DdIq4q8q5nToCZoLPg14WsYrrrsSi8TdUDCOaePOvrz431SsswuQRmD6qlzrD700/a9YloOoLsYAWtjqyepdi6sRCh3Fc6MnI+77klVOeW1Btff5MO9GVlfAl1T9tWo3e65GOwYaapIBz1izKHN9mhE9p4265GUKchGN6Maz2TOm/D9EZI5jTdzLA4kxSuCIQpnMWCDi5T+BPL/TRPGphfgIW4SsIBsnTZnq60uI2JNwYkuT3zpZYuUhc43QdDD69JY+dPr6fa9JBRLNeEreNO/4ZV7Ot3KULYGcMrje+gGOcScl40XihFSpl3zUdTs0i1Y637R6DkrLhXrhquz3aXOl2rap28vudxut5KlS1oo3x/DLHQTPQ+gWTDacvaWbQoPN2hxoxVO4dBHVc9fIr1JGm52CLrwP/wD56eb4RQHet6I5bWqA8QDZn1wfWMmKUbrqceE5tSodYdQllfZmvnzSsLrQ5M4yYc7R2Y+cKib0hcUcA78EKJ/i2wu8W1FbQhXQEXMyvBCuW+ZOtFLg9zqCZHowFpUyRUYBpvEp43iuLni+NVLx18ups17ZPH7PzVTiITQrv/ZIrzCOQLcjwM3HmY91Q+lhDTEN8/2tB9GEV+3/IIR5RDRFEkMnXjwhLsj3+HGimYERcViw9cf+hCE8qg6zJLGMRFP85COVyneYnn6tr/ZTolNXj0sM9jpnAA1DldqIm2D5PMokGPkYW8qCsiNiOZ+9uWZGZ04PECRmAejofl1cIyBLf67bxOcOa22dCg6ZloV4DHPF2dZBPWK/y5LKP8Lj5131zawvcXWkS58cWHaBi9/Ha5DIs6pOK6wz117XWoL9eQK0Pa+5RTTCYquZrGxGK6TaONsIKnqSFKo2qpMZE3rYDcOXTVvPa0pyFOtBOSFHhCygkISKpnaa3yYKFr8XBSVadxUZLjjodK1HmyrcV11sKGQ5kLVrBQNeujfR137I2wHH3Ka/qFY/PkIpBFK5hS+FPedt5hkFItf2cqqmQg1r++gywM8ywahNlIFt9J8B+CsxGZzN8cW7YBtttFRHGQIfDgV6822z8pfGu5EsP8TBHVn6xHqI6UKhwtZBXHQGDq2TSp7X0f9snbyVyNu9PDSnpZXo1ylJGOcg0kxmKF4JU7Is68NCaFXbYgqoGtpnLJDSTFRhGWCg003/8ElrpBfxWU+PPCDncfa2KvaobNbZ80gj5+f4ndCu2sEAb6B1DVOwJkRIifw0fxyyJ2u9e/CQH90brKJ+h3O/2AIaJLoaD+/MAAQDu2WM3faCZHNib48Xor3cgaonWgItmXtzEBYaJVDbwxF7Eurn0ad5gNZnMxSHgX2L8FNnm2PTfiD13X5aF+BO2/tY7Vz1fwteoM1Qgw8NfHKU3+Qir7vJcSUjJXnak3gU3tADv8/Ev8K8WPtS3puXLciDlEsGZdopx4SwkF7QWs66Tvi0Y5DXxi5IUswQl0s4ExHDQ18Ap5maH5FAC/fghKugp1XMxd+gRuwcNrbWxOFb/bXik/1V+5XxuqPediNqjI5h4veBg9A1Gg4q3bJdqr+xbXnvOKpTn/7FEs2WzBS4DFxvJs0Yz5xWQ09DeTqS7NGc0Go8GqYKh0ChSa8ebVwEVwjSp+iioTTn1MINcy4asHPsYQagS7Mk2BIv1hWIy1pxp8nZf1op6MDwSFhqziSmyHonQdsFiDCsMcyNFBzRsQJ2TWWyNkAQCXbjGW1cpQvYZBLAvRj9SslIE6VGiLe6A6rqk9KLtIdjn1BAoAypR7bFVSdw3cPKhp81IHBBphalqi7Tp3PR1VAdU8C3A0tE9vJwhAnA2SsI2XCmhGMIaP2yoX4jYSd8QHO6Wy29/ZCvyWoLtJ3zE4VZ8zaqNK/HEah0E8eXk7u4C1CM8pGAYjlMPHqzJruZxqdt+LCpNB4YyrpW0cMaLirn5aX3Tw6rsCneQcjQEQ7mUK1+LEz/QGorMAEyLDahVI7JwXRuU1FKxyLD5h5AatEVZ0jZhUJr7ZmEDZYBxJ5k99ufGoOXwpZSBNLe03bPaK7ksOO/5zh7lGspUESI8KcSOlCGEWo2ri/AEMkDFgyR7vID/x5CBFxMhb/5cJSzko7RN5PBYljFrDZCgRYZXdvVs8l8W0YBuonO91cvm4boy1JVnBmYUPRC6NKGNuzHJ8CQlS4HuwEHKAX/Ku71TEO0sBo0yTUOCfaOR69Eq43hMkax/6kK3kbsZbkkI+KW/gQ8KFw1xChLRL/4CSzqBwwzgxuhYTjA7op8jGQdVeKl9fmGJaX8jfMbxREoXB/d9bZqAI8gAAzlVaa51SAwejNevtWF+0w6us8nruTKt4Gud90OX06zTKRayvKOoaCmjwvi5kS8tx9t6buispEmFmw/qvd9EaJtssjVtOvpmfEj/KULDET68Ti5AoLuQpidkjCMpxBTqXCSMDtm4yTpInTOc9bYyw33OxGwkwNMMXkb5K7qWX3nyDFDlbyBrDuK0kFlMQO/wnC347e+sZyzvMZd//ukf1tEqwz46JVWV7mVV1Oee1C5gMD0GQpcJko5FbNXYiI7xidHRVMkYRJ7vm0bYiAPCP1V8fPCNZ6w5g5n2d6/05bT17TAbvjuw9FJ0o7ui5ejQBFI4rNF54qSCKHKp+ks2dUcY/R13+QT3iWZuL2QAkmV+UUzSOvtJhIA2V48a3GDm7er4PU8bltAtL3n5kt1NgdWmWS2zsW09Bh76rOruSVSiXRZjCst2nFE3tL/tq4etxYG8M7hqjx7Yh9z8PQ1xvQZcnDF7KvaxLgCaj04xEdet2mQfAitNa2dtKsG5nYKCrgauB/s2ZmQ3ozH/7sRg7sk2u/Xbn1w/dxQmZ1h1zx95wxbWJYgnGOJT4DJDjiCPOgf1jju80PTG1pZblysGO4Bn+wa78P9s/skwtzldX0VISNNbs6c1HXHLqSRHetBHqDFi7BGE6lHcMYu8D3rRPMM38hd3Z7VP7hGeCbYFghV7X5ZXWVXlFO+ed0Qsf+K9fEKFSK+N17bT9uLom3YoQWR01aeTERgXmxHQtUxH4NMLB2M+lSdqRUYBsSALZu/jqetHTi8qK7eKdiHbRrW+txUTi48G9hxI3S1iUoVB9ddbTcNNEh7gWxi2PzYmu0BhEEKRff+Cwl24lG8vTIioyivLr4ow/CXyQqH3BSilkXqGid7yjgI2bOEG45DKb/bDfvBfBy65zmePz1x8g7CjozaZuSa4x4vv4B1rkjaFeidNZvZTQn1PLqiPhgk20BkNqc/rOZUIL7vqMXsw+F5ElLkk1o88CZJUyZ8Eq1Ysap5xgfDrykCW7ZMuCglsEX9H68J4B+K+odZupuXONkkpTBEaxRcpL4lVqanjysX489evaM9cm6uBo6wmfDB8h81m0diOnSK8NBrNJmCeJGy+WROBO8i9dUnefbjJPooK1E9S4GgZjW1T9VMsFpncy39+AgZg9TEVs5LdCDWLrRl5xBWdfWDUAe3RqxP4afC/dX7LcrAiEAFs5hxt/ssOUMt0TmZrqsd+OrSfMtbnEkh6hn/3/IJHC2G+MqPeLiG+97iMq0nvtdm5lJWFJ1gIxKa5ReY/9Q6ZSvn3H1A8AHXBg/bScW9M0qXyKfvqFrwSJgiVXNdzLz+1INUg/LAqJD9fNz9lmudnp3GBHfurQC/81FTHas7hDg8rDl4DPDFdW01B1YIM/3rL8UDbpjeyeF9DfdY1bW9wvP0jUq85tgoMc5rCeuEBLxKDe/qHGnqa6ijnNgGFYMhyd3v0Vpso7vkElN97NRm6YEnSq4Z7GWPiHbBbk83LDpX17Pbrqpzw8LcEULtrMq4agbaGxtI3mLN+LnUXcEMnNtKKPPcScokNAhGcnTvJa73HVEowhY9gH7ioiV6ypXOxrccegl4Xbti835YMCKod84xVENPT+2nOy3e8+cfyWdccA8o1QFi5VXHppzicysfSLXz1ZsjeJAQNo2B2HOBslIQKKYeAQQcuEj2pWiraJS2WlNATEWQIOa3budhmYkOY1Xk11LAovq9j3joS0i5/GzK7eanbBar9EOfjOVY8Jl6wKm4fQQWEqpQ2KFkiWUy4iAUz9g188QUStW7rfe62YrmZFryYEmyxxEb2fYF+leHMlm1f4wAzexpUvaDM3YhSQ8osh/rTv26qgrcr6eruMDh7znqsLkg21QjM4N3nZb6EZXcteL152JRE3oMX5LOFvx5pXDevSJ6CWHmkxEglWoE5n/eujp/1RMcI+cadHjkZBdNJyYE1MgARzEK9PZnCiqOFjKJ/WxavOmZlJRoLzNBM+CD+hbjgQVnYcIefAqIDRrqvCleK5ELVNFGRly0MgGJyujUU/GZLJferG47BJ7LOw9coi4Gh3atAys0hokPw5wdDQetn6jGYAiFtIysW8rFTY5gDrr5vFW+UGsyGpg6wqRe6EBmsMXs0aNIaTe+E6ctwjt/P5crgBZ09PFoEBWfl7dOxYN8qEi2o5v18VWp61vFAZy+0ArHQ8tSGzQL72EK4KewIgmF6dme/mjX4yWFBbAHxe9p+e5uW639oTGI4xxkYf/xtgzoj9JCyB38v8ET3wreR7qji1wUEQ6lLa7OkoG+8OcSKCM5ZCaM+eVIBEqizDXDbsITyenl+wjY/23KKtnoNBKlF2EsBXuf4XbtPDqKDnen4sWb0hDOFERAbVxcdJKis+2fiMSPpbDcO/vt55Oi1uYhH2irBXWU5gWoHtVMg9wxw1SlC69oVvtuHAZgxvu8X7BMAlktUDHiY2/B0spFMx4iJpgM7AXXNK2yYum1NzUCuodC+vTZoOIEPJIqc2gLi0m8D2aX959nWTfxlOxf6OHeI41f97C00y3m0lfqCIhuq4g4wlakoY8W+KWk7u3UTbWU5Dq4RoqZbMo5dU3S838pIIdZQ0opgQxuk8vAdR1s4hH5znl/xDFhj9jXri6+ppZnE5h1H3ayNUiMwi/mHJN7ji8gfkBHOUHHDf2G8/OBN3huIQKvNh4BafL+rbVbSPmIcoyk8u4DIkHC39G4eHp/JuKYB+5QvyNGHAgrCCpO4mJh6I+/cYUxv0RQjZ7xKFby6/J07MLCm1vCYTTDS1KRXQcTGjrpO/MdpiaqdJioV36aMFTGH3I3FsY+Bsb+oEjyD46Xx+wf09nej0UnfvT7CDlS7GMQ0XPImabsIB6GccfRJRIArtf26nUGta01Z8V4p9+z2iCThETxi4FCMmsLcmui4k1bJ1HjKkAeKKrBKLSjiyKMrDxk0WxyUtB88vjOm4VNMmM0sjPBNr1UQE5fCeQuQlGzIYKRtiKd8IcYhPafWjrWJAeZM1z/fC0I8xwXi7ngBUBhrlGxg8lpoJYAdga/brtUa+N4NT3OcZ657OEmKqSM8ph/3a2IU1cNlvDtdTPlBHSFvinlvAsIVa0vrDCp1PMZctHKOyFHQlzCfPRwn++QAqMwKH1K+mg62epURuiQZ4XWiHXIme4zPTomNYL9TOc6WTaYXvgYES9Ro2ZDXGbucWO+Lek2l1TMfsZKkhkAMg/6mnCtiSn5ybQ6PMrK86oZ7ksD817IWyJ8LMVPi5fH/4yfadAUfERWWPV4e+kvc3wYrICkPNnnQF+6gVsNkGwzgBnE5+MtlxLcKykT+JTEZfo4RtdZIROuhrYKmSz+64b2Hkhdf94NnCYkWBZjMDyt1+0G1BCfyM6jiNwtDQ0wgDeH2s940VR96mn69L2KeUu7XHkDe93/sE4+U6U/lV9JvyAN1AtPfiDrqBdq5VOTyoqAr8rVP+vKnVhD6vutnggcNAgaYgDCQLSByQDzPlp19PcEWGXElG+K8Q1tsT0csFQUxtZF7xp19PKtQdcyWdi2c4j3OtAVezaWtqCBtedhpKP85gFqQElpAw6QwfBDoIocH4GrlvyTzcqSJ9DcmHYRb66qrOk71xmeyPM1R9IY1aiJmmilZoBLAk3daWy47yFS332hPzY5FAFkTcZ21EuTAFlE1f8+b1iZe2keSkdVc12kXFXrrHzo3x2CoiofiRaZy4mTH29kvh7F8CdqyPytO+M2UO9byclcp5uxE++IMrILLCCWniM7J7lnpqo61ngaFD3K+pRpF2ux37HeUFSHnlhZ5mRUlTSn4GJZ5wuHWWNEnGJ2L2WOfPvc3TS8z4/P2ealdUtnWnEYjk4a1jYhI5Uf/DOPbvrkvWqVccgSOc/I/iOwGVJsnLXItvB9CXm5hmSp+raQsBxQK/mg3teEQVJIgXekqjJlKvbieAoovufXiNJIiVS+mYC0DMkKqN3vJF+wQqJY2fzhLf028ORCd9HAMMMDsXwE/bx4o203aySR+O8wl/aFKOTMdzDbyicQscRot7yZRBDi7LQW1JBCd1tsQNZv2vpgSTMSl/5dDOSk6F4Eo/5WETQgg1166/yp/xPmGEdZXmPrq+TjHs3GAADC1LIfR1CUIEyD4u2Nn4O0fWMJq4lLg3tYqEo2h55W+SLm9OB8BLao6C1nmtGfka+i4HtKRmjufNoFH315P3b6SyZl+U3bnyJcZKgP5bQO4Z9M8/0pKHm7OwgExB3RsiInnu+SK8wn+FavUYjdDhJm72afxUGnRmDP7hApN3Tui4amBUC29F4DK32wTHTqiNwg4oeqLcWvqqbspfYwP7cqmScNSGZcWj5q/CsQLTNoOdnDDjoIq+Ad5YuA+KsxbryWQk1bXS51dhC/FH/FzzLeRLfNignsvOQ06kCj7AGwPZYAWNXQfYkTPQxKxtPge+XhmzhUGHKoLTvQELmaYeTpl6z9VztER3VpCrVUo+PKEyfCLGsJf8LljJGDn1QkjfH+ecILZWeVW8Vk12bEUnKP7CLlAV4LLjaZCjKoR8MFscBmd51Ez1lBVV7+XNTx31uo3y15u8fFOP8jAJLF2J58NMYQLgem4GR5eSLbzPnCo+DCyNMaFFPZ6QowJPetAMo5w7DLs97l3x9g5ogUI7+EFptOP1EFXwBG+E7Mmv0s6Y6EDCDpv339CPDRz8XNh2qYDAdfZy4pz1BhWlB6awe+CWQtHoLMHW3vC4u08q0mJ6050JKKImg1QS1Wse/914N8fWlub9WM7Te5c+McGVUOoC1oStMBDd+K53EjybXXbWa6TpwmFGhRZzSsu+tHpHX5Qxl3VI/UbPfVpyRaYDUMsJfO+zLQP2rbjKGIR+zgDA7I9OPLEDtHkKPNOvWiX7+vPoXieJ0Y5WUkboyHrw+E1V/YjK18PbQB9mfqRVZHP/mz5BSSca4Zwcs/ylGQfWw2HhnNAmsw2fQpV8DOD4kR3/7O9+u86vqiRE4s9vwasR+woQPrD5U00tU1EvqKEoGce7bn44danMQ2bYgOpiI/87bxBjT+ssF0BXUDxfpW+n8mZUm1YUEWsibPX9p/cm3t8as58/3Faff65wFMRm3ur086kvdIxCtacoP9HfLkAzRnzWI8L01X0oZ6wr0wjPKDLPA941ainxOzX/skqkpOa2wtU6Q8FW2y5LvhKqaPc691CiQOOBQLDW1VNAv7KC6HgLqqIDDOqBxzNbtgr5pEM80oALu4jTmGkURp/QPbe1bRRntqWf2xMPu7wF1sAJKktA5o+OVYkb2YV3Lcod3WrW1DBSeToWntT/3v6RUjKH48yEz4lBlKuHWglB/fOCHZW1OHmSGjbEch15H/Z5USL9yAFqeqT7DQT2ECPwftb0iPBR2Y89vYPceDAPcI+86/EsFQEXddFXBf4zhTrP3VKGivlJlEmAgbvh86sgEGSprRNA1slp/GGCuLzjdP+V/7Ht+IUmqsKkZaWTQfydO2N5atsRc4otAU5lhU77GpgE78UsfxoOQQ1yb7CufPbVyYHIKgELEaA6d4J6Bz3cNiiVEQNTo95ZF4QeIYTfcvjqqB+DlDORJx87s/+5F7zX+sxqP3L+dCZfVQd6oyEX7B3fa6mNOYH+v5GcYUUtQYcFT+eaoBqa32ZmYsPNEsByR/OUcoEhATeLZqzDXokafe8+ppEjvYLJEKuemZNBL08dDbJfY1y9nPwUPTvb5bvWiirlVctD3F7GNNjQv3LX9ozrZ+CTdMjbXz9apMMrKoae0f2BLOX6dCK410sx8E4YipNnKpuXNOP/UAUsinEz+DLuXYyYsS/38YJxupfmV5gPZhSOoRDsos4WfJAovyoMO9kJZBSXsT4/KGRayKU/i0N8IAbG8Oqqf69iHxEbnIC6fjOxoqFmOX2+YFRzMVzK7Uz8z1qzHnLbcM3RqRH1OkDj3mwsIXBntRK6biOUKuChTiK3agO9ECanXGsBV1ZGU1hBd6QYBC6quHqNeZw6Jd8BOV/qiwOiffZskl4t2b7jJU/tiIgSgpkyQHTP1lsH5Lw73ScCsXydlkhv4QVL2gdJZyMAAUAKHgrE5eYhNMzbeZcq+sV08jH37nNte60r+u6XtTe1SNWIDic3ylfZAbJfY1gvRjvwwJli4j0u516XxtFQbHiNwLXbMcIKlWQ2umFMJ7SxnQItOPrtSZq3kUMcNBFqYCX+CnSlQUbQ67MJjLaEfCv9MqP8AklQRM8ZwlJ5leFOrH6p6Y8TtzW4vriw50q9xoyUT3VBcF19uceT+sCBrRr/+wnZDeqlG7ayX1LIqSdkc/+gSGUL4EFnC1hFMgHFqSlGQoDJ4galbcBBkaf/8WllIQm/D1Y/4uV0gZ2v1IFj4e2hJvgB7IT13Gjg33uVv+mZ/oPiZWKYz4LCnuEbdiKOTOvzP4jBU+fzIXYm+c3KF6aseqrsKX+VIzhfkoZ6b37VLJqKLA8WKw0dFjLE9PePN1xfp48yDM1XCR8xSCkNaba33aN968bQNnsKvXDkZTtq2VhaJDCbegsG1BwhP2nrZTLjCF68dN7KEBnJNXzOgSd1QR7Z0cMo2kc0nJCAHe6OW8LN6UEf3HV+wkMpQ9cCnGQIuVbl2ZBaBmc6+vKRvGUZouXF2jB/ROG0XLxLTMyUNk3ZPatXtcPsrMggPx8EG44xCnoq+RLhUuV/lpsiO8pMP3dEnXAy0HjUtmd4eYadKAUQgBtyrdwuBn2F5FloYTmmGMjIS5+etH5iblXFeXqeFc24fGN2FDiyRLMO81q0fBM9D6WPIbjeKXGIpX/K6SI+h4p527jg5mGIdFeg/8pS5wEcD/W5Yvt+q9UyynC8e9L29G6EhwSoOUpbKeFAV6DuwnQLQsugzD+PAUpUYMWnJiInrPdWviw31X4HEUM4UbWY4e4LqhtqOP9+Zvc6T63SVtak1LM6vT4UQmDFXWDjjqVca9r4mwIs2SYVJ/K/I8cIfKZKKUO2632c1/ZWRVQsqJP5V9GCpiT7D5HOuts//EFuvkuuDukZQxfSqmK9TfBZcsCpegUCXrWryY8i11GDeLYHYi0YHdq0/gRFIr5mbmD4LlwuqQShADp3Ny91uDWmGRFbIGQlAitGCosiYYcjRp4FAcFq5Em+ca/jWy9WR2NyTWl4d2BPeNMRatqVF2BMNWwXLsm9XPUTDwIyx3tYtikobeN3GpLOLNLYqogFDzkBOA3kv12I4cguuKICAxu9S0okHu8WDk5TBubeXLPUXbPbsY7cnEHv4MxUaQ8YFf/tdmR7u7oaLVJd/1wSvX/L8EY7Vi6y//AD5CTbhMg1QZP0/bLTyQC5R1AsIiNcem7o6UarwPkS8s5ZWVadMClWDxyqCzv53YteiHseFcLchhUxELTpWTFzsYhlofg2DOjO29xVYV5LGu3qKPDEvG2j7Yl9sKRryyypIfWhDzW9ngPJWIwnEaBjn458JUQq9HhZ1m7ALyQg8fuBj6gUP0HXrbAYYwMF3mgHYjgvfoLoURxtSFUCn9B6dPSJmmFfLFBJ+WWp0QFs6hUc1wqp9m78hkIY7Hn+vY7X8YMfCKGdXfaaU/6GALriMpebb4exakSa/ZxXvQQfwkNL+a0nle/ZKPiintZOhcGZCkN2cC3+hNVJBCK7vDLFTKrNtrDUfdUv2v56uk1MM9C5ytP1kSM/mY9iTmLGQ6CktJKVTY5n9tGHzigq8QnebvgF6XMYdLSjErI3Jry5Xa36O1Mq8iOsRsQcXU/4C/8AatjRZwK9RRuDjMgfZYbvwdacwKaau6aL5RbPpNSVONBtKYWMgWFmO0ZPQuChkMrEevRtbltfX57qzPEvt14v+SyfmRgkU23T+E7zWZpl+q4UzAlsAF/GgHWphQRfSC0V0E3JYg75nIEiDzVsWUInF03QshDIZFEkJ7+WUD1QrerdpbL6uLuPwo2KuaGt3qt5QxlIQgCgDO91TOgxbSy4XAA4wL54AZEsBH2/qArc2yZ1pUMK2nEx+W7AIQ8o0EurU7f+KiCsMCAkB1vpbsBCC0YwUaeHEcQXe2nRMLko2IH2n8SjziD9X9j0xjlB7N20kWLDmslL0vHxxywwd4JiaCaOqMXpFiXgrd8h7abpiR5672Xu08BSArAdxtKS9UwBeHSHO4+byXXFJMLihTnBOLmjZIylpmOmcVJNX83sYSj2KO3LohRNwEsh/YhcWdFxMIzkKKVdxo9OxlcSUfXgKO8b7YMd/U4u836SLVyX9GNo8WSvWXXk892SCsQaUA7SgajGEWNuODMDac2dZo+Nl+Ew7JuOO/HhzjUam67C8N8DDwjNIswk75pw8U2ipVqLCe3J1dJaA/DIJwhmaYD6ox3okNyo777tXyu4XQm5j2o2e/lwcjqEazJFgF+xznt1zU0rSt2zAyU/NlOOPpee9qZQAZpAY3vfMcw4FWqo7MxRuOJFsMCcM2eTpTzvCERz7Xj/uaaxts93XlG104t+2TKy8rzI7HXCl4mjMcnqGbA6HQYvzV0I2ZiequOpa0O/SxkJ4CQVkTrZT/S+rI9yBP8htERgAbqpEFlTlQTwrNi0U1tpN0qJQrnq13C4B4sY870IIDw+a68k06PmA0/FIjSyu3ZSjifFhl+uhzcmBBR/A5PVQRkBCqCFuMx0Q0JIRhzSY9Zdr0ZPQuPgnsKKpDGmdlmw1iE1odNZgqNswJsblX6dHUGGvHn8laoCCob7ojvDCvqEwBF9OCv5OM7ARw8H56SP9k2irSZh2eWtbtpqHrMva1b9xcdy9s3jC2cL1XOclrDQxVQtI0Xri5nD/CrcVgz29Kxo+6r5ybWWTsaE2tNWootC9MsLOI8fxdvAO6XZThNEw7mBOm6VdpU2mUPVG4WGAfHiTsDhMzmx3hcsZM4z1JkEeY3wssjcdmJnp9H9GzztNQllzCxeU6khOY6WJsZasu07TwUhmx3uRQm6cj+g2GafD4eOWz8a1ffDtSngNm1OIV1ExJL6nGBTfraQbO1H5KiQ6bT0VrRk0YqdVooUEmTk+SbMPzDaZQVkUSaQNPLLWjyHwGjJ3SKByBjQ4e1Rj7bwdspuk6vkYQFi7c4xYhEnCcVsnkgBF717m6KYCqxx4mZZPoJnXgdqvgKi+MGqXjCuUa/ussXs/QeVo9muYQ5ibuTbj1T0C9gMkjwe37ADviEhkT7ODAk1GnLBIb/z/5PMET/U5Pq+GcpgdFP8pFhs38fVza9roX5FeZk9PSiemNlD3SCaDmY85WXZ9qD1GM9yk6LRrQLKV06NF6rnAaiUKYXppsaAhgljTUd+EmJ4qHpDto6+dh252OgA0xM36WIPB4ugHZYbbMxS3E/tVu0w+kFP9Z0v/VhDTIi49tkgsoICuwZOLpG1MxfNuMAom/hkvFwI6xFaqJLeETH0/pcIVr8Xw/OF6FhVl6GJglPOGmmnbUBzH4GcMWOXxvSGjkuM697NwwwHLyJMD2DOd+fqvzJUj0uq0co6EOaERbM/MuOw7LYZ24zvJiIOBM2cXGy3k+ILcAfQ8+yGNqQovRK8wCKoYo/7QaMdntjvznvyYGpfPCTR9+eyYBka+o8s2qeJ7qG4j8k+5XxxuNSiZVDiOJuvUXQKvHJqiJnYs5hw3qTl2r/nFuQWi9H9+Jvk0wcRHM/VNFr8Heo4BoIelufR7lTpyyBmbR3dEd4ydRKTx58XAU+0DdMnM8ibofFLR2L5jgyGtP2TvUF6Fsmt2KufW/ifAjQzhOWkHbfG8likdQhO0qPDumGGkBAQA64JaBdEW/djBt7MU+AutBUV2ouQbZvhLEJb/9OEFis3gW7KNhKO9yH/0IqMPkyYmPBqdy4P+kmzNXinyGxx7jC5QZ/wqk2clJHmkCxtw6igvOvHd6UYlYoAkM6SBs5uUKOrZsTBqtz3Jtxm4GPhnDJwXtyGnLNzXBOGFOS7B+HFOmL7dKYikJyaIx+0Y88dj6cM3ueAOyKI/U5+l7JRYczvJ6PteCvn5a0qlcLEnaKS1QGzMGqtdo20iqcdes7yjY2IBj7VS0CBq5womyFEKzHjdHnboYNXmoC+jCYAgPgULFbdm6B+5MIwzQTbwIEOqqMycmgs4QaBHL8CkSvBj6p1a69AzwyMnMfMYVtcBmbt5te9B+CR2L2pEEtu9W7pzEjhng+Ff1cudzC3PTTadZIbtFjVZE+JOriOCAf+iop+sNFhoz40OcngzGnfbOs6gQQ8XkoIxE4vVvboD35GFN1eUYWCT9Az5CxtQw6UGw2GcioxcqbVvv37sglcTaf9q4ShExzGqtIG13kQ6jpde2wP5aRO0Hs6VMf+WwoMsxsebK+te8Xr8salNCq6qQSp9NPLONyQqhrExDcBhgQkkhWnbdjPnTL1Y6x8mz1Q0bHwdiBpmvGKVBqGYV2JjcZ+keQNfFlD5SCNmUKZdRsqyCm6OMcSwdDCGL+XTU2+Ekp4roJEppGDZ6X9fGvWQM5WYjnF3ZpG3U0h16pZPuGlQFGq7QC6iMMGiZajvYJqWwDvNHqqcvx3HktWswObPXcWehKAq/K2cCKOV38k9KP59NAZx8Uf7TWNebomMalj3HwlKWS5LF+kjGhyWQ6Qkh9ONfDPHLWEzQMedBUrtAGvVieXM+hwgDkNFpUG1zkqAisw15rJpVk25wq26nJsbi4n/9GQGCivNN3dpDf1DtFrvMva3y9E6D6Dhlx4OK7QynMmuQljckOnW+O7huz/asbF7jrDBUT81ytWQweRcj/esRvWG4W5E6KfZRku5IAC4rAtltpEodUueCsN7iAJUUrwXF2NFU1GxLMGWpcr6MvhZ6qAgES8L4tMxn2BNOFGWB87bdDtfz05ey0yO+NnOlvbm+KJk5vMfCVyioB8okTyiKioaBFm3eRvSakcLTjXZcSsxf2FHPNk+hq0XknBc5xT4vJUxHQFWdMutRWdDP4MwziaaQqywTdAFKaHqdM8aRxe6KKrT925FizPCHZPatwjt4puzULH8aGVhE9C16NPH+O86fHOlvSI0iPJcgWLPwNKfDODjV5WMc2aKcDPS43drAI31RN97/cc1FwzCujZoFLvy8EzQK+kNeg2LSR2VYNTXJlf1Yycx1duPumoilMyVoQfbBEi4+LpBF2R2O1hsEJNZ/DMs2Qhg78bGh5PAtyZLmUCi8nez7kfpR1pA21jugdHnul8WfeOTMEh419iNraP3DyrA59Rq5kA171wtnuYL9h5hmahbLV+sHCeuy0nK57cxzJceehncrtdGTzDkB9cyVUKDTnCxiYR+5qBsmnt0agdzDMKFuWe+JS2wKKbAhML4/W+hAE+NT16HldLFPUSsrcUanOYzBoTW5E/HVsouPhCt0JmcfOXKVsjFbLaxA0djuyzKpAQbCGNqyoCffEcVBLioeZk6wRk/HlzHAUPtSlL/bPVGl/FABDuyT7hDUExuVNpYbmDxfmABintfAmcR2jx9ultxdJ8eKGKIw8hGr3nfvfDIfIaptLHVsSAvCXrU6E1OYN2vUO8K4L7IuwOKtK46XGhnZcFcD1pYOHhUnIyPQTxztfyYWPQPo0T2nwCMzUoCXEjMCbUq1QToyxMPVGPX4KeE9+6vYOqwdrVIIY8ZAOP3Fgia90EhEobGtepRsDqbQzixlovtA5XCPkz9/L+h8jO4dCFuEwv9LAWGZfaJmFQy8JJzoYUNuXSF9CnjmDxYrBtaLXu1aILBpehfhGYdj+ndt2uqfVs073eleNgnlFTVjJCeri48/NAiSrYv1Qzqd3A+ZrELOgoUzrPnXaahof6pk9YXgHIMzJiIvkRYCdt5VdoVa5uNCVZ1F10FAt2TAIkrjRDBinOX7jo0YYywg879J+ezheqiTEFQY9Jvvj8lOPvGHJknnDFFXcFwSa3a8sOfmDgxbWdRHT/usPr4tER4Ctjkf2noqJYa50d/2KXdPzoTjlrnkXHOlNoXHlY/PXPDxfaqan9GhKOWZpvjRkb1VsnGs87ecfTSKjszsWH9DLSxS+2bjJyIg1SwmQYsbZrXEuvbUOW3mdxcI3EXf9ax0xqN4LGvMYW0UHe3vJ57qzQfrWcUdi2BLkzaeCk3puZfrIwDlX+eS4HJ8cFDjodPyLTdVU8u6uKPZ8OUwu4UIBoTRjILkqj4CWYBq0KnIQo5TtTWDB8WNgZ/KWOBWLLfxYALi5BIMzdB2yonI57tehMLI87y0pR/Hf5kKpct7zkiuDIhLIATHCkoj/ApHKrPQQR1b7wHoWoIWN1HOk1QDb4EjKV/VeLKHzmnbg4X2nOKvhRQY6b69lx545bIlYuK4oM5VibExwjU4dapmDwybpg5lCGVotSl1slbH1ts833UMG0CFRI9VeJwLcbh8nNLc7EnJ8e/VZjI3OYQKMYhAYb0WATXOVjvMSs1DFZLR2dSRg7ch9+pNcf/QPm3M5OjwRFazI1AyFIAzN6vNttFDdgS4k40Tnh82/Xhc9ELnksiY3VUoc7lrsbDfiSM8OwGhmtLjz/4e+DjdgYg9NDSP/4zHEeBUuVqqwmEpd6tPfR27IyeBbxi94trjymm9Ru1H/xR0I2kiw9Xn5TAnDK48iqFCj7s+vyd5u3cW1UipXOxGLe6/mzFZd2W94LwZ0xjCYfBrNoCEYtHy6NlScGd2ktvag7s3QSVklM/jC52oVLPV6nCrlVQ3lb5KoCRXBooU952AZs7JMh1dc+QGYkHcQ5LKF13S3UR5YQYXXuXVcFVhuaywVpjutdcg7YSkT6YizDtM7nEMPHmt21g9cdlHSzmNsa2qJh/UfK8edX8fBplTzjBr1RKHauiGx/tt9f1Ap39rYYsGkwVXlfurzE3FDPIqXr7DI1a6ehI2NON3EjdsU9kYwYXiWaDFbXy3IEToJIvX5SiGSOBHZtC5Nn6Sw9jSJBx59VOAYiQM1x2IAV3nwJWJSk/AMsPE6Dzf1beelbvCN9Wy2t95Rw2iShbypIb7Pb0sso13WLU/NacxDNr++RsTWj0QlUA9b3RbyKQe8qi24aiif9qlihvadeQn8yKJ7G7gxen7lfJdAyHHgBTiFtPEOYkyD2XDtsGy8DugllWwErGBgPf/MHaol2fwNpWObr1+FMb0oCvbPpA2/W+OLAuJGB3CykhNLIZauUpoLAtN80dDSfHjSlsOFNFP0bVj82kG5Ch5zMRpKvPVq7bvjVd8mD0LDf5ozQ7eGn0iPhP487HuaLUsFcvZ7RRcRH2HQ5GvsMAVI2198kMgnwflsWcyWoVD4i8DkaJqXlZBwS+P6ZswcrHVpqOfyOQSJRKqKXx4ZohS115W/QpbagWBusmNJ1v8IBAaD0uJZinPkJTD7Y=
`pragma protect end_data_block
`pragma protect digest_block
26ed10d0378189ace48221a1c106991a8872a983b041f0bb787ecfe6b5c54939
`pragma protect end_digest_block
`pragma protect end_protected
