`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
vpJZCaXnZRR3heZlezG+/G07WEwe1VBGLZrQTWCbS/DPznkYgIU7GKIE43qrezIarZRXm/QraLZuLmikpOB/S+SEPcSYPZhxy+Y2K0ax67VQ37kx1piUJjbQ9JLI72o+BMDRRWB7tjzTt+FASXmRLeoDdnlV2/EZJYTdUsQY/q/5JMchdZW1wcxvypvdel5A3KHc9ZjdwBiaMv91IfUSXK9tBwWwAB6OtGXy46rLKHKYiDv6jIGSpdhiK9qG8RkEgWi2vJZPfPmYXp19mL10m5R8htn49wz/1fii6sSwSQcHUkg1UwjBzKTFP/NiV8zpF+zA80Hn9dUF5te1Rqx3T9TsU2INjdQZwL49GaB1XLss/4cOiQ+utpe3kAZ+yxuyQlvkRKaUdUXs1EogP5m38LMeqnmqo+uZfq/7IdXHcLSEqbYkd0zY8cOZO9olZL8i4XL4nZQC+h17ugkUHIR6EHnyqDn+glVwLKNeEWalmD2xvTep6o2Xomi2MsHrEolKoIxE8L3CUdhI6GTpkT4/NUSj+KKx+Mq59SZb4xdG7sTjCbl83/wleAx2cvpBQJH4IRMX3AtckhWPDFZl/kWvO2yDDLr/naw7J5ryJm/TQoqX9nza8DRdEJH8KgtfuxVLflX5g4vM8NShZFsKv1oyDqPYFsTPOUguQYn+KaKjagjaOu7nl7JkCa0zLZE10DuTqZ4FIfajN3z/WzXroKMEbbIDdNCDYxZkRNQAE7VE6nBqXwY1pDaNS++kJit7pxJwO44h5HnhHg0XEUUrvfVr7jGSMO0RabyqbpGA0TqI0bzZ5Kb9IHIAu4TOpRRBdBqvAiBOVptCS+4XFZcCNR32No4knuUA6zeTxFBYx9F/f7kmTnpse3JZagyfqL0/DA5mhY/UH2Xt0H4G7scZF8+hZeAic3s1Pff//qafyMnV/fNsAsv0NIU34ESe0HdvPbvBcvhpo9fv8O20o9SZmCej8xeVQfHxTSvjdUjNnmqLlOb8x3Q3IIST5nOvqSdDsXGYTUn1iVzvfkWLSOj1/yxgCKdQ4AF46JtqtCdbby58G5GoXLB44Syz4rIqJNfJD2ZjEtCVgPlNFsMaQSrZ1hrwaaLTkqCV2oFaMHTaLPaRWGUw3G7PeADm5VAaUo1OcGtbtpCiGbRDEKKfD8ewARHG4qlxMJR7fmm3jmI08xYF85PFMevrQZH0q38K5XF9btURlRr+Usus9Y6x0JBUshiWDh4RnQtaTzjV1MCE65TBQjiwryam3PXFZnk5aWgPe4Y/rIwCP+PEDsi07Kq3joqizxVEl7bb3BK/iS1LNn9jfypMCYRD84vhUaw+24QC+4MF5MGftFMyOmCYZMT5l8y9gkVAthx5HqVJkGJZ8IwlMyj1igzAE2JWmF3L9hYdd6ZsFcNxqOddlPLBRDBlkSkQib5L5VkNsHGtX4eodSDPxERvPKFNU4mC7u31tawK2lzzQtNOV03WCPLsA0doIkhIrZ05E15TFqV8QzBNDaug4ybFBFirJrqjdUyptHouCQ+SUuH5W7FHs7g2pyhBCpaxQQ6NCc3Y3ggM2hZcm1sLcmxQFcW+M9owC7m+hvORyTqFzJSV6VFgMjSWXScSqCKI1lI8knRMnsW8YSIuTy8i5dQayYBtMi+H6ZN5OXXs9WvN4bRHGEXA6bxDW6eGl0kN2kG2QPTWWSK/4IeIkPPtOiAw6u8WjgxHdW4vNo0pOkdK4R2rVyudcRSL8An6vNnmULthxjH5Ym1UXMcfbEK/BXqAuX1XK5VgUSsYwphXjyCKUrTW3ceIthp/xp02SyFU2TpVXi5m2m9nHnUwYITuF9yTMH5yyAaR0n2KDkLswNo8BfElOXRgKRdpjeWSRdymwGa7XTSBxN2ET6YqbcA9fa5RN4cRVp3jx/Pb1dqO0My+jkdWpyF2JrUQ3VPPltlH3jdMnY/YJT707sZtiDaUpRRTAaQB0yKPrq2rJMmNWrOwW1Ces5hqQL4Hf0LJWDdH07WqGidq/d1chiH1kl/KccatRtolqCgZXXR9jxqn9RjgyJrP43asFX60Toa05lHvhgO51iRkZ20gg77mdtv+470QXHPtVvbPnWqgs9ZOBh8CYZ1isAGpfoKsfrbJEx/Bv+yKeD8vhXDJ6xZo6Lra18DQ1OXkxojz7QAGWD1UKEBWpirwsSPdJmM0IlITRGjfBa4JZXp3pozhVXLcU8ABmU78DpdixWX9AjJJDE6IqTVEvULwxD8fawfJ4P6TtpcFh8+w2WN7N/UPXeqCIhr2A0QGjXptflL8bl4l08D0ityiE+TKNYulPj+po5BSaw707GXwkKDHQDWHRGkEH4ROV73Jc5k/d3ea1Ok1Q642+YRvTk1twdCjZmB4WKTQdCxIe29baJnbGsl97KCe7KryBvxJNStoJ72CNsPvdWWbt9nuv9kHpOHkl0lPL3wU0roBeB/Ko2WeHH5sc2qk9frheR0RZY6OuFpogfas2gOdc0jVqTXrLjgtjOY4R7FNaEyBqX8MEpN/0wd/iDwsMhvoKZU0DFfQFfIjGQ7yHVXtCwQGubSP/OOaaTALyrMD0fpjzwwFl+dEJAyx+GzwDmn8AI7oEpmEY7njYfrLjlkc7sB42XkVjMG3F2zt1aqUMV4t0KtSxq8Yf0v63gKw/xlhB2eEyz0GsYvOZzAxCIHF/go1Wpwk3EDWbST9EctRlmfAEa3AUirDWgnJ6oceKcxs69S/P5Ci8RGh0xfz27HOS8Htm65qDn6wW/++rXGHDuNFvfmOhKfI1EfAng5vXCpaicDX22Fs1XA1DMUtjHHsqWt4Pp2ZldABfX7YXrMGTxaB2iZNEFeQ2H7cdTPG8VJFuRVtU0Ya401g14rS/ipSAmMd2ybbSyCh/M3d0Y7Zr15fzV2ClqCn3fkU9wrD46CFxirvDTJotKgqzXurmqGiourkAa7wFYfgZ0PsMw96UQ0Ck/VdM2aV6vvhxIRp9kXCraxCqIZZI6VkufrfRfNLqI4K2kwlxyoLiY3Dn5GAI1VgZu9AH8NDwQAqVmylnWbg+nFDDgR1s7XJSW7S1Z1CZT47vpMBPRIetY2b4+AB8ulOD4+3nFbNe++h+bHaUcZgiwG//DNZUIND9N1vvhHi7g04r+7+/iXyLXQZS+T1aqDBbfYak7QeNDC9sinp/DxGMfl9dySasmo0Du0e4r5wRGcQvvsMOf/0Y2uuUiLSJdmiHzbVBv5oKCTN5aALSkASyB8LkNgTCWzytS1EVKL3WuA5ABtNtW0C7L0558w1xkbrM8ZrUJ2u/fapMyEbmdZE8Bw5yUhlc2qNDsNTpONGwqneF+xH2Lj0dkqGwkwmXVU8BN7tJ0uHfXDV+M8n+cGYL3kOUYOWeiZPBix+Izmn9k7E3IR4ouSRt1v9HFl/2jneZFdyK4IU8lqUCeJpnoAV21lxyNbh7vzJd/vH+OzDUuUXHc1S+ERVRDlgIBRnHPNkvMkaGJ750/jTQiUBYQILRH4=
`pragma protect end_data_block
`pragma protect digest_block
c0bed9131e485a411688794e1243716e685be56f5960b5fa6224e75cc5ce2418
`pragma protect end_digest_block
`pragma protect end_protected
