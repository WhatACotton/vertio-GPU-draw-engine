`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
wavU13abCM12pWb2bHqfOKNY8hCtexMJaToryr5RB9ato3BNrJUEGfpL584xY39KZBoOwEb3sRRzgf0MJRd4fJfpnvEP8sr0a9JkmubD/ZhBiLOB9NIc8hZ+UpamiXSLG0lIPY7drkN/GpTQIM7iUV7kWqZdqFE05XNYjtwGiOR9SoptcNWmAB/saXFkhlyEgL8PWftp+HYy+adRgaeIgfNAlcVF0Pr66/PCiN0AVNmpJ8PsOmHQ4KOwAzfQ1Zhq2xTUjqFNxQwE949TfSI3vKlSJBXduBeTQeIklk7xKMGtpwVTC0I7au51ie+R2lJyXZ64pN6v6X9zyrwQ1R1b/o0e680m+3yuGA561YetxFbvzKDm1xsfLBScv0KBeYKRE4rFxS02cheDarBJVPeisOgaX+q9QaYgKjfYrjtp5O4OYMhf0CCdmwTGY2rZ210rk50atIGkdrCtPqCMsKpSOuWD7s3cyasQCbOeAnwz3hOylBNZeQCrYysf9x9brCpXB2A5bmA11lsraQbNvwTV0ekiSZVXydQNgi9vAiGiQ2haAi4OwRHV/6T1zUP32nITPXDeDOLg+s9yLB156Yp5xOIz7o7jT32UAMuW7JfGuE6BRKoSCT7MXa6XVTC8YygoDxeAKLQkWK+hai/dEDWJogFm3CRzCE/fM6xtgwQUwJKZNemA7mvg7MdgHBSD3mk2Kce59ptjnPI0jIc3LVu6M3RUJ4bRvTaDKirvZ8zRUB0llLO/g6bhYMzzgLi97F6PQMXKUa+ZEjICFTLR9gPTKNzF+UQKGucvCDt0rUw5KBgyop+AzVh6WUjO8KZUCb2mJixBKH4PuZGt/ujMOitgixMwvLmgCjYkVQcWsD3g54XnavfH2SatKVdN1ocLqji3qlvdM6huetwHIZFDmucCz7p/w32/uyR71xYKUInP7GuQCFJ0/v1DL9LmFLRa7A3flwyk7j1CLVBsdRRUtAR6pfKPkU9tnKHpbTGt7GPe38fHnMyfDqu2aVLmzUKW+/p5DF9bCUxokp3Db30i+/b6E0OoqUVrIpt4FBiRSuShR2LOFHJZKmn3oAdv9H05qpHS3tTnxPkbylmbolDN4Z0vFLz1aX0MdWcVNlK51MGwude3UsPJaW/zWL0oKuhAAcFLNtxhxk74deKGLVRSTRdMub84UzDl4hmhEm1YVRn4Adcc36CxCgVNo5tlswmYU70ogWMR1NmbDy3c0NpdaXX3H4ZyiIxjHaOAeuSTdOxdk9tsScuZgGGvi6hLHQiLtqmU0kbQMPG1OMVO1VvUbV37Hs83fFYnxeTHon/ahUQ1hnBrwcQaN3luXXJkOCH28h1Xr1hNXtcXjLSWNluBlHlztiiqNKw8yQX6acMVE6IYQRhhEmxVQBbXDTcbUl8hctMYltLIsEEUqrg7cQRdbySn1gAWdSeqbwKImwdJD4xz41dl5Zd6ekq8BOYFS+MZ826nz6Zivqqs1UgfsDMzjqjCkYnBw8xo6qj+JQ2om+FovR2Slyo6j7bAD/hgfPkhcvTNJSF24KxI18qeiTnV2E5EdqSQCGaVzibh9+FMTJN9de3C4Cr5ZZ2sEwbHD2svnHVtWEV2l5onyn9xnfm7IG+6vpXL/uKmeYbwbOK9qNsqiy98OCNngAAgjF43tkbxmp2Cb/Clko/Uz/mQ7koOBcOH5zizhERBQlKUDM15+BJVJ7L7lQHgg00FSrWfIF08TvFfd90BadoJTp8pT8brisarJmQujyiq8MelMnn60Wf6ag8qYdcVWvPTgYOMot+XDUFrh4N5v2lKklyAAaBZsmxvx7PO0nyUXt0Z0LC2hqEVMrv/n9sphX6f6l1Z8rd2D0gjYeOrTKaQqXnKnA6NmSfHwgdBO5foBYE0jr77wCPe82KfAkxVxhrAu4Bqr0lHdqBoGTaejmD8KhuKcf5aNiwLepjT8K6kQXjWWnDGWMaznPkQaWCLce4pFWZlhoqwYja3T9u79I0NHHnZopv7Yn2+z1UEZg7JWwhpAeiTlhPkjF6YJZN9BNmkXfZHv5zfAI6mTvdx7xf0bvsJdI411YnBLDsq0qANnyRZDC2AHveiM628ZsS+5z+idWkdsYp6C3O2Pz0dehX9loy6LocfKCTjehvIOh0XR2vejZi2Xy/6MmS6qrYBHEgeDLeZwjWZolFP0Z0ERG9cMjapnTxxgIgLHKHfAi1+A24Y79FYxvKtw9HlqNmWnNH7N1zro57+fVfH+lHaoC+lNUo4gkSdPr1Jvf/5/vlKjTC6xzuilkYBBsNCNUK39tBsI5+wO++DzTQMbsCU78dLhP0XYWvchtZ8N6UpBk9ZUH5qxpK7WejKi9cO1f8m0KQMUWSZb/V/i3lIKzK5SqtygMD/27i+nY7IkatF/BuoUaX3F3DaEDjvVAnhOB3grkiEBPZiVqf0FFIM95nciQmtN9pFJPFl2E74qy0CtiJrRpYEiz0Dq/NLqG+b3EWdVvdIq5IxEnxt/AUAv8h0vRnneiBcG4b6qdiTEPvTsVDFOkae2rd7w0HI2Xo16hXNrrCqyaZnjnY+DsT8EvolufdYOnyFigUpzHOSG0+qimoiFWExR+ttpFT8nixCi2pgj59BSnW2Uk6IkmOVgPg8s0JmZ4RE0z/w0HLCxVeV+XzM0v6V74ucOA/Xc+RG3+I0j/W6h3NyTzSnkoIui1+kdZsexNgmM4Zx19Do1up4etOmlKckSewUb/PU7FOggmgpfmrMVqoOTDRy7uYpnUfTdxwEXb6JOS8YrWCpoXlsPGHV/HAiuIjlk3S9b8lg0tHjBaNB+smIXu0I1bsbyV7s5IsbFnP42VvkQ+/WVyN3mkCr5N/WRDWs0Gg6YGZy1WcJPa+f7ePrWUkgPlmhD4QptagBgaDiK3zvB4qXAUwV52mOOdYfmtJ7z+ZAS92PursPujR5paul1Ql9Qgz8kGO0eRjSuZp3w5GaD11tMnowSVUHfuiziwHREj07WfG/euhYZkzJ5Q4Wbnx+rxZ36V0pyLqaSP8ZuZPMDL8ORuDbJwxO7eGUuPyDfcCshmyvCJLnHGg+YDDZUFSUXNK3jHBp5/MbzJYcumzDC7kAAZqcS8G8Uc0RIsVfyZWrLuHy4Xu5URHhVM6xPIVcZhKM7sWppGpbwRAhsUw0DrjiyFo+uTtKQAwyhNEaXju1mBdiiTSXh4g18LqPiyTo84wnReJVUzTi1RsB7/z0K3r6c3aR22PqIcwsTO0t1/CMKfSSw3h8Ziv0uy4YIAegYUnuOrhRosEVfrBijGaMOvUx0QcXcWnOtsdX/G4b/wzhk3uhCIJzRCMtC73SA9j1CvbdWb7C7gwRKEyirFi5Tca1dHw6TXo/4/68KR1fMc3DebsquwTEfrQKGTJihWoiGOS9IuyrSqj6FgoeXhkugSoWcl0BZkneWq7tm4fkci0BdQ4248kiBy/0BE7f1AMoBH0F34NqGiAxlwYpwz8JG/aIGHeXSmwH7GeIjDDlI/9WxumDP+zVpR4WArwCxCnYYPndw5sTFrXn5+iq+LyIem+54zvdaBf8ySA1N7gZWQw6Arx3IG5IWVc1xLaEQ+HT2T/aoJ4MLHf5bvgvKyFGiuvCVHqir9Kmwcr50BnhIpSyzPi/+AdCt3kwD9tUAwDOS+lA59dPScmcSUxEVXbESwYlA0I8zUK2vSq0pexn2MJvAn1aKmeuOkqbTsgtvxuEKUoKbzSg8tQYopBvfMW+jvh5C/K4H6g0vz2o4s4RAnUIVKd04YT2nnVzEnisPhsjq+c7oCSAgvkxDBl8dELbTwqGE45g8YSbSVDZmM5YHnObnKBGT8wDwRQaKBLgpa3cffp7AkMRLmj6MS2ZqZRo/f1pr+V6Nm4gNRXWhk09IyN21+4gr1qSmLa9Y9C1/JN+sN/IvDuxwBnMh6ADYt8BRnNvrbgrJHCeQx/4+njoGwtqiVF9+ykMrWFgi6xtrgqztYMlMe0lvO1MA65nDXUvieIv/ATGxB0Vrd1fAKncoDcgaW6sa83lsvAzEOuEsAfUhaW/hRXtSGtJs3lpVoXaPOLA6+fExAovB59ULEy+mPM11o1ujXlIasGhnXW9fx1GiBZacQvr8CkK3mVkeaDom3DOhtBjIG8FEVTdJuZwaJDnIl8wgpKVkbKKuIl4gL711YVA1DiSwDxliWmZlhjGouxzgvv93bOewPxCe6kADRWrB72lBXgvtLlYU1LMeSGiyYPE6cv512z+O/rd5C5DI1ArPjuv/RLXn98g3Zb+Cq7CBTnGSVsNTa2OqQQjnxnKT5kX7g+lWD+kNgbIkK4j3Xf021W1X6AK29rOh1d2xy4XHntsMhl0cskkKGJWkQ5NeA6rXJYfCjS+W8p/noVB7oqpFxLWxlCOGnlVG7CBydboJ5fkpaFbu5djGJL6DhI6ocRY0kNYv8DlosFKHXR2p/6Q8i7P5/JCzHoOug08NvOjB6bOkxyazUEzmfM9y6yZhnbjYYNW/EJCBfaHnZChsCKpx/zkSHimGfnxsmoOw3WXmZu2Lzb7t0q6zaKCFOHYVBE50ghf0b/Ai+swfrL2K34R1d+HwtIYp+pnRUdnJIAp/qcD2vgX5Os1Y3uMmCjRq+46v3Z5z/XleWkMozz9kulomx3krz89cNYAPBzlejlFDka0igynYZHbZTgjErs5aq2lS/LJst/sQDWpQzVnnlEYD0802OmhWe72VtZUk96cCyJjsUfcMnN84/NtahW4rRDpt82f7i4USpKaj4DxLXmEW46AbL4vNw+2cBpgoKj+aOkcrI8fRixHiYW5TKXCH4hbJOSXxyeQBFdczlLwwfu+BYLIIqG5PbGKA5hopo94K5qO5TxAdUji40DOCM0A5VwLWMPCclQbJxY+Y2GlWtWmMtckOtibcAEPWlKxQ0kt2ciTRm40Yeu+lgdyvLF3SLv9XjL2epjWjFcYuriZNbYEG7ozGphTzPJc8CGPRCe/KMMlcZ/SMstRLncj8AEyHPFhNfDkdeMts1WxJAbjkLz0Hs5VCP5o01jr6giNlYPsCFHDEJCXUpWTBCD8ojv7C0Qt3/mbFehs0QcujtmtXAqBMdHfKcsjGxgOLABnMMhWEQIcvG7Ml55QlLEi+WspQ1mRvoKYpyurLxDWmrm5b+7LG/4jTwRG6ncvFd5dD6ADpsr8gdyabwnn8luXWk1lnTiLA98CGYxNDM6f45b7xnWdIfbsv50uscVxQYoXufS0aWNhpWbbU2B8uSWvH47o/mEZJUI0yJlKBlOpm+IPTuVUoCHvHLHMacFuWVPs8KzpyaDXsG0t3UPzQGkgnepD7gAw5A4oo4uu2iMJTvD9Nd7GQker3h/lSK7zoeMcE/2LArKvuYf4pPFIiVs7TnLPKOMDZ8JTcn4ZdgTlcpEtnmmm9824+lqITPskwcMUqUlTFH1pt9voO2acubkGcLyajdM2uTot2je+za1dMK+3AzhuLE9OjZDedmjGUI6IyFF+rcguedwacbQHv49XoM0bmatff5GSTMz+vk7SJjiq6sAqCiKBngvDUus3+imjCXOLj0sSt+gB+tbu2oxiNR/E/taxmzpNkFKKPWad/RkURJb2/B0V7ma8yPKwxoFatEuRQ5OZBYc0HXCbTMwQuExZ8BJWKMOd7eecvr8fOeXt/ylU6OT8FMG/y4Y5HZyk4ujvQ8M8xgcGcYkUqiIO+KI1hKQ0Klar4KwmbEs6R5ofgOztxhzEB3eMFuoN3L9TbqOiiFOosBYo1x3T6CPtrttB84gOQpnuVi246oAc246bvKMvW9QhcDPs24mFoz0/EyrOaWm8ZJQHBiVwwwilnKPTaiwCDeUT7tAvfq32Y79aMyyjEoFxZN9NXVmfxGRvtRaXkG4GHCgXj1GK/eNvBLnoQ0wG6CzP1Sp/CHPcMlwouXhHcqjkD5lyd6F4ZyBzYd3CHPv1ZOcFAx3xGKgT6ijxceU9jayyEv9jWpTO4IvY7BMKyN29qGfsfDat8WOqN31czI6YGnFRQmHc6209MyTymtvfM6OnaJAaIp6KV4yQwLHhLWwenRk4YON5QTrGZdwM1ZxrHW3JCx+ITyNexBPlMtolnkSc71j7m2DpwwMroO4QaIx4rNVANdPkrjwrgo/WxA6IVCSc3Bq3ENc7kd+9Szd1V1cPCn/CpPmYZ0bCqskI0wyHZFDWMnk4iGAVTEacRie7SqCzXK/1Mv2oiu/ShTZqL0QDIqZpjYT8SDgrKT7vZ94/c5Batbf+AB9oVgR0YCHrNvKhge0KgRoZrLd9M5nBUU8FMmYrSRyvJt3tjoEprvuwX+RYUjk4IpiOg6I6HBxMT9sy3CKkZWNnkHee8GFasdkyfgXEkX4w8VvGlhbYRKIZYWSYNZZkVyx1RtFKx5AeqNO7vIvbtDgsbG2c+z2Vvf1E45cUrSyUP8MUq43Smy5KcuEx6aw+949UR8H934f/mtJPLizwzGdW15vrlhlGhkP20e4434haxisenAWjLZlK3YZtGEHvm+/KyI9N/t6K63i7ZgE9E9PyehWwqLsko+5Q3GpKvUZe9GNN8vN6RsYr021KUXDQFt90I0sezB8HHwWrtWcRawDDT0TFNw8fq/Arbaq9GCpmbFd23lHES8E6AQiSkPHbQ68swVTi0MlEuiqEViR5Y6sq2nu4rdKwQFUkQ1852oXm6m9hNoVZlk0WWs3nW3QizjUcNdvAC0RpPh3w37NsSbQXi7A1C8ANdUDzExOhqc6cfljg9QRIlob0Np523Sf09AxnhqTmLoPA1aoZaNEeAAps7VkEo8MZfMpK2pVyDCCBdAktDNTyw2v28r1knM2hY8qDvw3XOcZ+JV+VvyEoyJGNmo4KRpGz3EMt7LIOyrJ6+ahWu9qzMb9lpXd7EANQunpxBP6Fn6V293NIGQjrsLQqZAm79v3gt3DJCUeNPmCxbfNfoFGyeuuOBEaQrWlBiS6Uu1lm+npCi+nQY/NWSVgV8CNVBgR+i/fzjT7s/7yYe2hCCKQlGQrdAjCO5j9HtKYatoGepb14H/CP30rblUzl7oDYjF1pRRm+qqUFRi7Sqet4ZFdUyReJFyVSCV6edpWiEKIQN3HlYDJt9lO9de7h2m1925xv5exF5GXHlRaUJPVeS5bM/DqTNL+QPBDsKYy0XaRE1JUJ+lgWtHF6kP+0P2gQyjOJRChhv+xxeGiU8+VLyu8OL0xMZbdCngpkhmKSEx3WLrekjzxn8GSCC+ualmuFq8CANb5FhDz3YKtYoTdYbLHmIls5V07IsziWm1l6Ui82/NR6fWkl4qx+n5l/ExWyjoeLOyiCj8GiT7NPUt1uX//ZtT/+NQn9G3AsrTyEjG0Uqbx5cpwFhhVaYeLKIIGjEoRk8ySd6GYN7udUQsC0z4JdO0pyfh2aEiYphLE1hFytqbZ1vKcfoll990BLNL9ZGN3P3wuw6zY8oEZRxRRKUOTnWRPCfx+vpp/5+0YEBBwfbxO0smad/J8HAYrmnTfqXnJODGvEm761bQex/zwDw4ivhvhPPMJB8ppPhw1JolTHz3EkFdoJcwyNhnukdbQJkkdO4OkHfI8FfSrKF97lJpwGajlj1thrQWd/G+8MRIHs8qBrRfppQmiTcIfFER7gGOOzD8Xwpg2cnByzdYw5kRH3rDbtgOvGLXMHLPCwdFlsc64Xt5Q9KQFAr77ZE9mDqrT8KrbsiwzRiXIrT4tiSezgKR54vSEtSWT+sw9tjdDJhLdgmP7o5aUdqKh6YMxpRxbNnpzrDsh8qKJ/C3pkjbiKO7gw107lzBir6Vett49V98s37lsSHYA+kp/5z9BQZobtfX770X0mRU+dKGauCO/euv5Tg9gM3RtpwSydlQGbpMz2RwNTyd/qgDgymyyuvbXsNx2Wh4jPPq6ChfgMovMJ4WpdZquZGaHseTSQDdpSZ7vt3hEF/fllTvx2tkTezxL1XXfKES8keLPabk4Dr+BlIt0pCSla7x+Zt0nRMHN+dgyzfoReSeRFN8/PanHeyiCt9PmX+R2GDEI6mIjKpFmnjih2RKrTIjnrEq9iOzSBLV8l+6+QTMbdsMY3lsBzpFBIjqqCFJLC5kfsuBZGvbWbOgprSBRp4n40iFcT7xhesePQgadrCvD/rxKx/CeSJyZPnSfGPaacPf7JaVLN7gekOF2O9XBoAXVjsP4EryFbrNgVkz1jIVTjR+S0w5GijBp6+rhRE+mCQ1t0DIIkLHxJuXzHn8cW+tXoXZT6rOjSKOknSAwUFnis5tYy1x77Z+aoq86+e0nR9avexiguI3+qTqy2xVw5uadyejit0G8KUI3+ZZe4ZPwzNGS/pkf8fWOFt32UUM0aVVEZZ2QBOqqYpP3n1dOz+k//zyPU+6C2xamPfbgz+4E6XbZxRqfUdTzFjJfIlf2Ol+KqSay0gnD+2IRPfraGQlatKhe0IL4dIwS3vfukTGEGtHSrL4y6waharWqk+Cye2iPpufsORGbLT7fyi35j56mruWz+OnfgmJuyWZGOsLRCFTbmLIoAfRP0nTUMOUw/3IqN3IYMysObRNGuxO8lNrlDrH3M9aYQikGaZVHsgApKTBTuS/MOz4eicC3LgQDykwimBf7r+N62VNiqu7RJK9q9NA+Xlp5T+8GzboluiymxC8gzBOwbfJoRi2P50y5MyrIkfOl5Fj89Z238TAML6QRQl3C9EXy4CjleF4GnoU45BAQUH00yJGvQ+2lsAhiWRjsjk4eYUIa1TohyXY450w6WTnFxhcsZbCfDS3gmHo2Vv/BI21+sZ+vjDrupWhAOrWXIjuOxFjnpD+6tZDaM3ceaIMC29J/4LhKaY/moPatgwPp2FJnz8QAssTcpLaGv3y2uKJriwT6O6RaqjcfJ6EwWOsMIC0pG+1mPbFFttJ1etpwKNkDaH39HzSc5fW5UWg/YuEVqIe4Yeq65OtlkoG15htIHFi0kn3BKrOIVDYHRenOFrpTQzwxZXsIGzuSeJC6uCVp1GDOzaG1gboiNEZUCNi1Vga/O2+hjoDtDlH7N9dVRGgYt2QG3zHMNxB22eMp5NCtlgV7+z/+Vm1Jk6+/vh33qp0GJs23U/epkAa9J91p2iD5UAmvqGcY5DAFwpNPJiCSPMAzrWG8afz2kmBRVYnVtu5EhSooISckvYncrOQL/0hlsgelMimryYLGVAteIeS09+nI1fC57ot4w7Eh+dZEiHQ91fa1NmqBi+Na+/q6kBU0c4/7yJIKkUHct/1vN6T8lzecWNhaoT3CZmzP84A2NgvRUjQl4bTRv9CdVmfbKtSHEMrMewkmSz9of1meT0o0cI+E/qZp6rcN4FBsMO02vKdqjOnSoUt84Wfzq7Igoy4TwbJxsgPjfZGWopUZ+EhN8mF3hLKMxSQxJnTEDTYWyD3wLqVVGUfBCWIFFf77sa8Tp15QraX5CqHw35y7ndY0fUQdeRNARxvYw+6iE3sS8M/BrtD+HAkiNSiJe2AoEDv4Ql1Tyz+TdesJx890T6QFVJQdtg6OSy0AmScuVgIP/hBGHupmG1vE4SGi1dNpgh8giGYlMqw6RtXzBkN7zEJbhggyAMStRXoKeHfJPmmRwiaM43kV23BN4x2nuFawabmjePrA/dRp4SMSQhn7WB8fHUt+hsw0O9S7g5HAsMBMC4Nh57FXeq4J3A0H+CxaOWFTYIqYYN5nOd+b8jWYVqX5rpm1rZIWmI1xDtG3g/cduhHDnzDhMQpcaZ3WDI1i9/0ivlQDkHpN54b2enijMRJO/qvly+y1rE5SCOiQM5jjVj04d/JZvMq2y9HK3BGYQ3B26M0eWwQM0sga0dDdHKfDom1CDWnIbGwwctMAo8aa4aFzp+a323isLQHbanN+6REVr+GM6lttpvuLFbJAI4dwAccRmwLRP7PND0yO1rIYJ8q7WH2kK/H2zPllqssagdhrMG9raD8pokaZbMSqkkOwUpabGXprl2sQmMXLdeWnsqpopmLQ27tEEE5ztRFMdiwBsopDpQoeg11sZdjPTqKfkcHDIXk0q5HCPk0604ULpnH802L1mCLTazEh3nAfKtOEG1NAyhce76SlHdr8nzABjsG4ZJ0f/jZQgrprOiizJEBWOnBh3ZU9MQizOnjrxa98ufiuDJPJA0W425zXWVKgLRXj+0XR0rR/81v1N3OK/HDVuPyMVpQvYJ4TZ+WlhzeLzIivqfW0sU2T2F6q2vck7T0yYzk7IYJA86MTLG6NNGrj70YiN4BDVtch9NTIPfNcA3DREfBtdKJkYY6lmBGgqguOpFLERIj7pr56MS/vPzI9WcawZ1Fx0GfsQ6Uy3yWzdOrqQk2+IztNTQeWOczwE9F6HprzePTqSA1Gaysyi9GnK4QRHVL8g8BHdE67d4AFTMNJMKLwWhybsBTFllf5WpH0Xxy2C4YBtIGQFEIRZIUBcNzfEHc/+6wvJMxtdraXNV8HudAqY7bDoOzPvZjnD9z04ftneXFiMtWDITM0qV/cSfTbXIqh1eXAa+YxwZfveMV57AfItZrL59qz2F7TmMagrq3yZiNdvYbJlFiqtbrvzmpJy6FRaZbd1q/UEmRrvwfx94BGOk7W9KBG1YhRDm2wdt3m2bv+jIiFHAbG7+DTwi6G2SPp+KMOKvI+Mb5bpg8sDTKT6jGsLhufFprJBqmi6pMUtZ9biccGwswVyjt0RkmiH/DNPYoMwbZ8pT89CnjuekT0smsm7jdRz1IXZO2SZJJVMdEmM2lVv+EKFfPjrwigTL+tgFZWsSaupPMWgAgS0KUeJN7rD3fgjELJ9uqrGVVYdH7uEFx38LTShIXX/iDGxyVYpixJxfmTMKxM3AQ7i9GehvnXC8In9jGHnJXvnQHRKw4SSWOs22/msWYJ+jRH59LSUd5+QuiVfcJBX0avE0yDRXBszekYLtiPG60CqI/4gxkuRCQ5T1OjapTNmXIZ4gSo6MD+xKHtkLvbfmf6QCPmGJLVofKWxNfMKtpCd6DXeeMGjDpDvEK2OKAoiOXZkRuWnbuIvxt8FCCrudjjirM/aF67flvYOitsgLy8I6ALfXYtfmPRzdYoOxnUB98pcWfNcl0eVfl/CBkSHaWyBvY9lV3plEUBIi4jX5xXQSSB+1PlzEG5ujz/ITYrmabEmUV0NxZ4sf2mzI0866njWRvsVoDO8V6t5TyCk+OE1180LnxrS52pJKsdpDRpBtd/NO7aQKg3BIk+jzG3b47B6ZvL0s7wIwsxkAMHhy/Hmys0ZQLjMV9IenHBaQz//gDN/YCb1cbh97m+YBb8vwzG1qLFvP2C9FfSz5Q6h1tEzX2QLjVvgh5ZWjF7+nt9zCouFhtGUp+J7KH7l7VX42G3RCSmME8nnkFx4FPVF4FquB7GU/74BaanQWVf9NKIzzWWPUhpsG+3FpH6PGrbq0u7FOfvYROqCOVrrNVxk2G2Gl00FkhjfkjsjO6Zz9bS86hxmaZnWuzj9SJl53WVdeS4ICM1vQLcxiji0+nJPybJetlwP4Gkguq3Ye9waaRh57IoT+IY4zi0ccLlt4osgoLSbPdXiNYqLOXhv/nHdHQZgj4NWwkmZhcgH8kIA4/TKmn92hwFjddOHV+NmayQ1bs1Q7TerhgOwvLU5n1UkdL1VsFbwImpOUFA/NhpQUmaBsfoscy5Ordvjojsnt5mmGtwMcYc6rf90B5ifTTWHIEZTBoax5Qgln89jgyBe2v5QAXr8JhFzPyYVfb7ssQNztrqpq1Txrt4r5UHZxZVz9yDHcrJDRHqoh8y+6S94vuq0k0Nv8EuvrbeXzWNvhhDTY9Wu09GRVPXIpJwx9lLdTksiCJmgCoNsfufvb4CmiDphNVZEyTjf8VPXVqHib56nYigaW0dLmafcChUMobplrBwqPXWHlho/1vCWeZ/UiEHZCleADWhnyB0KfcuvO+ftctPOgX5ngtAnRZS0yX7pnU+lkbazO2SJt/xlfUR7NONp5+w/IEG5t8gUUOJOuTfqpKgBZpEgDk3SjXsIbIuuSwRVjtPumksSwsgRmyeckxrep+AkVZgTjGaj4ArApqUGV67y0D3RNEOO+f06PUEWNI1Jil8NAvGbXPo5WI25D0uH4KqvNY00UkzGI9yorhQUHhvXAF5enckvG1CZ5Cn0kQqDtIXK8AIVHjY7oynwdd0K7nqhGTJ2pBSclRaLt/R7PoVvwz6DTwwTw/tSg6GqOdrG5SMnbFoUPnDICU+tZTC1TrFKWxfGn0ycF1SoYGqM1Gxms9B1TS2oCmJXxoaAtx1V9YJ6XrbfMb6Cb2ET0tJPvgMQVGRUq5cfOEnSNdjr5ttTxkFkns8RxS/2UQPfnd/kZdjXZBfcPe2QdwZcC5sifC5kLhhcf7VztI7FmO07l8/AJkFzjZJX+XHuZiSic8Vvfd3VCHbc7ughawOUveN/YnFZNVsoflpN0nPl2DvAbsNMjZ8AEicOMAUe0YO+VWVK03i9LfxqqpD4qYF9ibuj9ZKVW5cmmA6lqfGsdo1PaI/kS5ZhL2TalKotQ/U7rSXwjtaRrAX9XS2eelJtVJAOMpNHi5PXplPwOPvxjqBNvJSv6G413Y9ofdqIEjGrig7Ttjnhu72BnMZiRy/cHTcCu8WcrK1v43yMoMAfla/STexxdPQt6t2iJCWnmwILbeDFI2iIrP24Fn3YlK5/Klqn+9SvmPRLgtaxlHlPp8l6eZxurHiDxZ8kahhJlyEg8xRnTY9NVLh6UAvpYKpeipA21uy32/ZEnX0R+YTYHX0l6KOq28onxuk+XWzC9BeTr0VR79FIT3Mg2T2jq+r3eT1C9WgUD8VQ7N0Ff5oTSLH9IeR16rdn5Tf4/M6ppvFlK8LIMKdgmJqIMxwlQhBwc8dvREKqB9Msy3eIoyuNXDs0PCMlqVFaXwjkKMjkYz5a4/xlWtGsqbL9KWIiBzlPhC65c91l7zcLft7ti+8yQeYgRTFv0cYUnRaga0LoJ15oeYZ8gsp3yYOEk2TYx6woSZBmJeYO9odUhdIeN9mIAUOj/lKXOKRIBQmyxkoh08wrr4L18s5RH+QebVP5mHn3JkCsn4lTJGD259n/NZxFxJP9HqCY6Zz4xw3187oSemEdnpelnaYy8h3ds7iCpEI9zYSUULMoukeRQ7xQJk4pxAUF0GfU5MvUKzxyh8Gu69E3MQiF3nrvlO87XsEc9eYzXVG4+T7XBtcqGaAG0CK26XsWhiqf+SCKKLSTyN7nUlgyP7w6Ya0avJh8FUwAc0gRWazfncT7+9oMRhjlayUjm21BIgcKW7hNDZXUII5X3q/Ct7TsgY+CNtWJbzqihkvrT6PaaO99AKbKC9r5cft+lqEQplpRfqe8vfseAgLiImxZxGHzZGdQe+8AvxazLVnkowScANU0TxhRBSsYr8/sMor433yVTSG1nvnFAV5qfnnB+5L4e1sDgHQGcGsSLBDMWIE7DrPH21Wl2Fsq6CKEna9ZIlZ0+uhnK99LRKV9Jv5WJstp+uqL3n6xy0myQuFBE6o6v8P86iFn/sNIDjPD6BFtQ0s6Ffa9h/DfBbGgkJIWNuY8Hl7sipRec501D2stbSnmKIGIgqxDgkdzCWJudBaB2n0KKvGzXZ4M/hVm9f6+u8SniY7FPfZVf7Pici+bWGc1LrkGuYt/1TMIZzbx9sYDToSwmP9VsbvYsR2sAfDx5VNmHq23uGtist4+AVGmk9Tp2qMXULwWcH6rgD0TnybNzamnDG7vwnfJVmgdBc/X1amHzXRZlHKlRbdEAnNewwaaIQMlZ2TmbGy/bOPdSC6yRDrQwBXjmmwVN0/nEM8Rsyt4jNp6/6r+R85H+y5CvZezgYYbzZm3kO0RMv7Ea1p2+qxXf8WyeNnNRsfzU55rzRMswmjlA74mzCxF2/JeQlYUgV/hLV+U4zJyGD356w6Tod6y1qY8Ety+BJYL6v3APWpBr0pHu47za4BirqvraHfkoVyon6iPDwMQnOsd3/6+inT/8TdHK2UYBxR+wkFDAF27em6mePJSOY/8Fv2cOQaJu8nBh2AgFMsV2y+G5uePiIy1Gse/Txgdd4/XYObNF/iZYZuhheZ9IXjKw2cVf4/r37Tse3bn1m1tes69rQjLHMwUux0EUWpFWvip2ShCsCwtse8E+szhuqVZiokombIjhwRDctn7lSJVqFJe/bIyI+eANwg2aokEEUG9OR3vnh3/C1jSY1fFAlL0Ou02PPp2D5QEgvMP0Dod/O9pFdWq9dv3qBcSvcn6z+4nksYJFfLBX0YnVJPDuAyk7rvo/aWkO+DL94BcZLaA7nXGhB+rWNrd/MyLRIwyHzvRlgXFj9Dz+nPJ83tXMcs8cMPyOIABpQqGptudRJcGq7XSEZU3dDaUI6wA3ve8QNqB7fw/mcocly2I6yGWKPwjPUGZHwe+TThKDMGdih0ANAagALE9wWzeSx+7ZNBAbg6S6OGyAHTePJSInLsCxWeUkZ6NXSMxUR4KvBZMq9AyWMhK/djIl8kLlcxYlGopQ7bvme0Ggr3p+sm9c95ubyjuO54nW4Q6IvRpBuY7NoyS7iTLURaEMX47vlrhj5C7twdTHA1UZMvrQxul3YrirjQRaEn/tYB9ZQeNmsTRfJBwWIzErCsHERXLKjT83Sqnydl1Wyy99Wr4vQibKtymoRkdEkgLHepQNtjnuPyYwwUuP2aJWBdiMNkmTDymMd+2SnCPNVNvAOXj6LPrnAtiRVLkbqp6V0FDGfsirxup3tkTjEjQIxettshKHVhZryA6PIg3YL/Q9FCvjW2zWmdgx6J0vph39W2SpTIcBtN7DX+BmbMZMV3+fXLQHmXjDiNTQIWvv+PZZ85zuZE51bbBmruU02Dq3IYUOPKP6XEGvzZznl6Jpxb/ON+vdyB0bgG/QE4cTjqtWCowgeVphovtlRPF7ripUup8aGtKf5vfE9Aw80RW9lUjfeiOxgy3G+MqMMIgK9dXL+eZNRRgCPykdlYZy80VK+2KL5xl3B2z8KrduQKGFq9u4MgAHsQIp0TFFh/9VLsUkLiWMzJDDAa1HFINuvGsoFS+o2MA/qmEvXOxCkOcm3Z2rzbLFc1NvTSa8iNnWP6AX6lTffENyXVIzb232IcOKZKPPaEW8fJU1xJ/fqJbJ9Pi4FcBTukU3J491IkCIxcLrlQxzd0rXOYo1pnYBKsYSG9rq+X9qz3kCoV+mAdFMtiSlgLxI9RTcQ0qM0PaLMlVsHhl7KoNnPE0NR6IMOnFtqCgBEMO1aXDrun4y5zF4nbqoswTkh3cI0r0QOpujV8ssGMf0O1j4OHJxUHTer9aX0b9CRrggPIMyQ+I/AFr3lPoC8rIfPu0BfQEsOTGQkom8KRST9uWiE71nVjpZJm/o94+aJdz3OqvgSEBHEd549pArJmRu1SgE2+Od2PzpKQ6QAUut5sX60573IR4Tam829uQ+3a4SeuFb88Lz7YD3nuljgGtx824itykIvHLsyADuIS5cHnfItcJeoHb/luFIpJdecp/UBtNaU7w9vZjGB/OUHcm1tiDD/agzSc8YRg1FhXhQo56LNh47/VSGmM0B6TDgPBHp43ZtrxzcCVf2lbDXpZqKU0uMwUWQBVvw4VK3AZeiWRge88fQhWVh3DlZcS+7ODPYc3ZQUj4A7rDYDgy1QaYXSmRmGnK2CfuZjU0RWtXdnVRPnd8Qh/oWJO+aFEnZ1/dCpE+V7+XevX7UeQ1lcHlCLwMBXOkWY1yr3+K7HO52RzZY2wkrAP7u3Ub6MPwU7I=
`pragma protect end_data_block
`pragma protect digest_block
dff1f9d562f0bbda94209de3469f8ff23e6842b05f8e48dd6d92ffc4b55ab659
`pragma protect end_digest_block
`pragma protect end_protected
