`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
6mxsUd5Ptvec9ye/kydQGn4sDuyjdhD46N6/lozNCHlGE1/bFXNLd7jFz0KEx5TTigC5GFmXybiGkI2qS3XfG1Zp/SfqstFAJFainwcTtFdFiyfRfxZL5p7GCFj/GCUoIuIZjEMQqWQzYaqUhf8+nOjtoEBrWM9Dz7+CAacDBo7U1cYXLGgIsGVa5d12fX3wATvT8NDt4qFZtxmlJmmEgQCxatTaNwcIq0c1R6A/1rmvchOG7XD2Df6J9jxyKHx1hxjWEHf+YbBwAy7NVzdS5AO30kwQXm4mn2QcdWHmi+IDRa+F2V8NlPVJXMMoZ7+PzDhUcx5SqLU3/7/dhXEkN+Uwn3kf5OkhvhO25qgnpgS83+Ybd8zhuDNQwcojHcIUaiIH8VRXcryqSPpb7nvxXL5qqRYnOXKSxxNjCtu9FcdOuLEfrE89VMN4ZdywawGupVkKmDJjmL3J6V/1HGuLA1h+Qc0pnboOdEP5IgKS5d2WJ9Jie2LBZ6003fhvERm2ugdhj4dOmprYu1IPPpi/LsNOQlUAD1yekRkicBma3dKSLs8U8m4i1KnBa7hMYLc7R02OZxnUSucMkMzkxDYGlEWhMXcf3sbKYVc1MRxZ2upqcOfJmvrSxdZlhMsbhs3GTQpL502s9UjD41K/ugosG1WPqEZ3PMmD9ZOkRbCHX+2e1SD4U82ybSwzPTIHZ1Ucp/iiquPrET1W/8Np9DJKWzFJRvMow1XD15hDnRLpwSaQLH/8vhwODbr9tXX7g7vd7DIbis3icmtY2XxMNnAGbFilhQmpXfi6iz2yMmA5jK3pcdD7HfycOp9TpvkAm+kN0jtmcWzaGlqPuhoHZiHb1MFLb6NYdjl72+5oZMRWBodKpU3Dc39UgyRqYWY78u/RnP1YUiqxxjfgXBKPA3Ew8hXIG0nWe8zaac+yb68y95JLL0DQ7XPFOPNoOkzcgdsVaE3JVQNytzsnKhbxPoe000NKREK+sP6nG/AuicZ3qwf7rdxmO3N209TmyXQqkH7Y7cF5x+rbu+Sb5YcZbfvt1yIWuvmUB0DNYEggqMfY64dvb3QTaybOGjM12dxoSj6XdQW/FfPztAS9T0IGy6K2M5u4EMJXRXD0kSHSuTJPEFlyXba2buYKsVmgqu8qKND3ZbZl+/fUO/EGQflW6zENKWfpj9DH1L2Rbi47NZHd8wrIFOFug2neBojqKIh5xbUjl6oVogrCdnxQhKUAt0wticN4i2dzC8iJA5P9VAL0grl8/K4ZMOkCQj2lOe877aKbvdCfngBSqVcoJLYb2OQIozNhRRrWnw7Z70/4XUTb5ld1bFGPZeaumUVAwwUNupxBX8YktURiTJfX9NA55dgy/66vvuFpFDwZZuz/qLQhxIwveSMaSV1XTTBQT2UdWXe+jngsZlz8i7oQoq0Eo0B4AdJMCUWCTAvJk4zCc53J1esyDr7DGxc8dM7jgGnRbLMYkGlJAVb4SOC9h9BbvVxzt8o0Yz5Lz/2rPw7EDUpsNq5PWGZ2tkWR19vmwBIvSRgDxqS+gSqvCU92BxsDUshHe1cGzg6/bV7W4/62xWSg1Xjw8zqf2UktL89q0A68D6MgfAW1E9NMDqcBSeru65sw906Rr++Bj/tTRHiOHgCgnxCnkHbyCmPRBVpRZJy3WYlUMyscxzeRXagBNDRZta1x7C9rUx6lLOrrrK/5WXm8yUgC53bgzUGm0A3KGUw8XJ4rO9eGjQj/tJmX1qI3zUIAFgjAz0Iyxnt9v3j5prOnkpsMeGeKnX/5Qf3wsW8JCDFKVnL7jq7gfO/gk9HA5mekyfaQF4JHM2MrltmTlHU6MmUn/Id4T45V1saYftoDJ1Wcp4iw70OTBjOXPPWWjuoPzuWIPEM0puLtKpRdOwJOWe5QcPZEMUygen4182wY8fRvUFKHEp6NmsZVxWRrwFXJtDJuJzt3qc55P8QCNyJD5VBjuwBbCYuczx7//gFP3MBR7oxXdH1POb8p5qn8DvEpN+2nNfz1hyceUJr52m+inTfiTnrJ6zNj4bJKvxyqsuO71mtQ4w09AVngqBWKw2wUS9vKW7SHslCdIf8MHw0wCr4ag9bdj2Ri69ybY0/TmHsinoPzK7JEOyb1CJMoqJZXxUdqVsv6kzCX+0AXMrPN8pWpy/tOtdhRhnLjag5nDseCb8KSKbH+5lbs0TQLiYCvq8AXkJQzeCfmf+1p0FxTCOiQWdV2S9gV+uc47/7+dFWUEFMFSFKTeR3R/Fv0xbrW3gbFwGJyXAp3H4zjCWUbqNC/0E1g1w5W9J0J+n+zl3A13+BxmhSBf/561Bl+u/UE6yATjap7xMS0DOYI8204pjZHEgbU8TcCpa4/dYZY4YWFzRz7l8metrGZ3zo7QKkhtn+uCpexRTjRJ8RiINUttBQ4p5dFyxnBoLZPz7ulkxh4GyLvKgPvCZTXUyYgF0iGBbrcaHdIMVPxkjTOHwAlF4gKyzULy5YeKe532oqOkThZ9h6MGYUYKvAqaZowaS4qRgVvgOpnHwZmwZaC8MwSrAyEXpGxtBSJiDhw6UsAITBVgv7St0xOVaBb1CZ7obBCvEn8Wl8BemFYogS0YEiELd8qwOEwTltPn4wSdF7b7nk+7nKomUMH25A0lW7sRkhqYy05M+/Ghd4ZSvKafNIE54qYGpPZ/fBa3OuaowNwyRkq7AqUlVwOeU6azRhTAEJb9pvj45GjHvyqRNQdVSJ+nwzY8MEilPNZCaCnZaqndC9B26VOmQnhqnC3Ddv5xPxGZQ4nriOm21fqOEQTlYhPa6QeLzeoKMOr+tiyFOkkYhMMcpMw+1O1aheA3xakgQywAJ7a0O4gD2hVo1i8dcJp7yZ3KmvybNjfik4R7MrbS4mKMNZJMAbpVr01ZoL472C38iRpKUC6tQ2Uv/5asCYDdMYsibgzbq8XkZ+xD/WCj6O866MUZNCp2MmlwFz44LFl1bPlrMFiqiarqd1cSfLXYPzyyhppW6D7XJw6GshaQm0EucqfS73ztDTVGATLsLS7Z/Tcj1sEYPLNSz0KzLWhLHTP9y5CAcD+t7NR81ClSoyH9Xf1aA2D4FSPR3PWFIOyEe0U7aRIIt2wbTVyrHcFghXNfphjb6FM/dEQu7w7dtbp1z+5b0tGIlDxmAWo9oxY7FcczWrDKa5n7rB2fz3n3JHfGX2V4t/2UsGRFwnZwooKshdERKmiFbg6cQXAcdqLPGTWnZawqCOYj3wYYkl1C0ACnFZHi0EXiLpxMGMh5/NduF78srXjfh+Gdqp331enntsKRBwNFwWJ/QbT3Q2YL6l2m5vUgcvSAQ6oZam3bHPezwSHDO338LwA2moVLcjg3aIrVYhnPONmALT2lLrBx6eMXSXJuR2Oxqm56+WkZ61N2bp+aV0UIBBr22L/ZRfaf9HTeR2A73XQXbnA7LzuSUpi53nWr2tJoN7vkVABV+S4WPEIqRoSBqVS61RrqP/hM8YncbOZ5ELhZU5hqgB7IGD6OdZbl/SEOyD5ovy8ZR6QwahZOPzZHmcFDC4qap1p+20KvrBAg8oQckj/5WCM6zjxBDQ43xLT3xX4MLB5wxVmTi6ylx7+1ByrD6qXY8fwglHZ6iupfI8m426yEl6ZZw2iPE0rhGTgjcK8AejPR1/6obsf2Ys88a+d2+80xLfJNuCCZZD+HGjfMKbwewPa4e2X7i80C7FGk/PPMz2eG3BtLa/tRugieltheexFcmIip/g9Ch2N089ovtPehytjjp/yTwaPZyySRPaFHjACLWvMf/tgNqte9QYzENY4UzBljX+RiXFh9nWi8kpWwMnmBkCTGSQE5rIKlqHnZWtDM7ToCWZpDVn47sJZhfk+NEYcCIjRg/L5vXbHRXUH6pBBtZ724gIq0ba6MxVdfNmH/0LRqgCuOp8pLMCxPDZow/xTXFc1XqODeui7jAytA+GSUiLS4xc5Y2zyy6XNkD57vD4LkQ9X3VhQZWEweJ8xIDG+dnCI61a2vg2S9uHs7UcBrE0xbBY3ec6xRsICXfjzSHexVuD0I8Qm/xjzWFZbp5p1gK7Xd7Mrl0ffy4EtlD8YgMcCGVb2P17FzbS0Hz6ONyphtXhxWbs7jSrMkYUE8tzqEcae7ldiB1bwayORn+T0wYco1qZZKmPjzeJ5ym5moEV6It8ELQOVHJnvFc13T0SI+/Sr5Y7B4UpYZTvlGvS3GnZvH2cOLEW+8oYzh1Tj/8wLIimnIzvXAXs+zybPm+hKm+cvUOuorVqzNs2wde0s42Lp+A+wYjvCz08NSF4T4KoEGhdwtBOT3kJCT5GMHBM84G700z2r5vImivPGYyWC3PuK8qAnziw4pRI3ytWZ3r9jOUth9Seji1srAL3o2Ymuc09p3e29IXnKi+ZZn5t7DHODe/7AjCSh50VqHhyOhv6vJOmx3AoTga1XwMG+E4/ZMRsuUOMz+YcSB9tJXC2gwSCsAI5RMDfKYTihFRUE24YRkrQ7gka1WbLehgiJq5wdrq67XfzOhadRHXFqHWKmob65ZaZtl/kloZ/IVp3zyQoqC5p8OcsBR42VMLEFexw83nJiqn8ze6UpTl4TwdBPw4I+FUm4tv/MWg2NRKY5yQgX2v/l/heUIMhk2fixIcRXbHcCuEBMRiDofuRNZ9VCQfp2u1L3V54yi306vbXLVWBlhcX26u5VQK67vIeKxS/5xmtttPZL2fEn3kxYB1g6JIyblzXLLLuLjXKpelLlng52mRzHFWOmBPRzaQSkzjofVm4z/xTENpmRfptV1AGe89UJz4neMRT2zcxWdO5bpzNVltVifHFSjti7xaNBc5wxhNx7lbp2d+fRdvuIWHbDFgbvpko7jcxLlEAbvSQ0iJcUbHHVw952Zk9tepF2UJQPJklcuPwTblfDUV5AKrJesceauvHwoYCreCJH1HQ8OfryUg9D8hYj+07OQ8+ufggcV/tY6VUtGMC/LjBpzbYdTcNUx9+yRgqSzyKzpHtwHMX6qzAz1zzi4H1mj6C02R0PGtjo33tY0CzhPVtWbVDPDreIwgzP+O179FFaSTWmqAYILB+ZpwnBUpUNWveyPcwqHawtL2rH6shFpCfORcP5szOXpq65nDJ2FMh7XHz8ojAZFxA188FTAAj/xPJP7342XahAqal2lbdcbT1HHyn1o5JfqjqW2a0ZBh4pGYLLkew9FkDUuo7crod7KM3w4YR7BffKuJEs2HnG5eoDdioo5jpbQCcNaifaRKZGRdV5lCV6zBBj2qSgOuiJowbBoyYs3X/TOTipU6WFkjjzrhpbVMiGtBQ3eO77mMkWzozVI9v/TFePw5wSi7da7fuLlCyfKwUw++0wSKFNxnVpRjJ+48hgybQ7C9V6qBfNF+xXvn2fy8Q+qH5+FWcfGv0/j+YW7VU3+MS9c9JgznBgr18+l86IBVhImXMIwPi+VqprzEsYiMpn4i/l8st+2d7pqTlaWXjuUSvx6Lwt1tHv2CLdOuMGUa2ixYg6aQFVP5DJob4CAQ93+ggO5bxXAIK++2JKiD4pMvqROdEkvLOPElX+EohAbaykKCI9BKSS3ovrL8cGS2hdWTzsrxljno1rPOt4SBVUJsRX9qsO1XO0oKb66d4Ss7Z6MLxAL/Tw5ai5d/eKO/KIH7C9e3QVmjqPkDc8UWqw+7ULlq5DpJV+y86wCrXMxdfKsU9oeFIX9wA9VpJZZWukQZlUpyGrVnWxC0NnQD/wecVx3X1tQEKnrGGRgn60iFZn0L9e0L29AxHhd87cjxdgXSukFsnUXv+EWZMBIwVUlcbBnhwQJT/rHDV766XnHF3mMlogkt/WoVpW2ALwd2eafBPV97gEYB9rGq2AzKBszWfUaIS2L8hCzTN8dz3K6GKUN80aLQc9TnheqQFQ/QKAr6nRHSyrrkFukn3L/w5d+CUjx4aFkez/i+lxCaTYGeoxQ6KiTSh9mk5CSkK2oQDYrLrp94oP+z7GmJodo+nRNII1OuOmpEkWEyyE75P/2FmkIkGisNdEq2CUyRaQi3PSpkFL+vzrUHSxeZxSzX67oZMj3+1Fhdaj4SekjC+HNs1jlTO4hDsMbtmdSklRzttO2ol8tGk+uQwT3q1DwFoRw0rlvnKByw1BzexZc05kHGCzHpBjw4F3YJ4Zjv5veYoXf3oS03/6L/kSQ71CYVQT5rW0ykkH9tq4viSfTlXzJCXCdaJzIow9YJr5hD8lYSDSgTxJkI/PvGd8SShU4MbrYglu1+/FI8Z9iBv1Gok3Js8dxsx+DHueCulbtRE2oGkZfVYRZz1CRk3jCOq594dxGc1t46P59yfasfeiv28Rg6zdURRgovc74V/jGNCjNVYLf4Tz0JN5eYVjHvdiihcp8C5p3bEYf1XhrGI/XfLQpsfVtp/ACX2sMR+KZHQBY5+2TsC1FioZpzOO5tG42UhNb019nqlsG0pbm8j47TSQGSihx7iV8Gj0/h0vbuYVshi7jBeUaRxqoEDc6dnq4n9d/NMpBy3EuzI7fSoybX/25ymPyRHv7J+uy0kFI/9swQXKUYh9luFPVBC4ob31Vd5V4Q6jaC3M0xDi9IC/j44Qz5AeW0ao7NEkpEqFrBkiWyqZMXe3OWT2IbyyKy0W88IMis2aH2MAjmSfb+OKtgdvOj/x9CUEIio7I7Oviq8gdrxcQtPFbGrZqbdwB6dcyNuptPaTmicV0U2hsnQdh1V/CX7R58Ee7B6okGFE2S78O96OatdmjmSsnwjsVwE24DeT0yGtjPJ6qQFe0PUzzfN4vYzzOJfd4wBuJWLCACvTkQ1W883t8XgufQi4bzsEq0eYNX5Re6bypFrHhNJeG4Ut8hOnSR6E5+kIL5AZHjmiqfCZzL27IBkL4/oQXnActzSXNvNatUaQXi+IDUJnu0EoFoawTBB9fh2XYNeBcj3iH+V1qdNOh4xHldocXmH7mHGiQ3oasRAipkjy1W9Jce/hQ2kWUaIXWyx4DwlL7KmJu9reD7mplBeULLZh34gXrs1SoFGfq83ICoPd/4+OvrlNBXRtvEBj9CTuhlwOzLYkCMJrnyTDNZoJn3l6wvq7yHyncg4Dh3KZNlr4IgL9lehPcQ+XYX83JGQn1HuKHI+jtfVlDUNQFceo1vXkBr846j8VZC1GihHPXCpPvzvCbfDXjWuMLaQaZEgAqCFP//1UorLMAxiytzkAJ05VqXwqp0xmSLS6gbD6k9Lqt0KAXjp8LVDuqdrDyuJiTMH0HufeBNKkl9esZZcKs82f3OSDAusT2WmrAniHOiFCmUUA8/Yuy+lCKiJlGepObxdmgnWkRpZ2a3umYcFSuBfo3aVB/vSlWB3p4y3bAiPRVBN7sBSiiTC6hcffWyHkry/1w3nlFqeX25CDnN2UZVjY6LWEG0x83ovTuGPJ0KtvR2nOEy0oJooizXpreCD7wMduqp5PIxp417MlmQJb1tdmVj9hRnKlFI6rlVnXU6I/Nu6NXq1ICIsEzWxZQeqz5k8ecntbBqFOUD6sBKW2bLm2gAofgo5l29lzyKm5gvfHKmx20fiH4xZUB9BATFJMhssml0XNCAUs55jo8WIgQ1oDvvddLqBTjPHfd/aoiZLsYbNa5xiY0g2nx95V35AI5KqXFczRYVBmM8kSGv5DMeRg5/4sFswS0MU2wDmyIZSSk2kUFpaQQSEJiOlnHdACqdUg0aXl4SdIGlkgkMWswhvDXNWLU9aaVcKYfu35gnKCKy6wSnptJCyIGxsAhDv9T9m8jNXeJ6G3lxrmldC7fgKMiZeff9jP6bfTcvLq43b0RfcNccmcCXipokTYfb7iQUI8bT/jDt1U+U4C5bOV77KSW3bIHLTwZ6ISs4KYP14ruxYN7b2A3v4Ia0xSuZ4r0zMu2MhiFCfIpcMMPzSpk7TYoZdnYViv6uXutKPa/OmdWpD8T8Hn7WFv1xdXzOiFdOzfmnrfAeUe1XWOT1xVTUpWT3o0FYzz80c+jDcUbg+BSF8w63Wc01Gz2nhgKjDjop1f1fG8RJYHD9LtJQFMkIHuMwH2hbbdwlUFoS1ccT8XXfIeVcxkIyctJmgi2UL3QZQz6Atd4u1D3M80wto8NSht5SEfcLz40s3bnXQ5IapkeaDo/+37em7hSf/uNiLPxX3oFsQonlCayWmSvHiwQrSZwXnBC/tHXU/1+umyP7CeIDP7OhI8jWwzuY+kOvyaelogXzT9l8DnCZyuUKGtgF/dygTCvBXJHUwax1Zspz8EHsPaTvPbfDLOpj8D+iRs6Cm5j/dpCaAcj33KJ40Osgs7IK+Qt+LRvZXXcWEf5gmaKmdPrutksZ0ZERT8KwJda2FyhrfFWtCtQxCB7bdwa6NmyJcAQyLFWgCfW7R/BKkKz5M0K5/52EpKnJet4NiH/UrEbtF/wXaAfY4ul7cTUYS0ogmomRexSbLAcKRrFIuSPiZb5j9FCJ50p0EXu1aGBOgzp8vx8BOEplyvHRjrS+4Kv9iXoRsx7542rs8Dlb0jyr8myqbUfpcydIShQRb3T4418WWz/e73RyOTmzYetErm2Tu7cictpzjadkJgD82X7DzfUj1kTi/3YoW6ksnY26iJ+sXyo6roE/8TNr8rg8DGTDhvH7clozLNQA9q3RNQiKdrv+OzvCQ318lGaWn0vfH1uOzPhKIhFHsxPqqDCNL0yNcs8R35YFU35NkiRLQadyC4L0gqUdSe6Jd/m+2WXHhhNln/sov4VU4yszyRDrlcWDZAzet9TF/9Lys0kk3AQk7gJTEUQhxmRJQ7v2QE9XZx8n1QiebN9PNp7X8TE74tj241C9LtdHTHGQeB3sFRvh6vHWNHaoodHvvPwZ7IMIgN9EWtxVdE4SuNije5l1Iva+MKtQE/DjF1JGIZUzDBKS1sDRX4r6DvkPcj6+cpAyfqR2mBegCJunz7m1cfq71sMNmw+9bedu5z4fNBQBquwCk9UtC6bll+XYaA0+byRfw4Qk+QlgVyfXnwGGw5E6Aa81oiQ8TMoi0KTiUl71bes3M24uLeH3zjnzLoTY0n3hu2t5//7Adxc8loe4c3Gz3GTjZBveErfrGJiGS5nyquxRGI9DYAiUxW8Qi/kK173vhnX51dU+xnU9gPL9gAagCfAElmahTtHuem7DERIzexiLL51NQ+n3FVL25CKF7uFRvQIz6tUh23kLFzicFL8dScLf277y6GAXTbOoWHEfS0ENC2b2FMAm0pyQsJ+xQASDQ8E8cu5EshBqNLeAhlfjl9GPzjhehOWjya72F634jz2Lo92zKxc3O6hi2mEmRBfubQ2PeAu+cei4ZN2ZIYRQOlkCszfUf2b2erd5IsZT6MtGpeqLxanSqWfZCAJxHDM48nXc4Ct/C+/06X5mvRUjQ5PueEN4fP/MxZq99wfrIn1K+jg5i4gM7na+VbNuZOzzfmzA/zDeVuFqnVX2Bo56KS5w1jmUoMlFkWV8RlSVtuPf+qFk1zk++D7INBkwJpMrzwMbvA33ZrWrm7cB8m4C4TGIsIiNdfG6GUFgVhbQIHQtCWC9suKxuqw+lg1o62swoqddjNVGOCwgImjTgpu7T/LaoryqHNjEI2Hj+tcDy5M/nZNVYLNmlkYpjojrEglxShJh9fBiI7CAMtZxjFA5SA4WaCsjVxWXHqBbP0VTVWVJq3fr7nW4MYd2TdpPrQigWxrVsU78e41ccsHkLbUDj275xVhHCKiyCSgqD4g7H7Df3GFebgDRNdll9PCaGe4DICSefnGxxy4Vv4GQkqiwbGyJ4uEE2vB82qJJIAZ+jbW1Tb3jcbV2fmmr6xfH3z3DhQKtszgGkvAperbFyqROKqna+rMSldhQhRduvexjJal3NLzOZ8aCU5kU8mYLLtyb5wCeJMjmY6ls3VXUh/13d8DI25FeGGLSlFUyMDL8vDQTNUx7BAqJ66QYLVTybU5oHp9NWvPjSo0Wvzbn5XRXKPpgvpli9pyKyA3BzjZ04+6JYJ2Dg4mYT16JeJTKlqHVoPOR2akyI77l+Mwqe68JoszJcjyotAUI6DW/aBaUQrD/lc42I6XS0ufLlfA8ebdj0+/dMwiy6axfuS4CvG8mDy/C/BpQFmajsuqwv1biWOKpdYvUgLnvPT2bdeHcqo5/XWplzsBHIfYmGZ9Gh8cfkBdDsgEL8oEDUp9jKIqNPHblAnce8A8NppQmk9B5mevLW1p6D5FkS8fHwN4aIEO9JJwqpBaDAeTj2I4VvH+GUpa0+Ma1asTcY6NTOwkHxPeGEiAAn4nE4E0j6XXMiCfUlO8kbAgHZidn70Qcubo5MZXeepQM8pRg4Zfuewoso1vJWhqUeeyEGuxQDr+6VMC6M7IITqJfHAzifkst1codSStMdXn/KXLpolukvzAsX4b8dYjnZ0BChX3jJcoX5MuILwTXrpMiY4pofxWP0fROIP1lEq72m9u3517zmg3oytGIbF0ZpT5VJrjFn4q3Ad9v/Yc9xT3Mwa/Nkwjv6J7dksHp6u6D1zNfLm5FJPbkJNMm/2zuZfeB/Mf7oxEqL5w1cMHsekBzK5SEXjMeuilVuRuQ3SOUK/Ql66Y2/vrMmRT5q26ZyKU9TcfNoXbaPFUJ8IK8RjtTL7ubThZzn2tPDcVLuU7D76F5Hou/j0oGDyLXwx4ThxZoOVnI/QyuFtakxWERs3q6xFCIf/+I90xGBSUgcOII0oU/XcFn2oXO0bxitpMnIKY76Qxc2a/4wpRVOVmGCoJ4vd042lT63Vg7v6X1qAmm7nEfh7IHqTcyFw9KNzJntpf+/VQR42aSpGDYUkV/5HVas5gf+HtZiOBdd+E9Slu6UzxNNire6nvUUZIr1i1o2k3iug46X9Jla9pxsk4pMqLex9Ayi5Oo66kPn7OCUVmzlLIqrk/kgsWL0kmM9O8fpAzC5Kl01cevg/+YiiGfzmnvUVOlGZIyysSNEBfrn4q5ph5nDRVVKDnaoP/M2PulH5EhJ6IfOISKjyYH6mKoKa4w99wJZruoOyz/S6Yg3KERIHa08y3lH+rX4UhmJCjoJ8jXZ5pMnl4hb5dcT8nQoEJQQHchWr8MvdlknBUkT1Nyapp40VFdveydswwEjD3saT2i5vbk65+lGXLVnOW7eTLJUss2r33APcQhM9SPhqPhq21X6kUQFHPbZ/Mn10sXpdLfiu7+pwjAGUZA0VEZMV18Z1yNw9LNDU+5PPpQZachJFRrYJKuZBCUjTRNS6Ng8vS4wS5yfhzXqQtCsyE2GhoBgAbdqCubyyKC4gRfTQ+WVCJV2ZyxphEYuQxql0KPnFZx7O6Af0opVVA9CQjeY9HIBQl9gmBlKU//fL3edlRAieGQGPEY/bG+YL4h7djxA2tyduZDGHnUlKUIHP8AwKw57J+TUOH5Erc9jOwt3AfxYdZIJ63GOtdUZuGo3Ibb9PPCAwjXaAiyvE1AJTvtGrmzuGtO6aWubZl+cN5DCHDt+oE/REfRaOerCViK81tMaEud20HzCqQJdU+AWKuo/V52aG+MPT+bST+dVyng42FdjPSIJXW6D6chloGw+/ZxE+5VUXNt2b3jQJJ0LCDjFML4GZ35Xgqf7Iy7Z7pzEpoZTqqwbBMLUtPEGFEwhLGBDNMUenKR+VZNBMvV0a59BkaybRMlg8IrhuV3ZNwDINR71ZeXl40CZJpB3QHPN+Ayzod1N14BV67LXhAVFgD8wcKH4KrhsQkx0MEft60uw+VLPQ9qN2yMcSXDCq8IuEwhOCTQmQpMNmaGRQRXI7ElyB/BToCTcvAd9dUqaAyXeosa/euMs0uNGan6qJwiG4cVv5jGi1fQa/EYn+mAqI5xo0LBQBmzbPOBaR8s3f/jYj2wV3tSXWl623Dh7+QH0AZANcyD2G1XKszb1qyXoZfQEGBT79SEY1nX2txhtnuSv9YTYaZu+ZFgX+Jjb6Bgv9pda4XZH/jWZGhZxNr3kA0QeGEZcE640YZdozdobufbCU+1/hOC7ofXgtCFEZy8+/a6iA5L1jOvdcKGkBufHbFoe5AwLfGzNJs3hMRguc1t0vCiWd0CJPKzwpySd/13aY/f+J9WfIpyt39oU+eCGZ514KEvFgroZyMur+A9fQTHohppy1m2pL57U+ZCekzBBiw0eUbcK80ifoTMj/BdFlepiMbmIkoKLw1qkkbSj6iAJrPUgswGt1YqSMqsozNYyJArWjN5oPsTofrRWTP7DL1YVKvhKWs78gzX7XUaHzUCHaKreokJ1jr/iV5pr/0pHnygpbr8MFHvz96b1WqJmfJseLit8poMZcjA7Mm+acR1wW4bji95WYFzim+eWJOHPd4xy4ZjTuvNSQSOJ77cHord+G+9JmNtAAQ5xCss6XInvPTvk4Obna2tmOCaAF7ZHU5F+TtDb1ur5fbEEkuJhdrxRTXZiPmSDQM19yMC5vWIy2L0fw/0eCxAqBK07Ao2qGC5Vb6z2TVvieHUJHsw2c3UsJuMJWgldh6RVFcwHdV1AHA7fhvSHTuX00DhywO2jCbnu+B51dgyg1gOPKg6EXL24YmaqofTZI01S5zZMURNdvQQTVNJv1NDwNyzx3j27bN1MkdOckiBm8rQ6dw2Q9H/CbmtDpS/9Arq06CHHoHXbO32KVuLWlU6GkFCO4JutAG7eD0Vcg/nnJvhREze18qayuwojHcuN+kJM5AOPxfTQN80SZjfF3esGeTIaOTJKtSu8dVjpSG7GyieeBJ5mXISnhUmh7H+11aZNYqJt971mceUmp22Lsz5u6opGBva9D7qxRufVRJjZN1aeLTKyLpwGtm4BeMICvkb2+3GOBPVKG/NUMKmXjjs2eXhpNTCwCXxbUXpSsP7gLjkf/fN//69JsIM8rk3VtPwlEPruhzPdShV1Z6bB4RQd/XJDu7770IZAL6yThrIXauF7+tLDD0vW+V07xTodunWhXnlFwCeG6hf5PbaZGyPI8fCrEXGYEEVgLCK0aUHhsuGwCI9HnErRmeisleOuzHWJ0QEp6c6rGqY84Paw8gROv7DrOHrGAP7rcwM/Olxooed53qtXYdLmuPNFCJX6VfJrytfAR2ZxwIAdvto+tDc7JMRsem1JGvuOC53JEDI+LW05f9fCveOgQ+9/bigPr3jePlgYnqqZ0qn+MMnQJbsXnGduBuMDaKJnwB3832tl5MIruKVKLwKGHCqGpFTTDLs99tKMxPKnEFJcg8aI141LDIOjOvzVpAEYpdN+y1qZ7Ks5qmr5QKV1DAsZ4NJL1W9Ke8F0XuHXt0rc7nPlLPUuzroSvTVsaO3AzosjNzmNNN8Kph98+3/FPuTe2PEmVYTBsYTD8U/RUeGlNS45QYBzW033dNfm4Jm4EUR6vSYS/H9Gl4jB+XUTkIaUScNusUd3ADs67ZBQjj1GgDwVkLFbruwc3eyKXT2GLSaBELtmZRojTfLffplORDGZjUW1LORdwr/6Ra0Hhc4zCRvlQsuKV59kVGdTX/5NB1n5IVJW+RdkfhPYZce5S1Qumvp5zFl6UeOZMrWJEHGB5fNNLtQUfyljtKacMvi1LTtwt4SFZ1qzBVGzMMlmXb4NBTigQES8HKBHhaRtv+mAPAObqYOFXwzcJ9h70BqcGfaf91MjgpLmqLTV8t6zAb7Vcj/EBowH4vNRaPujTOpupFhnKlhQOJ86eimlgNgB+s74DufRyA8RlbJ0dnIelpUNGJCYbvlFSP3mvbseGdAUiWBHsFNOWpA3kB7bg5LtLySfQE9/ooIHDEcN89zaNWcLgorPUrF/bR0lvCLXuEunof9tnGULKYM5Jzpsx5IsnGyKl6TdJqmr74CYwe2PeOrMefxJIRaGc9I3MFdVSsfUJlbQXRwCZlRj5AZBMbK/HkG6yFsKsGhe+1WifEyI2C3CnU+qZncBlIitJMi98MeVYzylKEBLPWOZY26ktHL9bqpDX11xkaKbWnH+Pnth/D3LXsJGcAIEcDDs3/ERIC43vxamecutQJnH+uHS7kP2nKrCuVNBh0I8aAddsWTd/ZWLKpmMo9aMRZQGbVEGUPr1+fhBpo/0cx9UNJNcY4GTS1S/cexEFZZckPGEAYV3WLmE3r9oZ6Jwb3Hu/tn9lpWsycMq7CTTVTAFvA3UqgzfN9DKi/7aGu4t76SIzs/+90TRpTZi367GztklBFio29ODyOQO/lom0coLyODA+wLMEviuf8bb4ttphtdkkCjABqIvwgz8OcUD8nqgcnjLCn+KhAngEdeIMzM343qdKA87L5XBNRg6b8qt6AaGwxF/GjbIialWnT9NDAIWOP41se2vFcLc8X4zyL8AUAKwF3ncSEqrNb1r4HmbdqG/Pg1gVC4E7NB7l+m3pXJD0A5SeUaVXXbn+2WSyum0ruwAry97lwBIkfiL3OpCDZnsvY2Jrtvd73Xk1jK22iBCJwEkynI3nyA+BmuDTpbhOblYAaLy8306c3RV9uJuuPmJU5STLF8ycLESTQsmwbTgT++dvcQu1OQ40Or2iDwa2eorJgLAZL/XmTpv2O8bTe2T58EYIGSB9vZPRFf2r6jWBmQ+pzbTorOkSUv/fyZLuZ/mk/OXZ5ukndMrl9wgnivbz1EB+xsTJqvZ4kyyJJrVf8jHt5hna4HHw3lz0yLiyVx8maB+JHylcVar6b45sX6VcTg3jl6OZyaQOWXtOym7bLQNwkVtg8x3STiYNxro0ONcKZh2Nkm+PuRMCKhCJbC9Kjklp/ANAiuzBH+PPtDH2ihYbJ1p16KdQjwaDzZLcJhiDjSuBMHi7t+b0azeEMeU75YR5slDd5ZkOnGiTp27pIi2Ubvh0ebhGS7En1bbNiWjjkp1BgOJY6nqsg41G4RYFRsbYSBN8J+CRNsP1+cp9LHbNl6YOwnk/QzVMDD7UApDxy0fS/hitHRP+rK06uHj2DJtzc6Tj8zMGhF6xVWoKM8OQBAKWKLyg+IA7KJLQo92ir09t4gw3rJfvQ2l6fuEaMAMtzWyQnvSXDEoEAebjvZYbvwuV6uqL1nFcAakLwqmD8QG5PjkLzDCi96a4e7OSBMHP59+5sDsFPbvVJmYA1HuMwXytmhjMAKphsI9Vmrh0tqgsz4QDAwOXwtmqWIKWzTBf9zT7wC8skO6uy5v0EK4BMY0m1UscB8POxMJa2UBsDtx5juSHJszyFuce0JiuncWLlsOP246+4rWRQKtV7EwQJUQzEQWaKnl3hgIC8XgWgoEoTDGipxchl2lL6f9tNfoOzu2eeWA1arNrD25LmXOEC8tWzwYUhJp6f0rJySmy3cF2CbeJJ+HRQSrkOWy0zN3JJ1UOEuD5ISMcU4d9mNaFaIG/PG/Nmb0Ta5cyjPHtNX50
`pragma protect end_data_block
`pragma protect digest_block
5a882689e0c92e92c0a31aecd1f143fda4d713e104fb296ab8e6994989018f52
`pragma protect end_digest_block
`pragma protect end_protected
