`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
H4h4Zukmil5cEYqCzJF+OeGWwh+dFzAiJR3DaoDdVEolGDHcZ8kn0QyU2vo6dsX70gisHNrFaqHtmETno+6Ec/1xMSI0gnVo9OC0okMpV2W+UmqDBX5jxR0NK/p4LZlnqoMditvGq2FoIZQWpII+8bH9h+2XOYc6p9ntaQJxJIguAJfEuNhhBw9DdUHgXNpg7Sw3ldob5xbY6AoYbYVrTgo3heu/N8dNOF5aXTdMOZQPMqPOIcyAv2f/OFExRqw6dapnlOUHyA/p125mTd7Lygz0LZvxQmugPfGAc4xIAODj/NWxltD4Wk15/eJ2EUUhPgXjVRB5X3SAPXYQkVHI74mRdS6nBscEEkwECdMDfofeYojoDtIiV6YWD2K9daAMr1RS+KU1r4yG7rxF6MHKJqO9A4mA5jk9gNxdqWzF78++AmXwhgGsJtHFjE94/gN/rgxsJcqb2M9q7tzCxgsxj4wfTjfdwFbTmVi9xFZcDef/ZzyvJruYR/P7jIEl+SBupYidM4bv2arbBgEWIqjOrd39dJ0AiwmyrAPXN+h5EqMg9Jw123kDAm/dhfFxN60y+271a+7NV+3bi2k1gHGAbW/wy7GkphCeG2NqE3HQX+zkEDWnod5lQOHPz0/oYeZvvoFFxe1WRCCfuOGQMGgLRGvJ/bDMpI3oG8M91ZiJQ8FpQuA12bERVEEO2aJcIUnnpkWYr+79rXgfpLpsJYOTq8Vfwm6QKtvjIf8h+7Iu1LOvk5l2eLAAOzPY0XYetkXpNZvyF2Q+ix5Qi35iFhQ6u/vU05JD9jWEzvivCCqeQmWypqskrIsVbWQ6fnc/sQQnXniI9/p9c/FwSeVXASyoWdvr3dY/+kpFGTf9P7btOKoRrXp2hAZG3rLBZS2Idu4XAoL1CrrucKyPWFlNBJ556/nc3yRsGk9tYOMlD1emmFLhVQpXYh+47/IXTxB+AeLVZDT9x1c1S0SxatJGnkhEF/fc3QXdQsrqxoJhoLfoStxC9jF2tDF/DFgCTdn//WaBnqrinygr/Uc1lphcE1siW3HJt3078y6DxNtk4h5DkR1sg2K5Vbkxz6K0LYNOtK3+2Y61cHeXtPr+tHJsbqL/JSblMIRRP1MJ9p6nkEdcj6nNKxDN3j9UInJEWU+v1B5xFASsUExEG4fRCFwiehYjnihARQswqhB+VGNfxtJvADgCsSmkwJfpcjDE3aSuoSi49YVmkmdcPLHNkegN9ZW8JuqPm1oI6HoYeifwoECGizyCzO4YKxuDoiv35QE2hgW3pwqn/9HDC8gw07xoeMaGtGzfjjhYyc6g7MCNQizQZFn3tbv6Z1ppwvKNtFBsnEgZJJnrraG7R9KjCbDc3vql9IbIHfKW4AfloqkOjJoTPVyZ04t414oK2qaXGu+tb+v3Cwnf/RaY508WQIGOnU+3nsPcfGZWh3RFZHTg8etEWSrxS9tumoFQbWWvh2uK5Rs2uiyS9zfWnmZBmi4QbrAnZ/2834I5bKpN4+6NLHBxtItbWu9Cpt36AcgjVF1Cdo2TtJbLgKEU/TVAujzQEU8v6AOgV9DLKTxJwiObaPjWEKkie9fRS51AtONapYDulrb+L1qohdKvXJlf1GDbJchFuDsLgOlOpVQu3tqKkJ8uqkLeu9hKotqzOeYNJ7FTFy/EG7/K/gUq9SQa5vRsww7TUjPh93VXvgLMOG7782dmAUe9QkK+YUiecDxdBfwJX30JgsInJQU8OXpu/zwCsjiz4gbw8cUUOJn4Hwg4hwHgb7JBgLCReWUSOvmguiXpGxip6N6mjsYtOo6BrGR0GSGUwr/1rE1mUxTkUaVIdcTNzFcpG4KnhkMdEvO5Vd3CUfasIg6sfm7qlVz2adJqxJ7fmjecciz/b0txMYaFxvseSdVUBLFVQtrQFlamhEF2YvZDLeL+lMkmEZHDV3qPQtF2OyMgbHK/6kTong8NyLabBAwvzK0bH8B/mprqhHXPNxSI+mx8O5gbOiwhXGi2+bC7g/TsCmWTFou+KtFxxatBmFHQPrUG+MG9tWEFAh2UESzyh9oHfRWnSGEyBGF50z0LllJL2+ECKAHMAzRYyEfobgJlNasIHPK8ALPSYZLrOR3JZkRYqVq0qcjmDEmVjFYld+6Ro44BLGk3moG3WaROl/1PHQxSHOZYwBmLjLd3gM9akgkKXXfDpRoDi4LhPPRYE4po/cVzptprTUndvvMxDlEz/j4IFCrgz5M+ZtLRSKXRgvrzZymdq/L1tut5dQ2flR7/5ewKpmYhLr88nrbveW5j/LrAVCEDOMSpqohFNJFJ4kQtpqkE8VwXmeX0/7N0DT46m6BoxwtmGal8zTsBAb9gQw0yyKglvkAB8IvV7R7bmQIeuHii/wtmfEX51zMq3ivoa1ltwiLsxmpVKJ3BVcf0KgbZgxn2ZrDSEVJvmetpnHEoDQ4njWbt7BFQkLsrxJeHsUZXWluZ3G0jCDRFHoh/3GOMRlakE2K3NfVjE+pErZ8jY7PwzXBfjtZtF3j0tKBIQve05ganvbqq6XDpDcJTsSqPSRmq3u4rxfEURfB+B3OqiDTdUVVMSzSCb5vWwjCVuy2BdOOyYJWwTdpyPQjPeSvr2CBg8CqRhQ93RRee6hMtMS7pBu6WvX0cV4SrbT4ITpRBRnovJYrLhWP63vIeA1npthJ5Y7ci7DhTnE2hHJA9JcKNzP4R+8cI2p4wu+VuuTY3UMWKefcnwv9uMbDEF3p4eY3c9ZbhWPN8Y+KmEr1QhJwDJIIuXyj+RUGXWgwadeHvo2bZti67iN1Xeg0+aNb+bRPZgHEXM7bmH0x5uVFB9IFZyy+n4/vEiRTQySDDfnonaQqZ0a40X8swBKxpv7y7Ie5bVDxYejA6BGSbOeHH7WFNvKU1AdO2SXLMtXiszEFBmOx0Iow7xdVv2pbRNu8iXxPmOP0vn4+ZiWNf5bTBKgwvpnObtx7Ue4WV78fcv6xtoUf3CSat4EBx+epYiaHvdjMvBm8PSj9+pT7CwlNpM2yIXbZsZ7UQPKImFUtIgTynM90wFcpVI1BXNjWQbICOmNNK9bJeFAHyfidRDJkDaAHkWzYE0oPbxNEeUDECHOnC4jA4ghRNpZsuzorNEdEYCmgfSyBugkM9rtc6f7zYO3gi1a/B8iddDBPy4IOKkWCn1InO4tydOguE2TC8p7MP2yeq4QB67iUI1myErdivkm8tJ+rLgtzbmLr1Lj4xiPBFCYzqHxQ3NMPH8i64NPmujACir48xiM3DvMCTNi3d6F5sLyxxQG4H8FwUXQ2or3PsvJziQUcGvxeJdwlrhC7IZ/aObl2tKqaHS0LzJgYonaXgws/JKBOaYnKiz/NzuFGNpyi+WQ7WMxOkUP6GubY1UUZ0iUb8g+SQ0XoVojT+Dpe5KyvuZk/aMnkyFhkUM82NN2uOlF2GbJUY1hmR1+4PWnHcEFQ1EWFHCbp4x3G+GQYzB7Lb04ZGWXZsgbCUQ2HioDg0G+5CsGAL2xpqDKLnMYR/eYfRRbvtu4IBO2MBkUKGByCcs0Fi7i4yhmB/n77JB2QxeKhWPe1ydIPcDXbs77JB9Zf2WUEM7mD+nlBAt6ptSIXKUtIFwhNPJdzvftrWqdOEAccG3/pPO04rBZVr0UX8NlCIMVFmKKvw4VCPUsvuHDFjfP5XFwkx6ME+suNQgs2Ur4iBRqWj7Wt1Mg5jNIVg5XE7Iugg4wVdh26+DVQQdOaDM5VslwhBIg/cxE4eyQHWi/0XiijRO+xOGFnF0XLEkljVRah1IKXuEG3OvRqkcGgvsOb1Hi4HDFvQDvFuKOaIoGg++ur64y2BkGpKV2N/Ou+coIebl2aN5jbMo8ac1SZGzgS/TTX8NS7rXc7JbcMh4/FPCWMIT3ni7gJ0RZ5DN7xdqImrx4e7RjrWhotzGt2uNaaiXT7B/AuB/FLavH0excip38qzXIPLoyfvb9mTEKIk25WtHg4/AGumCT7MJUEQny/3Bjb5q1Mpy6b0KVDjP+5FlGFacSz5VLCNG7Rio1ukuli+whgtqO48IAHwAI0Qb3RSOFRDODERd0UNZCG6W1aVqXsCzHBkD64d6UKR3vADY9tEz74/G+lp9SWn06wE6FxVA2VMHto4n0YC0CsoUxueZGWp79nifeNborgTDPb28TqqR5Xp1Qstt5UiiyCKgA/v9x5MUQ3muXhLC3EshODO22Ze0ALcYlrNmeff4qY/C0MAjdBgGh4LBUBCliY+W05tpo6MzFkqzj6VHISDrkT+nOMeQ0aBhc8vfEt/Lz0DxpMuUMmUAq6pPMUGDO2xHEMBpHmyEncFnNw4PsiZzIfCq76JCqKpIzlXjzDU8rKzA3XvNJHtiI5v+hmV5HLpchFxsX2XlVgqDl4kMOS/GJlS8V8jQXNVPZAKHKI4RyVcS0e9BGG4SyTpsK4oPIabWuRbdkN83lDH5MNiwOwaR12+WZvxbQU8KClN/Iw+HWZUg240cxvy8EoDNE1W1rsrohWgNXJSGC13jEl9G0MkYKaOkWljxWzGipb9uBuB/ZR0g+1VBPKHrJyjgCDps20X1iRrVoB3VXrz2gqT2jL0bo0Pb4QNqPoTBzSFLgTLCqqtST+9wFkHUrTa+s3qBMVXxYJFVRRBaw5TO9xsijNzMRqSnOrW/8/3wz7TbIOfmH8FYMIKOBCDg/Miur2Ed9eXy+8+62XUMZPqauGJsBE2422U7S0kouFp80XKjdtGzMuvWTYsgG1SO5mZuQJJRfRqfATdN51XHsJGhkKUExh48Nuid1sT5harsuPCkYXPpsZ4EChzb9YiU7nKnF2ARc3YQANSPLGAEHcPLalUe0H+LCwCanQsuXwu7BR/3HtBzjwlS4m79t0ERN4vp/ILNEReTls+A7bofGlM2/S8/yWlV1jGwT2GEw0L4jzOpbBU54rvqpXt99yootthKY8Y0AyedVNaBYL+aJBnwsalTc0v3bIyk7n4q/eRp9odsd3gMKZX+PW6N7L58DBJiWWQoFfsPygmUw8IxuI8/qe/s1YUoMOQb1Bo+uPbLVwi3IGokoN0tcHhaH4RnutrwNJorwKHv45znC4VYUuHN6++py3hCU+zTC6gla6sqt8FlMQD92yKJlsPXK7qv8vkrmTCniwdDRZDg+/8vNAkmzA6F/SuQVVngjzQUX+OB7kKH1UXeMqq5YlVQ6PA9nTzEFuOTCreK1AS1Bf/IexakmCmvRpDIhMzMsm9/CGL7dDNjLZTZ+yG4IYhssxap35C7VKOCP0LgDBcBkuLhdRKnzQxg2LMBFGeulQiGZPz2eObaVqrPnTE+/SoPTwt8G1Y2ugLXFD2rvz4WV78ZqGOZNbT/AOWBR0Jymnk9RjmFt5nvw57EoAGagFtTfJCpN29kb9C+yD8hP/SqS0wVrmWkldhqZATeFeRhRqKgO/u21ZPDIK7pU/YR6dcr8CTrZmaAa80RGbHd5eBlGQorF+CaMtbRMzAI5qkJm9bRq9mkrt1vPoJj3koVMdpOvBr9a1O4VGXTbI1FswTm3857kvmnMbx8HfrH0us+Lrn61JO4e3GynaIIX2WZfFY/lgayKJLiwUAVcSZeJlz01FxDg5Kr02iSg0uv2dfYLEqpoSlqCFvU6lkzQJI8CeW+4L0XGmYPFY2q+vfkYI0hU7QzIee+CfvzRNETOIb/xqNGK7TNBOVdExC71RvFBZY+ImOdQBLG+y23mvzYG2OPanuRcxiUEmSCYXzwAfVDgBZCgQswfjr0J+kyAzVEl6lytvwUxoMQuDX1RTKuQsBPBYlqRUJgeZxgtZVinMsy5hhKlHyRPm2UTKJo9b0L3/JYVYyWS0wvsKPHRqTjWgeum/ovGSdWp8BC+2kuFeFr8xA/zWGqkRHYJgHezVRF296KmJWewNU4dqOcG9HYBaRirE5zUutxOlY2/VnB0ocUD3YTa7HRk1wOnzv1swwekc4+oeXr5tOWRJaAlJZV6ew7XiZM8rt0ZbO2FYh1fLUPdXRhTivY+v5/9gTNumuz4c66zPMJ6Fmy+XxAzo5LiKw/qOwFqu6gHazovd3QAJu06CPdezzqZ/5XqxN85R77wY6VCpIZTL0HR/zeXxUeDd6XMWpDPiWDsUbUwSuf+r4dhYhkNbHKj2vLukQKmRreNq1u6U232vBZdzs0z/biX5QJJP+pljCtPHeekouURflWdbpuCMrliA6/mBMeZV7CGB9xrNSEdP3GK73wI2zWRdwHJ7csWMlnEehmuvHQlfE4mRliziAA1ehwuHMIEQq7x3O99fnWs8wit6tMkNVZBIoYWj7AXaeo75RsgxB3xNrhpT9JRUJQlMSsHH5b4cPbIUhWphhtGKei8OIrL6HLCEKk3H5kGTvxbSlVJ5eBkv8gdNqUaupvhBbUQUoos9PFBFvnJIiDtJYZ55YkrnSRGI6w/7EN/k655mpuFrD67TCV0VxWYrPis5R0ux8FqccXtcTN5m0iETBG5slSnbD2JzLKUQJBsY4CUNUNGW4VbwIY6mSzXOyRwlVIQzHvrMTq01LVo3Fg/lAX+wcmhjJJfIktOEs/llKnyWPE8voazZ62z1Iqd/FWaOY1M+0yZawLaYtFHWbHl8JoTZG1aNcFHNlNUpgGRxaFEfyzdxaB5ceHD31kMHznglefZRqTbMZMt2Yo4RyiW879dVhj/dHRlppljA74+41vGP4KKbbLd3StISPrc4FrBIC02lGNgctUC5NWNoSNHoRnsKJ5cISHzhhAYkVpIxFfjiAAIolflyLP+L1nvRy6qG+Y8i8Xe+ms3NwZsiXnmUeFqK76lhVJzIryigHtdRzTuHPBntxgV7K6CwAlQBsS3/y+mDV7+I2cPusEN0zmFJ5BLLorxf8XeEPh4DP31gIkkaauFSiGSr8dwMagT66UAVlU7o4uO2rpzUx8EPd90WCvvc/GTDpc0NBrBAqp5Nf/a8LJJcir8CSsJyfainBJIWjQ1pzL7IyTHS2XkBRar85U9u09C6DW0yTxwr4UtpwubhhzWtY8OU1UDXdqQMZCkHAbxOXhRrD0hUdqzoYv2apdVgfE/8GumTtkoRukt614x022PjpGRi/bfVL0h2clg4Y7/hNMs8aPMStzvYvluuKPKUtUKYavTO/XJ7SFx5sP41n/pAfkPuFG4bIAhTDgHsRBUsZXIeoc6LOMulZ70hHTMypgKjvam3vgVJRyFPTYENPjWrynLW62CnQSa1C7J0Qed/XTMP7Snrxh4STeTYWUZpuVzK6kY//eou8GxCSSLyyZoqFfJ5Q9ysGpbu4NB9iQgBwZO/vh+gYxs5cZ2LXc5OEltXyQpTGZkHToG5EGDqgSjGfoxS33D9PRc+wNW16yaYdvyaUkVaYxs9TIfrvgTx4MUsMLP/cXPLbiirKBcMMuvOdxzDXA8BmR07BdzWAEfHQ1R+u1QJQOh2GRP/KhzCb4B3/FDDv6uPknn1OPug06+HnVuRfQLfPVDZhfPPdiU7pSw5anrcHOoNfUXMaQx00huThkPnP5kx2HlkXjQ8ZI4YLCdXo+5zUMU+mkQ0wLHOgJpRosFGd/qD1lkZKyA/0RAcbuOjU6ieny5qM6x6WgGctC5kyGHYB3ajWwiXH/ZLYbLdhEf6FyFa3KtC8BqrDJzlbNDLMAC50ObOHwzIQ7BjsgtDOQcAPEM5Ygi4dwEPb3pOt8cBdGvs25SvGApZZBf6vlLX8VEqyCmWNF+YAXnhXXzIUONIOzEzVX9CclfmLxkXqo5e6GGHZgQg6O+SK54LbFtAgYYgT7WPQFWhlN4Cl3PGtNdYkhONOt0B0FwH+vNA5pnnB3GtHO0v0LkQqw69coBWfys6BgjIkX1h4qElDqFKOeVXdb8n6XiuhxzD8K+jRhapqfld9opHLDMoM6e4Iw1aqjOqakTxb0+l3JyoY0bUxaxHzY5DQsJK3ztJfW/D0DgWH2589usxe7XR+XMvswUKj0/g/uG8Mnsca9VsNA+/WZXnq1b6bgrPOWyUi0PMOqzmz/B0HHjGKqCcleSdRVqLvf+44h0d4hVamTxcyzmmdfllZLS6db7osn7SjRDV2B1qovEesSbr0P7aGM1DU4I5jrGOjRC7F6E30PwyOrTVMNijWLdxnDSfbZJngQZHYYwC+ksoLtYQ1JZ+OXdoUMT/QmeX1yZeUlIfoD10Vp8QTeaOyoxGS8JsRru5cVeEIQW4VIz2js5haSri+ubxnE0q02+k6dWKGpIUzlfkVEXjNCS0BYfxUXPgjbGqZo0pFdY4Rh5GgYBXKo3K9WwVOU1G3DG5qyi8/ardrTadBygachZAjykkTbZZppz/2NZesg6B+PKf/dfK/PYYpR5pEAgcKiCOlBBm9ycEhuGXK2cIQYE3Pw+zrEtWeFcQ0+sMElLK2f3jU9V/XpP87CroeI3sze5inz7c4hH+qiZtm1h6I3YBiIpsNRZonyrU6fwNCBTeCg5iE0UQSNyUXl4srAC1soIW6PRVPAzNmeAVq60vvrkHuQPRzN6QPZKO/Ke89i62m8/2SMx1Ptk70D1dgf4+dhYxqmqD9tlbfm92wz7UuiVs214eWXd74QWQrR/ST9paqT/rJqAp3Rp0KC+D3F6A+wbkxOplKWGDh5nN16WiSwaLA3/pdimZkozbv32DcZLjJ+rw3d4zIEeMgLk6QXEL9QU2mhSzXBAlfhMkPHpKZ0HtyBSeDlkFXoeExH+vYBjOZuV55PFlXePufrTjl9m+/0NyGIxHre+bHo2UN3uqboNIWDo7ONvn+B4Qq3qzU96rIQYp5EZW9EiJ4uGBd0tbd8/HLyFLhdbkze1kYb4tcgkOInJ+Id9t9jjj8bXBlwyf6qoCEBi7UIZC6OBsKT+MY9u4bK+xp4Dyz2gl1xpYzZFkQzTURmJWFhZgGzWrB3nyRFtZkBjTxrZ3WOd1TFjrZXSqSQWcCzF06pOLZj+moROxf97GiOqeLrC1upmSoOtYxiYbsuoIj2FbAu1gOscPDRRSp8qTwwfpmf0Rtl6Wqf92cwthA3zbTReE1UpRIZToxmDIIq/JcIW80eX1kqZLxWvBSoEWdLwERt3Qh1BfFwco8HeuI4O3oqoULx2xalW38D2F3Z27pbL+eFlNweZZs9+KTGlU3feO21wufxZaMhsMgJYbwvTBhfVMp4PTcJK89OwG6gPcG70YBSS8+L2QIogUA49iZrr2F0cOR8Gah4HSXhgXhUpZmYN7+s3fxMuZ6ZUJfuapa01aTM/jS6a9YL6L41hihYM2UQFgALFdKW9CjmbFsLuoLs4DMH/Bubi0Xv04Z2Usp7Fkz9ttwkYItGvLk2P36flSAmK2wk6LBHT486tOJnYITpn5Wijf0RMDeh/zApuISMgnDTmPYi5ziVWuHdWfMQm5FhuvR/MNaGeJbiIzARL24Ud892gHhX9DdMtQ58SvxuqDzjGHaLb2Sd0/cyOGbJcavmuMt/PQGCfjUiMS5gm85/RH6ZA+Eu15+RGHaxcT7nNabs3aUbn3cbMdkSSV/8myGO/ICpO49vYgPcMAue4iIkJxZZaflHJiZTs+0KJhuM74Ydz+vy3ChnIBV4nL6tbaJyw7gBJ7Z2OhA8gBnJt5o8gw/GwyQ5tG60CKu3xTJmQ0XnhTk+JOmSiXaWfEUxPZcW27aUsawOFa0hzXhT8T6dS1KhzxmfsWV5wcawV2XCEX8ziLb0cjrMa8MiXhUUuHFOfuHYLlQussKo58om1PXWqcuAJs0UnnTveJ4+efYyz6UOwvrlM1s0Fy0XJG9N1WN5sjcAXFq7BPSb4KXYn5pARgvff5ebSL1rtCPfuF2XQNp+2JqfwIPM5TsUtSNvYI9P5atxpC+jlwhKSAPuTQOCbY6xlK2bZcXRG1zwEUIRzGKL8tO1dDc42eFV3H6lRpafDdEw0psSk860VrHtOyH+vMxV+pdMfIPt4jd5FusTFzhOLwuJ1kF+JImpb6baay121vVjeSSLAwKU/lLc1YG3ZXWvAkRfDJKN8gGos9YD5pNMroARrv4/7tM+dwMdP3CTyDfdA3nx2lCIU10yi7icN/DrAr45RpUGHvpWoqh1+MnhFwjWh40r+PuxZmKbZC4IFW98PFHxdnQIaUH4XxHxnMpJKnuQIG7yWnr+LH+NzrEo2uZfV2xlq3QGoNRanUgVXUSqVEOCW1+BtdVlUzCMA4/pUl3C+FYmCWMFjxqCk1web+elceybcdAD2eIfhM6ZUekyVQuLPVxOqutiSDVHQA0DOdCvDgBDr8/zhCMts4EZjo4/kjjVU/uSCjJjn0VpDvnSybUiPoDclD6CyF6an38+goLUbZXwnG87KCIPSeuWxqunnOufZalEt453DPdILoVAU0AIJzPU4MNOB7IBDirekydNJfTKW67YRSX7GTPDGgR84I2MXRMiitcLHlc9iTiA3y3843zudONgftUrUqZzD7p/0PJjq+zEWiP+Y9BTdoXwGcE0yN3RhrbORxPHjCYnnFdF8rAhC2YcqHwNjvOum3IJMd0ZV+lkBPK0ERS/5zxHHguV+1e3oGx1XB8Yo+i12i2D46lOmx74+pNYAUih89QBpcGaE2cYYa3QgXpbH1mEihvnITeqV+QoCaqZfz3HKWyw5tlD224V3bwvUeMFPFRARELiSU/ylXbfjUd2pR7lfAd7XUPkqMgjmeHRQHrFDs/jHEzzw+CIZaCMTxwpbVuWhnbCBtcVsN/9Y9wNr//WLtzYch88E3OfvRjonps3Iq95d1q0uJ7f/NLAaXkKHFrXas9OKhXwpzfIWBbBvU/ec0Bt5bNXxw6sa8Uc5ojMfgu8z1wcws4RNmkrPV2ygd/T+MGhIBMV2L58Ak57itnMrzuv9yTwKxlBYkimRFuxSae4D0xX8GHrARt2n7iHrRtOxJYAlQMYA+FOyiAPdKIHMQEtacWqv9G1TqI5xosK6slw/imPVLDQJ3dw9Yjdyd6Z9EvS/eSjFBDqP8fQvDwMygeMIPZek+TGTcuIXwIdqHSWSAuevC6lwZKhnswEzDXViB8U7FBHxLKtsqZcFDPU5862oyLDUYJCnRVWUH6qIhLp6crJmz+TW9avOi1QDW4edww0QgZn4gbjyHIwh2SQQWo2ggO+RWX5uCJlMNF77q30enPeJjxIcdjWVBHsHzVVjSgYcVQI384sBDbcLQsjGAnvlvKM/T6jOX2rzkrqM3el7DjLsbVsVFakJp5eXyTYENJ0Tnp3RMiLmuxFwLZiNkQuddvN1vlYQP4rv6DQFKWz4BSL2F5imoeQ3uv8p9kVrXOOrkmDl+ZtL3C/2uD4syx6TZL99425bZmcHZNskLaarZBGx3xP8Haq3Lb1XwKv4Z2InBtuFyF//63LSUm+2Gi8G4JR1csP046Kkm3bHQf+JY2o5vESW4RJZetrJbdBLSLoHmU2tGP5nl7jo3JeVi6ay/DRZ5y1SBRt0Zp8+rrFvuDhd+K38/6J9KAOfaF/T6lmQY5kPijZ5HBErtU+FPI+yaEey3kItifnijWcPxqVq04lNr1zChaGIlIgemAM0UQrmY7YzLoeFmAD+QCkmH/9FgEVR71gpWPyjxRNLZWACmq0UZeEphp+D3KUyyqxHvLPeI6BeCJRKDwYKWGyLcnHktSbKVAgZENw8dQvJk+5Hc8J292iMY8zdlQgxAaWzKVJSCErBmvXYJ1Euso3JvSdIjxwOnXSpu3wLCBlaup3oQcjwS1M/DqLwNS8J8BSAo2qxY1mHJarLWrE4Ck+OcoahPhadTpd32KhDsJNiTHqAx70xMU53+z6r9tznWrVK0hqkT8czIpBGDSEOgZHjK7HtFHitDpvMe+2028vlureBVqMGjXCjn95pgaImqf7k3LL6Sx79krWyiBZjDOZ65gk9q84NJ6+Ip02Sw9ZjJYDry6NPRNumY96IH9l1sF19hz2hCe8swKb+Kqw0MCeAcow5DD1Hvyuc2psgS4gujDp1e/aFmYNo0JJqiWYuus8RXzOnC3SgrPCLtcTBXi8/Fpr1EVuAmdOqUSiUAzgbBpjqvMmwxNKI3Sci0PVo7hMvsn5f8WRRm4Edp4SxDjoKPLl5U8KmGBuW48q71ZN+yhabuVY3WjhCWKiDKUV6S9WEH1rc+qGI1SGmxQO/qnM5ZZtOZSowZpPRKvVXwmALglnnCJJFUr3Nf14/EW8nT8++zk2B2a24tezmJRhkLSeqz0P1dIcV2iwdKL14LmWLxDszyRTcvsCHjURdQaSSVLG5Yg0al4Ajfj48A+HrTFEmBUjYdKVINlcT2R9xf2eiozZuwMRZ6ukOH4xM+7PBop0ITJZDvTUsEivrDOi5UbbNeEJvLOu8t/x5rwOxVREFVcQzTRBkWy1vj+Ff4RTiJtiCm5G/m4XWgqI3sFOpZ2nDvZgsbTYG7sv/Elb7ui0nJiL7vflqCvm3J67BjOAaAMrlb9sIwp4CUq6cg7iUUpk0m1GzNCY1FJa+Jkoe2yF1zKlNPPSWEyVmLCoEZL7V6QqsFUU/g28LefYblqvIBe1Iofs6y6SC6pU/wdF5ho+ZT+S3oRS+bS55zREc/m1oD0dTECZcCDnIo1FQ7O+v/XyU+clAbHU08Dv5XQ50vcQzUcV5pDjFV8/JShPFtFzfjZ77mzEoUtZQOSu9LO4V2vKqDux6T7xLepSf3Xu7bZYu/ctriOw3te3cfATclNk+ISFiXrXLR/pbiwZ5HMavEVD67MKwcrhokF9nAE7r8KMYqT5ssajNaDFaGP6eeYt74zmS3LO7V+A603PoFxtx5h++DgtcMkGhhmuGa6NmkBIPWBzsthIqVoCbNS4yXNKuR5sHsDwkUce4dL6GCZLt73EshNOdcL7eUGrdRNQBpdMVtT8wgxUdm8T7Axw5chHtEH+xe9vpJwgpF9IsDuXYd5aNm+hygufLOZe/hC99+nGoOFzbpRLxeEBTi6fftpSjj1DyqJLJaqeF9ILLoz7hgy5SmWSAPr5RZmjfHfQPFu/1atut8JvCW44cVNBlaJ/1SiJY2NZmI71h+3KW37dH6piJ/wNfnccleHH/9dGHcfCsNg9rbasZ5JGuVpYi/ED56uXbccd1wv4Lmu+eHifQVIjYgHS/kdZjsWNBj9duP7e8JTRqEwQ8LzaZPHju9Nt7CGOJ2jdV+D8hb99P4syxe5DMTm/TQ2uD+W6mQ0Sl+hXHRei57GBayJmKeJKjLx88jkDLNiJmQ5T1OGXNRCuN7BVsnB0z4PwHfTsZHkeL2nAnhs6DDBlsGty3buWK0PTK+ssO2+D4sIrNQQk04wROxM1PvdwdIyYtqQ96n+q7CrbWrYxd5xNXPZnEk6ABntKHLncNshRzCz5EVF06fM+/N8jiZ//Z99K1o6e8sZXmR1Q00K9PZwCuA1z8VhuxrU+5vHygtPeiJVO4n3DDQIg9jnmI88l0QaVZx+kI9hjqXMzJinWiQyjiAiOI2RUoFGeiPqNmFjBjLsWubYF80MAsKBy11qFVaIUPn00ARQ94rGdC70ShMRXk9UF0QSMpli+q/KSC4eHK8nq3OOF0hbLJP+cZ5tSYxpSiyyEKKJccp/pMfuS14cRXH8SDO82vaUyxlBwJqm1J/9J1t2usLLRfKl4w5dz53xQbhIOIQFm/5Y7bai6vyeEdmskUaIEsUoBt76Wbb0qPiicOjMmtLODsYUwnHFpHOBlGoWKJvBJimhrNNLuMvkF4gPE4M3iVobUTElTJuntMAKK1N4ETY9bCyPXaE/VBqAYYVGiA/Fr3CgpVIHNBtjUvr+nCqiTOyB7q/8rc7lotd60kdvJmlQzb3horXdyl4F5uy5UTWLhcL0h7Jz/YPZR7fDBMFblcNBgXbr5cbBhbNF6KoVQSLqM3/EIxzwUgF1wGlNDAQPzshc9OW+1LF5NGUn20eNgZPXDwgikXQbm7hPe/UWb+gmoHTIVa/PCvnRNdsee1b7NrXr0WSrbcw6fRwi4DpEflRVoDaZgCk+TsCz9ZrIUmZ4pAo+U27uPgx3ZUbs0YiIFrZ9I4nSBXbkuCTi3cenT9MM0xa9yEVrNoHT4a9m7anMnSavQZG3eTLtxObV4FPp24T3lf8+9gM0ByfNmS4PB+sGCDhRKgKmumZ6y1guXIUCM7SYFXYgEZxVK0OMaJ6BYbaBC1CzAMgoRm/tmgJVseHSGg2dCpRM63IEoy7SJfR11qCMe8V8Q6tjAjscQssDw1WgYufLPSPWLt2Sc3lGZG6cJiQXj5lLIEnAFBIfMN0BMyXrJJVfd4sgDB848pkvfs/MS1E1Kzr1XGcCKNcc/i4TOZdmr9N07IcdybJVH/uNtjoy0PSEpKLiw6lNHsYkWdkNpVNwP50/4mwUSE++r8uznXgjrMKkOeoTPDK/5AzHzPNYQSo3Va/tvnGjmubE47M3gqmv04P88eyQjBnZYGnsqZnks/BfNMxASVxvk1z5U9ftfP5jmXHplLwOJHpNE8udiNjWkoUD3TjEsqON6yui3zaslLh+5UXWro2EvcXNRPwXB1K0kWLMlaVZ0oXr+jFKqulUGVfIX4qjOMh1S7YQDd/yHvzSFO3dBPDVe/syzzKAmcJg5UqwB2ifFkKtLvaB1UhfZfQpYq3FjDxwF8JOgPu+iQV8JOBBVGpVOmM1C5LyA1JJQbwFbhIiwjeTh4pM7vNTInbIYkXs/iMjE6bdS6hJErQe7FFFfnP1nGmtnyiXsUOV6itMHFYA+E45qgdA8AN48PPvNTSWoqOoWmrq9aRl1aSnOTvuSHKfan621vSksMK8BO5nqcxKs0AfF9hMiZr47O0/jRXNfZUU0yLiG5VNYi/QJcFNxTPjcT/NuS+o+fkJFA9CwAyWJisEcTo8s7fY0w544cdYGW3GpyGq+nZxVo2Z5zOR8AHaumfNhbNy3Nb7/fmOOgwhX+GDdKY/kyzPvv+a2mye2WM+hpe7B1DzaRpY0wcXryCuiVU8FAxEB7NKZHxK6XDn5rdNgjMk/x22nl/+kyQZcjEN7uiYi34dteDMkmJuq93a/F1/qobDDN0CPYVg897ioEm5ecqhQU0ijkRrg7KyYvx3qetzoOtm0izCFLkdo1x7EfqHQ1wz8IdJLoy0qZkt/SOAv9wx7l5kxryoMDYiLvS2hIgIOmwuY/mGe4BS8lUn1ooGZV4pBYgIktwhUXT+Zh1T3T0SzAyXRJv76vCVeiaC7Lqy5IcvCQF0CDeLCQx8VHtS7ACrHdihFfdWk9xKZgW40jMp4ilLMGOIEcJ9hb24MGaNBxgzBkhY8tnfOToAYSrrQQERfp6I1LJW8U6vq0OP2/bWC5bf0JYsdYAGHWhRic82btoMq7hZvsrM3W2Z8LgC2rVATQ1AZ4ITw3V/U0ImKfA+4xFq/w2EaNtKAhNlovaQeq+XZjU/3aP0Rn8zQRLuV1z3QbMhi2f6ju41q5atGYo8L0GR+TQuH7qtratzXj7ve84g+VWSoi4EMJpDVJQHG0ORyzGs08pVQciYNDv5db4qHm0GSG6wsI2UV6SGafsA5AU5bMNDcsCFcKEeq+CTKLYaGm8LOYQInt7irE/PSff1xg36ItmMkh3b6tJUz77THM+SQfUOrc6cr0tRMLAWyNW+SW8x4tRo7bPbfdFK41rVM0EhYT56pmR3pVMNbkRJuNUseM0Co3j3hL7eTiaOgkNRwJCA/01oiyfJKrX1dDamGAvurxbMdMNCEHg33NCufBGK34rQl8YosLG4DJtwBIRq8ZjALiNOlZBtVPV6RVcH36jRv1p18eCrqfVP/p0Jh+NhsXOOVf/00hMSmU0+OgV73IvXiz2TLh3s59h9XlfAGabOQtMpZuj2mmc1oy5Q37uAtcf939vdXbsAm3mZfroCkbdSGiqtKc9qk7qeU7+t2s3SqlPljvmP4MnUvtov9DBt2qvpMKihkmsrpuSxzPU71HJxsmVK9ZGrcQY4m+aKaj5JcUQfK5BUM7ik1NXNqdwmBC5vuk73ntegqyu7/1VuktAa97IoDc3DjgsTM6RxOKzGY2QzyA7nDT12HbY/VMwFkW8D7+herKujccayvb+C5G+voX2U7aBBm+NGsa60UyGbqM4uShYOel3xwiVSCMURcJH7Qzv1pq5LkTh4VcpXT4HSSv/lBD2lDJUm68A3yEd+zX8rRBBU8H7Rp5eDc+qITy8TQT8w63yHXw304YIAikoAW9u8/oupZK2mOoNhA1LiGTr5PUuelaQK8PWI7DbdhZNigtk5DkOTy80ylQmhEkbqrJC557dP7RnlLOyLp+dfOzSWOl7gYcd6HpRBzr+TDPMfDnWftXHhUKqMoEHQgqcxegflkzqnOOO5MZlKogdm31QpGbRJO2VvG6O2gBNuA0R1rj+ejLU8LnJK2fsX6fcp8hdGhLNCETjAYOP800QgnIaLhApKg7SUg8v04px+1QYJx2l45zeMVOZBEAoFX7uLhvDlw69zmS9sY6Hd81Nh+IVKEsFTLtFGMx+xZLLWC7hp7j3XJi4D0U4qWQivxsd9O1GfJ0ZjTO3VQBL19ZDtiXcE+WYq99wVVoIdhWM5Sk09xrEWahRpdS7baPoIzgkBXQJYVng2hb86gsQdNGFRkOvHDBwNEChOp9QlvpvbO8km2+HT55UMd6a2E+Ze9djIzNR1xTWBKG2I7D7TOBKUA4RAw5JTGZy7TQ/kZue+fDwkK1dp8x/2Eq8EpA8qQNtTfLxEDHkdO4+UMmQQ0pvYKit4xDYbUNsQh5cHJ5RFLMg+1tQvzTa3re3yxLxQx3Wlk8Biz87jdFTbdxJQSbro6bA8EjWViwHdEROGvJTxMkhWBsiteaLrvAVmxyGUY8V5f+iPIGMQfU6nEmTaDEdNx4cU4uej0R46wz6cW29wRfWSYZ0TJrLKhGuyWimhcwYMS6x851xZVCi9Nv5CoA42grJJQF7j7dFs3PmlkPrkaZi0XHhaE0ucoMdfrw5DQE00g60IV65GIqIWML3huozC8U5fhbwAvVNB9eq3kfEV40CWsw3a9AF8QWWL2XgYAaBc2gO4nLHKXEnSyKjX5dAQPjH4UhE0NqQW2FxYSz4Q3EPDgy/AV/bNNS7iYG0/obOtlCqHoHQW//Z3K2gqKbdCYA7PAjNY6iUY2pbJfKLxTrc+G/8M8NvGipy2GoS3taY+1rSITs82bLrWXZLfLuLNWnBFgnvAg6/uTo8isssnA+gfwMpCc9EqWCS69DkbWeirwe4XPKcOpfx+QTodzSvWQQfYuW6HYq2gKIVwBAG5U1rbR3+SY77LaLnthiv2J5641Yb/gkd6vxyWWIP9Xnp+jXQ9yC9RqTDTZM926rY6dhd8Oo6hwOf/snQSLhJWs+SxUHyDI+r5HlmFeOuiZNsnZUZlnUa1jK0mgAHb7UvLFInP8Oy8eREOBzmfGjfeDutHTWUTSBf1L8UwnHnqwD/HsKHVSZUIAOr9y6RknYF1TCbuuF9vob9YKjrw5BjqHURJBrCa+inz4J/i1wgs3pCsRkme3h9CpRr0HCdOpFzKo010AQajIAJpBwztvurgYa4t/D+ldZ7p612/K4eDOcUvPNCClK1jycPtjVske3ySv31QX7rKl+UqJ77BgiE1kTBeOVczIjLarIQAz34dO/s0xTtBHIzZF/SA6JPXwGkZqn/OCWxV6P5GIZs4HSDeexG5MlOW7XvgHVC+q36PpmM3VF6kTBn7lkKfHW7lZyOI5ca7YSIzGQ9gYBsxDWc77EW2izQGROgzFZ7nJpS/Ph60M8O4MzZ1+bvGSLbcOSZz6X1uDqr60dR8Vi2Y4coVglR/vMhUnxdFX3p9pfaFdQwcukXzK+DWStcMsRoHPaXSQslvJ2TOnhje1A6ajPn77R7lI4XqKyQijKWZd9a9IETD4MdQABEEBIO/9DUcC5SlysxFpiTMZV9DPHEaL/RBhoC3ZoLhCCWPgo/v9e0EWUhGwCXBUCOFICLhahKD/GCu7k0i7jGNT6S+5YcIsotzI7IoXshCbiX//5KLmM9CZK1q1Fb6xjP7Op+aFhrAQEn/XDzINkdgSoDMiiAZCBNRoqH2xir5zT3VlTt+4blv5qYqBkMdEMxc/kAxdVQiqXIVBbjuxXFe2fM4mrBVsqhYQqsfAlPiiX2A3SabNs0J34yD+0gzqlG86yMnuYLjuDk3ipmqg/9tkNkZefXw9QvIhSRoReJY6vxEIUX16EBe75TnW0uiZxZuFDA2Io/ioTsfO5BXpJaYj1sLWY2FXVnlJG0smdcliTlDIabLxQhHJaF2elLB8XHv8ZARSirJGi47UmBFKV40t5EGmBjnMkTVXdpqkVUt81+oJ73HUYcBTkIipL7+QB32pogmLGStnfolv5mHxr20UvrgOtvHJSsR/QVbbYwUtP3xc75c7Qhuge6FIB3DkHXCRCs0UACkBpAkKjC9agOFWNBbytUkNvzZSVSX+02a4oq6gtDMqYTZ9ttbK5xu8wcX7Hw0X6oKUnLRNtkO18zm8XyDOxb7ayYaUhqb4BOtCx/akdXRJ1EPrWGfoisJCthXowEEbYjYxset5hSKAxj6aMMn3VAQ/8fGQi1u/tlJ2U0R5dx2cvruLP4Qb3zr3cGatTMmh79Myh9Yp7WTH9yHGXG0ffCRZxZ+J/qvgNo7uF8jxGxqCIJHJX/MYlFEv8XlRRkhnJhouiw/QUR6LvjNjszzk2xdBz36FxqMdKjLli8ptRbclqHCkZIT8FEcj5ACRlwtdund3i9BSxJ0q93YhekQ/zTwUYhvOBE8k/MSQ1mLh2N1nedPBVVA2syTYsNgCHIKYbllRdZRoFP7JS6vN2myqLMiWu3AKvkg4CE3Je20RhX3Xf6nBzUGm6NMBKukbWSVVwxCG3/9BJY6SlH3u/WDMOMwGp2ZTEBtoTvcxMmfp6O7q2bgGKt2uVgc8D70QT5rQlcm5cRLmHqIw12YpTR0m0yTvC/b6VzhgdSRw8/XuM4U3+MLZpgllfkriCf0SW8DGNRFbD3rfTBqW8UmYWXrzmowE+6/AyHa5ctM7y5Z0aSSfY3LUJJhfyOSYXW9TYjxVxshESDqJ9ANPcsBhpVHN4V+nijD2bYlR84KSf75f7hMAJKmNif8ZxfE/G1reKO68mNkX1efgpcKZlPyf41uhFEk5cm4zfh2MnSOOwrFx9HvEZ8UjBfvdfrp/BdItsRV+Go6Eb3TjtQGiuXvGgY6dfdAAGh9q6+2j194UVkN5huRguGwoaYVPJhuDoTW1o4JZimBWFRklyDnnxWaFPRBDlrYd18FKgevIc3oiZbIvVqvyZv2wcSw3NBWDLmfxSkkIFzqbAprOchvKnbC0Ld21Dc/fram0AR3xe+K2axOB4j7BJsZ63yVY8lWWhtbUQcI6llkv0fZON7/j3iUiaJqI1vjz8QTamGhujFHsrLcOfPzWiAH+4AQ2Cl0IlaoUM2/GrvKtSnurg/0TF+V5XH8/5fYt2T1iz9Yf/fMkAU7HNoi2JADzWZJvPoggNhSdxBBZI6gn4HBNEwgyioBtC+fwwByVSYt2wS2LZ4GWeGv0U6oTrh+SCIWVMox0APv/CyfJ5otrurlbcwPTtbnyvM9RTcBKFmj/I5pX9zot2NCAedwzcbQDUW9WGXWhKRvkL5QiZA2S99KmqG9sUyPQQ7DI//NSw4azIaQDhEEit0vs7L28VF0/X7O1H/z3ez/yV/5IEhGfUBuCIlfrlWiZCDGuViJRRXrbjB52YJ9H84kUGOivoKP59E+252Ll/cXsJQ0z+MqQC7yXzqnVcL4BuzsqUb5tTjMMVd6evpsZISsMlKgZqI7TJ3VCyiUQqfwtLGdir0DeKuHJa0fKDvhJ9mzsVDyN8YYphKKfu6m51yU6Tu3sivCU5HlG03R6q7DUosKugmpSeLQ4/Fkevx9BF1f8cVzcUoiFJ7CcJUwZf5E0E2k5/2+4I11VuSpWKJyDsT30WmLc+MWiHKSufipeDrOUnuraVr1k376ylbr9JVtMCtfY4m0xSTDApSEhTGjJJnDTuQwdlflfy7g+HYBUSltWhfn70ATTj55NUuz5rAY0UO7SCkqoKoQe5N1hTizLhE7PXOll5uZWfLA7SPXraUngubfy9JkHZb36g4GtK9BpUgb0H05t+xvwnVS747QkhE4uLmcTeiJWLzBtEX6SBrhrASSaFO3upE8lpt8/HmWbKiq1T1L3bKFEl5rDUBvIW6cu69gPn78lfUeOcgzVzriDTF/ay499lABoPdSf/ZTKtgPu2L2fztcruXUm4yK7sm57Uv+jTRTKZQ72bG5g+BgIMVaTu6Bxd88vZqxqwunCXPKkWATaMWXvJeBxCAfPiTs0qsZpaXbNFkPO4edIDGmQGDSGYUUYGII+SYK/CXztES3nTXEIDQAx4iJRsWSOJlSFQ3jmc7k+iuCwrx4iwdCvtDzhTSOOYiWmXOIfE7CO/0V7lxWDutuNePcvqjrJaIM4PSmQjv3y/yQvuvHddlNiM3KK//a+Enj3L3y5FHpILRO9pAl9XLFrbBIuWs2Ke/2qjbZrz2LLWeNsJ2y10JiXbXcfh4ALQwhK4ZxRxoAA3swK0n5c5pQNdcCRlmio/FFfQ2cpuiIeCyI94aRmIWrs9IvNSrDn1czXQ3IUuSLx4VSGLHJ3iFT+P/f+2g=
`pragma protect end_data_block
`pragma protect digest_block
6ff55936a0579c35dcae2ebbaa8e171f574d3333b3feecd846d7ee1987506a40
`pragma protect end_digest_block
`pragma protect end_protected
