`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
f+lOCsRi7rucy3vnlEizV9Q4gF8aJajBd1NVDW2zylVHmZ/A0oSDpvl42qKa7e1CW09RAe4g5tSJVkW4F0p9vRu2yiR0zosRrTGUna2YbplO3GpMV0txcQBiWOJn2H3tJSkAuhXQWduxeVHhWi1rx3h2/1Zchzb700bIAHSqQkLLKaScV1gQXf6OYoUODD8K8iFGZtVKWnfl9RGMWQUs4JkowhzVwbEUbBkskbrgUunP97G99lC6Qloa+Ktr4pDogEffsEwgbTRV+I0lkdydK0jipZ7MJ+AmvcWYcOg0xBZEGBUoSXFqy1nFPJUlJCkcY7oFclHz3o62jR7cOAdzl5WbjK6SUpLbRS2tCpm+p9H5GmUy4tHjEqq80SMLbYb+bqIJVVugpsiPrTRP7VGo5Vl/XGfMRwghh/BmGOxXfraxi2XwDGtgvu1T1K6KQuTbvo+i8IGtsREDIaF0sqRdGn2P49l1foybAF/xzAqFj4/s9/a9rHS+E3VQZs+dk7tZIGtLlCzobfkjhuheKm7/8YgyDiGgEhPlRjDt10c2sawlUK2EjtQUMINJGumIx5kzJOoF4Ecfb6MIOXy2UvPRJ2R/B/nl7B3GmUnpuY+SUFOCurxqTcdKnsxf4nSGlwkH2qV2gJzzFuOnufQHXay8Eml+ySg7CGJjkLjPCBhj5LkifRyoqxd3Lpp1tsKp4afimqU5f3az8l4cR3W1AobWxqhKp+58qjAaaMRPhbvCtZIMk67Z35I3QAnlKdAaWTJIvZlEO3vKj/WjR69kVP9O/GERgfW72WB1ypH9qd2feLuGE9epEyJnd3R2g67kIvHgufnBAjbUHDwvFBZRXElSn7Q8UvrALf5pAFCJfY1eWr37SgShesXYl0HFKcMdu/seFcnA5mJvlIQdPTWAJn+UNNdXtihuQwPL5gc09JiFzaUrl/lcjUCnRRa3YAp/tZnGPdlDEmMpDsygB8dODI8eVR8gr2L1aUKAIpWSH/iLli3UCNZIhX5RoyJ9Xz5u1xKigBA6LKsHTmAJKNQkN8/kknNLY794+K54iBJ16+at6SwTyzY2BYoGgQgcBsiZvb4R+jYfF2OF56jj6afLtMn3VzHEAayH0CQ1YU7smwgQF8DON/k2CU7SlBISBRi+CMjg5ws0QK+VicAVWbsNvHPOz4brB2Z7evVpP+LxpRvKWwlYF57+csk0L2wHtNF4Mi+EtqYs5unSv0YYrLhOWpyd9+0ChDq6EQRFARXTS7mgNN9Kn17hQIGU/cEm8pBPzxirPfjXIv+vBrp9yoCP8GBe9Pv+/3sAZg/LkX2BUU1BTYql2BhohedA+dNbWe9gI5y9V17fre/7pEUgAu1vKRj+LtND15kB4wm2qBCqnVISHqG1SQwecDk4C2QGi+nm04riiLCxQYQCHL8eQYVfk8Pma7ih5+dd5Ektt4c6gjYSEMTDb0u2pdOR1z3Nfwr0Lx1O7e6Q9y+P+CPYWEiUFXH/RZbP0C7Xs+tAxIWA1JqcERZo6C2fssfbsU3ONLBPNt571ZYzHrWm80PAMVQFAxVxKC9TYKqYgceLTXmlyERQcAMw6GfBprl2hAz+kuXC7HlIrEliiw1/ZvAN95UlNZ7Ek/TQmBly2s5UM/1YcSqjFJMweyocwJWywbTaiAfyqgd4Z0dCJHp4Khr0G8qwc31NruXjg4A2IhEgIT29BGcfY+mOCuXqwgTmxmjWiG6aBK7VxZjUy0tLDiVCbkQv8f4ZX5BbwXcmIWoojvs2Df0PmnOSrwcq6B0dPtE9smNck/JxtpVBxPXMyHN4TjjMbIKDgeNxvc9xx7vvS7GdVIxHUchTAYX2yyQJForzDRfLlVPl3iSB8tYwBBiC3edrkuFqzQlBqdVUQ2mlCCMdziwrhkhxrQwSXvMgcmNmoncvqKupq8nGh2dI4VuiB5F9nQmHppJayS2jPxxTWFzKfWwXcclGR30bEBOqFovzmPPNgqRc2a2Mz6GIKrPXzoDQTbANq+b1FXs1tpfNyWQSlW53gzUZ6Wd5DdcQtmLAqbh7+OtKEhSaPNS2e0Z8nlMY8Q0eAphsTNoz/zH09Fum41XR9D5DxNKrcyUqwP4ItW9Ekhd+4AjzpZ6XIfF294IKNft1n7oeACeFgJ34YEm36rLE7hLbFsvC1prsFosieC6RnbxohDgqgy57bXFu5YC7eewsaypuEvJg63dup+FZbotuG6hnbzwOikfLV8ZLoYjul4PDkZLMsCzAZJ5cZ1N3+oO2IrTFH1qvwAo/sw7Mgzn4tHmcjVYEoBhIYOAWh2VEM1SpaWQxayClqEB9vqeka9drYANOyb+XyS/vgpKfY1JFeld1Mo/pPsHMCgtJS6+BJUWFmE1PZ/LbUFUKe41WT97Jfg3pqd8DL8240t5uDVkWK182yUUBFbSTK0+PsVMzNVUC24KgoODWqYr2nagG2SFAkJJUGIm4JS9a7Q6F/JbMpYc1Xk/36kZv5nvUdA4ars2xjW1VDjbB0rox15q89g4K7hDA+04fGHTRfhqQSXny4W8aA0+/7urgpnUKPQJr1poPSFbTu9fjIPgD+7XeX6qOMwwZs4fm6Ld7IBLa9t8BewQwuOJSKhYj1mViyA8dOCAWVCN7Cqg/KYvx6vxqYogZz0o4+u7wmPlYUZTjPl8J1G+4P8M7Su4uQ9LmGBGHtsXJAaWrwMKwvmN+1ed+FtNm8kxScZbXD07HQPyoXa7rDDDUz9udbbRllazceI4a5CtwOD7ahFbSF7hYV/87g72efs+Gshsub2ZXIt9MHJEFZoUczUxIjKU3pienU+TiJ9Uj+9BswY3B9Y48xLS/Xt6PBGLHouVAYMCxmygXz/nMPCyxBub8zMTzCnpcaRHaRZBRagCgw7kPwQcwKlQQ6OaNwRH0bFo1tX6Sh41dKUykSLcd98cAY82WD8HG2StFhaU7nX3uGgyNX2aU1h3k3hyB9SdO7faaBPgSY3OV7lfDfvusixAOyVPa3/oWlGnmuXDhsnaJZDyLBxCkEKcurDZ+LXsdTJ9odtC4mvy2ziT9AFVTWaHRDgWmNghgNlVLWfc+jniUwOULinIU8yEF65ymn2pexvTQ43k7Q0z8NuYcwXOlinyMMF2PC9T0D1lpHCxLGXlQmQlQ4EvQkhC5+Av3UcJcWmXQ8W1no6PcBoiBhopCsE4RPfFC1y6t5+iwheKxDpgQnE0/y9kKtCY4utrmXk1Fbu08vv1hCdRnZnKCEGuOvyoclDYPCziocDTki7d7dQTmjlHy6QZV4B2/0mVOIhV8FhNGNCUO22O1NO48nax+G9xha1fcx3tGGTEnd8zgJdsF3sylY2gpLzkKtLIDhFm37ngu9rFu5nur+iZ8ccQCetqrGOlM3N9EFflEQgNKOWEXwPvzEHUihM1O6EOHxGGLEZovixEoqKR8yrd2rMiRKzkDDmjCH7UL5UGIwoJhOI15y/+FezS3r16n6Bl29BZuJbuuP3ZfRqEHjyAHAiLfpUN7qJXDxieURpgx2TwoSz1jHuBI2wblw2I8s0+2tV0CILi9FsDr7C6pTqit1OlWHFwjL1Li3vPR5E34pk2wzEMx960CNqz+AjEkDYkrE/0gofS5hbzMb+qbR3tdgkN7CglKSa2nu7EZfJ+Hcb+kJos2yA3ZHmM1KNimOLZ/2SpZahSdLsokLlqcKsyPwQkXpM9zsam97yOQ2tw7GMMfU71vFUL9Z8AkX+dW1kiH7B0tcu1Y8gg4VPUNbUwjfHX30i4iw+/J/Sh2BJtuDbHIbQvFwgJcTvi21tHHuPUf9pGzR+rY3aO3CXwlzmJwUx7nsAwzGau5K4BckuYb/gp30Ia23RNuTc9VNerLWjcAHkkaG26Cb6xmkWs7bSBxYbflPMVx1bvGWim/ZavxFSCqIJI960en+EW+hPOpxAIeGapUxsj9qC57Lnsk3u62IkUVnOVJACqCEqkqsFtU9fCJ/9TiyXpWiA8U0iZ3d8j1swKJo3xIBmNGuOOA6gXpjqfPIJREOPm9ZC1SlepvNtdp8ZjbNgGwz1Pi2Y3SInob09B3eAZxCOv1lUOo8GNfwghT+pXWUNRFD3xrbpXK6IZjriZPHh3Kb40ZbcF6Rfy31wqPnbzP/NpOv2Q8hAaG4IZ/yekxzoKKGDjOOHt3E1c9LtprQp50NQE7Xc2nMU3obHpje9LYnLzH4AW5JPZLYMlAlPWlVN15Ow/Hbm+GsesAK9MKCR10Ujy8PqEfRsZxsQLSHcJF3Yo4+g7D9cZsi5P2UWRqt6YxiaAdJ4iw5SCwWPRRjnspaaQBNPCubYEByX0o/BGtHPdlOnaQf/hA7Mz3FubYIfn0Zji5kcUi++FgBXBDOa9At1MRSzvP1r7CFr1nScoIGrbFzCWulRr37oboRZjOKO6Q5FQob5X/6rEI4rWgUXcE0MUsCsx+L7T8URzjAIvvTcYLlsdfdPPsKcIkeCXM1wEPhrdogUqaWy/ioCI3D0DHG8ZNFTLICrGB/Vbkjuq03QsTuSNPz6IuBXO3Xsl3GHTusvHJekr1ILJLsb43m5ua5WPyMsfnvKJB+NUlVed5qS59RbGNg3CzzmIjv1gitSRG7NqKaQSaGupqGGZVFaS2QxkftfZUwZ0aKpeP8I7d1MO7dMZWWsEb0/uXonhBHcn/6GNyE8DpuomheQeaeP/YnZOoBEKldoDkQA4ip23sq+qjwum7t0d4ZVejkcnjBLc+VuK4/CKOE6flkEsJRSG+TKL7oSJ3wuR0P0klNxeJb6DnC9JzRoD67Ksxpz+3U/FTrVrlJhwKpgLU+5loroOAB13SHcogClg0bxWgxt9ym89Ti+X93zd8yqHvWpwA2/5k1QsvkpLvYvhoD+6gA2exBxC1uA83ejt6LUj4N5az2BI8XqobIfp51Wze7vb3s3NfLg5MSjLSYPS7mB570tvy9IcyL/CAe6i07zkMNVSzcE97EzWT7Un10RmRIi3doclcka9XbeeEHj3Pl3zghlXAsNREZv3xrG2quL6P1Yw845wZCmFPnypffSYmkK8TnWuisgWfoVBJkl3JrIyqKhVedp3GKv+s0nkLoH+T4RRq4X+vK/eHH5p9oe9w1fJtNeZVA6WICFmOV7MWU9LmPEBZvaSqznsJsQJU5nhVjKdgAzuukXpVDmMx/+d/rLrfVCQHEx/MtazxIJvKD6fkQqD4glzif+XkVeivMbqcIx2E07lBFxvvpang4ZPgxscjOHMKORBvqWpHKqj1US7J0Ngw1YHMV192/Ed0buVwezkEmT7s84Qf6lYlqWGmEPoBLw03M5QjIAp90VCssDvgu/aRZNIWYIt5f0//Pd7HzzYnzK0zqBQgtTGgnu5SUt2/uja2vsvuWsScmNBTJZcxmGCTs4hrlD7evWF2Bzr8uUQlbQMO5RY9MbwfoLaBDMraBdM4TjCkxQYzOaimP0rRn3R0Bnd5laXVi6PuD8P7/yADnhKf+vZ8HAeB9gqLljAoC7bNSt22Z6lF69Y/Fya9B8ZRIMr3cKau26duY2aBXVmG0VPZmGkcP7Rm4pQ2o0+pJ099rtOCEfZo5+VMeLtgpJa8V7W0sR3airwrCll6TSFWsnFGCWRwzBI+f6pWXWh9kdqF0EZuUWelW15ZXNzHh22X6RBrO91B03lvCmhbiigomo5w1b3OZG5MOPUIiuL86VyPtgvX0QH6gmOpT09nGynz3DnnVUepyb29NUwliu1t6VpyUwou+/pBNdnDTXOebiA60wnP0qikKoE/meoDsSgD7fOMVclziXSNncsQVr1kv4j0Vxm9a1YsHxhZhMP9F05bVBrivDKcLoyM1RXsAV604VXkW2Iz87nFLUXZFDrNzZHojLsuNuTYlqtWWEPLWEoBj9MCCe3HI/iuExWO0F6G1myRFJy5r9mh9uQjo5ftE7d8iJ2NQ0GdL8b/uzZ31VK7GoL7qr9uq88j9MG5FyyMnc7X/jflt2yQi2UlIKUs2l/3zer8btzwcZhx8v3xjrKwwi4tLOKX1ZYcYSn6eOILiAY0Hj7G6xSZghB0UawY1JB1syfDeziqgiyR9zmFx+F0CK1o6paaUMBGvCttr9MRxe5pSza0i56QFwO72/LHbsMcKLI69dxbFy9J+1N7qguDK/GHLptXukbdZ8FySlG5+2kRwxmlw233aqC5itTz0+uUz+oV0EQNQHlT4fNorHbtBSJBfwVpUzMrS/ysLpXcvdmj7Qx7p9NAU3afR0/QDHby9xZ8nIt38HcYOG7eCS+WFq74mXvZRPPWxRllcChI+1oJ4KHndstkIwqt6LH7s65y7jp8DXRYUprCaBFyP30ewKTSXnF3Mha+FUjyksW9QzC7+vLF+EA9eoZhsI6zHHdMW/9iWY4l2MxLFk+IykyG64P52UAy69BQA8zGfLHFfyhCgeoEfp9s3njqMr3LusYFL0zK3Ek8h6R0Rr5X4KyQupTSOOMt2q5VNw3V8sIlFZt2lxJClfWsZGL9goRHyEmTcLRKkalUQXnSTumSb6TuwJ04WuL4vm7Ff/yk27+5IP9v1pP83dRPfV9qzzExXaVNIhJARbrmzg3ayOS0hQ4cpcT7ZJVekRwSO91X0j7+KX4RevxxgCCsfdI9EValcx/p/V/bXcT1CB49OYGH88+YnIVP934C3kKc1fLNLUnfqqe9MJJpAM2/x6NA2AjG+9gFQIE0qzMCCHhAJgaQfcgqWJ9LCyAIm5hDt8rSw/aiSkCBIcnS4rsgwTIwKiaRFXzieNT1a/RIDxK9fpwCQ+bthR6g+xR/Af7QhXxAKtbj2ero3LwKtHRcUvWrPHTfva1IZPjLa2tjcPFITx1NVLG1WG9DBpxSsA6MysZpWG795vpA1kJ4hYL0t7pSTSWMBSXlm5gKpN5i1t7WQZ/lf7p8ZEUJt5G7bvaGXWEsAqOuTseC18Hrkqc3i7dS2RS74ELAfZbzXeaSV2yQ9Mi2r1ckDJKjVdbYAQ2b9rxj18hMZL+Oq2gBeBWk/UDPS8b0ov3a6W5tjDDed1NKABxgEFQYErLLOB1s/SDmCTI12Nv/JPJ+3gn3pWsAaVf/EPkYUGLeF66c3fifit9wa4reJVFbRcsNN5lOo3EYXwBgsTeoFvw2mL6zswtCfxA17CaDclJCOSGNMDYcT//SPP8MaAdRaxC5EpuaryhKxSJ6VN3BaooeTeUMX36bSdhrbj4M90o132zGa0kM1itobU9SPE27ydNvtC6VVDErVeYDwuY3z8Se3PW/YavK0UBcL6VPhMQ1ScbOwHMbQYSLeh9Y+WFRYORpK4Eb3sx9N4QBysBNv1EaAtZaSBNACMcirBUR1mWgi1bQcWLkW1AVlXOLne/7oXlYpBhgTDh8TjFpl7KF633F8+7Lc9k3UMHDvEHeVPu3G3Wt3KB0WWTAYWjR4MEKoCKfzXFG3rBhVtGd61tMs9x+jdWRnPioUQ+DWy+hnNysqCAUdH3SI9ahhyeOt0A9xenZvR7+OVwep8DN5U/JImPrgl5eHR/qplQ3yBd+8Ia1gOYPXFtc0U8BjWcMmgXpnyMeqJbhx80FXQqoiA6svufUrTRM1y6Jv7xQ7xG39gwJrUzVfk/99HTca3EGp8PXkCXxcJmb+hlK9X0cYRItuw5tPM/K8ORp4DP48XWWPqT2lUWK4tuuDbrY1PiCdApwgBXYu8ZPQ5YpzsNHwgZtA/z1rcDaAKVnGBWGxalD54PR1S3L3lmral7QrJPjQuUfRr0xEn0o5qYo4KNU0QspZIT9XkW0t995uozRIMS2kPrltbOickUZZqz6vguSF5vChxbRw908kdXOVEk/k2FNElDw/z/k6J2b+5ljFPR0GA86YVrImis94GaNRCPjpiEM7cXwvBuga22XJiKdQqx+2kiGAVTW7gBpAapv0rL0lHmma31fxcyC+FjbGo+2jJjUJy/a6+d2dawJa7SdPzu109BDqlHFfxHonz2oiEYmDgYyF0O1S4OZZ+4a0Q8yTP9oiFnGuECXpV+SFyNQme5jEwupWc+Y9pHy+992Wxpz7bzc03jtlrdVIuXNKw7Lm5cY2XNNODSMdZjXjrre3WQpfSALYVKg7R5iXiXm+A+2hV3kwBcTa+u0niHEa0yPPf9I0nALiFabwK4vp0CkZznzV490LwryEHZBDvYZB+ZmBDhCX05040DdNMqxir5WSEk40GhijxkD905G+GN87LTpRX7CUz2q5Uabd7piK4Ioz0pB6gpaOBCdwF+koP12G3xABOiQhsbU43qVEHBYMz+raQQDIUFhJDZm324pbt74MXVZ7qHGk66Kq7+zD7Y3m6sMd0IF2Y9J1UZ3L6h0PQ1KWmOfuGAmaA47KbKSIb3H15yGCTGCjYC2YARvbiqB7UxEvjuJf9e8qFQTGJibNDZg0jmm70Fhqiud6xaNZgZfSkiy60HJ1CNwTxVLOb4tB9yM161vFnVxrgK8GNuTNIIvNbEU0fLgxaxengL8A803UJtk5bTA6urmZQokIivSboJVGt11BAfeeFGdml8zZtzLHx0+Ap2V6V1Pr15PPM121zbQUqHY5aLZuYTOHlkOTZO2IuiZJhWYeb299I7645PY0OqnFfpgeEUZLq9s5Y9hjwExu2Ioq9BmpJbJHcGHoqGjh+BPnqHQ3HSDufYAPAB2dUYcoA4XOmRcHo9rigt1jzQVtoD9Mn/a/0GstbArnEXQFBezf/RArk3bDrxQ6haEz3xFJc5SWjZ3MIk4xKLIbLrnpgq+5dqIwB2OdM8tfRYRMfkN8lEE7oqsr5asvCa6I5RsM/fysbYeEFVyszT9NMHnTzd8scGJDDb4u4EsmJTXBClgHy3jxtNLMVHnxWqmseXEgxTVWYRqJJ58EDkgj5GtIGDQxJEU29t+ENPX8KLuDdYm7uVInQdgATmYCXg72GiReyp7FipB8CTR2AfK0SuFE20+lklwlQD7C7dzl8l9cHAA1rVyvjKEmFbwzam6a8aq/ITSKYAbI7YgGPyffBT5o5DkqNHXsAOxilqnAtJBrGmQ3M90tZdtKck8NOuKFEETDI5wqpqXlsjnCV1myidDOGmMUWT/7peyoypWMko/cTbIxKZycaSYekXadcnv3maSByNJ4O7bSBsm1JjWLnaIXexGiYaXAD7qsBdWH5SgEcfGbLsKMaZLkJ1C5dvozQHtGwvpvug+UyRPdmR9c0EEn5X7vng+mdRa7SmG9YevmZyHS4O/cNvupUbrHodKskqFY67NYkLyPDIwHOQj0KKg+hkOXyIapNWcCf9EieEWkf05WxgnNSj8lSjdTwYdQo2zHD9T1ieisWf9j2SJvs5YMwP02MCVXW9icvKFptqxNmYWJo+OtuINvxE2Ej3zQ0V0rYupGCO0oBeCxRzDuL569C9VlfIj4lL9kD/HwFbUDdMe0IyVxLA45ABvi9T+8V/CwjYetPzCVkg5jwvTkbQSIAltG9C4D4GjS2zTqctCoj0BTKpHDFHKsw0svit/32S0R3g2EuMcehGF43cQ1OiXbdE840z0/DYovDiUqIQxpph5KOSPeghE0S/46H6FNbzjYUAGxh/BB8FE8ARvN83ZXZIhSQizhGVzVnQipzwLktTRN2rKvw3+E9YzCGKYFLuFWM56gBuwgRGWcWveECjHbdNJAHt+MZR6llpU+qlPtUHEjsJ2Q3HDZNIIZ2MEXBtnQUK52yzv/1nROFgv0V0a/YC8y/iD1fxXkTGslKV+eDrwrPQ7VOcWBSGgOM4h7MrOfZVxuqN1wjohXD2+eOhl1xThmt00uHK1hIZb/MoxU/TA1jZlmaFAjewsz3kULjp3H45wYagHpq+afuV6C4DpY9MtfdrUNFTzubscZ/z3vPFv9rRQfT9xXE7Ih+zBxLKzfjP5zoS8NfQsKECbaHybt2NEgEpfBEHdtiLbMqwehzGCcZuJ7efWTnsz4ceAdv9nLgZBl0hUrfgk0wHuwHk4rxwdKkLJXvLaoQPXXmgQpFQKL3fRwv/hxXMI0BbrjA8V7PSGiftkAD59/TytTp7Rw7BAWMiAqCG2q9MD6aosECap7gQVzrb6iTjXwW7j5zwgmVIWCOXY53wYdE3EOfvVLjZ9oBb+1aIqTG4NvYSFYtp+eOXFY1bdrr8tBeQps5SsmQAuq0oon3d4i3zp8zT8hkPoRoXplmDLyG2QlMqg1WM3nm5N5nDJhy0inD5D96D5au0xN+EE/iclPmIASPYGZrRXyV2Jt1vE6VOS03bW3aoI6Z17gISi39vLlgMp2XAfA5GHJ5FQIrhXTffnsnZrgyVBDyH5tHYtWmLyDhd4tiuNsx/v2R44Yc6DfuYiwasG2E63xlr+RkOHnQT+/J+SnpRvIEtGg9v7VGMRyxpHSLJxoe9+wdOuc+ytRvMw/PbTcngy1LjUCitrGL35MtjOWevLnZ1vmiPB0HLks7/use5IUw1fm9BWe1gKox3Wx2V4oCVkW3SMcA9NPBRJD86IlcNrvBYFqfcVWWUFRAx02ubg4HMD3FmN8gLxnBi6sg93f3pTm0LmRNtLa614IZBV2n4pfkHzeVm4dvKTXQ7UUTGobTHbOhPzSKxodwQ8CIzQGxpUIRvUJwFTX3QpuFT6BZWJk21l2jgbMUj7TcZpMQ4XG5elcXSl/jvbuurMMEfrfuRYEqsxVLI+GzsCLR3RGsG7LEC+3omtj4D0jIE7DYlt+mC74ScH6umd12RUh/+x/DWE7TgW85Pssq87ktMTOR+zKay7d9G6SdTUrMfnfkuFWA+o1+gZMBEP1QmffpFwPo/pK2FZDcAfkaKXZE32BbLLq7dsQE/XBCLUgiwb+JfehfJ4zxvAWFlq1x1NnY09/vTweum3IKDL+xZRsTmDR4YkZwjq6zHc5OGd853QME9takjIxYl9KnxaKxkBmrIYyzGOT2n38Kj8p+URMh0H4SYcVFLzlM8qLU4tn8l6GQjBaCDyKowaTdnxKWTrJthamvQlzT9fDhHHO45wpD9vk/q++6TZpSK4gteHpEaBni9pdXhFgPbo5ZFWbQQ6Q68ZHYDaGDnWoWeidXusB7gAnSDxzJWTkXejHMruioNHIwc2IwJRlkXqYno4W94UD1TDUXM7EpMppWKRge+hABPXt01wLYPAHAYTX0VcnGSP5t5RG6CV6j3PUCB+AX6UilUys6th30BpBo8qBQq2FLMqsGUOdEaBONDdDlP6tLAQaWnTbg/gbGg4tRL5P9imty9VJIojhQ2zjgJl3+qlQ9iiq3BnU52POa53srGtB+y5KGHfnClbibNB46q/TzvxVAYhA7NpA9sx2m825cjQvMPSlVINgEpiOoCNiMIeRxhijPXRQlnhJtJKiS0fxvSwOjZ6tb1Ahr/qyWrRPIIEKolpN6tA2FGOYDz+bdiEcrO8dCLurxA7YtFzcOP6CLMltx8o5Qil90AkdlHsQbgwr/t2cyke3TS0S0OPiUKkIZtDUGObB1yiD1GOLm9ouv0vo7cB5o41pgh1xEaklQcgw8gx+BcZ5pBKd3bR8Hq+46CLv0stgNVNgFo05zwwwq9h8kD7acmz2mVJD8N2Tmc1qHLNwdayL4yOynZgpoo0L7YX0EL4MezqfTZ4OkszPhsZugUVZkYtSAq/08l9gxJMMXlHWzOroO6/y2Ybygs5+lWvDCXCpnIh005AN2CJ9VsdSshuZjIbZNbOAhDCTJu7u1oDoqymNRkaZ1NZ+8U5yWXbxjm7225s/EPxqTvFTFhlwpeV6/MV9NurK5ZREirX0lO5TvXsonpSN6OCKF3PDQHfMI1sRuge7F1KHfBFeCzDTtSriCizgDdZp+SetI7f2T8ZGhOvLtRY0Hs=
`pragma protect end_data_block
`pragma protect digest_block
369efe7638ab6b5be914d6e63657efb0d0ffc3e5dc5dcff4129f524cf3ca7bb3
`pragma protect end_digest_block
`pragma protect end_protected
