`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
u0g66kkUoyd3eq/5uyAat2pRX9eKT6O9I3+zk51VXGkjIMpcOV7Kh76N+12FmTeWjcJZJKa/1QbW0ZqxFoDzpngGfN5bYoZEl2fCWeO1WIt3RJS7f9XzZKK1fLsozoyAdJGLGIaPlAUY4VuG2de0mHOaPEakATESGikdiFdhOV9Ffhaa3HB4qmTqUNNxMq4O7dggkGkFba9Yx/QdgDKmUW33Wv40Kn2mFgXRskIFwuYfhvPfvgvUFxPhm0zqseJBsgUniCYkbDFl0c0gDn8SzUnxTV5WabSdIGZa+p8H8BNC8wa877M7MyL3Z5Q3IeAtwyknav5tOBZKMWio/WntMRZyCb4sVpG5a/R1fNF9Hgs9i+NzBm3Mab7VpM9RK6Tp8fASxnuTUnS/VprcKoOHRDE9uYBREvEcc++EK83lFhbsYmoZdFOmaF77pgcRB87LHFYl7PPfvfczXRCzh75aiEEksbJY2DD7shGEoHXWhUZzLHeW/8OqAjaVLd8IDa3xNtNM3L0BWE/Dbog7K1pK4Lqv1w7M/tozzVTam2rPgvxPjzz0E/4g7clsXOyxhYna0ftXEwZJP7ioR7UmFiC7gscXUgKTue99ZmOkIJCCOLOb7uBiNxNTgjtv9lyg4D1C8WCrkkslMkM8eeL8mucc9ge6xiz8xDMUCXOo3SzAf1FI2eqDw3j4LCOVLZ5BxTJAEOQBW8KWOVy/9GfiHRCp3Mfckjzv6vaUPc+8xWv24+Bxv3DaNitIo3Li7sKlP/Q9vYZgrDi5juNTJjMCcFpapP5UtkgHfb07e+2Ku/ihM5zMonFJXVJ/jlkjoqyG47rpbVVnkICQXF4D7ythZGQyJip3s69HHDhG1X2XJhZCBRCgb723oJ9IL2xByF0Vk57rPXqV6OHcO+uCCADvxvOPNizxbP58OUrSYz4AiM2JduVdSr9KK4qKzbaujxieZXEOBSWyBkhMsasS5yKIRl1xuCE8nSqlxxHpR02dQHONsi9unENWfN9c44LddIaPyky05i7ykdHrM6TtvWkAtkOZgAhFuFGbwNarSjyIrSBQsiG0HL0XTbHeUJxQauZ9EWHCrlZ5mTnr9tmOVdphgbihYkYS9a41OBiv79WHUZr7v9N0KBr3jMaThUeaDGMFOtJ8s+uWzvWf5ZBCWd2EgYFQx0J8VudDc3arMsPEw7aifiHCjx8utHCOFHKrX5OiVERxeawlYq2qJkVPs09copAwIdkPPjjVjghGD9jpqUAppUqML6n5xShc7Nh7I4UnVOTipC1cWJYrOfMePX3iFasw4me/g4k6BQc3z5+tg9wjo+Rle4x1eVzZun7SRAAQ/WH2OO3kG/I8+wzn98yDYqMLF4hyx4aWjs46yqmKyYQVVM9XsELahdxD3deAUzn8FsVtwNV1kularktI9uifVwFkWT0MPdyjudyn+neg2J6qR9WI5oI/r4wPWJ4xxmzGamQcosvmGOZUUbx6Do5ptkRbwBWNpgequWQ+gdDfA48YzQAKK1dyaWZHCw4xeFMaNe6vm1jObNkHBNyaIlY0d65WMmW91WYA0PIGqGRPn6A0H7SAQaInEixrtnzjoHDde4h7SutnqXLqqVd9xcaQaa2IXgX4olOLX59KDh2UgZAV0w9LcYsOV+S3ExWvpq88Ct8YyP6pXipeva8ARi+VsQBydAu4WRXbJkTmtktZkzdAOBAg9G7cBG45ZkOYzSXWvVD9MoEzlUVoUkL9Q8PzBwOXejZVXtSrZ2u3wD+oGaJmya3XJTKJ1ky6fQ4lQyQcwcCKtMJmC2Wp2x6n046sxC9S8BqJN4+8d3QJgC9pd8ypudI7FvcPE+BnN7OlmlgxDxn2uBejrmGkIPvvyJn794yIyK9/0iaSndXlWO4c3qpXk06gftd1gFZE7gM1hE9FSdAHkKx1RIG1gKfUtu6MevjyKDbkdMwIWaVkkuqn030YolklZ5xQzAgE8j4PHv5cJOGb11aJEehVe10OTRhojD3Gc2hPY/y8cQLAG5M0TeprKBlVigduyT+LmU9qdLUDepixJwRcCVDDr8GrmFaXh+BPxXmCMrF1GmTdCTgo9iSay8rErGM8lCXQEWRJ5dsPvt/YlG8QoPRkbTHTfZ8QyyAp7A944Vq8u7fEScL96XeGJOQNlXEJgpBO2hMIg/RiX0M8AG9IlweWE4Q7zxjRAx8ouYejtqEK8nQfJr05kdNolxXnOIAoq9xjH1CfkgQonp8rAR6H9JXiP9SNv9qGCecWcRqflR5v04c6gqPztuMel1JCAsfnZIWrmn89Zoaa+WBf64EYxhVPxlLICiXMOWEXCiikJpsdRDmK8+me303ZzQ6Mly6cEljDAvSM0S0MF5XxWI60kC55VxTAgYFlfV8IYdMOpQrl/oz07bmIsDwSed2j6AFKTeodAmvCdxRrUdM2w/W7/spOnMq3jooeuzuAgyNeXVsFOktjiAE6BQgXkhsP+mUfMee9djsBoXku2rPuFkimvprk9mCzEZfW+0d0foSXiPnUSeQQtZRmA8K1wjyPgl5TrG0vHjshZrJ4eMniwq8s6+qJC6sr/yD4xcFftBzPBvfq+lAE/W391sXe83tG03mfaZRewXrxn6Y8Gz5OKf/rs7dw3NrhAPHLNGBPTJGAijj3JUCQDzyrelLLektqqot3RLnCERjdiXHelKl56zLDMzbxoITpFPuNIEz98jNQ7qsmNKwr7KOi1pVvCh9meuccmXlfgTMU0jvK0GbPFfkLPu/ePHEV3RoHExTqSenvbbEtgKl7wmjfSj6PHCCKWQb2WqvOoTeMjOc2FpCfxUkSVgJVFEFfTtV1zGtJt7tZmklumJxUnaiDdy1WBZ4FWOTOvbQrEniJI51yDj1NBh18gJZ2cOimxgD4WBCuy2so77FH4YeT67bgPDu0sIDPtQNztZRwRxXtvThhV7MLRAd3u+q0655zNTeJr8mC5fGpt7BUhITsOMR371TRyb12M/y9dOBOEhaQzEo75HFmQbNqPjMMmGAeriV0yWsJD4rAeoUKHdp9CTYldiaQUUuzP6cKcCzGXDgYIzfvZ0r8048pK/cfVkIYvTlMtkCQB2IJoBDH6RMAHvl2HSyVVZIB7+1uYjbFurhpgh84uz7Ck03nstMlKO3X0CYrF6zL/F/StiLDcBTrzKI6BghjOZq3hhzSaW1QLHAXKUm6qe9u+NvaPJL0eaeKASm43J788IMaOU8/Gqz1xiUAMj++yDdNBjN2QxP2WBItaI/kbZ6SvQyo/IP8+J3OKL5cR4+C52Fe+sODOGOpWsRSARmcE3WAJR+ueFLnWuYQzqPVz8GsphMFWliux82/zuB8HeCojoS1TYO1cJm/KmWTq8pefaBjmgp9CkC5lw/uDfOC3SK8z6Pa9IUZIjcMU/fCZPOtikg578BbSKV3HYslYAs3S20LxflhxuHJJOBTcTgvGtnY4/oOlFKxKv9odSp6Fz5aVVaQgRaXD9AD2oMXY/3Q9ltVjLY+dtRDeWlLyNqxGSVGix4031ddoAWXtj57sCvdFwPquVxulcrUnGUu9f0i5QtXH4k7101BV+gIB0mhu2bfBnCXtnpPyiVnl2sFo8kPR4F5Q22qviQtNk5HS/LzART431ft9WuKxLHRoRMKKgUuZj0f5LMHW75P8alMZOt+1VM+XA78cqg2izTeqw8mbSExCTLGpyxt9T+y0kZzGMlICu0sE/4Ym5xWFLmCTjCDu7urhuvZCJ+MRabl3qbvK+8AoAJ30NCjIavMCZsYa9et8W4E2XFvylyJ/PlPYG8nCGBBorTnHWVfUxQx8e1pJXx4RwN1XkhdA05H4FlESFvloGfkdNKGFiM9oBlJ3HmvRDyaLPCJl2oymrrhPuetTzP6jtqlFJ6TCMmF70Z6aD0VA8a2tVopN/cdmPo3NUNb1nRGjnjERZjBIIbwAKnelVbPvj9LWktGwWcNC7N1g1EPKLPkvEqT1JgGUJsv/8eMzQzqixaUO2eF5u0R+ZYVy4CWeh0tLD5g4SFEJy+GxBhOt2MlEjWjFYEura7xZSfhDJFkiqr3prwAd3nQMP4OToNGqrkXwbixjiiQ/HJt8UDIssGGZ6uFB8XagGkkm7N/k9WYIxlmzQFDvTY08a4+FhHS9e+4hKB+X6FR0vZj1yfyIcTdE6xwqnwRgkVpo8lsjdsEvRtkicBaypVQegByw1bCvYsP4wWQyvk3EIpbLibAWhMo1Obz+H4KQdil/MtA9DTL8IFkd8Y7kHBWQUZwaEG1GAvnoZsmFTNoc+K6N0A3FlwXjT8Tvty7XJi9WfyUORzvp9+5Kd9IuN0NUv2jex691Qok22R8IJYVqdXyAJiKIGLHq9E0Nd1XS568AXqoCsIkf9EmKQDs7UU9rJToYdnbW40+f7kgv4x/oWE5BjiEb4ejE8BoMgVg6SwjXqmLhkfEHcCaIBadNuQQxeRdiAFxRqL6fT4sIL2GR42MnhSY4o/rS/s5i4myhqVq8YUaAnSB69pG2IH2NtDnW2biwG1fJIkMWhChH+T5RQc0BhMUI8ES4jWoLzL8EvV3lLMk1jfY4itFwHYHowRMJvlG/DKXmNLwkjzYO097gF3yL99tkhhG5pGAB81mjWDrleMLNk1bOV5G4UJwjoLRR5ugmm5Yw3jWAR5q46sOEw4aJh81orm0HK1dCvXzZiBbDm4hNHzaDORnmlhF49P38qaW4ktbVBpvTCxCs+tcfdgMGqExMjTmkJL/uQhSfqSnZgaKDJO/bHKzoFlVDCslJJjxqvZZFH/D4RcxMqpHJ1nooZ4rvifesIYHwhEJbc9r2wEoiuxdCy5uiLv3dTyiq94eir7HJW3idRlR2LGJonIYVBRiFQUNV0KeCqTzCsGFcNbeJhLSCeKzONoLRxKsESPgQ4gn4qLf3Tv22zQ27gTFPjwiv4A6QP7y7089umSykKXq7PQeivV69WIS7qgUhd5LKOAgRhqF9z7Yme6TL/bu4L13DwsbZF5IhOEOPnDDfG2JIfpD+GIToLQL7AKaSMpFdjEAtqe7Gd1g6QE8Dc/gSHO1/G/QJX07yMCnZaLjwMAcD++daoiT2aFI5jCqruBLZLQBpRCEcDvd18LghG/oajih33Jf36dE+0+RjLBYT9rKe46l4gaj/klCG8khVaP41IKfYFVGAWoveXt70Yhpk4hYsanN3O8ISiEyveW1Yep6eJM7wqq8cCgnvTVK78WsTL7an9SU91utW+Et0iorh3nlLERsCGezanauNFPznAtl0Dlw3ZJE5zFKWRBn197o5McYKSB+Zuuq+AywGDONlqqNdamOdF0kci9ymkiq3Uw6T442ZQ5PnMpZ0Fl8rKP1I5RIkQ9sRV0FVy9FhSfN1IKBDKSd3tbc8Zm2q18lbYDlWE26exgB/KoaRPL6IVI6sLjTWlKK30pHfW11d3BwlEaTdsxdUWHoZBbbQ0Q7iRfaADVH4SJKiPgohtUJNDs+YqMzm1VoHP1e9oblBreNmE49BY866cGnjldePWZK6jkAI8FGsILjuz5VLXCCeRy3oxDCc7jrBo6ZXI1maYSuYvS6F7QiB45nb30CIyXdlkSNn+0dNZfgb6nTnTSFTSatnhsnV9ahW9H62OEni5jwR9xMHqhEpkiPlgb5hY5Jh0dYZCzzrE251/fgka4cl4YZ3V9FhzyQ67UyHpd9OnRF/6v56AnmGIGF+BaohU39CqA1jk664OehE4Unz56z8zqc9O/C8gi7DcFhocgiLp3FbuhyypBs8aRp3jr/rwDIgqOqqUWLWoD6wBNH2zmEiTOf2JYfCDTDUACEpsCz3Cjn5B8rUvdhXr+/Kiha8L2u8uhQ8WRmEy+zPHjwyXeK+xhPnwBDJlm/F+h/F3jOEK7jbgkvpHAkwCo9km+Qew8cEo3KkO4RlbdXaF49jk7r/yyrCa8C++9YJ3aDMMvWhez/tunVr9/gN0sBrtNOLl5tnl1+n2mHz0z44JkYpaD48Mx8AGVvO0UdK7aoVZqWoZrFe3sh0kq8bq23ONHI+wQ6Lexk+TCXFH4YQXwrcOQO5k0HbgBW8bKnzp/rCJ7gH7X43bAvfMCPN3hyFY6bOOnStz/P1bWGHgDnAP6bXokqAGryU+q1wJoWAz3FJMNrob24VAxCnYIn6JLO7gyukpu2bL0wUbK2A0jaOGGBydSYTZ6y9cUbbbyNE196rytPoPEcAwdICPgqZdPDoc4HN/tkZ5OQqKUqvQ0EPfvSHUDd9yAh7W3ZpNiAGDVVT4h+tf8J4r0XoeZtDM/bwsFWPacEYRT1cuoJbgvtWQ3PGIdxJhKe7s08Z06QE9vEHCY8M+HNSbn/gt09y9Ad3vinwICC2mhtCscgqg1brt/35nYkJjTr8pxmfir5zfjOqR8bqfYl5QiECmklULYPcbVfQIGYsTXj5OpJY5agw5KVUhAjIGNiK/6+buaBs94BKFufgl9EQGYW5GlAwWT8bWFkSq/vh7mlxyCwQo5muL+y8Dly9qawp5fZfdpVKV0AQQIjntVQEriLJDpWllgX2mCpJ/VGjQDBRF1V0OW+WnB70yFW7Bff49N/7ap5KjeA3KHkB1W0MX8bZbmxW88sr+AAWndcS6HDDW1vqepmZOO8ZpyGIFwEyxF2VfosWVelJ9FCXAxeMs7TYWuYit671lg/r6339k3S0Fn40cD0frv8n0jzNozyIYTVzxBYOC7PSV+Y35HNqGgpDMHoakAOH7QA02YxqBDO9PaUojwgg43gpFSuvtbVpnEDwJT7hDX2u46Rw/kKtK4ETy82lxv/xpZRvR9eiihVnK5C69122wR5Kcheb1260fFYDapB72p8RfN58OoT/+lUpGhqJGP0ZTNF82qqe6kfu9SQOx2fwN9/KKZabAxSF1B/0EkC2dfdiICwg6AEzH8XyD0VaLWq5FLOQHiWxHNWZ1ZF01wfWk0NeoOaqMhqfUocaowK48ndUkbORE3h/l7jody5QtJa3f8sDfyc1uYQGJ4uCkk0RfFH9p25dEp9C4q/fxt7mDQblJqg1mAqu3E5oIsE3g9lz+hcSHs71bauaHoErJdOsBCo19v6XrSXOLFDnbDUBL1GLcc0sEAS7SRbTpnoiv3W97cVILo/vKZGSBZnqpV6rMqLl0EaWtidGLutmOr5v5HtLl3cm2u1h1jSR3kPglWLoX3zBJPM9+O4ZSTsHpBkmkoXFz22PgPNuf0GViszPTut0BQBjm4XB3NrRXq6pKD8CU4hgeBpc4F0IH9refinhNTmGbJvnRcL+SGud5p/YPixu3FZ7rIvbQWZjGSZPOgsLgVcTn+rozOyioah8lz4JuQpFTvOWJ/WWgQEK4b4lkZfv3l0q2J9k0SqiVNTLVVS1mXDXfFsiEW6U2uYNNxFRfoqwh3gLz2B+Y/23H96FFrDlJtl2Zh1WqG1gqck29b5SJmg67UhASO/9Lhma3F/e8VH5KKRUDlsffXKQrTwf8yqtfc8PplS4A7HP8obao/qnAojNDe6B4YeqaMhClbHl1+zIFwH6SthsmOy1EG0nutZmqzeZKgmUqQL/8AdMBNzbcnzxT4kMM0E69ZP3Kbgt8fV2PK+MLIVi+WTSrCYnR2RwwZXShrN7KsdkxpXu7Q/PaQTAONRdnIFySBKEBHupXZlLqS33tQdRl7IVAQ90+6KnFkf7a5j7U8SZJg8YDIqhouH6Mqb2/B+5FmNgOcx4UMhkZjD3drR4ujA9/LpKAMNYqCau558+IwOCsxWVwraSnzGytW0Lif52XmvaX1zPmeY73Yko1rkR+75Cg7ti7Pp7T/CHX/mrF2OsxmseFrWbEPyYakoIuwtq1dI1c8Ci2mRPM88vUYT3PjL4KhfchViA3wJgYjPviaELXoxaX1iohBZBPZEmbviHM6RGoWGQ/AtOlsddX0HUy9Qryu2zjgwa5zls1IIKOowoIz/FdQ7qlKuFum3LXd2Uj88Okk6LYCZx4bZMZkSxtXGUJK9yE0ooFxn7MosX5WBuuif9PaY2/bFYIf6tPvgMS5h/wPQHDmPRX+s/ObNyagMrmkPfZ09yjhNaX3TxWNJtrwgmzAkTVxxqFb02Qv7KqteGlhlG04tYV99RdSyhNGSBcbw/IhFhh2oiTvHGjIBhDGcmmIrSwQW2/ygrW+0dYuQX4z/1Wius7AS7xu7nKul+1TVk4pbw5lgzkU1gTN4Scn7pq/uZpDvTfC7groRNVj7lDGO+V3+9wH6npE91x/s9APzw3OOEExWkqkzt12qecR7uj8zZXUz4GK0B0Kb9Xe3QGmst9U2mbZaui+DIo07ZG1ImjHmtMbfsEKkyBlBtVQibG/A5YmglEAAYfTGs8MAOhTWdHavKWWmVsbrB5MQ6wp/1iedapWFbn2QY5MwunImxVzVtjiR5m25ucG9nwTzuBp2zVXhw4Obi5TLB7h8uz105iC9Gpi6KkLWcQzryvJsA98Jaeh5GoI7aigk7stJziZzLot7isolJ+J2B8JAxM0TJcSeDbBRx9Vx5k5IYX3dK/PGfgI5sVUWufnvv6oGtk8Y6F25Qj6KVJm5vT2RaMlOwnzv0AgWAGgvQ/ec7EHTtuOqgdoszpIZ7pOc03jccQvIAbHnLTR1z/63EqI1B6tyU8bHijM4CczFj0+vKX1qOqm/4TLDdW/d3LJ10ufsyI6WvUc8ZrhZMtEDXS5X49WPGuupbK4zbvdXP+YKt54yYKIgZ3dlwNpu3ZXj9RyI6saKQU4daq0JZU/7PKcrX5BuDnefZoCmVDbzut3yb60ddN+oee2i3efeQsG7CjQQI11wYb4xuwnuywLSNdvCC/J5WfMsr7egYYmCwacjhSXRJyhwwVlZ+R6BWQ7q9y5haynQm/KHRvrR41UF8urXhG4GBIigfuU8utB0mNNAdNpFbGN19uwWfAF+k/THWWnXV7aQc9nctlO+KzC93VwmEsUmasHTd53Z//0TcPLrAN2wq1C4x1uOFQpH6crAUKdPT4oAAJ8/2+ovveycCahaiaSfRE4uHQHL8i7KfLCFACN0EUs9e2eIrMtHtAeMw63DSx3P44oqCzreN9ugtUXzKzAHE3rpgATGStl3KW1tAf0iZ/sZ8ypudhgVOu/kM59atAE+wJdyIpkm/Ika3dMPz0ehb7oNVAZq3FpKQj7NPY0W+q9dAzScusWh7a/YQl4MGQI4oDz+0g42IbXafOayIbOqYhV/KTejaFMR062JFV2fAIy/ZhEhMq19kiOMwnPzMCtu9iYulufB+im1tgIvXLdyggaY6VlowQC6AxWQ6Imvvk3iCNKgjJYEngElLyqWxmmAG7Lf2UDLYiz0JFaIDiQxn6fcAu8HBVcWngwM1FHH8vP4XjGKCl5mHZdfbMyusvH2UK46WkEW5sKmPt1/i2W0niEQLgM5NmafTF/mdglUuuhKmlNrLMVRzacX2N60NyNkFmIxCUDEy1+USWAEgrenWj4Kj/HCLHR6L/juP2arLHbFQlcKCKmnGFSs8UR1NRh/Fk/eCmXvYxcgwWKWqzJCUKYcnh6LyHB8FIbYoXJgm/p+xVnbXbNLW4M6eTM2sjT+nx168wY8cDHGq1w2L7kcx0kb7Lq+RjuwLiQ8w1lsAgerJZK+zzbLuo0/zWp4L15DdlY4qpLk7larv+pJ/X4uIMFfDYbFyYU8Dis0U7ZUKmvlnqTups23Af2GzJVL5wbAsGWkNQX2R6A6VfAA2K1fykj4/1AT6YhNCm30jpUphpktCpJzc6tgo2XL6fwszrvkURe+Mbyz69PKGV1lXQ3xnwRUurbaAuBLnJb3dKj0I5RsN4VYcS3jgiovjDs7O9pTSt5ysPKtyM7Xo6oJ0E9uSJ0aQL40zD1gwSSt18yuh6uV1wh2JmNpwlWOKBqA/IJyR6dwojHtNFbPbdHxzuY1BHxyoke9tDa2S89aosWu0tHIc7spMXrabevsawDhDigj3n32FlHSFoJdB7Oe6Enp6g0Zi85a2zbQz3RnhnMFwUGieQI2voNzMhGUCD4d3gu6FgilrXDltjXCAhFusmBBn0bfukVmhxFyQk7tFGIYDPV98H+8jNVwvoMNY3+k4LLAmHKvh2W/9LGSwxOKnhNFtT/7tNpfSke3WvXhMafReoPYEBHmGbTYSl0p2EVBSXrvgSqd+Ofj+/AN85ua79EucxcM+b8dqiAUG3rtTxogJyor+UP7U69N4oPlyQwrkfyATXDINyYdiuAR9oDJLKdZ3dOh8n1WYEXRvEBiYmorHlSpjHe5LyB2UA3osDjLRY2o6CYa/dRHaVFJlCiXm18Z8vDSLZY64PK2iuXWs41UWTTFb4QAVC2kS7R3+zgqnDHObBVHUrVY4rOGYAzN5UyD3ge+p/tbgGDcWghHucFoZBMAGcZlOnxg5Z8BV06hQ8p/Vf9Kux+TLhApv7Ma/tcvg2iCz+5vEGcb4xankgC7wHJd6Xau9jZfCC7WrLWoqxg62N/7vUPK7Zgi+XvvHDMqYCIzholEG0/8KsJzUt2H6K8ruerbKtLcE1phyMqe9HBlcRQDFCiyzSMMU4McJx2NcQCO/5GjUv61vWDAS0rNyYbvw3Qg4fi/a6hhgA4X8GrYH4Usvx/qVYIeveW+v2a7qV+Hv2ngdTcXYMykoiF+cpfI5jRVNTmpgAhcQ1nc8sjTpAlxy4YD+lFY5jpr5l+jF+KzZZ8+KH76wAXT9611hsRMHfG8+/YDTwrj6JDbdixCtWRsF4cfR2v1nBnHrbwsje19j/07hBquiBHymCimT/KPRTKQIWh9GTpyzUhFuK5ftWEwvUoNd2ZETO2E2EQDYk2j4UwCrN3XB+9LT/2xKn+d5E20O4ZqIN72IbHXC1eA5aiXxIzz7PmXQRWff/FM45XkRWJJPY89FUgJyufUvbSSrqhwh8fqTLZlJf6aWlD5eN9OpB3v/xi9lMU8eX9YQYZt7cqSXF80p1kkNaL5ahp7dsFq75xL9z8x8zRE33CTNiNSaODHSN62QJ+lCcoNm5xcu34uzQVlcOgBi2UePIDloefnW54AEOFkvFCf2phPrduDWV7s5uvcx/nv9xzDubOp2zafY75huC+Orb6lFQamBuMf6r9RTW8ZuSBCwQgcwYEISDeEDU/L3pErUC8weWzf13eHW3FlJ1P3cJrhLTXMXfKWF+ys9tlczU/togFvRHmZKwzJ6mmqLalwS7OkyhgP94Qh2EjepI5HtSTuZN3ivuM8r6EV85O9lQ7fRNKRjLvcoyQ14kXZiF6mxW4gQsiN63ZQvb8S601bs4GYsxdiJNQLP4oqH1H7I7xTd8QdDbr9Tq75Y3Jj5iJpqH9Bt1wNF7I2eA8NO1r3fTq1i+dWoHGJwl0N2J7Se6n/g4QPXBmVp/pQiVBwU1L3FtTqupQIXl/ucjgH0y2Mki2nYw3fSlTCADEHGJgsG7+91WakIsrEdwLo4+Oq+bx/Jsw7HLubHqSrFLtyjA8C3f0Q772/pJmIeQOkh4QXAoBu7sFn4xxYWw4W/dV0rQxX0JaSFTD45g97/+FwtnW/Yvvy5kNLuUfAbxqBsFTCJH8Cm4s818uxQGJXh08KgqVVbw3EzX+Ic6oSJytwSUScTynnPloJsVqYTXeqOE/8ddJMk3MGeN+GGgsP4o7t+kcd620WXA+oAZqHKD3K6EdKrXtiE6iECMJQ7yw2mFlUlwYozpUh7vlJOEZ3raMcbu5w7iu5Ar/AmS/m5NJmOEvhhoL1wzwFBrsZIH/4KeiSRumMLnyoCkyK7kC3/0qdCM1eiMH9KB+OHV6bMRv+cKDo7LDSsk/dmPy43h5wPQ8WeHk72H+55CmNrDBLZXm26e64ob1er4Rr7SStyyEmutt3AmIFmGrApym0cRLp32RBix/MFyfWkT3gMqIoi9j3yltG62ddLGYSwCUeIbgJLI9z3yOgE7uey/djxMGM4BYC3suEA9mHrpAVomUYZpEt6qFIDxqzgU7+1BO21qLDj0/MoA1GvEXqCDJgqa90Xxd43B/Lcvho2No0xU5KqXQ522v5/BdT/WDYWAMpCIZVvIVHBM2GVrnsftNb8evzoDm4kVrNC+iZD6popu8y3C8ZqVD3JwKpdaERXftTE50UBEQVreYYv7HVs/gCIQG+FfsEml/kkTEPP1agSG0YUmBmddNpmoP9zgNMjh8elM9ugcCnT+A9daacQA1IWIAZQzYpQueHPhi1/lX6C0lmU22spxIPrnLMO9xG+nAV1ApaX1BrE23bQsiS1EN2rB1jPadpsQLLSsRhbuN3AUCOQDkxclD2wI+YECG3a9+Bd1lvXXZoKIYfc/YfRsR1rb3GNCSf6ij+s7e8iTPRD+xpdc4BxxemUTetZ4WyRB1IEm+TXDT5qOgIYfUoXNdJgBL+RPzBP8jfJPXCzYWDCUeCEgwY6nOzEcJzHt4IeIYj2FVa/oJnHCQKbnIIF1/Sl8TQXA6cII2W62173EBjqM2JuMZkaRbLWWMWUz6Itmeyne07vPH+LzQwQmUQbefHD6Bk4CCnAnfe3OqhXpBAjzW/zbFloGv2N6ENrC3SqIaSG16oi6QETbTXTaOQyfxLS+5NN5f6nYO1Cn/giKEoEs/XFeZuShLFR047Jd785rkQ7XTFW78gyLjG1zcnDmSx+5a+e1lCeFKCGG8B6dTOl7uQiaK87kdrKVZdUyIeU00o7Bk9R/oxVp8m8It7dHBvozvO5o4v8avMlJQODUjIYFM8ChQxIJQ5kdYL6TcEOGuGbHZVrW4yC/Ch5g3Aa3bs/2mJ0gL9cDagwSsfRmwn/X+iegJ4k19hMnF6mVL/hXuyrWEvznxySC0QuFfQ1v0YKs0oUPPTEUnBZ4vS4tEEbLdww8agM+WPWIeJYTu8yERMx7M+ZmMx2l4NxlbyQwEfQUzu9cOggV5druHpWer12qSZJYa8EKXe0BQ/Ut+cNwkuMId2UFnD6Thy0ribpWUuSBNOiL/EZDm4FGmC/+54b7P+xPDAEencE87wwuMpffZsj20tuuM0pWjYC1sm9IsTc3Xp0U1ce8kLgXC9mkMvZRPhCstNARVHnTqMD7N+hAQl7NpzKxMjwXqwNy7N2hN7HCOV+Ou3ufFpK3f2PCgQW8Xf/0qQ3zGrW6ijp6fVMJv7CPwjUh0zDPWro0MSVUVBzYNTgHOj382DVukn4NfdbicSeXJIkZ5RlPbQWiC6KVd9ISRbrw82leSP3qFuOx9dAGBNjt/yD7Kf4viqSJsrp8RJG93SuYjQdcQRT3THP0VVMT3Vm1bBQkKvjdLzc5uZFcY7tdZ4rEyFjZJecnd8EGMehUHFYS3+zsbEZB+WFVx6e+MrwKbcndutIne9V/0ejHJjEjgzNUn5aYfL1tZjy50cC5z7npQnD6BBc/9PUzVPlOgODUUA70CZB4iaySELkS9NLqmPbHY0s0GvKBIB025tBxzYHjDPi325mz/cxrGRlIgkz+Gzl53CGqICDnUSNLSkvqxoIMTdaxGwwpdMt0ocA4ZgUtW5FHkzragbVX8DxNeVPBRDaldtjGTv64viJ9JA6bNnac59Br+zOwKa5ivdGil8rzr5W02BDsPbqfSsXU2qqn1WjPe1OyaYbZXyy6kkE1OvhINoqU280xvSzh2BXaVvI6zESGPPC/KIGR8f2u6+ahP3hWu/TfqdyP2ihRCgJaUL3VFY2Z/qkuGSAuUCQeoTLE7Oy2CD98MjQdw7hdgUXDKpBGrC4fKLes0uJLZ/1GDYq5OJNEuEUzfn/DXgneAKvK79c7OQQceal+s+B4WlkaceMuCSJr/scLLp0jy6hJ0swORdiRBWefwAQdGszq28779YauA7Q1qKYGZ8UzNHKNWdz3uQtFoowxUnnELg4QJ5h1QCprTsrRiReQirnN4jqoSbDCy9jdVN+Qap1BSW2WoOod387oOcOi2zFMnEMwIRYaNkjXmBj4dMh2EHFjnALrhFELimm3Lj2tG8Jv43R5orbXA8GgFvFWqYmyV5xmA16f0J/sT085MT5/55laUipjoIzJv+STthp9S2fLN31EFvsh7M6H3t98Ylk7EC97o1o1PYSljvUK7e7KpASTll3Kr/HfWb6UBiZaOM5qRS7acNjzrIL9i5rhYiFbThSOaLoxkZNUxvKELWic6Siw+utd/XUjn6DDLk+ikFJmtySBheLF2m62p8uG/2fXTYwpK9wFSTCrtkobWi5bZMF/IvjJFcOIugmpVXWxDvI8HgUfbuS0ERQuUTPAKtarF8VCPZr3shoY6Zvl/ror6X7NiAiFKNuWvFIAaCe1AkOlrWEykK2ikWbmcs+pR/ed6kMdlkPx8RD9cLuTP7/IurdWGKK2oFmcB2TRPKhuLTARK0gkNjBx2dY2ciDcp3nvx5QgO4aTTVdrJBMWCeMIA15JrQAZddovkZB3vadl7mOiTNNGxyUfcApGs6bsa/hlqcdIuUOV8vHB89LxwgTyv1UTGhTxuA3IGoALfNiNRWwUvGBOCJTXoi4KSQIELgQwvQDf9t8dfDxQyEytg/BnVlkZIu8lXOns3YpRS7S4oGe/u6RwovvgztojBpy+ylbMXmKClJjwJCgj7TnQtgC1AB16l2KD5iSErymUi41kJweimhLUcitFRuoPV7o0cjvsGR3uw7tdM/AbKh2LNgALjiq+4ZcuTfQ2F44/1JoNnvhmc0ToZl/teZFIeFMGT3qdSb+zbD9LCwOrf0+wonlUeQjD2bFAziV7xX7Df7lVVpkTx55qWLGBTrfCMmefZHV7QhoRbUcy49v1HFv4rtro9AbPxdYWaOGv+vmC9tXWKaVVPm9yZULbQuuaEqlrAF/zpRVjKEb2sonFmNHXMIkMOcYfdNnJnuPIaPd2u1AKFE6ILxKEqqqnq4Ad8U1ApMhgwGBxn3kLtEWBjUnEJkaCSI3eEDxpxVZDKu4zeT+RcNQ0rH8Es8JpTCfui0KP7wY6r10ZAZpbC+lK1PYectihNtoaENoCrJ623Nkvmgizw4mYXpgdMUFNPYaCKL37CAG+DTnrG3nujdh5w+scGi2abGGRc0Qeeq8MrgXAHYleXCtRoFWrp4FIlxzTXDqQXeJKP9EBaQ/iN5DczImi1kAdgj/keGITjmEr+07RL+ThWFBw/L3go8tCOZa7kjuUsbL1MvRN/uFA==
`pragma protect end_data_block
`pragma protect digest_block
9c403c291f38e86f3b508b23cfaf861301b9e2d0e5c674650629ed3d5ff979a5
`pragma protect end_digest_block
`pragma protect end_protected
