`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
V5ugosxNq9Ov16Ufg2KlbW5HQgyqlGDGqf8k1RQ/gq+7VNTpxgDYq+B++Po7VuXXRSWP3/3KsCW0Rx3ku8T3okoz9rF2on/eIbz4oLZ6uWr/iD/wux7i8kyO8V/JjwbAgQfFimwTCYIj5yTP+NLkyq7VpjG49Fi9MUXRlNEmIjawS/tyYib6pP9qR2Tc2zTrrP+H/XDUQPS7ief45Xf9llgunakqRzSHPxYCi4wx/Gfry9j/HxfPnvahR5/gawiwUFRH59p+dKO34f3ra9VH1XK8qBfiaYD1ucf5Nvsl9GMA1z14V1Itj+ghvayelIqrxuEeNIKTJ2i+vjp7zEw2UhJ/+RFOoGHFW/zwTfrtMrDuUYYnOw3XUYUtwnhmllj3IAo49OuWMY/APeHm6gr0TmLZs9oNWuqpEAxYVYEZPSYzEipHCHNqgNNpqgNnN2CC2v5ic70IBAqgTWXKWRQCAwbFblUJLWrWzQR8bZ83X5S6CFPFfj9LJLc1gl9xAy48gEcFDuUtSezxO1c3Rgz9b1kNUQDb8cGAyyY9i71zFr1/GoEPXKuRT+LoovrUxex7dWPUnwRoVxKK0g1d7vftyq1fvGztOgO36bNxTSsgMCRIUNX9EIArGqEOqreCXWY/UUFH70bYiq9QVXWi+1v9kN3rrOhe/rGyAkol0MWsKxTX8zbPpii8el7NYH2LGG3OMt5yROu3emi2vu+Q0LDZi+Cfk1jeLQLM+xpEVTxmBmJTC5TJb0Cryq+rEjbvWwe3O3KK4nkSrlqFSH+esabEFW8Yis2sKvVxhwRZQ6v03nNBq8hH74a2DExPUwR/ljSlenS2K/XXdvWn+SOfcLIMvGS6AzSGilta2CNIdEdX7PdkKUeryUH5hpcsVR1QsFPmuCt7mrO20X5T8vlAJr488d28GT5219igVvntCm1EnZmTjTgGTQs/XNcHcMCfzbMYIa8OGxfEqOkbefXlFEMC7sa/azsgkoxbQGNmZNRgMzxIjA/dReATgL3enYxGUXJfNPCX9c5RpEOXMwOPbJyqNXA5Hh7ieXXA2HnmJl7haNJb3W2ZxXjlcekZBi/H0QQf7mPgHKrvijyV88hcd7yIBrl8sg1HU1VSfEtLIAyRFjSvXQm3Ce/l4HBExMNX/wO/GFMeifoYMU9+5gKr+8SbVN+43r0CF0UYn2YjsJq2N0q4JrYTEuoJSRdCuCuPt7S299WMksx4YQunCcll7nA6peNQ08oEoEYHkjGzvTABkOQhPoRGlLaVODeg5htJJLOiTu4d+u03D5I88YtS2nLExuhgp1Uongj8XOF7XT7UjJ26zgfgSDx0AqZ6vkavyy5GPkEAbs5SJZPy0aZEFrg05+rTw8/7iM6u8Km7nKcZDQVDJFUEkOLVIMl/OUPunkK6VM45Ol2UnN8gW3oKYeDXjuwUyd/A+kYvLkdEC3CixMZarpHEtu1jMh44TlgKsaMTlnPBjngWug1kw4ZWpPW1Xy/tKf1nUbxG9B0LUrY4GKhT8qspTDV9uzUIfvZ3RQ/ffoprbjEVm8BNcOvIx9n/+a/UUFfMYjfCy6EG4S+kuWMPweYDZPzRB7pZtMU2H5rxRBsJMMtmIYpLWQ2rSOu4I5tai0Vp5ui/N4lqhxw2a+8vff9WwBSCNYafK9Ch25KuGJ9MUh67717dbz6/f3WYWfd9AIosC2IpvosIOTWLlG37fwO0xqaig+fKunT5MbYtYwfmGVrsg0F0KKUoFuNjZd6d2z+xX24D8e9JcmVs8E5B28zJR4RM+/0xS4YYTIWAlD574JRQAL9EQyfYRQlzFGSvD7HAldjurMM38DiCv0jyPJhwTLZDFqaq2y9UGMXuOK6I1Gc6Dhs1gv8JDBQoG3n7Eq2496zypclrKGWhxiIfnZM1EIqtJ2rSVknxLIzmAinn+A4J+YL0DiwgNM/IBpQMl+VzE90BFzgHLXcfIBNctcNuTBnus4pFo/6TFxXucwy3gi71ZNWlXr3egB6xqh9wSayaHlKH6M0sn1Fvgq21ZUhl/T7wzr5WnFmfu8nW4v9vE/Df3FVtMKT/B484ieprOf5z90ak0MmcfH/MZ50To68xH9t64EDpLSvNsIb6fTXVlOSc69T69bNqk1gaGPeU3R5r49QUVha/UewM/6qzIy7nfNW6bkFe5vFuMQl7kD0LrQzIKkZdMyNEwORKUijYfLCqXW8orNbS6KYAgAfRdGTss/LgCVi8HnUmh+6Yc7Nw4GYixoMMj0ZYmIvhFKjd2Dm5OWYXmowBUGH3WGSsZxuIVe3aPFNmMZNpTs1J//hCUjx/+hIfwYvAS/fF8SvhIKhDcXOUW/8KHFYmM7bOMYF705JJpJpbqSS4Coue7MakzodQZJ3EUiZ4Qx3Vn2fx7HihxydYmng7AwUb8vBZCDTUAh7LL2oy6V4IUBoVTKO+eSjxHDcOr9pTZhPKekAjJziLnmWRB94EmvN7pV7Z7IM3bK1xuCl7w84fDkfZaAs0d+aVFkQd5Ax0O70qDQmq9pJLX52cfmtmRJ/QPnlsLGzhDUIHKbka062sFjTI2B3Y3lpc++iFnmLWjt35LB1HEMZK1wOvYaqOjvSP14NUxcFyEsBVZVt9YgsqMfG/TTNeUv2I6lsavI5q1nA0ou5UvwMNTU7pNIHnm8QJlVc1hhQjGdinl8rUCySmVqowmFuF6Gd+FLlQEfa78z0ymq2VyeoeMJ3WxxBsg5qwFwKqtUKrBGQeg62j4Mjv+Bp7jhwXMP9OlZcpayDWPM9ZnVIWkJYlPZS2jMF/h41dSXhXA2okIviLLK+dsiEuOgKEaT6sV/ezsugdeOWKXXOvrBUxaC0TSrzfuwWyPHNmehMUedmQZSFTTndPXIsboQtAuYBGDQJfJYCw833ZPRACMuaotav7fnHLwJ82jtFSCW7Sh1qHl7A4DXhJulJ3vVDYEaWNjx38iHMDluGkEfbuNMZxAyFahuCoEEnwXrbeOoLT7lyVQxbeov9y4863Q/8SGKAWImUR9umYdK6uXAfCOeCzaGpZkB60i8mFX64Ov0eD8kRlZFEp3Xw4u7bdJh0Wchx9q0VM8blR6t2P9cBhxLSm4EoWVXG2Jrn8LlBen8ybH2Iy85AAHNY0JvnCrxiyhHTAfEzpaJ9ggpdFEvwJF+gd8QAuL2iVzkF6RAy7YdR4ide/e7P7sbO7x8Xemv7v3tvIJdSdijRPmcjiZ/aO8yF9Sq5JKcTCGvZVa8t4cp1V944g5fB1aArYCQnLp4eNtIWb2Jf32e2z38AJ1Ouxo+G78lD98M/UTyPBdnpm6PL4fEnkB581cqR/NgCsPQ8T5gWLFkSp7c+ffmn+FLoSEDXsegBr7ePflhxBbJW43q/A3XurxCHhd7H4fi+nF6g3hZLtCUNZbCKnFi8RhFGCWTiiHgrGQjhjqDmgiKZqEFSsFYPxUw5awrZDk3Mq5/jQAmM3opavNiQTDzyVBHtKmC4Ye0LwZFw882jmwiGeC4NvqZhi9vJ5ULUTD9PgKOPDGrQ6i+fcbGuBYxMvi/cC5p5aBhNBNWW7TuCSfKSV2mRbyyT1SwRXsomnfb7xdqnUsmSiNhgcAC03gwKVAcWINKkQ0F366Ej/yb/UKdOLQPt42EnGxmy4EcftL9t3NeMMy6k9ER6gr4MM6reuAJ6QfflAFfJhxLyoI4AbnksMFj9JX/+Inpmgi9+FP6NrfPTxf0fcrJKBIijn59dSVD60XeMsQe2xKYfWCwtKaOoCfuQWorD0pBFjDi0eg0h8Vdmzxd/RRFFi1YFIu6B7cZWwY4ARyVUPv59Bw4/nn8GiRt6XC17GF03HGCs52HqHX7I4K1Ve/zo24J81b9V5tea8xY1xSc0sQ3aY3XWsWQ3VfFq+JifwIZpy186gdXRfo/6qTC8CzglzekLSEXd7/do65wlEDbUTUM3uWFunrvHs6amElKo51o64KD/aLnxAZkW7ILdOEg/TGk29OZSL4r8zwFPBMAV79zlVu88BIcMZiUv7+OlZGxEp50PyhBlac6KSXSN4acJEK838+rOypnQpCNQzlbVDlwcHcByYtwuJ/lx/JsiHgphKIiYx87IEAHNOjpwznmq0JcC1NY1orZcE73zjqa83+2nWKOLcO7L2d5G14ZurORD8N1X7smOXHwqp5HFwhFqDBQwAtptc6D3tF0y5c+oM49eiIJ35HrCOoNroX6lfoj6W0Ze8pQ+x+ARUbjs/bJvoL4ePdkHV8LgDVtA46dY1QETwuQdGNpnI3WfTRlbh2r9bUaIaJW2Pg3dNmv+oOivdp42houa1HYkN8TFmpunWkPLZsKSrYE7KhKiuosbigLwxxAPibzDgBMwVyWiJLrz8KnjmBAQRUqaHbjvbqIF4hSYc5oVWSadKVRNkvy9LliEq1SU5hP7L1adIujILiHOMfIe9TmNGycgq57chcZpB3cKoSP36muSSJjOMVbwBF2Nuy6/DpkHHvA3dKxi1UdtuU0/VHRZWsX6Qm/7R2QfUKv+dsVWd7XN6nLxQbOtgeQFRKHeLKgTxlusEm8iuOA6VFj6cmlivP8BvVmu3rbNnlDKpxlFYbRPSJgcfSAtbu7hgAcAmFHpG0SjRMRkFUPYZbTRaffwv1Cw/+c2y54fRhOj5krcLYxbi9aITpaEq5jxLkjW7iCpI1fPsOsqYHx9VjmLdLJ5pfL67u7tmoBwOALZ+7um3IVn80UH7W4phuj6gIbOws9C606Zw3JgSdmJ1DYXNM1ol5b1vsvJG7LJUa9jFzzq8uD5GXtrS0L5QvvuOT+KGjSXSQqanvk2mf+SGZ8z7jqdk2AvXT/pWaYJdePk0Hnm3TX+LbnvinYBfniNpJ819Y2EVAF+m6m02jpUAtFDj60yH+NE6vlxW1HOvZux38bKESJr9gwh1Qy0194L+FUmcm2lPyfh08Oh2cYjj+J8S0jsmnqhO54wekg3ebnAT6ajLPQJd5frSZfk6ppH304IgM//g50ZBbJ3doKHi++3d2BGg020XRDAsVNV3VOe9I90VP4sKDhqg2IIcqRZVDmlIERgpzEQNdknMz5tdYMzVY1OV9jgBzr1MR40RU6TEUhfkYiwgC3P7ukBu+G9fxoo4FA9cP7H7dthkrUdcy7lmGR1PvbelRFE88iPYPaZyoS2aZkAI/+KXmVLD+Zk9drOAREM8iJevj77HawGBX+KJD8IpLKXioyS55y48woWA6pxliPLvmdP6fu2VNcsCdNzNHFUNR5XcnTnfAy6jyVODPgnSpXW1tDY5QLZz3IxFgPQ6P87XDbiTDHvpqe6j6il1y219lL2DjdyJSCboOFhLjWUdguhWh17QdzlRR2jjRuTbQtcBUiJbTcHF4Fye0W5SAlnNmwFF94Zqpe+9uAABZ4mOsbn+3NsWWVIKx11T4tswziqNoppcR1ly+7zAq7YqJWTz8bOORqvHuKfGiewqj0r9nk/GoYHl6ivsoUodnDZMUEEDM01wCwErNMybuvqR/UqYiXI3YJ7bCaTIc7Giel9efti9D5ySwSys5k1ZQJbxwcT2Cd/8gfgPiYAcuLtxsUPJIGNLg1O4iOU4CEzHVMzMOkxNCDB6N+PIB0CwrG+4SgEW8Hn6RZqlpPEFBOYAMD9MbZ++Jg+nY+/fSsqFX24jfsfKBXu/9B0Nx6FKN+nA848rc6RxRFEReRjMbTXoGeD+jF4xGf5aOKByLxLo8CRTH/JCoGXTGF1Va6mqAPp0HhmwwDTJJIzmvP+f0YDzwnq78qCWo8xPwxQIIYYrV459sOStZTOSi/sPLIrkVU/o7iUS1nmP+TlOXwFiRQ/AClLEu8mLtRKmDCo3xeryCRBeXP5l9DBJfPQP3XiIykMaTY2gEDqAdJ2chVaqxOaIfePHG2AhlQRX9dOVEhGQcgA7DzAnHVv5MI8U+v/rPcsqQkytqPlRdykRXRks/uRx9aaAjgC07cYmTKaf0glxBUc9d+GjyudG+GzdGR6GTJ4yE49mGXW9N74ABXSYXrEjx4V435wCG9i9V318gDhFJgXPhimM3Isat8GgcgwLUCzy+TTJKnAPvR1BAnsCY7C6Ab0GLHpJGAVUoGRPoeXj5IzpTBBa1OBODrVKPRImBVeQSN5/IHGqD5g5XzsGIREsKBv1ca5bSo5hQ+3rKBxG4uEgfLOs7iPhS+IbXSII84afwYBscCPdG8T7gRgAxZRC5iDdf7+ags6vroV8grvcEYqejG3IFqLlGDPwCR5MGDBE8wv80+FP8E1q4ekV7pj+SRjqNmivKCHSb/dTOYhp4ggkbsaU9Tw4kH7ChErK1AAOcz3M/G2CksdcenUIViHLXZtgsbI0dLZr5BoXdC3AjsWK6AtnZnj2+ZDBN9cJQH8uKYKFbBvb/W8q3gxmzRSltBY//EbOOxZtE8GDlTn/Dpo3/1gAGBQ6G7q7SvlZ3ezJDV1NX1yLfYB5j1tBiv+Nvu8QK3sz7vtC781PP/QIXZXxYUHNvLdCV+9UJq9/i5fkPnfRz+SVZrhDr8GM17RdniCoPEyaqUpJWwyCWath7jap+FJ8bn9X72b8qTmVgmiOcBq39gUSu3fEE6echLoUcEppAoBD7I0UFk3qBzLxt15ebNTe7jGbsUT1PSl/JvnH4pTGfCESvbBVgNgRYAbbx4OOF4jVzial/1ECGqQS97zCnTyY0leboz+hrRJBxkcIeQeZfoRo1YOAvcCFtNwxZhPXlLk1ALPCivSaZHqg8eQJNUkpqfXUhhhD/H0bKUKNauZS8dLIYfZO46CeQU+Pp6u62jVj4L9c3eMmXSm6A5Z22MjhPn3X3yencBwdYEJNkc6IYNAr03CD6wxmrsNyQoPjOMlOBcdyi2CXpkEv4CrYt76a0US6PoXBD2e52gWN14oESk60cJ+jmUP0NHIGJIh7iBEXjFf259a/PHU9suTe5MMURqB3hmJbsNIbsC0Ox4/0+9CeQPBQgIz6eZS54q1tUiO0e/lpeBAOKpAAQQLZFQvpcsjA2H2sdWzjrPvwzOcrsiYVHHjU0sbvG7F21PqKYJd3X9BBpTNbjaMrqW9UC/nBGFRdwk8vsSPZButw+5ro9e7JpjSX0ZQW3SLV2BtOz0Xir3mIK8hv2f2Z7rynHmydoVfqaBdfHzPa3l2aM/5L8/W1zKCntcyfTrMynU1wnregIzQQBik4fzAHL3ZEB29shR5T+se3U4Upuz2WVwnzDWBwM23YIZCEeAQLK/rFftMm2sePLYj0LE9TSLrboIFLWZaclvbCkjhg69ouw6ojuzm2MzO4hTx0uupVr4EaHJ3FhwXvEyqHcEhc3qMrXgFawnfEwnGaPWrkEnAcjzUpSlzhMF8iR+oeq4lnf3D4FgtDWEgBDrg8f42G485MgA+mvoZPmVwOfLks7GzIoYIzaDHoGn8UTg1ZPFtoaHQM2j6KK1w+evK6RIAgjsH3CYAU+Lj/PisiRotCiu5+LTscf74xZIxKCVaJaTwrQGKNlhO9r7LSSJ+TZv7sJaK7chmv9A7EZY8fFZzNVb+0YnQDieWWRFAq8Emz+iCENQ7V0Nev7PQHnA5kU99m4at1UU5/0JPZuqk1n2sKE3NFD1qc6lHXYeX9Cq0/69rNH2ooYjmo2BIEY3HhBGK2dlU5NtfQXiRS/nKqemWN0DNXff7GTFPRDoeE3x48GQ2K+JOG5KGH9qak7LCbLJVhA7+lLngxW8DXNoYis5bllYiw3Wat+uqpi3dyG6C5sfxolCaM8fF92x7uU+4N3u5IFTyebATsbI07usZvwYBY9lA3zKpErq+pFiyUMCbjL3RaVl6AiKEdMJncWe4KcCRvnYG9fz1zCnp9G2zwwH9T3z94OtDdTytIhSs2wFhxY0dkkI9nZcG20zJ0goMxwj4x4IWQ1bM4oupw9yrzBGy5BKwQLQQG/Lv1u/M6td0I5NfO0NcnXbDYdcChu6FfHu8WXZNez0K5XldpsqaNCBryHG7FPQ4zSRkiZkR3x3ZUcrVSyOh/dLca55XWQf43tXW2y4wJWpcAuQsk9zOqVVSfy0GldkRKHxAZor5Ngd6XJtwC3eySaKMldf48etUnMc8ZVqDTxqSWDQZs9SOCoFxSKCfsHYw0enDozb7d3fdlXU5+4Ei56YtyN1eZ5Y+9S7ly4e36m+BBPvEQ3CRJv4ykiz1G9CopmsFso8lUX5r/6AKmeHLTIHQwHHLrysZOyrApaE+G/9IOEnY/7FYw4Aogna/C71J0BP/qOWUzcXr0fXtA1vukk8sBATUailnR7ETL92yTKuZxel1QDaor9/eNmjuXilqKj4kq1novSiJ9TI06gY0kMqj0jVR4wop/r16Sy1KVDE6SGESi63P1URWxP5MzhJUv9qYlWGZky3zdBGoyfyUCVTAZi9UH3c8/X+9t7AtQ9kasYGMXkYFKIXHywe4U2T4nlGXlW7v6pelB4Ojnnhc7vB2opBvHVZMoQ4zZ3B2Wj9PPhJBCWk47fI0Br7ieWgrs82gNEmTpgwjX/ZEEDL87Ex7caWaKYN2t1JoCYOreUWlepncF9AxIr6neg3spw/coWW40H6A/Xb2urE9DGh0BMnIOvO9WEyv/BUZXA0VTrV3gSD3z7FgVrC3oHBJZAPe1z3A+V9WXWQLgRIutLMynxqyu2PFfi/6lwjsbKU8p7ZAkDL8/T4Fr0qDrKVE0pvYe52mIpkj4KvEED1q07f3Qz47R1HitKWgegPz2BShlnn7TvcZV8nfElHwGFTsTFbV1jQsIVQwUUS019eaNcRi1wrf+VPKZhr4nlYo+dr0MSexmpWBV8MVN8NwfQS+mCY2tsH0DNwzMgxHCYbl5j00yZevRT/RI/2DJLiSiXZRdaDMYgkud2gSUoSEpOwMKkixvstP39M5coMGbOpR262oFAa9BDce6kY0ZX0g4yPJqjH7idun41+a1a3ceUr8TUX+cIoUjLQVFEQNFOQh6iqeMgrvaoZ7zbBDgEmoeqM06vdLOM//BfNjE2RiMZ8wzVQss8UvExOnCaVa1xmDpwIg81DcL/T70kd6aYqLxOCmMQhwQ2I45j+bwUVScV+cjUZGeVBVaT7uDsXnHC/Mpr49wir/dNcFq8BvGC3KgNRZKle7J+VEzUk5auPRbGFFmI/mnLTeGvcazd72rfPNiO89vfG6/dgCndAwoRszKREbic6XW6c9b7dnxhc7SKr63ZC8WBaWeON8TiPBeAqf+NnjQ1k5EDF/0ziHCvT74ct/jZWzlGX/Rt1P0PO7dikL1Roy303jNto8fPRNTZM1gEVd2s8Rqvi8Th9wje/353OJRL1KLYQo0rhE1+vNbILjkqFCwyZfCxAI/dDt1vHxfCmutYLwX4gEGXXdnOuyiWhU7K+GqolTUORyH0+HIehfa3uF467cBkSxYG9x4pS73UHFXvbKRce92sCv8ocJB07UakN3M1lPcNWlgUecWv0rIvJkkYwhphifmsvsQ2TQbRiXBCqeDOy+2RXWI9SWdeCoCKZluKrdMhPr1cbpCMA/m800uLXFd9Wd1vd7UdHRbM7Cx1KHRkCHb9DqwKPWdVE46EUac8TGxbyFGAqxhF2tTWGbIvTMktS0kJyE9g5iDF12gULxACYQNk4p3t+mlVLSTupuzsCdtR445ZPG4ibzQS+9xR8IuhUGGvtu4knPXLVXeU3bnm+FVja55OB06lq5rOKXv9LzB6VTCjVPZfilA/bSkGNKLJc83nsC5qOyE4dR/5v6qi9nPQf7fGYBAgkFxPI+FL68BjEOLsvcSbShrA7MZH2CEfbA69yruoZYM3ZVCevX3Q3GobTe1wXN2wDzRI+83DprHuHcHCElA3Vo9xME2m7OVUbEQEiMUQ1rAvOXLkVvykrpsn+YRO64/RJ5aPVi1vQmUJpRItzwiqiBJUL7m0tyrGPglZWyPeznfjjAeJ2Gm6IY9I0/ZZk2uQ0NlwNvKTzQj0j3RIphYr2ahKKdWmYSV1TA8YCxSrA2VuUURmAKyqD5q7ScojYIoBwj0TI/zV8T01fipKxszmNm5K4d1rjYFgeMeP3VPN/s2w9NAAZECCpBggRkIIIk3FS4esYP5izEUCDYThQ2w0FsYUwgpvT0OdOmZ3DHrKfaLFol4N+4K3hIHY2PZk4k0GYFZo2Ry0hC20KCc8GOX4IX/dx5mE9LSf8TbX+ElxCsdkUJJOmEDDQ2bZV1gPKYe6pTRKiJGDjEdUYeuAa7qlqF10+fNfjF9lezgho1lEC8dHSnjODiq1TQiqyNItylEdFWzxbCgS19Ih3OcYftYLYUM4iBb4oLRdgCiValSCjV4oYyXxXHy6p0uJS7rbmFjdIZLc6hfALZkQ9G23gYDEU2swSaeVwsEu9ZcJGBnnCTWkX33s0Kdz1dUJb2B2tLIZUKmPIOsgGDDyUzD6AAn/pv1P6fzsGtUGXFcnglaqT3q+EdW3xoa2mz8uebiGx9NREqOdQLbHiEld4Zijjf+wTYbJsAtVth4LonJPbeHAHYv8cQe+gc6JJloc2uX5pg9ouYWkPsnoaYnzDcU8gSW4qTDl/Ndsihmsq755BdgwPxljytCgPnSY6AiPhSKMwAM1e7U6QOJxJhV3JU+Ay1Wi3WVpvYJMt1qpVx6GZfSRhkLUCMdB4ZbpDLx2O9SicsAoLZ3FfQK0Fgjt9EV02y+rAPe9qMupvJLLZP5JnGeFSX9gcE6tYAj6OTTjJ6BTRoaubSZVX1fptoYtiTdJ/3JW/R/YL3RabUwgh7Ms4V+x1tyDdaB9calbp+J8m6yG481btL5XcQRcs11o+JkmWmx5QMLfXtoMz/RVw42bdqJO8oRPhCrHhr0URAqLquiVHREwB+tVYGxKGocgxwWC8eODq2a8W0zTrvE1twWNbqJ1LY7137eQazpwvB2X7W6sDhxlimz6nPTCKSenhdGEXBzjJ/YT0ViX+7MS27027qxVBumx4jqgpqzc8EmrahllPDx8F5nnen0HRS6mdj8B71EaRSzwjiZOcawpH0Zfc4kG21bQR9o9agJXFODnQNtRZ8q9MCNmsu0qp3N/oRFlYwAb4UKgeBqJdMQpSro02SNj2gAez53qHjgUX2YUwh062SE+8FSzKRyMXHDY197KiFWq9RvXBKeWUSlv3CV2Fpje7mBre1nv44O9CH+YBDM7vPHiYaoFc9UHaQI6hOUa/8HvHzf3LpvBZfDrCaP3Kq2wDGfEOjv61/7+ex1Nd0ukZ5TmybU+AYk/p9xbJAEagCR3ECQu545yVCIfqFu+OKIHJ+jp4PP5SnYWgCYYtdyRvL+knPpmj0dYtYmj0XTmhGjZG3S5WNs3FxPLWr6XCcwkdNjprBLm8cvWg7GEkJa22WjEnJh5O/vNKyXKKeKbfDd5vrP4BiOxxubf9sCVJxrGkrF17QYYmdo+LaD5e8gqNQM0FTZnlAWqBRIRwHuOTgDldDTVYwdKCGRG+VRql76FaVAol2ykCxM1inaIpHYRkhieGtY+/oNBtyEzITJs3zVtacNaOg5+C7vyWMYXU5XjpnHCm4ogES8CebHSFApyTEvem2+MnLqvcEdIkX2w4qTWCVTC4T6n86W6/loLFWgJoZcxV8y6Q6eCxhS19ggWf0trBw57DN6gIZf4FepzJCEcbVDytdqgwJ4WVKXaFj4lDJ2MPr6jcvRLbRSTHV6MvEX4vuSO81aYkv0LryUJxVbdsPmzO0JVzxbXYU2Ydw5r/G5o0VaxtgAM3hILd4TVoFQKmJKcrSwo85H9VHUig5jPmQKDnCm+dtsUdzAyRYJmzVd0w4En3ijn52vX6Gw+A71ilGwyP1FKFxzdUTSHyrxQtlvWOH/qlCVlqiuDq1G5T4xxBQ21UMQ6WuzOCWUZme6M+o4vrxJLucLLJ7TRUp7DCfVp9Aa4rsIFSxFtNK7lqwnsRr+b0ONhqbd3n7ZQv9L3LIXvRKkpFJrTQUY8EImDrUxqvHGEN3vdUIjEwSQ1N2JELgWMJGlm4GxXdGEY3uD+X7sDK01Cuc3wMNhwmewL4Z06nK7xrOlZWmDPRVeRwrowem3uDSc6pcdg8pdFkFirp15pI3LVbtH/SE8x/Wu8Uc5ZG1coFcIstwjGqaQhubf7kfKeJBJwv7UT0AfenPT1/lZvScsLWIQVkaiprmbSl7wlbTE8l2bzCFVyVRb+V7C3idXYcDM6Q/JAp8DfnXr88xbe0In1U7mqia2IOl/8r765GQ1V/YJPqfb0QXug5ENwHzqQ+1JGVMg+Zdb7DXA9xYrqMAGn24hiXRilD14FrvAWaLdHTTySxPSN1Fel/vc0NvpD8Ct0rfvb4TSORoKRpEc3n0uT6pbKVqXsl5igZNDei5CCXY3Vq0Iq5dPrYyPZSTXm4Z7/6EtBgbsuEELawtO3+xDExhEWoldpz0RmxMOlmPWqXiG9875oyuIk4zJH5OdChwF1i0Cz61k/7r/zmvfGYzjD+tsbVkQG1W4d6I9OgMxwLLpixvdRRrNdbkKIOnnk7C/vXunJ60QG0ltAU3AHgx0TE3tTq/rFXEy2b1cLA7Ul+sx5qIuYNcr2zOnObxlE0SB2zXQWhTyW05DMgSolxX6GdiouDWVVVxRjOejTDfYgP75y+lx9HftGbuxyDHpwjDCBypHgDlLE2QBLjQhpMT3xzi4ljQp0+QLjz8rSh6DpW727LBt1524I4ZKTOJlzMUqoK9XQygE5//wX58yZtCqTAFBtIhKGpqtcSeZvCevgnXoCt86IjFzVqRI0w+Ycxkarh6tFsos7uuz6fcisfaWWKWBZaecIRcSnQrITzaAjkP2WMujur58fH2S8tnglvoDBAc//d+eMyTzIzyPPetOyZh62M2CosGlPKkNlSWmuQbLXijCrPUc36BcqDk3XiHSv55UR7gR586l/87rETQTacKGqO+awI4Dp449pkukk3fL/7KXxL6cSycli5jUXWQNtbJWYu/lB019TzPQZhKPuNmaYBLflqsgv2WUjYs7XzUF4geOGX8XlM2x30ai6fJvKvAgACBWD8qOj1m5Vs0XLYhf/t5iIJhza9r2VEruzziw/D7Vkh6hGbEJhjWV4XrkPVgh9Tg5jlYKeUuOE+8k0ONa/URo8e/WGM+OPoMkGam9TTNfYdtL/75W6Okl/xC/UaXd96DVx/7ogaNyasQq++UNSYIFnxnKca3jrY9jM9R3v6qfRM3irQay3dA4rEsLCillUZLEkoAEhv7EJGWcxbNxWEEtuMfaqur6wxgkvUcAlNtpAqoiGLNelElSOJBGd4ekJ9qKSnrrWskNhvHtK0dh6HsfwnXJ5MS/NJWMffkL2LTWlL39aO3zeqW3NudCR7lTsCLG3XaMIYgixxwMwSvDIXX/vLtZepiUngxSViXTiaAiNlMGTGWc81dihoJWC9uXlhg+EzGTc8dLYC2oWI2seWri4B688Zjs+NXStm346R3oW99CSKzcWuD3XOf0Ap/73R2W6biux4ywsLfzHG4RVmMuIjGuBVayIhMkflW49ETnj0+DNYHnwpvXDBg6gMAFWA7Qa0rgHPuc93+rg1V90Ih79Tm+lQcvpUS4U05JY2Q0Oa9PpS1uUFnGAL/5PsOUIX1SZkcaRzghI9HInB1LdOj22MxNyB9rPz3cMBRmKrtgboF2N++f7zxFGXmUpLx/kMjWoQVncHsVqlpRh4NsKRDI+e9ncX/APE0SGm7/741C1xfwVHHZFnqiBLtsXyp6AKViJwn0M/L/lMW01+UAzc8ZNe74J5C99Ve7d/+lITDhxgz6w/thkjYBboY66Jk+J3NWTiY6hEm1Bc1gH/yZ6S/qaIE1rFMuwNTiOrHmp+QLt/bIWip4jO1Ruek8+Xv+kQOdkvBfYMFm/BrZCfr73M9/6Cd2ndKotAkmqH0eQWiAD0g2JMrLbJCXOpb0CCHHx1r4uZZoiuHQrDMFzaJ+sMiysUX+ZjaGzKrV4eQxpgVIk45Pl1mEq3ae9RDGv/WxjOJis8DTPoDCXlzeoH/l8V3djlilJQcglFUJU+kTJGEO6c/JRxX/NIzl4LJGryxatvDcJ3FQO3yApQWd60hbLDABmhauTI3aqOEGAkEgccgO9AqhHamuHUMLux5cGJYDSLFPeqyDndgDOandfhvIKytsYToFQWBPt7ExWf69hta29Izb5PgvRYr9BDk1uo+fMVT/dFjesqdU6qlDhlnWClPc0duU78SSy6ex5z7QNsg6raohNyUEmgLUGatG2VpARVHUHd3YiqLlTIfDTgAzg35/h1eKfrXv9dcJMoVBTqCpsvMF/gVE8CEi0eRCycmqwf4K30d5Y2UB4VdRXZACfFOebiV+nBxsi9I67VnvA6b0Sb12mFIL7+GVwF2Px7dnFn+cZG3Ts1u+x9fjj+tcT29F0ELd0pLRTyLlm3vbHM4hGa4xEWzoBl9aNK0CbTIsHvAhBsqYlhVvc4DWgdS64WkBrEKSZ9c7ToYeH+FDmdM7yrQkutq2WdnU3Ty+7D0RJIkmFV+stSi+CYK66nZNp1CFGRiShgWD6nS9SPvqKtAKnEP3L+QFC91BCI1thSKmCeUvvrP0eNI+60lw48gvaYm4SR2FC5T0VtegcM1Qgl33Li6tLXgcmIEawo5sHxNDTZKR6ciG74tmRLZzAL7Ia20YYjVZtrsajb0AqhJq3tqnQM1++VMDWRtWKtbKr/M/TIRSG4Sf23X1xQROSLVOaGJuN1hIyeW0/7IwHMQbSXaJN5tEIaDUvg/ogoA4GoYCaN2XbIBUbK4uS5b45vuk3a3idHjxwE3WWWXPjL1KqzFFOr4piFw8eLdXEHZPXg2wYRoDFlzgsd++2oQs3VIJbobHHiiag25+vOdU1mL/8KX/eTSzPUdO4U/0zpqcNvklD77cSHty8hbWZ8b+pe8WdDXwIvZ3uZKZ+89nYhXGJzIP1V4aTn7MCfIdV4I1IvMLae6YJKppimQwBTc4TEVdHgQ5HiHJupQiQp7GehT+Sn/qPiCX6dIlXEMs5cLIUJr2hisBOCGoDnpqHaaPpzjFfuxbhZ+vWSDXcyWAerEdd2iHoHvw32ztcQPolwAl33fUrX+RNJYltcbrOvWK8lxp6p1GOZ3iH85gZJKPiknRdm232t/bLUALa8QrnJ/89NaHjGaawVzPnV3XgImmpgPQzpvE9nd4OjyXM5LEu6kpUOcJoLGzGSf97+CWdfe57C+KWdeV4ueK9UxcD39w280bHdy5wHmgMDlgImCzsid4uGDozXxV0rMOAeXfw5EyNFiRwT1qm093NxeoV3w4bI3l3kIuENxwsftLis5ETF6uQcfj2AD/FXL87NeXPqVb0axXCCSvI0F794SQ2VRgL/FuesS1iYZeZ2a4qnDPUZuazrEoCImOgndTa1tJCLOFZ8XzBPglaD60xReMos8W5f1JlhNNNkiC2x/AbGAh/6cUSzfKv2otR0zmL+8uKTaiYSZEOhOCQnZyHlyCAgwKysluWC7eCCMGKUOyugoFvCIvOr6AwWbCYzD8Hkd2pbmBc3pQOIcZM0djZ329Sw74RRsKeTaX33+am9hr/UW29Uqqfh0jJI/xETgWZxG54ExGKT+0Qv8XOE8YK5hzMT0aOiiEIRRjF8u1sajUKSTZqMA2MaE1cDUx/mX3so2KnXtaNudoCk2Kp2vTThf2WGjmcglzbpbht55PcOkJXbTiURLZ1Fon/gfi7iQp9NCvRBshiaXGPfLjp/xxJlruJ8jdsJvgC7Kt3RTJJWCLhdnWhsemRXPC2GBnb+oAw2uqgHcZbeeBH2rFuM0qO+CQOPh6ONE+9HtSG55eYA10O9dG6QI1e413zpfV9TTMkm5GlIZSslRDzApv9Dd3NjhbU+rMANblFLBJeU8A7/mThjHSFlFhPWlJtH1XlTD4S2SfjOpfFYrR/3w5bE2ZQfqFoq5bx3fU62JzOyxrFmAyccxUTdC4emxdTvmlkTtfVXHm69D71Ma9RB1z/jMzxOUB6fdI+gIG8l0XrFRf66jA0Re6WGT/Dioi6Txa1RJe3OmUE7ozujNcMYpb0ZSl9J8rxczTNJpu8qG5tnQXTeTBdElZ/l5EwmaXxFAFfD/ytRGa5Bv4tUvWXJRhOqmgAoPvyyDb/yW868CFJnNJW+6GIGFH3xmJUVFMsTUCtCjvvQFzG0LRYxkqWLHITC65Q3ik8GBYMlZLYw82/eb+ypY5ThhdjgiSO4ZZQ+u+0zMhBx8jjMRy2LTgFQ7X/GCXb9uXGQhIZ4tY6IVrgRlcLrI7L/sumo0Dv5Xr2QB79UlHMSjXmCOHFjnAxxUdi2+OFyYeVH1x4nWu+ffV+TwScTbZdfI/G5ZfmEtwEBAoXQbtQRCfuaOoxxDkR9tm7kLTwtK71r085oqyp0CuU+7Md4/lijwXabyfNWgRoWdFPdu2EjwRMDLpfV+4Y609fdMuvjomCbcaMM2ZySTcfJ2eLdPY5K8GZpXRv5aFtOy/9nSD+zA8RcssdAMOGtxC/+hwJQMoXf+bYbBocTh2Q/eV8usnLe1GIOIU8+E1xcP48Dzburcr2VZdkfR89br74hcHd2ZM6zKpqGTxVzeo4UvrmrDfEwyrLC3UeSNftjaShyccSplUd8TTJ+g7xjI4FFfOIZbXR6jS4wKQ9zToYf3G8hqK9iHnB4hS2zFcCIRXFIw2bLiDf36zXfWlmC8Jhrrvgyx9YOzIQs7o0WSc+IcfE9jBtDuAoYuAzCAD6jzawsfqq687v8BtXfDd6gAbnld91mpMCYXbwomyJJ0MXZ38usbd4aO+BGq7Cq+lv096MGxAkSeqXUEjilDSJeUmg3FBVL7NOFKLxzbq0EqYfn6z9uv08g7i09qOTEox/LAnbzjbOCFD/3NjX6kzjHs1gjWi2mjZWTYQdxdhQyWMD5dcR03ywcR0JZJ6KnkKoqiQut4sHLLWLoalMYzaEG1Hc1aKC9JqMzCwcAa5n8Sy8DRJ/VHEM4HlZYzwkj69cgKxhQXAv7CwjO4koJkS2TjHh0nlxem1OayPJYvOr2YqgKwviuGoIsc2UP7EMy1jfiB1grEuyL3mauAukxAz9mT/S2e/+Bpt7EZesZIryrtcG6DmehreDuG/aWEUKbcUQdm62YwqR+np8lAF1LnIlEFriAGDECUYIyXQ+TlQru+6PZgA9NMNts1RVq6ujUtEbbQziBh0EvhybvspiRUVScKZA8niMTtOzcK9YodlJyZygwY3y4JjC2+ST3oKi6DIyD1DYki2OqMBAp6fRcsEGzH6oUEXNr8udfHXQmE/2myHZRUBY/iMSTKrXv6zdILty3MSTrC1RCEZNmmzuYVzTjuqyBPy665BeXnmapIsb6LCPh25A1F5ULLBONpGh8AFqUKTMxcf5dc/1DRuH8k/l0mVsqJaxUoEqbT7pdCAA6ViBcs9mNM2KiRdAsguQBuwPobwdiLS3cBPYnEZa00XANFZO5GAGjcMK6QtFVKnVd/iPpLdBDt/P7Do818Lzaf+zZ8a2OR/bGpMLx3BdQ5KVbubdYFck3ztJ7BYAAqN3fo7Y5we9MnnK+rYcgJ6qm3HLy6FnzAZLqQkyJqNneeQYczyRyVDelImpjX9BWoBzTL28uQuKmYPnVXc0VUqE7PHEUJc8dBouYsMhs7bWLOgTVteNYLMzmVaxahD1LMcxTXcqN3kn31HFWupnJUjVl+6nF5bEIva2zblLc/3tEENk4VLpBsyO4byhYZ+L75s0D3zr0WcTDsIEz1gJUbvwEaLwDLW6ovbvKulDxjPEGO7OeWhX9Iah9ARwpp65i7X1ABJEY1Kkj1ezqJFmKIXDgIevKO+macH3GDcf3+HjisYVvuYyth843AydpkWiAyMGZpemrWNj08yXaratSmJI+g4KvQR2sA/bUIMaC96vubt+10GNZLMklRyA/qsQa7txWY4RF4rqI9WfpyMpRKJeZHvgp7UtqZVR/1yWpQ4A7DhYvj2c/iHF1o/tK0A2fLo0Xd46Y+QfCCeqFtoMSFcsyq+6u1xAi8+wM/9/Yy10tKMPxfJ84FBV7Cr9olFBhMyl2Qy1XAjqts76LLrpdmcO1QroEJXKAYMYdAaTndX7ojlCRKshMlahGr9TSf3L/eN8FGJ+mF62xsis3Px7UDpnvljAjmZ5IkTMMOF4o5YHqVpOYZ+bJoVgCcBU/EpbrWNQen2KEGLf1wnMQooVLt+yEAT0ypk9wuHLCVqY/2myMTi89DY425op3VLdyZtktsJ9doDzxegq3mILm1zV6bmceukfIF2xtb5DA+HZSZp5pVfPcTjnmSDs6a7W/MwhxngVB9fJ3ipI/t5RNhp4jOC3RBHn5JUAfWF7YyUidy3HNGqJZih91i+sFNyz5uzEaezfbHI7ALnzI/0c8KMKYzcZnGQyDv23hrO2yA7kXSlymsHE5FQG0AGbfhovdIJUEOLO9RI4LZF1I1vBi+IiudpFESXi/DXwQ2qti/k0nw1tIC1W4odtxBPWzIruoPXr7386prPucqjCgSuDf/WhhIW/7211+WF+tRhDlLv0VCiw39YSbRVRnMWjUGrNIfY5uASQjVG9PM4KBoav+SRUspgIiNnbsO02gXxB+uv6ui0Uxy2fDx2dZk/0Ex+a4HCJD1FsJaE8k1W/bT7ORpVH7dNBQTilXzRREQ6gzRIYk8JzbCW253MbFSVWn10VjlE2xNlFnN2xPIXY2kqKPZQJGyknQ0rb53+NsujF2RPSoin1/k34G2oNaeklUYNceyMFrYQ3vBKpO6eedmExJojdB9sUwrBpn+qIEfL7MFdH6ymedYbnqGl8oyNXPRx5XQGXJ4/wDWwHZIjxVsIdEzvcnAIlr1cItiSu7OmDzogWzr0WkDQ2yUBCWGEnp9Jy1sBY8hb7vZ0Ct/3OvqKtK94DHje6KD0H9iS6ususiyKcFJCWkLwB20GMEyMjOyHE2iNKAa/LMh/7q+I4oPFOk//cCsvMzL5kUs9+7wLURfsRICSemNZ/PufWmcTV+ghqh1xBBYDnTu13eztmw/DPwjhnHglVhmfUuxSJKGURKePrsBJx0l03Jmp/iMZ6hee3Zw+zTXWjvAwl5Zs7QxJgvJlRwekPEzvvot0mlbl1gVxu/lzDXqV0EdJNXOMEV6wzizlyLTdJ86AZJKQD+SmF0r0rYT9a6GEedmVJ9c4wuYgYKg1JD4IMh70Gjxhupdt6u11JPSKB6CbRlMLmpvq4uwPM+xWF4Rsx5xH2BRaqO3qP2y100+1iLuj0BYxGEXZKKTi6Zj359LRNZmjZ/20ILfsvRhyid9JlOcTTCJ3wFAsnfpDWepZnRTyuS+ybzZhV4QO9O+ZBRrQpKhhYiiMoNCzaGRguwS6StggrOiPoHsgtHsvwc+bKoPlYqD2BgH6k4VR+qWecQxk8PjdN+z1vxCfjSmSQRnEB3eP6noYw7Bt9VOup3nDaWKRLvgXY6/gCFgPkNWf6uxIEmIDbHHAwOoN73bdQebjCMgkFAz2wB0af/MSiHD7c66xNZGj12YBg9bpWa0pMWTySHdX54sRt2CbmsmlvUeMVAHP2IVZyGBg/zRaVgJOZ2thv2cHuxIXRgPEHboIkRU6OdtAMTL3gYnmoy1tuWZeY6qJhBvjWMGfUgOAOaH7auMgjuHJZyLYVmtG1zHk/mTVHu1NZ/ZXAnpQhQgYAz2fjojyvEpNz3OKPJBzdmEow0YxI02VaZSQbMgiKTvpbqiX+rAsE46nsnCynCWZsNc2CDvO7d565X3QkLCHu1kSCcWvOCFnFvSRKWtgKCCEYFE7vt7Xeo3uhaYmvYKxzJAQ9JxB4sb2dHZ+TPGffHN1oNzQ/uG9tPRBdR9Pl//auwLCelRI+EpUvUpaQb1f7FQh9MQcmUtZCHtnhscjdJ6jsRX4rglEsDpwWI8WPD0E2Gm6P+SYso884WMWN2NDZYBVY8ZzphkmILv0iJq5mGBBMeq/Nx057uHcSEgF6GCxfJAVwBmzFCZmaP66ILNuuewbeqU9zmZ/DTILPr7vobm5xwP4rSMzKypXk5aLbjnfPSsnWfWIJwg0l2x/lIPVVy9MvBeSHY1CgLRWY9N2uf/YqY30EmeUgzOnslGDvcjf9nl31N1MzNDh5YYhi8tfOeNGdjcIEIcR4ezm3YNhkCQ5XA2fPA2mLhLTUCPejKW1um/iL2SVbkafTzWnJA53coh7lTBV3U7NCQ+7zND021vBxpr0qtKih8Z2YPucs2z60wJGG5PDpvJIqlRDQGl1nENC5CJULnSKzFCxw/WJ5EUIcrEQN34BB418eASlcJK2h/bZU16nyvEp6wahtJS76vtDLUxwRSRuWLMaqUQDwOASaJhvv4H/y/jBLxDJHrj8lT4jQGgrkq4SQMqrT0YyJ+uEk83ED2lpXQ+zmnmC+yjlK1QbFKb693Pt9Bl3T0gPynZOQc5G7WP/3KYp6OD68ECgVxi0bYq9DCRifU3ZvU5BS1aMDOjDmsR+23hrhnuiMe7DCdcr1aI+I7mJlYzOj0/boEAEYv7034hhoR5S3AU1D1uNA/GN2DeOTSKq+rqVa8OK0klfudJDiJ+pbGdTMErNqe59hNBMajHp2zhe8RSOmL9PxwwsE2jW0LZ5vYcumyxJDz5Zfib0eIlUrsFlvkN6mCMNXvHHSXCqBAg3tFCwPX3Fb03hdIIO3QnTslqCce8RlYYblK+helaEqEooV8pTg7HXTIbxww+5CvaXcaa6jtFnviaj9MWCEeKINuD4I9E3opTJytEdVniIvEVU95DAr97V2k7eh9OKMnXrLKVaggWKnhEkKy/N0QpQ4Kwjs2WiqjByTzDbWzy6afnlt2J1AAwDASw9e4ls8UDTG6h5F7uLGc/fH7BOsqQ3C6C3X3og73cgO+kFcUF1vAhVByFL+YpN66ozADqSN4AQB7dUCt4BtMHYbaM2/5UCi54doTSBt3tj379g98Jw76o89tERWil6sRvo6FZh7EWhw/xELNMFkoIhaPVbwFz9zUipqnR4NuB5pZ0KneZWR3uONacz5HjjP39Cztf+vKNbN2idyE/Cu3QkMvWRoImz8jNFahf1KmYYcAk+9T/u6Y5rxwLwlykGzhq4TmwnQz4rMfIlK1Mtay9ZTOI8zuRKx+B+RmUG7u3XUkYwS30lxU/KYz94Ks+4OoLOPvrchmjhAkRa3Km3Op0YP/OqHm9wq816o9OXyORqpxSxrcCZVM7f9R7ScpBuodzButhprHyWUt2+Bz6Ho7iPauJEWQbeZV7dEdHpUfvxuDMDpUMd3NNfMrMQ+b6Kpklu0H/37oB/qgUMICJbDtY4PARqhsfYsS4PlrZSDj9ly5zlSNknqQFcZqlmxCvSqWir8w4akMVfzRMBn0MqWMM9lqAc31yZod8G+F3G/PtreZs/kiWMt2kJRXv7dcGt2kdfdb0JNXCYpJT0yvpF2djp4wkDsT1h2wctJ/wFZpM1o49tTm4gNcgzGZVRlreKBbuUjbuAKGlYBL5Ejf9k9Akrj2dowAUXGFSqXQFHwZAkI6zXqZTFLw9E847AcaVtRC8QaXjA3Pmtp3oRpmFXtAOrEwVKZvLWjdoYRl/Gl14ovGWh9q9aJS2iiNSdG8wS45wqLJ17Ic+nNeuYyJrXqXnebhia4w9EJu30Uhj3yKoq1lNrazAachZvQUEFwzy8ai7sULEFwOCxOxNPuQfxLFlKHhbduS2cFneV+FVj365X/zciD3ppqCm5uDs121BkFoQJR5S+jXteH+/WJ4XUjq4LsdwcmQuadGmupgTLcMSC0uSydi5GBZmf3LNMEiqyamRkfepx1DORfY6t7B5ecUkWQCV6xGCvhgVfIaOT0A6z4JXiTOBpMVK2rfQ7IJ9fWYcQDJIooKwgu+jZg9lIwjGlgCTJzcBpu+0XUb+fh91A/0eTWlmCilQAOkWQhGY5Rd1dkooAnXyIl3eQp72lOdyjIqyZ0I+0ILOZ7Hgt4OQTToXAVwGayFwCYw7hG8VTKLPkX7EheBi5HxoAFikptx5QMPFD+lWasp0DDxmHdR3lZKUKhEZbJUrtHRCCFD4DSIbg93S8ug9uKWnNmuUOkh9sdyrYNoUHQP/Pn97cmxZrka0TrOc50gaMrTjM+IJ+UDJrMacH0zAkkGTYDXlEestTatYBEeMyr+ymiTKEH4GR+UGsj1C0SKizk6lUOSsfR0jbUnQqOirzvk5mfbylV/e2LP19328M9FrMhk5vnYVjCLmsiV4zrVxsInjGAXhgjjYfmmYHVRU8Ft6q7TDJycv7tNcrXVgWSMwbefO7JZQ7Re/1WclfYtMTIH+US5Xnj2SZCjZEdcp/rZsaSYFGFwWu6KQq2rdFGht0vn2R8xYk4PEUYQiv7WQirDRCATFDZlP7A5ezKOHF1QzSpH3uzLu13uu1QXeI4KFoqD9N324wlv8BjoBGc4iqPCS6zBl+KH8l/koGNn/DIyNhrboK0cvt1S72bT6NA5pttiZf7Djsn/PXbmbRYkcQ2Rt08I3+UVeuK8fGf0h4DoH+YbtOEG93fzxZUva6NRJVQjaKrVNrATz/NLXtnzBvDyl5QOqyGcuzepHwsHH8VcHq/nio5Dc45AiIlfaEmUeaQP5hTkI/z7vKjiPbWDbT+ahS2GPMWjONJJpOh6QwJlxViu1iU73/kdATV2/S6LuAAbxjidSnlKiopc0B1VI601ZPrIUht8xw7Pmovfqy0/xsrV1yfVezeh8Jsy04XVmYZdFpidd9bzuKAKFbdfg5eWsBeVEazrDGR8AbcYV+CxRLHYf3VHMODQVqtLzoGBqz1tYDvCy+Ey+1KE54ekTnjoTWSvNWLO3pxWNP8rCL9jidGgLPdcccnJT70Hfu6zvzWQbLo7Ny8VbWnkq5D3B7bYvZDUsJsF6CqTZnb8fsLjA0d7HqXFN/YW+hUJ0zlQPv7UOOrXMnZTKiiqNtO0cTuSAwgBTlG5/DgxxOLK+nyVDrXBnWxsd176dnmNzlnteq29Z4AV409LQHyLQU8Mq3BfKdDklNDiyTuttvYFzJgu1mL55Al/FGFv/n+YWcF06juTOPBDfJ7JD5itRnlz+3pZj/9+/NRROnhlhkaY5ix1bGmM+OKx7zN46f0tdI2Co85eqXE9xLpBRT8EqkGQX8W0NeJMbnUoBZwYfHyIFuKBWd7F8WI8tQbwdX62zCjr+hATr07kOc4zcBWMHEgJrHhFsqDW9RdXzL6IFo4EKH8+MOu6m7x6QeH1Q4hyYkHnhSBpAA3xYZqmS0ixJGVvhgUdUeDUzxXWQaZnIxun0wb6rpkzULIMLnZKOmFa0g/VeR8kXDKQZ/0dMcb97bEE3+jIwyRbO4QHymeSzJq1MnEynd6tjce28+nMeSVf2oQ216PMFVs5YR+ctG8Z4l8LAn66cnCVUS5jpopLCb/2CGRJ6C+H4xZf5XC77QwgHXx9J9TXY9kmSE0yvhy9JcQ8ub0RsfVQ1k5EjHA6fdVqBnpQMPRPASbMm01srf8LhznGFkgiQoltwreBGZc/qlvxonqsP3TpIV7Q6wPp8DW/Ao0K+KF7fplx9hCmChIqw7DPYJoXQuqTfGPrm4WjuMtwHYgyrDWf3tQLY2Or2jT+/xKKabVicBiBq8BDfCuJUQ2TxVnOl99sMJi1p2OKcrAmzg9xSElAQwPZpCkQerm498KBLTScdPOURsHjdvOb6s5AHgIXlwJNV99xZVgJb/ekj5AKZcDthibhWPVZL3AQ+Z69X7BZ5X0T+X3ZOL9bkEWGOvAnPeYyL60Wg7arew9LQ=
`pragma protect end_data_block
`pragma protect digest_block
5efbbf7368a2bfa7784e5f7eb48edd49fc30bdcbb5e30e8bbf286e3e58353ae5
`pragma protect end_digest_block
`pragma protect end_protected
