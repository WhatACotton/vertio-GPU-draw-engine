`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
c2ZrtO2VlGC0hI7Vo3bCmPtrm3oaUir+rCX79rie7tADuQUZv24YOwLAlcOrGQ7PXB9bbZY36hf7XAF83m4WpsGUZETp+ikwPWhYwYhpBUW2uw/C2ln9nsXYI2nY2q82W6o+BZLm4WP+mid+xIvoafhc8mpGDtan1+4wQePTtv5PEW6SQaVb7EOcOn3Z15JBsgcvg0WG/4RsIPwcJioR8jLxWJ3uj1VTqj2yzD4x+cp9d/NpuV9aRnonMakLkyzSUfQJkHEbmeNVYRT6TRwQGJ1e7+bobL/m5tOdHk+R968qq24XkLCb+AMg00FLlZEwVj2HD8UvzjSorbwX9UPQ88z9OuPbwgJcwWOWR2tDwdgpyKPjvGTVrYVW13ps4qaZUts05+r+dbwfpIuTNFqE1+1KvFvRKNDBJSXNRC6JCkBt/Oj4+1ko64btvK+KMyivSYpn/4ZX17achFah//N+y36rrDSQwxO8nFzlWVX3d6HjP7umxU3QHhnINvT0eA0av0qo6FzeMh+XhG1tpn2M/7ULXmf1mKAGZI8sZSwqO2zUobfglkMuvXDRb/BhrgsotDOjSnsYt+n1oFHN0p3y8dV+FQz+t/aar3WdgdSD+Xg7cr7Xr70wHL4PcGrizaK3dUEBcWqwdSDVDdTY4US5fVPi9PDbxzBX35ZhNL+ZyaOXcIsrw4zXWqvPZ7EthD6EJFcnAnoqjjgV1zim9TZ7okovEyNDXAxnTRgCOV64CS3w03vs1thQO5R2lUGwYwRZSQJbomc8UDD83c/IXyruIBSRvwIwngYUiAJ/HLE9Z759L/ceQ38JJVv8Xxmp9BhBldM5R6ufF0HhoeFdZDVGcYfEtr7EOnXPW35X6FtLYYZXiPDCWtmFBZkMAjMJR8zHsiqbbCy+iyJHAk3h+54oM4RhMW19BgI22WXIMsc6cDuUaSPU5IoOEMFyLlpSWpVsxinGjdAdC5eiC5+Vkd1isQ70wJVlLhl6a+qTAjK6zE1XiV0AWJHXAaSt/HeudajbO60XyZeMca3w8ywbAfLGowdpbG1aZGbJL124yndrSJ5cHMnYtCPIlTIi0YuN46fPa5NmunLR6Xn/KcyKTWbtp4j/7n74dOx24tP3YkRXXii4/Krxd1DVr+nERcPrla4+3Gkgf90i8UTes6NmkL2c6byJuT+dUPHBc0q/Sx21+PmjMS7JZpnpUTc6HBkBdW9MeLG5wYFHISjW8CWWT26+X0oAfUa1f6dxeqdNXBeRryonIxG8WdR0X7e6HzHwJl/iSa3O1IoUKrPK6cuETXTpKmgp6HqP9Uc09muuIJoqSRnE1xFOV4Uajk2fFebBG6bAZ7HRckaPg+6x81niK8ku+K15/XiF1MTDmpViAn58beQI/J4Dd70ILUIefYeZxWeHAuVK22x4nMakkaY2QRzAUiP7K2l21WjiEXHfQaiIXD65PEvNZ1GdaK2UP+wDrhZiUNeMigKMVb5wFEyxSMu6kvK5uUV8qShZaTmhLAR7jflclYecskaCZY4YdsJT9OaG0zET6MrqrSzc/Ow8qxH6CvUmPZ9mQs6SaTtKg/yVhWMUpfeIbQhwNGG6hkGTaxwT418+yGVaw9f4/g9Crll2z5X5TUfrF6mIgazNCnbujFiYrlGBtOQ7wGg1hsi/xIuztjiexCscvCgf4aKiT8+x8reZtvU+pWLfFD9w7CEf0mDylKyoKR5oqRqo8wk+BS1M1NQZONNNlghCSpFozfSXoo1vpE26fT0/z27JXzaAb4lH0zLpoHjL7i4Z+/uYGU/49dsG5rHSlWPwmNrB8ex6vjLU0u7v6DRLrGE2VcT02E9PrLSnSCmya2Xn5p56ek50lVt3uBcitJl2hIg9cODITKSahVzVzb2yc12EbS/f5i9mw68LSBQQRSbQg0rlW6uK8tGF0I7X0iKSl07+t2GRiKl3OSO4DGzsYFyX4fq9AcmbD0KnmnyeFvEDHO5V73dV9ocJsd38eH84MbF+aFr54foFhnt4P9wyP8/P+pNo0GuaaPytaICZ0Y1qG/9bOzbOnRDuDA1utm+hPHrESTwlI/Zt6On8j3ljfnRP9WkxYsBmTW2waTsZ9jotnTm3pryTT+kfEdzhlFNI2Z+fidVw2aDZkUHU0ay94PWBg9NegRVmjKzOu7C1IURZV/iw/tIuV++Nm/391IjqjeAxkF7bTmQiZLE2+uwzVWwevntWPqjSLFSZdIb0W2BMHl/CjCNA+KQvsIfJdjx3ZtVkTnBxYpi7ySUBrqUDeJksboKNEunHOMc8uoHjeFhSkKQGZXKjcNKe6zJUz3lOECwfV/NTMjb/eqR0x9YqPuv5fophcH6Apou7SK50sZ52QAeG9VmDBwnlq3elOKzjDxXiDcZ0ddlZDQHXOaJmKb9taqdcF6kW836rR6YqGcwkxc44CYvhCgnfqGpDk4oVUu9GO1cQwX9lyc27Ez+7XGbo93kd0NnNMRHR7WxQoRFxX9EkFkV5HDIzu841ifMaa6RlVTIsqNvuUhssQRgBK1qJgJPc3zNOPSoRHAg+fV9yNEsjzNEMsnT1DYxEjEPiVRiQxbf/43OjkvHwdGx/gRlSDRx7Bp+6/yik6BnnEB47JCAiQjTegPMLkez8g8iRTkTTBtyfiOgPFhVZB/znGBhZ6F3sYmoeXWwPgT+omU8Wq54NSATXY7Fn+IZb9fbMQTjMTRq5vSGE2ePr4uhCO16A5xILPLi4kEPi0MTgZuwr9Q+lYCU50ycUyJR3bbdjlLXjMobIWUR/ZZ7PyJaw0Z4ysQjEBOitZODPAL7886C07kzsDtDRQe9PwxmOfLwZ26ouM81yisfffhFnlm3+si+9hr2Ep213T+cDp8ec7+NSgmOdbn4nJOnFHy4Pbl8wnfYV3JravBkdf2SGnCU+56USHEIbVvVxZOGVNM3XK4zW8bacC74BJMhyQbNRbi87v/RMOwQ0VwQ6ssoR9Mt6AT01u+P3ljaTNE6zmXJWbkgBziKXST10OiBecWZpfBwitW2xCrElp0duf53hl7S54HSQZL28/+9Ze9waylA/equmH6WitDjh6JLPsLmeJ/bgtbGFEgxW8HxW27IQYDH5obFMOzldwFx3VtrrhQhwtKWFvqj/4ij3Qtky46xZQv3PUhRbPPxykuY9rcnK9x7TAWiqNb/3P3Fr8YIaYpTy101lXVRPdwiMSBFc/jJ/w6oUuz/FxunnCBOarLqSPw7hROYK7QctGkRZfuX8SyPMj+oa4Oe7Jwg2bnLNuJTuuQeHaW6XFeweaes5WU/HqXhFMmj/iV0dJ1Q7wSgSkFLhlKyVrj68pLx7CGDKNhE0g1MK9GFDPNRV0nkIBJEeGSJlQlT/8SOqbNqA0EXHhyDnL/2bsK5WOBDYq1+vaeM9OiwcwsuJj/g79EDpvW0cp2iQr8G4StmUjjJ4hB9PnPXMTVJILmD0J3zHD5t+oJyogaluV3QDTofy2f3KVJ1ZcRlK0hqH8MKO6AzyMeL4aJnt70DySj8/S1fSIbPfhDAAtWVlXmAq+vB1nMSxSWFdtgCgreDLfrlJmCV9aAmrjxhJvgzslZeOSuLmSuc2NmheG13tVDm/xQC5RG53TLzdRh6Egbm2lx7Ezv5ioqj3j6gBooKZe+X8rMByFNy8sbBrKyf5FDIxwFyVtJKsDaasaOpP94AItNqXxxkq1Ad1Syf359Jtdh5Gmkh3UGR7RAGPrMF2VO8gxXKyw4FlYaOaNV6CSwwqHXZnTGjDcadp1flg+5Ci1m4ga+x2B9/Xtuj4QDh35Cnw0bg7eowR5JMNMy+GMf6/G8P9DJPxKd1uSU4pg5wK+z41rYvazQ300LXdwWrFu7sjWPHMx4HoxJTS7g1V2tZXBCGWZb0sSWrnA+CGtsnTxGtbL5eAUVYtUDkuhXI9weA3eVwFu1JW6LBOm6drLiw/HY5AmK0555i/dBqCU3fU3e/yy5+bTfv/f2WahF0/2k7KD24diP7XWY4PoeRam9StHAckG0hSwOgiNS8rMIkwj/TdVCC+BhOikZEP+vwJQlZWqvq/XlgezpYR9O3rgfuf4n0dWtRl7AIzvfbK2VjZPuRgKyCTjV3azMcGfmYv9RymUi8ZeQb8fKD2TpOEdJtiYdIjzjtnBhptkSVfvELmJnP/n9CvIVceb43CGDdOpBg42lN8fw3yZcVWwxoiRbRnj2lLY0U//hwT0u3vm2tiAgeNn5Bk2MxYTpaPlHyZX+Fw0/pshf+PAnLPU+u2+yjjrnyfNx7X/0LJx6Ij3Wzcq70xNvHMXC5NKZv/a/M6vpG9AwqU4Iw0O3eWidoc7aTRXGtftxp5w+7or7heTn7VHMVclWuAo6PzMvt8Qjkna4+E111LZ+jmeT99c7nYIq9FB6XF+D3sxW0AoTFaDa/D+kATipCUWvarIi9xx27CVdErIbGA6TrzmVjhepV8fgcH8lvdQI1+YZEkHUK12HIGWZtzyUk7fSleMs5+cd9MZjaQxu3CY1LOiumRG5s0BtPOC731Z7CJNi/kjWJBiPVACzVDj7PUDyEjD+BK1MJbLnqnpmhzp6SQewsqu7Es84XxpQ3TLjOvHPzE3Nj9CNRloqN2ri47JeyH7UM5JdbOjKUINygeTtb4MycKUPUr9lRfE1o52X2vENtCV6MgeheGYb8KMTWPPejYDpSbz3Btbie6om840stt7ePAq35ABaEBkzK9hZktng3ecVp/I1Z8MlmKcDpLJMtHmVMkyscCr/g05OV1PZwGDx11veuv6iRRrW9PVGl7ouKAs18OXmdY5DtLdm4MNBjHC8oKbXGr6andZ2ZCSzbdufq9RwUAJO5xOmCsHyvptbAdaYsmUvo72jcSdL/bTCH2inr1Yj1Ia7dOvs4lClwb75pesZL/BnHAqQJ+VmIVoBtSQezm5nJcg6myeankmHFlMOSwttc7ww1AHBC7JTMmZrJi/XCKHTrvbvdSZSSSxH/iZjDSZKNrKCEcjfoLvzGothZNy1WaLFPKzJo2M9PXf6KJE9Bbzq24w2FxvEnzmczTKjlcFv2+nCITypqxAXQ/QNVgK/rCgmdenydPF7Qs3+1LXS0r6Wp9JaZLeaYMJiP/0kGADmaaayxbnQUpFKQz8gFdiEAAtj1wnRzBHXlWDH6ZOOCBjctX8SUkklX7SI2Or5bU5pq6QnLpZgwWIFB6/IuEEHcf0scpQWZ5py75TrGLeI2mPVy7yM/ajvZNMimh6ztm5gkgFVIcoCPEOE4atV2Ph6fr6pqSTwA+i8TvXjROv/oc+IYPHxhuJSBTIxSdhN1K8vvbTGcqca4H/sY30+TCC9Z+QT5epzWjSMD3TZTSEWdilKiG+XzVVvKkit9+ZCXhiyIw7+znhQ5lU9szwGsK6K7FCpDDHn956XLkQ5S+bIGSf+l+TsZUP5ipaUF/HnfMzi9JY9/tyr6JzOzffv18VjtF54TbU8+3q7mGk6dsqRjpQWw87kW4n55qVYIycEk/bznZi44uI2HnQvIGZZN1hxNWBwNbBQ50O/PKwrratatnxsMVyKe6QVc9ejF41kSLmj1KrpBJ5uEaal+rjOl1mw+libEHn52v4vj6/uOok5otU1Vf6q+9Dl3kWt9Xrq6fNSsZPLxZ4NaD8EhoUlXwJZRKkAukwYHQUUA9Z3Gk0ugOnzcm7zymHkr9caJwp9jKo1dMwrhRCER6ZmPcE3hK/xwdrgkfoQC3/tXKCk682LfAezpA8jgK0pQCAJjorIyzwJnqO2PSQ8ToZX9qU39JmLf5mVV0qh1TaXxqQFIz4UC+d8svLqAwv7GTDOCaPJBlfKavRAE1x1DYU281JW9MQjA5eBrEAesw480zN2JfI0XaycG337nmXAhqO0SHKydUPrTFJBgw53aUZzpNlDSmalsaqY6LSG/zyawDtdjUgZ0/R/zkYzr54GA/FeYDN/d/fA13VNtf/EGb21DugdB3mUjb8hQfIxtyMwQO3/tpi+HIoCN16ey9yiHhjZccb1cyjgZYe5z1jhykvugx8pQm6nMtfXwg1yHpw+x5Dbwy5HRdVLHsvhbOK0JX50N2B/tg8c/q2Oyfl7A2iE3XJW6nbl2aKqBd3Vtpi4948TN+ZX2+A4xrMyL1UzpUX+GcIMeqX7GMQDYtCAdlNLiQh7EH+9GgoxTJgTu3OUnXMh4CBK1IL9iXIPnwBmr3iLJ4alFH2ODz70aRdngKvvVFpQ6Y5TA/FUpL5wrlI1Ky1i9w0EYY7DG1m82rlolucpCA/t2XL2C6oT/mgGuDR4bh3zlCIHiokrd3Hr6eGbIgu1mdUVfaEIDpZ6CDZ/dBK2t+xBv3jYUstH7uwB6uGcL0wLKuZuxUdDx+rQh7S82STsifeMGYd9oEnbQwQ8UgkPT9pR6v0jIQyxVKCrDrq/1y7rZzI0LZJbW4X1xoSSAvEeB11o3jAGH4eFmcmBCdhyO/UMlMnrvDSmml7K/bFoTQ1rocnGjeC0zb3eI8zVad+ZdL3R2c//L7qGwgdAIgrWCr+dWHEVjYugh7NL6SAlVlw8dZQaFCCBebEN9Woq/hqAdWICleH7eMcuM0VH3VrslK5jiDjzGC1nq6d/Xbhk8r8bohpPQpNTaXnXSqoaOFBPisZXdOB/IALKpZbmNOAcQ9wkwd276WljjWK+i/uLDqaKfJG2fJuOd8Tj3dmmAVUMLG6faRNghz1jV1Dm1wrFDq106r7A52I4myMUkXMYnsX4DewtsjMvbxATTIabptuTDb4RvvgNum93aYGLtUgElucza1S+4XpZW4nu3hYqVttGa4oXOdr20S0j7ieY3vjsk25HXW/rxBYZGIhrIJ1RgvCNAhMiWkyVK+Io11EfRqrL2zoiThVJ1MxUWvlJDgciIpkMK0PPc3+SVAkJ1y0G+GgRVJ7xoa1/V5CRiVQqkoK4WaQtDsqXoi9LcAK6NYWjXUPopOUugsu0DCCD8TthfH/2CXIxMjbzWzfZBHo+ox/8zzj0sARIyWpUP3D8t77BN7gqXJqX7D/jLVsS7Rlq5OIuDJULEu1J1Mrdv8iVKpg8hXYuiBImm1+NNWqKCW/RQhV92KBaBEzY+uFxVmzi/y1IpAXb3aCL7VuArCMa7+n0D2nu/h2fm5VlZUvEmDOFxtb9+VcJr1QvQBiT5tm4C5z724gBTRdg/zRfVXELd34BgqRgG+3oabibpRLNGZPqlQWh9a/UY3FY/iFvgX1ZQZJpAXyKcWeAXb4WmMPvFiiXJtsUA+iaJtxDYuZ+Zxgc5hq96YG9BAdUDPqhZ8oUrlsHOnurDLfWmJ3c/iwsY0k1RobX8PljOVO9mHWXS8/+w4uZVbltq2aOq3rgbUInBTfLFoIMGqbvQvxtCKIClkDGTN8bc1R2LDoTzgh+z7nq5KYNtAY+JiQKJugWt/7XIeL4S13gV4rLW7phtaq9wn+r1hbeFjMoU5LDRajgw/jIJgt1YVzcA0HO/iRZG0sNjWRrqAa0Cut6L6wVILo5/GyTZMKukhzJSZKeo2Ey2e5VHy9BpIgXguL9QfDSKgSHtCAxTVTniMABCacwPHri3qtsyIZgOCLnc0bZ/YCdDCo2w/fTFU0U2llVhRNJ7do/+kpOVhdPUWEdHQ1KxXm/JbsQASQSwV9CQ3pvHX3Pgn7sleBVQWcfBp40XouMkYNR+HIBmjyNHEmHaIyYQYX/4UKNj3ZrJRCphsGCEcamt1OHoJcBPDw3udy5oeWEOi7JuV9lqE/i5PNyzhxGZ6dWOVgXCId6SxvHV+SWGmmdtep7tGVrPvyS47xm3cMNe4Fm7ld5plg+KMJovGnmudo+d780xcCvpto+Lgx5h2d78dcZ1ZySxR/gh45Lgx5RTX4iiG+Ly4XtvSFr3e2hYse5bmGYMPmbQHiyU2TUvue17z6YV/P/8nkPmny+bWeNGETXQYMMKZfvhdU5rYHsUmEn2M1zAtu2UCODakXnvVNvF0fJFiB6aBsxf6OoiocPzfhiM9xWaHQmRQjlj/DRuRL0MCFsEPRpNlyDYzQel2fja/AWbgezuWmb0ScY5witG0Tv7+OIcOayFN+81qrPAgvoCIxY14KqHsDILp/6VIFGO9zDLHZWbp0RGL3uT37WmPKVn8Efi+BzhCXyS9ITwUFxEo2mjOAVvPmSsZajnkUDvd9ZKKrv0ct3b2sefjkenAhId7aIR+eW1OsimccwuJvzvMM+2twU/pSVTkg2bqEaPOsqJavJmxxWrDtzrwlu9xBQV24slpDUHpIh3PSKHXp1WGt9HTapSk53Kdku7qwbuMj/LloeUMjw/O53dy+0eBMSPYTPoWlqFTmW1WGvSEJdSqO2l7W/6cO3YjkCDgjaikWCvc4QxPrvMaT2tLmFt0FpQcNLrCGjAilj50z1gsQuXlMYV2x+z3TMaUs3hrkcNRbWCae3/19uZ832N1q33QhZKfFNitkkxCa+U45Q3dNhVgxoNjRNaK1xDg/t2xBRIXD9+nidCyunEwNTOk5JVZY7l++6068iZg8ni9hZu6m1IjFmFVo/5PkOkp72RqPisUum0X4aU2u/QmxBe52izHD8LszHORSrf9KoX2qgfyCiJk8Q09KOYvSCJRRD0O98qGa0I5KxOnqE1ZCCbEk8Ac/vnCNC0teqYVrI+cwJFjXZteQie+VqseiqasQO4Csk5YchvSb80D4N+NLzTjUdPdL/iPcI9rufqtRngyqgC3Xj8QJfRms7oYXME/zW0sAToztIVKvv6GxHf8GCbAyn8G1ncznXtANwdQWGuC4hAkDD/m3Y47EIehSe5455qVu9/qLxp7J9NqE27mC2U9DBokiyulr4VI3w5HoyHL5blPVDWW/c8+bHsrpEIlAFOT9ozTC2w1c8Ryy0BxvXfoR37eXypQJykNbm++4N8rmHR6ISd8bhmw5rpXoD142lx12Qkug4fpCzkUD+R2QpWmHEW9usFePhtiPfMyQt5MaCsb+H6fe0ZjPj7kIf9tHmxXdzQ499hlKrPPbPH9Ml2Xs2CMC/FJOyrEikWSdL0H91BpHGZ69WgN2EuDQqrRVp+FJ3SE2J4A/WP4PRMP/QGKMEcERCAROB3IzFDEpA9JfLLYFoOeE5KJJHscVIuhgFRXlToQhHpR23iVZ6rq/5JIv44+A9TxJlHZXJF3CDYM6Q7+Mz9+SrwsBKOUWsnj56Mt7TiObehp1qWiaFbzaPTFPJZNrB9P294LYub5EjgXY59lBBg2NM81Xdt4+Clo0BAR9UuGudwKuEWvZeTQPsdTfm+515tPCjp8L2bqaSadmGbZPdN7Lu8lKO8t6NoZPTCMl4W/NZJazwUyKnA9AxEmjWDIK2o2NXqgSQsQSvHbLULlhywT4lnMw4SOfSayG0Vpf+ix9aykGzMgQZR8rpJVUA/6h0ulgFSV1RBAw/XeP4xsA0t5W+QlgRVzJ2jDJOudg3jlvzX9qmVQ+6ytPrrnLGd9p9n+I4Onh9SAA1HvN61zVCfvicsdnAYpXo4oRosrqDG4u4qk0pKJQlGsWlYPY06TE0/29AiPNcaWRhqlmNyYePICV0v1LxPn1cZFWH55Qb/Ivl5HnDPH4Z2d/yMvpwfmmdR2xxnMSjq+csRjejv+2t6wHE+/ekbZWiiqv8K+20D4TgxXfjMV0KMJ4l4A6de/h0oWcF/4LozED3Dbxn918coIn9XrxUrrD3T3SqOLvd1lTl8NyKmJ33RL7rulhlsYKENImX5f8MGa/QBvTQkthxg8wtyotb8+47vsFEhXQGz5Y8ZzR0SPKqv+hFoNpdCtv9Tyfx+HpU/qQjyHIL+cIvVBHpiNHe07QpRNY9jVQ27DQ2C9nSHaWhp0kNFtwOEJv5/jFmn2zpIp0A+yghkDpLdwCN/5TlupEcAPxFXpE2XbrXLaAH7O9sKJB9CIylLK0baYClmbPj73f+v4vlIEobnpVIQV+Ri5YJO38zQbWOwo98Zvjj1sMos3D1yBQjkDgtgeMl7fm5RgvdZXujPP50/nCU7XmOICbrb2TbEtjlIBHg+RFWIGCxEIfYpQGTmjSfpzmAe+NogWTwbRLWnZchpuL1H2mPmdiwpQ3FcWRVt4GF5jRg8NYeAaGb1Q/XZXc9zEggTkD9VL5KqckVxj/n9ePEoBPT+3cI1UXl3GUGnqUXWLv03fH4n+ndRDAQSAXFnLYZx5mce41e15nD1vEOEvbKhWNzEHWflLakf+4wiQJ/EK8v49ZSNGJuRnaHlUkQIAZqU/1Awge9wKWLu2Q+14IBmx5nSlUeupu1HJfwoqoO5z7DZ4zp+p3kpItzFapOd+Hhk3Ra8rbyMdSTCk8PHaFUUKiwUUg7reEWsHFXxZA9tMP5v7tgKkncfXOoeC4Rztw21Fq/z//iacaULzRjqoAbsT7zQqcCB4v3q+Cv2pL/IJnZseL4DAdB8l68qvp6YuWkwAHQbkVTr4RClmPQgLk/QaNMo5g189bBMgG2KiorFAaSUyZRyHegCnOyjWL0CiejVkgFh3HPP18vD2tWKuefT8wlsMB4aosBMfOYxtWv7ZZmNaJGE8p1uoWuLPPL63mjoy9r1o8/Z/auhkWkR8f++dhdbu0Stq3OQ1CHsl721EuxGUGEug0ggDX/UNn14tPKMM7so7B7D7E4T07KPWPibVKfWBliOK3J0GncwVx6g17TD5ynWzOCJDENj5eTHqRB27REf8gbDyTjU1Sb8maeTttHo1J8BrNDyUyisatw5WkshnpCxBLOC/K9UwWNF4px31DgBx+CC988sHJwxmODeCS5xPa+H1eX1tx6sZlkQy6ZOf6jyEWWIziddtP3Xj3ct7z3oFOFXotQXsWnvLmsWURzAeqYfKt+81d8+75a9IkBh4LJjVnbZaj0VGol+ubsXs5ZnLWyNWbQMnz/LTgnjUybntNhrTb22u5IOEaVnSUUN+fKsSs/8PRYMAI6YPezun/hGdtjGitWs4McOI1XQffwiH23bNa/Fpi3QNZRE8SmScrJJ0MSZN0l5cI9vuS0PGagR1JhN1yQCiV2Up9mu+U8ARwU9OjSL/WLA6aUC3/J+FdsRE1T9d/SftLgbDgtwZFFhpBGEEdoHa8zeDiG1fbp8ZMJFwHTmlwOHIL1XKk2W8Zn/9h3Lo0CyiC8WvQThHVNjC7+RnaCEgfWGUdy0HW3Y6tNiW3Pzu4xtBnSpJ3sBDIzr2XI6QvzC1rOW2g6uwZsHuVf5qZcuccmEr4x8n9TEUzXeTfocyOJEe0/yZBq5GggyWGRJLM14/hW3uSWpWTXGQNSXNIkOzsa/1izEI2KtLd4/M8ut/JOWJABVotg5dxKxCttSQX441D6qqAp68x1gK0omz73L73YocPdDor5u/R08WOD/YiR3lo1CSGIB25mmQCOJUoMtXiAnV9EO49SZ101XenfgJo08hlHKkmICcDm/kWkqIDw28YX/Qt5rfU42emmiDXNY2TAZvQZhqQr7guNLrE721HRMTMmR0fAPSshK2Rtp+Zl2lzw5BleE0ks7AVdfIpPMAfH1Yjt3RtUHOULLtIpqEBD2JUJMY7tg/ZEC917evDni06QiCZWlYZ6/+HIOVdgVcJsUDCNw3OUy9pPiPdiGUfL+1G7KyeHPRfaIfnI8AcdJfQqaHQpL8IUCAFm3x1JZ3vwIripQIXa31cHoo7xKZ9ZYkCz0RUY7z4CIe8pEkVH0nVhO2vUKiKWkWZPds5IOfAeKkowATKvEKcKT3gMrQoVB1camRUVAkmAZYjmwzP6j1706sa228YYpHWieiGkqRigBQfkeU68G9GEs6mLYrZ8LPO6MvtUeczt3pNkdf1nnurh4RksUNRRv7PQ0wwdA=
`pragma protect end_data_block
`pragma protect digest_block
58cb5dbfe99e59ce746b9a3d066a43f3c37f926990e34e682c7c3c3c26b4b40e
`pragma protect end_digest_block
`pragma protect end_protected
