`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
Dd4mIOZvDWcTuS2imJB29ezG93IwJW5wgqvXZOMKsX4nJz/rloN52dJ1mvLGBaDELhjXIs24Et8+EgZUjARlPHh37ECzFDSNfUsTNoaRoC0Mew94o8K4i7UIi5gTknbjAwyYGONLkAARuoiuXNwlkIWpVv0f0yhf5Kb+D/Qoagn/jH+8wtaMOajk92KHqwwyd0l4FEB0xfC1GAOiA6/UMS4VStFoRq2SsRe7i7KMhXvye0lFpVH/I5be9fWSNlp0w9WYdlAUSJBH1ygs32O95q7/GY4m+8K9LZrUf4dhH4BhegSo6HgQnp2rC8XF4oRjClM1I4vqjHnh9nsbAnlQzyRD4OynJTfqRaQ4eIrty7oK8quNM8iD1aKjn9cI4mulPLbV+61gIPhQfGZcc+i+LonGGSdd25vV88gLlBVMnxVIoz78jPGC+B6F9q4WZISW0Knz3+iAs8S3TQcTJfCENBUq3v4YKznZK7G9ZHrED5Bfdhk0AXVQLC5GqtmbMTY07RG3gW4Sb/ZrvTFKFjo2p7F7M8PPz7z3JbuVcGuwRlG290MDapYVDEeCEIm+kDLD5sk7JCUflWhSKCG4sc5R3zdpL/5z1R4yGXcKJzh2kJh43uz1oO/Z8EBGjYgAQj0/iXDH7m3+aclFyANUEIk86EfhQF25GqasqjuID64WX4XPz7cE3pzI9MvEFBKaOdvyh+oqUJivUUdZ/gIz79Hub5+Jf0WTStcqwqKg10U0HJqjJ1lV7rgy75Nhf7/BwsistjtHtauPQ3d8GeuB7o9P13sGOGuo8am970KDR/gP3JuJqlezebgLm4EBn7RiuEJkl6RPY65qCOqwbsXuLS727l/SS7HwT4vqcBjf5o05SWmx3aLe2oGVUu5WtF8Qz/0u7n/wITKIOWIjKUJm3853/+UOjyYsJat0Z7rHKRgz8hJtygqUVgFwB+F8H3g/wlEt0jIsEaZo3b7pgkW/QhYXCQS0ufIBJEvEHAwoNy1rkVBZ1wqVb++gywhoK/tfOMeNCEByNALCXWTqw84PELO0EBROaTs00uN4ladSUZcsLSs/Um/4IX2P0S3Wxk/pMneSBu5vq/S4QbhTOSltlC9KHt1ItF/C8l16tBKE/JKvCdnFhxwuRz9rtkZJBI9lQYpGT+BYORVNK491hZ/bgdcf5+oUI0Fu//hVOX64yyW/WPCtcaFx09HPK9J8/ICWvBZRQyfncDTmoy9sIbm7KtWUZwgVKxve1ZzoeXl1oqysJlTyyHbrrh/DZwHnIGzUz/XQudkjAx2G6TwyP2dkTfY7PUG1v3ksUKMFi4GYfVEzM6aJNzfjF/QT/w7x0cYvsEkWBE0IHZU0fFMXTvcm8NW+cszHR+bX8t4V0NzGxWhVjADlvotLOw6LZg9t/0ZodSVsLWxzLQJ++pn3r4nOrFc8I1AsvXCQDes7kG/cBjaa+WSDDCRvL01q+te760nHt0a2d2U9zyEtLSGg62JXuft/VxV6mBMGhHRaF56jNiDVXtsigFB/ONfleeTQdWNf1/0IJ/ap9/BjNUCNCgCSsjMM7tiDOraVnINIKfxl90buYuZUiN7vC3Paezpo0FOHxCYFEsOkOzhBTO/0DdPgq6XJ947ggLZIDzTSS3lZOtGlnutMauE75b3WwqHsqAaMmjTqhaD/iuf7A/xYHn/wzQMsoImj1X3mTuaKjfME0RHiQEto6I4x3TxrURx8TZ78L/E6630igIz2DXHyRABDnGTii0IgsTY472cKyKYNqkCaZKdXJ8+tNrMyED2nPS4pq3EUH24NF64MeIdOO+sGpF9h0QHxuh5DaBOMcJ2CYGLEUch80v9DXFFI5C2ahD3DfTQJQojc/hwMZNTb+H3TylCjo5ZrBUrk/UfLaPWRTohc2tO5+sK8TS7DRU0KnX/8CAPqFcd/jePm4OdT0rUbcDoc85okEegJru9K7WVJtsygHrmIFt7zLB2KLcveTkz/7s7TmDew061DJDqH1HKJNCskV4cQbGDlaLoNBfNs2AUDD50yW5dEh6V6qwwvTCMuzNSHKgK57ia+KpTUE3GQcQsEIfnNozoNLL29KAZ0ToTl5WsvLynt0XpI7A+5mOnvoalM9AkUYTbWqOcqHEF/5kWLEl2VlgjyPDE6P4Y2y3yjQFfqXLXdlHpDAySoWYahXA8v+8vHzbM39rsrNe8xQGbbWrkWL08LSlze8azpSSiFVUkFyq6GhXIDbMJqeCawsNYDfr5UoKkOYKvBW3EDEEOqVMCh2BgueWqWj0priXmE+vOzuokrNM5tAPzY+VIvW0wf4EIYpeIiufVcrdvRnVfrb7WmlmtdWkOyBKiQrcgbXL7q73egXJvot8KwcQXymfMS6SREE9uQ9Ux3g9Ky3Mx6vRxIZoyBYdMa2OkbjjLt6YE5pgc6y30CUsnQg3Y7809fmU6EDE3GOaivwDUZ3/1gYZ6ejgrPvFcOt47scCKcgyWEAwS/8PKyKb52cF/RQ9dR69LgHeq5FJfrFelVNE1HkyQ08VuXFozJzyJiWtsWlDQpgXQrOE+xZZyLR2ZdujWvgkE13VjlySFjVovtxPDtHSUiVb80sS/dxxd2Adpp46lkcxeB2yfxgecE8BRcuWRdjeNY6U3GxMiWSgkQhfjFC7hQFWVZG0IptNp158FB1PbBQ7boRrLcR+kULbCikdsrkd3j7e+QHqahH/WRsYvcfnZFLDqrJXHoP5h2jMOtFgWMqNA6oZViqsL8PJvhqb2eURsY/YCOynKEOPrPxPuFd3raaD7AClSABgIXOPGQsrYhhwKhc9l/0NPUDA0pOcL4XaLuRj0Yme6Fnzteh7WZpQhuvZktatb+Q2IsPUHuZWLVBHQ1Er2hdElurAhd6rGB3MMK4SD56giYqbEO0bxzSEgESOfxWYEmBtI7IW7Gd84LZe9rkjpzgAyc8sW0eR3y1Ms1qCzF6JsI4MhCiRvjL/QMyunSj9D1A5OuQtrLHLg1ATfOz4nbiLRkXZk679zZfayLxUmiFZPrGnKbB4bl1kGbsb9i7ekGips5tMSfGc25JKmpwJOw4TCTgdPgdwqIKhcf3xGwCSx5vNUOeZgo3R1UikFWPXOd7EKfRNSMdJL7CFjS9iOFxCUGU9gYNu/wjTTf8gnZ3EZSDchr1QQ3kAGnvxwYb1B5v12lVHZ3fCF8K1U7C5Hys/vt8gxwMTsLlR4zljBU4HQ8uKi5nsxtFyVknRcuxqRBFFPMkmNSCo3jB398zN4L7EfQHnhi9uEKeMT6xxjDqUnkbaom9Hel8aX/bJm0ZfUyVRAOEPM5OMlRUELh6ZRKANnb2g4NJB9uLF1gxvYwRTVb3RDlbJf/rO2hexjt7Fky2V9c+Q3+JKr5q6x6y6bHZyXhmdaWOfKROtqvUDxzJ7+qdhvUfuQedXzom4qPo4rluNoUO95bur3guSdXfI0uyPqLkQFLsFcF/pD9oInwyS46QCrhL/nqExEEYVJp1APwUvq/3oRRq9rqPdQbS8DlDEBZn74iiiWJsHhp3T804tJ3I9q6TYpo8xjgb/kuPGnrphWHOHhZ57M0qpoJ9SCPqT91wjDcYUKIpr6TmK+EgQne4yLSiNd7DsYSfGKyQseYHhaXB5SW69Itpvlh88djYo3ymsg3NkWDWlYkC6KvdUsLaP69hemwlHzCcEo6McS/rG0OXz1Rx6fb9JM2JLFi4JUmvkzNS/q57ejSk4z0W/eGeZd3hs2r1cqPEUej8erJTcww81XxChbJzUcT32qEUdMIJu3MkjnaYraQ4iPqSOyc2m+msmkc7nlzFA8qTaHGUVyn6Y0TftgqLJuop8bdPKHYJndxMCetokOFzExARmVV9DY+PUHz7u0BUdwKeb8uH9dKezFDNL7DSGhn2iBwPSwrqgNzx+Q0TW7FiQEtADy9FwwqcSQa72j0BA2KxFxZ9g1aR97xz67suqLpm3ofd9uHIOJJdA7T43GWlSp8mEiTABRXWZk/xxy4tvWsoyphdXB8g/xc1C2M3v9qRtXSxlrftwgBfymDHNKbAapIGB6NGYwndSKOwq1JlinPB205dl3oDvaC/dSInV0fURx6rUU9mtpRhUH7N6LcZyhyS8X+J8LyGCMiofDD+U2d2Kq0w3+mVBZzYAWPK68s5f5V/AosBQMHcG7wbGcvYj6eHqg7M0/l7lQ4NerftZtNEHVLhZoHiz5aq4ke/Ytf0lDKDtCr0NTSuxvhR2b/2uTwJSBeCZOlwwcljdIJX7j4f6uBITQ0/29UODN2q6chllzYIdUQvjUewLS175B1gWeBU4yqzuPmE0BGHK3p36HBmpS+GdY6YEBApTrtn2xSuDqBX63nhP0hmRzoBhDPJ9jdCcpj8BVx7paiIMEehc+ZxdwmNNKODIQ8BDywND9QtyWCsvB4pMQh1WQbpcv9+I/7U01BlCTlbfhHRpbg8Zicpiw77IjFGeeswpvzVZVn5PbsZ/DS16rfkFukM8GMRxYaiMCkD8UGICFz2mRMiDNvWxqO1l4wN9GzC+Wv+QG1032XqW6+/evlXsGD96MMxXnz2CroWB+cS+IxlEH0hRvXrTVMAd0Kbccw+BqyIeXCDrCqgneAPFpllsXT+6uq5BAVfoMnQWIQT3oI6ytw4gemcHhhDxd/qenvQypxlUBY9t6J5KV5dBmnoYO9ULX6G/yOG0emBO4FfpdMi5EHe/n0WFaeelkCliJhlQ+BJObco60xsJXaVOaYZ6Mp9XAyK+ydsRkTr91GkK0qpERRGjJHy8a5DqZARAoNI7TVUJg3WohQWMdXL5jpqFIDdimq6IwoHb4MuhGCnAEYYChxQxXXZ3E5uwce1jR9XW5nvQZF7gFg1wxbETZsuMZTJe9Ki4Mf9YQjflxGldW3QO/CF/yqQozYrdhkfiui3HQ1sd3b2aDsLvwRfAPA03G4POgGe1wQHTmcSj7ZcJrQR2iZXx26kLDsLt9qSXuxdT7ImdjCY6nvSmVLP9Rgc2arbkY6cyuUWZ8nk+xvVGgeRceH2tgcARE/oirm3Gz5lQjmYJ0I/PpyuTrPz1d6wWPKvPjlYgOG8lfwQTW/Tp+CqZxXSb4HWb0EZjtdFWzEt/1/nfq9RrQjVSXwkV62Yoer1P0FF7V5bEAY+xISBesEQIQdVhtzwHE1FHO6lmO8w4YtUdiPoK82+DlRIAvfsuu/bpterqLIsPD5Mp81Pj+RhKoA4DmuAQEc3Pj/pqJjShop8pK2cRxq5sC8zVUb6zjpK2Oa20iz4qw8k4oJbQdwvdSGD4DZ7YSVX21MB+DyuVQqJbWEhGQaNJofr3xcX5M6j/uVJrciBmkd/DJGk2ORhW1wFyhsRvfXutgrSVanXFgNIVaYwfyQseQQF5ncOyq18Jol9V6PeoUcPhC3pymTmHmjzbFkKi20/0ICayjf+NgxfEcOHGM58Jc91KvTUkbTaP4KKsZUu/lFsPa3+m1kbW0c2TxRrd1qFkF3K/UzyDGOJBkVkyFV4af7oR2s2Utc+lbUjwu6TxcCOihDyDYkjvx3BkXF5zkhS5aD/1Y30/6tSyE29MOk5rc/qI6FFrbvdD9THZMnX1Ge5pok79PTvAeRV3Hr+Gz5H2gq95YmFuHKkbtTLdKyFojhrZY94hM7SfOf9OOwBpq22gyMK8l3QOX3N9QUcj5QkkTW4lxgXTnp4i9uwpqtBhgFfynAIdf3NtzrycKq8Sh8M0olEbz4wJof72tZ676HZseTSWhZGB1BLFrMFgTWLwAZlzHxEsQw5BQj3K+pWnIG2h5JKi2HyxE1WWu5BsB7OlGonYCLMfAyWr1x2yJV0wMEI5yubCTbQUJgQTw2Gn7eMGNuSJzr01Nz3RFWi2kw34GRFj4qcuu6sYSrILxq5kq2LqrkHqjhfRDi+vV2sDCTofjdRCe2k8AsMml8k84YRceDXajTpNVOJD4R0o7J1rksjOXfaAylRYL0cVO/0B2TM+TPn9vj7Uv8AqJSIq22iSGsmfitRj3TkVOA0ncmJWUfmPgAaY7qpmCnDdH793JMAyzMmkztjQ73vcRaPRS7HL2FbcRF6oACcgFZnLl/YQF4scQm9Pt7J/6VfKWRfORvNYym+JMQ+c/iVCVkbhIlylj2/oy2rcQN5OZAbtPI0dxmmYVq/6WpBRNnitwV4JXXJfYo1By5N3rMNSbq7pVuUDywciuwEAlnatjsFeIPq+D2KCY/ZLdNpO552M7mFEmFQ/uVyBbJrE5r+IqYiULfD35f2BIMMFTBm3HLR+x0H0G6/3vrJ8AaPsnGwcFXC92W1Ugczvko7R7zZX+tTqMC3M17X67bscr0keGxSzYZVYPIba106TZXKwbFljbQfhmX/UW4S5lsX+6+ocCNCGi+pLo8nfDbqzV2IFq3OS8tduJgX9KFrivjje6140DaO4LC7OlAC8R5guw/zXWDF29Jm1YmAuH5Bcwlu/1EL+4VoOFTyiXXXvKNEbVF9Q3vnAsPvPbz/99Ypj6dI8HzpE5EPLgrSF+ldCsVIHd3opi9CrWcu1UAwW3SSAmMeWudxycYKo1Z29wP98JcWdXSEqgUKXv4oAnmiudYG9A0vaKpZJ9RWXjdyTYCr2bJ30CqKv7QlvSijkbMJtDe2xdKCamrxHh8IUchZ9j7Epg5tpoyAAbjJ/+ugkuKRsyMUgwFvEenkQRXgAcGDe6iDVBF7Tpj0gHjY1sekDk7nu+WGECs8CykUf8KS1x9j38WAx7Hmg5j6Lieddtja9Sts1Zvd6ggc8t3YQahC49YHR8niPZzu6en5fA23VFLfOhBv2cNF61HhnCtEm6mWJaPt3R3OfmzZl1BdIZujNmFS7QK+jaYqQUpElfTjTOi4VgY8Q4VwCKL/kzrdde4PBzHt6335khuzb3QtpoX+/lsiJZYNlvgtiX52RD+uToRxpuzsOb84HobSuQko89d8lIskzjRJhIu6xX3OW4S+ObEBgHHRrHuYoW4uu3Wuq0fcxWEHFI16QTE5VE81j6siKYo5GVlww8YDrDeCjlAjOVLf93rGgHtR+RCmxPH9UfvdDr55UKJHJLNpGMUVtknxC4iQIktussMAWSK7jySu1FfPbNDXFs3lJuBVPY5CmdeUFR0GWyQ7e6lG9C0F54FNYWU3pl0ZxarxO5x0Hp8AJe9vyooHgDPFbwc0zpMZR3huwOrCZGyPZCloNgdyn5Obi+b4AkdFjOhrtW0YE8yUt+hXPPRFRTTYxHZ1p2jojF+mUPlWSfZK9nx3nlhFVY54y0KsdfAxbdbHNMQHHcwwMxnI74t5bUQ5ig7TVaC7v7tk4p/AE9UQbR/9BeAm7KkWq9vnQvuCT41+qNDeBIM/AXpdmeE9xRiJAsTc9aj12jWtDFGqdKH3QLUMy4b+ILTlRulKw/JZpkocjKxuiCDkWfWYulqj5mnl90PB4AIL5YbXh+0jpV6j0TKghqpULR1eTb7OA52JlHv1dv5giO/XNFe8lYaFKvhD/Oh3JBbU8IfOacGmEkjtsNcg/6MBziGCWAT60huGkBgYQ49fUPuOduStxgFzH0PdDpJ2sNhSVQpIE1j13XRvo8B4zbp02BW46cMY2q8koj9+mc8AuGxQ6Q9S+nmxwx2hsHWjAJf13WWNHp0YmHvedEUqih4rCYTk+dNCglj9UMXG+29wVwdJU+85NlqHPcPlTXt/b1Q+8ArBfTs8TIJQfTNsRE//BY67NAVHVSGnQByiCF6WUVK61Lzt95fF6K6eAD2WBCAH6GyahgrWbEaWF+ledIUHX0nK4s+shcwf7+vqlzMgXF/I1I1q1qrmX9Q/CEcARTqBnMD46cNYQpVYBEneYaAhH67YuaMWfbLWJ0cYTk4vN1tH0boH1m3RpP2HPsMxfvtZxsmMeGnbKCfX0FpJT0guqjYTGkNIoMnuoGJpFoDnUmN2GZd4GonIhx24aD+6x7tS2blgdKT3wbhmVhi9r9Mr9sId4CLtUSqjYnpxlQrGNKkmzH3g7FvOCPgidQo8o83QLGbvAmlGV+rGnz3i3msS+K3nvnmtCTmdEN/YkqIkWnggrX3alf3OM7eHTOCa/GBCNkJsQOyWUsYOEi0/jsa5y4DgXFzEI9s4Vgfse9Jiwn/j5qOxEk73I+dh/NKdqS6vK2n6E+7qj+6Lh3WwRPUTs5eeb6nHis5dU30BvlMBia46/QP4Jri0ZY0WojvfnbRucAnVK5zhfM3J8gNQZzzTp83oZH1f8sw+zxjzRsUFYK1aYoRHTL3fFmvaXbTbNNXF9JrzYTH0MXFFjOmUKRKGjyLeqf4qqByX5yHEScFP17tvuzKQGZKacqmY2Ctf9/sv6T19THCreMBiQRC3Mx9m4CjYDqhRU0UJ8cJB76Wk4ozFqb6Cwn7qYQeqdOkPikOHCGIay7P3vwsAljE1vO8GmBJRa6t0BEut56kEe/OJpJszL3QxsaOLg82/ScjGMWmGpnFyN+qTIBirZSECt/XjEyvUL+KFtoo8lg9WdXGr75SGSkY96w36RcYrwkLX1aIx5lstitzC3v0lNErSC3t6LDuTJmxmZCz7eFZbkIqEhjNElUt/tkCAONm1NpdlejKMWlV7Lux/x/a4lQgrRp+Efk4MnYtA10XBSjA2JSsSus0Km0WHBw9rGjJGMEdS22i+8GidHjkrhwnHNbp4R3k054l3A58ZekNrfQAcqOXWgBh5L/h1oNuEmqg3l+tJ4uRJk6PaTGdQmaMgwBcZ1tV/U47IhBsLhi55Tj+l1XrJjHEDluSwv93tl0ezL2PFxiWVfnVU7DmLYeCSEL+k13BKlhHn17rBme6G/mVzDDjB8EYog6jP1w0OzOLCsKJjuLXNDYswJy7eIW7gLizD3fPD5+JRvmm3zyXdtD5XBMiobNiN40DEFqOG2LpO7iYqItuTrfp8NAql6yc2N8QsR+3zKEif2b/iDn4nqq5lwoarzqss3chuTKPXGOok+eKOnAod0XEX2GYNViv3HFT1HHpLHrULEcwZg+NvxivBweC5RrTRCz24j9/jNe78NGCF32RiXfd5X2eeBbwlPD/012Y0n7K2OozF44ENVoCCMAjnnUAp7hy4OMEDXGZV94Xy1id1AuhHut6QR+9NTPs6qt063Z1pzJakTn3b3DeoHg5GSG0rPjkHcn7FgZrBReOlyYfSNq5D2xVoFYeGGklyLJqKZePztbmX8e5YfmWi9b0rD55coGpi5vhsQaDpKoy6R2+/ctCVzaHSiPJWmKKVS2RwcplHyBz29HMkZptKWlRMWg2orAhOlIn/1ZUlPkQR1Ql/C6SXzc9ah2eHN6JPpS+sbHyGhAtJzZvXTZktpBWDQcqLwkb4S+I3Vm1P3MpXNu8rIOun+IvwGbJDDY73KIiLMt+QkC2sSZFHcyuA1Lfs6eYq3QDwVlJthCmNBNe0f+vaPZCvTTIKeWj6HHN7A9vjs1hvkkvhCco7i4mv0SdQm1dfaVJHKFvNDDJrhUbDEiTOc+L6zpqgh78YmRFzqS24XOajrePhvCtVcHHG+qhxTMhR/XZyTJfwnxAAPVLqnTwxCJ2YeWf2JYpoJRDwarmmNF8MMjp+yWP94B+CD0K6y1QYttlO/ymbFc1Zuo+1GmSOlZbFv0SnzlWPe3a1DQSZV6N/3GKTESWTWoGpZ83zfZplZMREfMkuDs3aa4aE9ruqUnv4YHaOkMbg+Frl9/J8WaCUztjeLMzdL9asTKy+uvE3tx2GSCDr7nJiOsejQgOt7WtEtq24/6l21OSI1V4nR92QWpAR4K6neKqn1gOYO3fXIArPEjAdl1nfq8qmrxsEo9mOFTSpsgCt4nTAQgZ8sbCwEDaY3dhX9Pmgmc1sX0cTKGeowzFN4JSOiSXXcsaCYKLi+hOS9OR66dsc8tNXgRLYGJ3Qyas47OMROsFPMybK/XS6NjBnatQycBt6qNT5JnTShHdoABpvgPP5oNy5u18UVa95VHhbc3PXm8Q9eTDfdzdsihUSTsEkAcpqGSdstko8IFaRLwF/OtHjKMYbIv5ctQRH2ulD17XD/NNmicsNx68dM0BXXkpRNcQxzgAjyAzBi+LXfL2n49tttKndyfXmz5mCHBHpO9i3JLXXNJGfy2URX82Aq2Ews060uX6uDqpu3dMyC72hl0rE/0o2Db4WkKCJxiZ3VPhQPsf+NCKkvxp+5+LqkHFcqCRq0XVcOxzlBYSPkQmHfCgjB5ETAlUZl4lOia6jT43ABliat+DynVHPlXn2QE5VOtmLhPJ9ZcNXcF0E62HEBARj+E4egq5U66Oqjes/PvQc4lHaGOHYiAUrt4e13yvDg6yyA9W1YVsYQOhx/zTFe1hRJxr2syrGe/rkg32FNbJ7cz9IOm1wH4A2iu6PpC23irfY0CdgX1OviXOaj6KnKgDuczizA7xeT58HbS6s4PvC97ke5yvhrcwU+oKfdpcOVHugZFJf4IwiNwjQL4VWla5IxcfJvu28MBkEtSeWWuNo/1CL42Otycu3JB31CA+K3tBrXJDjwiCsw/jsroRbu9IArQcEJsjucUj4FA5PfxEQ+AGIoQRNAxTyScgtO5sPCwmbnSIipBrx1JqWJj4srBqMF1a0/q6T+SfXQTtOarpkkHHzOnWMRZrxCH7XZf/ayVBO3Wvz64RkVmMGDg25GLPCWhX8tNWVgNfeQaHUP5Rqp+h38IQ3rTjJGozTKfyZPVYC7qOb5wfAR4DTnzTIrrkVWmpllcQO2vU7s6NqKOvLN4cZH6vSaNXLhDCKPSyjNyGTVQcdVgd2iJRoSzRCKwU66GWrDEzJSvl666pwy6V8CgdS/B5AvsbRKSC/FfW57Cu8WJY+oezLbYc5wsn9DCUizDHZOyZFPI1UL2rDsuVc9+Sk+JnNbwgDlke45+izDuKNn1oI6FzSg/T7Ka1Sz9AknuIcHp5l96+dS8eFXArG8PhAcnzyXfDIKPR0yH3qi4mte2DIP5LfUi1gm2PM9RKrPtwQE1YL1YhVLJcBOpdt6ujiIWYdXzPZdNCFXcKsI7n0Ge4CAnpZ2Z5iyELwxVmK3xnaIDEy/qqEv6J3qBRM7RB5NyjIAXZG8BeKe+QTVzCGwoAZhH+VEX6XgCJHcH2vJsfyKZzVbQs5tbbA2hGtez1dZbGDmYGLSB9aOi/Xz1h+PI1YRpi6Lg4Y9SStkPFMFzBUUvk/Y6tOtvvV1IITWOgpTfLrpkLPYXPBqXIcqKO7A8lfmSM8Ai1IfLWmSROhVTJ5PNVk2K5WNbI6Qh+4f7JaSS3PqyNm7Rq9kGO7rsg3UizFxBQv1rk55M2Z0k4as/UceDc+wSVJCpKpwGAL9iPMGHBek3Bv3+YSxk4y7z+uOrFPOnxTYUydnhthpu4lAUoQ4ImPMnkxQRfVTUgsxhdH65lFqsIm06hc4Z8zuPCCnCmuhpl3E7+TVPZ04GISK2Hr4xHELRu1NIGoMEfXe3UlAf0KzbrRRTq3r2hN3Erw6L29FsfIy4lPvtYxbAfB/mWIoN+mrPjg/MrCbNSOKQJMawviRJd1AfDPUPEqStwI5EpKS+iTxaQUkSJsnyNNqRIAFu+EhMyvDm8mazB9drZ7nmO6bPC2cw2QTplrBb3ptdGpxsIHOdS5R0nhjNiqak0h+W2L4r0/cUye7awQ62Elahf0vgU8ZZkXfmB5HJF0FI8qUWK5UYF6anpSazvsiWvR6tEBdgT/s/m8k48XsVWPFAN534xoS+K+ptCE30mDLzMyl3u2+I9U7CO+wCKQaR2p569lWG+ehewqnEfVspxGKGdJnsl17HZnjAT0r1f6eWuZE8JUQ+3Mw8zdoAkLI94oAvgWf+Ke3I4lIWhi7iNKMBA1Dq+XrsJ8n6SkIWSXGJIL2BCEXon37o0Cug9RE96G/GUK5obgEhTnBG5Wm5SbEWAAA5UYZhkRvstdOhOfD5goPbL5lUaqL/wtvfS3qYgLuy5c3EwbGJDIvUIhr2wEV9Di0O0ZGGdqDJbCy/acHjRt/Y3HTt6h6ekxguNXc7nMSrbu0efgSA0PRf4U3qy2pHo94bSeZkro5uEHlCiq+d9R9c+XIOTBmtrWrvtIA1QO6qRh38yRvwwlNXJk1MNziXNRxLH1JSkylYZT/7KVm9binq+JiFEgIMnNINhKX2A6pCJty2621QRw6WJDxViFO4LuB8sHhjL3ZF19hp23HwvEN5gpXXlyHij9nxSkdDIECVWaxW11fi/UN+xkHw2SluAkNfDIYZrojlrbLMQjn3KXB2M3NEUis7QVPUDoh9NbFn5t0I3qwku5BpJLQIqe4bjLxl/MimIYX1XlHHmn/rJQv+ru0Mu41NnXxUdiLwSzUIEgpGyIQwca4NkDXErNsdSmAZOwVsGYjqEh72RMO1EsQhGPwzCcDNRFUUrLHyKuHH+n8pG12oHPYMoQIJgsj89XByjY+HrWG4grPdadbMCqcnSuUeFbMLRUGe+xkZuTqkVqostFycLrgaNDFDOZ48+aXgk0iLd+Nj4fHUM4neDW6TAFRQ9p4zQKLj7AAxf5qJYTKwvgGUKaRjt58Ibl4B7/vgkMGycVDf67I5gG3/Bhd+TyyWzhl/7FvnUc5TwM/GLSr5pwucqr8HRv1mBTrcKHrPS0Gg2QBpPFjmPylfyIiWyIyBqolBvEVM0cTlAQFm1pfbh5dHbDemyOESyQWrZNA3fpeCfUhxtm/07O/IvQopR4Mr46KkR56UB5ZK6c6h/HiTzl4lWZoIrEHCsUAISWSa3sEYzAdK+UzpSuVJ9pOQyYJLFNgbhhb7Di6XqJ4r5YgtvSniEMhCQZ28lzoNrC+T15NIaf6lf11J1QmcuO6wBSU2WDM2r0aW1e3Dg3bKks6hnlSjnH3cw//mcNMczsP3Pr+V55QROSSruiIJGyyHViFg11EJwvnDaTxxrLwlb+ApfAc9nZrCpTXd+yNoxF5w4ClfnDPIVeC0jQJIu5scZLKT8P8U110mdPbY7n5NQLBv2ZZw7bHdDhxBJ56S6UCMorHaJZEdvroxFtIYQO5PA0vlsMsP3K9XAIRxSf0uPvGS/x0V7WExHvw7sdYA+nbOz9qel6fFXQJrbugwSSzfNLurgNO5ooV+u2Wa3+rsjHkzaciI43Jbd4vBEzqW0r4JVbEA6DVdnciNYw0TxdZpFBOnzWBLuyku3isZ6pJSK81+aPON6JUdiCIyXmf0RrDGhrXCtz5Iyq/L8pJfT+nkshgSDNBbiJRkZpMqMvH2tTBSx0YMgZ5Fx4ZMUaPYxekCgbzIBLeBhJvsg/+gcb8cLgwxoT+Nt56VSrTkhq+5O0ejYipROyz4NZbCAx/D5qZ0RwYZnfLde4NwLby9NBtTMb6RJgvJA0/paLFKp67dBfyqhiQ8MeGE7WcVm3ti0xV2NrMmmp1NbNNFun6t63yPXsCPyMfp3UJj8irI7J4LLMH/2H9KPfcYQjQ5iBsCQlCE6YBFbQzeANk4oOw1NNumpxFU4HUflKTBizA8uzdpUv1b7p1VaLMicM0L2AG1vBPoE7sQlWbqqwaesq1kTlOqOR2AuixnQkdPZ1DTWq3Wqe0g71VJAXL+uPyRAFzN6aYh3a1ZP+ZiAnLRUNS6MZh4MRffvRIRNdVjzQp3V45uZ4fJhwFoA7DMwIju3eRWczRqNl4tSXWvt3wHqk8DJNhoDT0RTrCgT5Egv+PRYJ5bIJHp0AqkqRaszXrT0AZK2zCHPh4s13MVkdktnovQkwTnv+nQRB0XmcTN+5ehBS49KdTfBtrOehEbM2qy7FTGJ9RuDoqHNbF5cx2yOnUuElypqLCXgd2SsbM2OYSSOvCnXxFSiRHbuG7xPNaHRTeO3f0Wub+J/X2HPnB2dFfMYwIntigPvA69vn8oweGo0/wyTdCGGZvZshKYor1Mg3tn6iioPvTvItrqEjDC2gPsiqgylve1K6+lFN34EKLtT4KYqYcXD6b6ly2jzfDV/WwOOlrqJPA2glMhfDMcq49eKdsAHzgTTjmDrCEW5Kf9i561PHi9Ztfx8EQn1GaOcEZiOZLxykOojsgy6RB+IYnZ/+QzjQ7Ue2hzk/Zx1FgDiPl9ufkBnPcdD+kbPy5BVpRAo9s7UcnUgSmT9rmxTLYrD3lNaomrQYgS21C9xfs4OzV4ppdzTiqLQXgdivzBSSrkh43KQCkrmiHOpv2fTJeALkK41vFx9OzO+pBqJRE980tNkkUGfSJ8vZ8VRY5FBz3dwPyzeMVYKnwLr6kI4YjocvoCHQGeZZNdLY0OnTiYfEoCV5SQUb1N2NDMyXxRf13xccv0CRNSCfDsUGiz+c/gC1CM6E4KJiWl5TakI8rVY2jEfXl2Pq85kcWvC0UoDks/Hv76YkYGZj262f025873ZKeiWkWJ0DEwyh/pEsGcfcsqDBLGTtnqV+vFBKHYMliGDzz8bVe0B6nthG9Q5YIoLo/im0h1orbKbC1bPol3wRcrhGZ2uhO0ghy1ttHiuHxiGCEdD4kKqFkRvrATmVfF6xFatnqxYpK0A5E65lwvd1AvuAsjrz7EaDAd0g8TV1U38sSIVLKg7BaOdujCjpAZhk88hbvIqmJK7a5b59KaoVQCFcjPsaUDSgd1pKpczTyWvtmx1sds0Q2UAXpkhxcqNpYh4q+wDgVV7U32u9lkxoVGizKfy2dWbZehEqLkRsb8yee1SojbAd0/SmfJMoJ9xVZwumZDn4FfjDMcwQaRrUPX31hJus+kWCw3gUrm1YAyedK2ZnpEzidXp+26YrVgWEOQip99hlDcPa/n169Tu/mkWtlsjxnZxqoXFzoTGwZF8aIhcTjlfteTAp43oipr8PQXjce37Icj4JWsZmIv3eGjo3eucuLKxPNCB9sub4nUz/aCQpqlJCLQ/1xVaIAoD9TqfiPxzAcF0eiYy4Fee0vnfs/P6PfdKgut8wtCSAAB0Vd9zWSlzFhetuZttA5IKx2dFJ5gNbhQ9KHqeieJ72/keSixOFUmLqTXMdW0KNFR1ucRYmJYahyR5BXnnp+cMihCnjXx5VomXjMDbdlgBbFTxlwcG1nkB3wax5jFzxBfwFZhrkDM0T4DudTD+sCbuTqgmskFQ496fnQ8GeMnnRm5JT+wIB+MM47coFgK9oHA9n9372ay3q4nM0vWeftChgoooGMjxes597jNkvLHPq00KG0hocFuQD8SpOeVWTaXY+0XACNXBraCAQAVCczI0+Lhacfza3Va1Mlbks3Suxd//+t2WjCfwVLzOjlnVYbln/jru6jzGV4hYCG/lY3YyYtF6/PLhAhVSHol2m69eXpaKYPrYG3Dn9hePGp5Z934yEZIRACVGh44FxxDj5zVytCjypLe6w4yczl8+1VYgHHvYhW82q3KXw1yfVmE4UpNpMzOyoda8+dgCdFvseHAEsiguSwudm5WkBm7hm+CrZ5pwTxiYokOPcv+y3UKEQw7STd/Kf8Tc4sXDeDVrFcxq/1XEZPse5yM/TqF+iMEMlHqAkIoDFXepv8uE2l7S015bxCNJu9VmFZPhZBOJU/tdZzB2RPLIPqBvy0X57cfTGUdkdCA6zcZtK2Zi17CjYZaBrH7c9LpbQZKic3Pgn6vIKPCOSj8ijm0n1CUxvbKZI0BXS58VuHRe8ntlKR26Ul0Nh73dqQOZHXRdFfxQqC/Of5/PiaoAF7mcQ1RxhBT33cF+sPEkKmdTrDGcFq7ZypC5LjJwlzMTe7soDF7UtoRMpIRMZX2zVSbFTjzEf8xDtEvUIJc+9vv1cDQ4r9W3rnRTwRI=
`pragma protect end_data_block
`pragma protect digest_block
55204e8ed54197cb4e713f7262fefdcca84f71493936e9c2ff8dcc105ee02acc
`pragma protect end_digest_block
`pragma protect end_protected
