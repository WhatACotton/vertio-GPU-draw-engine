`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
+BRE+CsP6uH6sXDblkXTOZe39hI4gLtJMHvYjnbZlU16nJlhWp/+LQswn+5SEcMOv4A9XJY7rj1xC3h+1otYath4vlW5lqg+S1qcEzm8DUS6aS+MEqbkuW2+89hJRnbbdOkksbXHswaSX1RhdwuPROPb/DXCXhAUTljQZWaxbrIFHpCZ0qnaMXPOjkJ38Azn8hiJqQqpafrPJbbuFrrG884ySxjdThn0l/262TPBTTjUVqOqNpKucvwozD0s0Wz+xQfnEMDck7FHtWfM3+CEU1cZa5J+DWfp7OLowrmnJYo/9RPZPNpN/BkfvL0my9jFvKtr4zsV9+SxfOlPBMIc4LXjwUuce9PAOHybUk/NsYLHbzxpQIS7Eq2HJCImWOLRzGdl3lPBEE1zENfxUAc1tWq3dgt+eHVMwcIR1pRtl7uUec+CSSHUBLHAw+inn0xHp0gF4KzDN0UBYxOqerb9hrNNDhmePmun3cWM7WoUMpHxDtewDH7rwvglfEJJjIOkih7WFeKxC9rdouY2/tsTNR+jBRIiNPCfjfx3OFu8b9FHNQfFIKTioDh2xYZikFvaDBDR2NREhkfhfNgzrbd904I2pVpCTbU21viVr6RWRQy0k6W4pEe7PJTtta90KlabdRXtBkrPQ6weaTUyJbxHDU6AVY0YDwfl5GbrdRkyqJlluLvnJUyGexO889vP+6pzuLeIA9rPMuZqD18AZd6bLUDezyt/d7Lk5xPoZTPOxg9yDCOtYz2GwudwC7IsrlG7hpNTFTNaWS//9W9MSlnAHsVNgb3Pjp5dMyRgiYqa57A2x6sEcToQ4LNbnSYcZ5+eHMma9Zt6I4+XQGN2umDHET3Eotz/P57MkL6GKjFBQHUcMTodiJtSBsZ7wEWc4VyOt/PbXwbm9WO3xZDmHoP6rXfBvqptk0x1Zf8jq1BesowHzxYLlTGdjzm34+tBVbXB8KVdX1BpIcFs4NZFJZip0OeIuujXgHYRQFMvJA46GzVb4HflZy/DTLX2l1n19RQ5lLG3l04ukO5v5IC7sa/g2q/4gYJAnwRKdU5Djl1NMqu9Y0223zmrX3vXR+0HreVnJOCB2EDDUji1ZVjjG0O3XsOQxs2oFjMGrJMoiF7LN5QEjKxDaB8hHVgVqWi6ce6mk/EXcYrqD/6yuIbObnBWwoxfki5FoMo14aM24rf50v1uDuJh8kXealHVa26p6fX0ipVVY3YH6pBApEYopoqEeAepiTSl4q0TBm+MMs94MV2d0JyZ60fv+PKbs9HC5pJl40tsuMU1/KQWBg4OMQ7INxXSuruOocVb4FthDa05uY7IYjRdAfcZjSMMPbqJPwjWrmCLLJEGZ+T15Vyv5703t/4fEgZOUITljAi9GNmL4tXPsVqD5+BflNxS119+RnQu2ToXr0Uyh+9+MjdAclRug8ql1uFKyZGDoUGrHmZ6vRTb7HVPdReyDY8NEaousqGRqr6vsmp3VzUp4WV9XJNcCSDcKkB5AyvCUYCBAT9DMoNqwf9VAs9fUhK82EETfC5E1cInz4044uL5HIccQ0aWDEkvH7y6pCTtlsPRTyHuQlsM1QvAqwBoNFFQ6mF2UHHnW5CwBJaIeN6QDzepBF5PwydZwAIAPmH9EoNpaFkiargJv2XH2lhCTLQzaQF/g4FeqIMpzKuGzkNjJ453tQhDe8Hcz2+hmUZGxte+3/xWwt+eOmi3nJJzZ+H1G3FUiLTrDc0L+YvVTGiyeTfXEo71X6wezLnlLuGBPAX9kH8NP6QzBgb6r1eNL9G/unasseiDkwCr5X4Tc9bPOd1USKDZP4Q2JHRANdlA4M/gVr5MCox2TbGaUnPnOnTQnZTvs2ItG0SHYkGI7UbFRHnL9x6Y5YbC+nmVQLqpEWuDU+AuSYEtfsjdILVpF9cPd2Ukmm0LChLo0sUHABud6qVYU/1a+eTgamtSJbSo2WL2hd0gBOUtR+1lXwTUU0gjvto3w/IOP/HkncIKNDCVrXq28dk16yWG9O2UuOAku7MD4jF8cIXvh1shU+8SXm9e8maMwPM0PYDC8nO38OeGfkDHH533o9gM15DB1Y8tEefNHay4Z7jkFou9M8gGCtugV1gnPr6gAIOrfksryu65Uh9qYfdUZvR1Yz/4YMWRwsFXv+bmTlRNnWkulSsH04LVyExtVKwgrPb8ozatCiaPGyqp64Ep1pcIkD4DZVo8Qv7AEkXBvh6freQsdse1IgcREa3QnMfnFJgNlJfcsZbIiMZu6/X4tmgZpoNSyTi1WLtATpsscLplvCTZqpyTFnBnqaWVpWcViQ9H21/JcwUtjG2s7r+lCxHQgYFNs5/LSut45E+wym9SQpPA+nZuncgqVq1X/isFSbFVR2cpB+Ea0P8pGOmiEYrhXPjgoBrJ0m7sxwiWQktaLuuTdf8Bm1TZ02ooKri23xtg4slvNnIOT1hckMF2HaCo2YSmGWqFMnww6txP0gJyKMyHTz7kcCAby2sUrFmfS8LtuUqs5IUFboV0fDCr2sZoGjPx1dGFfVvsRSEm4gz12iAPWHpy4Mizesu0c/D5yHITLn+1ceXxR0bauFF3X7v5klrQzK/I+dI87Gozv04ABzqrCOPUjgdhbc784pXddCk8fQv2+bzjZtK1h5/YM0TyOdywuV3WuA3NzjBBG9D8Vs/mkNgrtc3ijrdbZ90BR7FNdkeGgMdvbPYq1CiUu8AOFkxCBkPSWz5ns9lQb3CiYTYfOWdmt6X2TrQAIIKK/7c2iY71AI2dO9kaHZpZU2UzZS8vU7sm4iHPf5KOqULJtmgGB9pM3iS2pnX1hpLo6OVXWNqJD15CsWR8L1u3hJSNCS/2v5IgaeKfO5k/6LK9J/A+ou5Xy9SKgLDVE6swrPVeFb1im/JeihwCMoR4efOcz+YB7S7YdWmLq3Xzsm/IxbNHMDaLKFhK8CTb1BlIXNEu4us0ZzIgSYqVksKCiOl650nhylvCJafVwfATdEE4nc7DB30IShK3zGOjVqyxLPyp4pMnp/oY2o5pmQOs9e+4xJstKv9R3ZZX4AjhoT16sK1cWpjjyA3tp0ZQ/R577v/XyKFE5YRka3G+eyGHZb49Sq0JDQKFbhkI8tckZK47Cx6a6QLKTNiKUOvJHJnq5reKAffiqu56YesUgX/3g9gc6h8S19i2gsBx8SJoau9/5oCihIwwCrYOPKoEIkwosq/TwsoSqkQbRPa2UXYYkJgrNKHTofzg8iz6twZ0B48R3ZW6Pk6eNdqEv21W8NhVCANc5z3DePukc2msHn9S5QE5jtwqN4UsUjOqdUsY/zokY+/N/hJCnQMh4ZjkrfjmpQYojAv2cxVB8i1TvCreYyeya6mT1EnqvfGT8YFT25imD7vZ94Q+3LN2nDsemS9f3RFx8N221Sg8+WnAdKWIW4VMx+y1y7/2Ra+WIkavKErBHHSGJDLxwM41w0s6QIZd+Nq/HnK7LWzayBjQyqvp30eVYtFG7nz/Gzjhf54KQly1+qXoGUEPyvUxOOO+YrbE2kaYbUppL6C4oXPvAZBfz87RW2Fyu7J68xy1XvzyS3uE5CpkXWn7SS47bjTxJpFFWOiPA+GytuSjDGVkKvybiInlwt3Jxjv7Tukcuph9DyNeETD8pUjOn1lfXFM6CxBNralsrMhwb/XRyvOWjhd2H2c59ttC9HbeGvgQRHCrI9zGbr5awcUI8mBwgIdvZAGlLzooFdR9MFeF+Y/Ed3OTYytcp/zTaY6wJOqGwptdc+7rapwB+m3+PoYBye16iSVWgm3EKyfWz1vek1ODFPs6zbIpEQc9+O4zr75lydL5U/yKhXUeVQW+5A2mNNhSISFMOUTQh3vZyKFAUTx4HjzyppnTxIRwAZ2N5RhNwgkadb+IvF+2A/Xdo9y8Q+2fE9l62v41r5FhR1X1ujKkwkunN/BMAYVINTGeNxGA/vNuXo1h7nTPgWtZ3gPT5csHY479b3n37wgmWiI7bS1nysDPL+8PrDZ4LUVu3qknihXHBN5DIJkXU87OmA4ANvDCGn3qUcz2DSAmaz51wdtUYNZpv3vnYvMW9wntd++IOR3dCWZD8N58wny4447HKmP4SEsvwm5daU60xImi4UWXcG37WWcwyeuDARUauqf/d7kVbAaAa4RQ/pzyZYBcHE5+Tt37dXV3TZCgK8kTUs4KU25kFTiKOUc5HxCCRcMNtLzmypk3caJoH+bh6vrrnQAZqszr3rLuLDqtglPL8eZrdJw8DnHxD5l9Ll0wMc3RWCswxSKaqVynLLf8C8SNMFXWEdRppGcgcMm8yal7cEcyl366VDjsy3QZl3dSKqSUD/JqRJDkcXcnuiW4eY90oiJmuDFZagVnCnOENI+06FttacI13ztx8ncZPPvXpfuMu8SlSBP3btMuS/ubhP/94GdNsCcIOWl73Xt5E40rgW1IHqlmSnEFEJO0ceAE7nRXl3mLjn63b1TrqZ0Jmeox8jMbu38AJ5ExeMMgTHXejuPtkN8bi+MOJolUX2Qlevmq9L0ozwrzTbaWDO13EyZVLdgBbRg7KtZjU4bDG4ikZuyNsuB+EwwxVf0jH8Duko2FRKLyOGXHrrbTKymMagZmgw2fAi7yqJTpbZSiiuj9AmOM1k5TVZk2VgtbLmZZ3H4sZqxd4GF9IPI0TZAWczO6m84A/pUIPhjXW0iNVVcZNLC1cLhhZZb4VBtcpp+sY/WIWfO6hoZ+CmkktNdOjFdxMZMiKxtolVfMowPEs8Tq4OihbDp2gu/fdcuspMrTupHVlUhH2ph48xYmTKQ4rtSO1oYZgKTdSfh7FLm5mV/Nz4hBFlBeDvhQSxLhRaIu4vMaWQteq82pnvvv3aQPwguynWkPTQs7CxA5oe0ITkfnO9wIY0AvZpHOSAdiHih0ZXW/42hRcBtg8FIr/hFDEEAI8EAPkINJfa85uguIQEFc/NmaovlCC/SluPUBG6JV2NWmqRst0lNktAfgoa8zubK8DGNcUoe/ocCLQk4wT3UPSgRsmgrRbFGJ6Pe3wCgEHeHlMXmEFEMAJZfc/GOzHcXPQTOc7IqHrzOhpr+ds8WaZ9Zaj4TOk6ph1iwZ0tMJw9DoG5+cqKoKiMcwGR4oQRvo2VYyAWUuvMYrBYB+7Zv2XjZ/Ap/AK2VNMJjXqGTMnuUJyfovcyb1KbgLEulsYs277aROrMt/mewlBh4RxSA5h5lzzKbVlJ9z8aqZ2uEkifzC06bMSK6GIzobzsF/0+a3peHFDpmELv+iCE3Jn6ZGRWSa7Mn5Bj3s8gWv2OydgmmuupH5cfyFw9Edza3DmyAr7OJ9AfAwvuX6nGUwef/kyWibRPiwSTnkiLGvn94+CgHhaO9As0Qm4V0wbVVyIvHUX+7w+pTuwFgdzqZoJ/ssS/7BzJROoPR7yrpr/2GFOANcSjs/+LIlBx7cg9fr0ceoGnwsSqDKxa53pm09GB1rskCaf5tL7lP4LbeS9mEy8/nc5HIP9IuIbi8Psnj1gD/YKcS85kR49at8XNuG5rQAZUDsC7K/6A0JlvrZjueyLyyLbb5kkgMu+HImMltfOA7OiNGZdYHe9OHkC48+YH3a2RorpiXCI4CnEp6SCsjijYQ1S5Uh/N1z/ZOhG+pkfUfMQAc+JF9GkK4T9gIpkaqpgae6p25BtOiIYjtyAj7Tuuf139tif95bCLaVDSkTnez/xJqaOxz6e11gjdyCjjSqfgk4ZApeOukTlh2V+R1DsjK8FJZIDBOW/GfXtWwA9OHjRCT5whcyRhGk0JL5WMr4CxpLS4lDJkNwJP4VLWIk1r1jcXgBv7OkczUHO1j6XSjja2+bBH/M5Zz8EH8sDPoK70mALJf7Bts2fJO4YXrtnUh0ZrC7kRmLcXMlOwGEnkwDeyDlwU0BJzrg+6YZcOa1gFx9x/V6/HRI8sO3yREDXgs+8/lggvHoJ7nn7w2rCvFQhOSQNTEgxsBKcbbFsMbAAgrj0esm4kQTZSgFNGwyJsQ0msvCZViq8f+zKri/5cSQqSPi6UTd5vibJ7Xo6xKK3OHHR5tDMDlZOQcGOJDUciyjLR7UoJJvWKSeEznDocsNyWoYuRcX+jWvYteaug0NxAsPKHYJUWvFvKuAukc+Y/uOdLycd9RCwzkWx1RPW++oFkuHjoWlXcDaHNzFnF378Rd09oZtaGOdXubMk322B6jMZYGrxneLfTLTV6gWuJcDYS3Y/JHlzANtlnf7MnhRVZMW8kw3LJX1zpEyCETl5Wv8RexrGZRJRA4yn8QDgKJWvqRbGImIlR0s5794wtquB8zU8/VN4d2rcBRktuhUc8geTCiTwVgJqtKd0S+Km26wyx6MEsglu1m31UNsxJUp529eu1v18iag+m+lrBWNJ2p9MeDHcawKgm4R0yy3FxgWC9FipjdtKfoW7Y4fFusGcO2GjoOKGA71t4RFsYYFybiGdK2GoruEd8tc38ctdbq3CfoAcoI4cy1LugA+lBSf+4H5bqtjeMITzZF/SajIR8tKbdX2zPEHQ6WBuPP2+3g5PzbnbnD4Fp2z2MEnfah5UlpEDVA+fyOZ5W3jnkfRzi+2B3zy7/ooE0lmiYy7Jss7lvZYaHfimc7QInhLW1O8uK3DBl4ifn0M6He3UOVNExUZYTTnjQbBWw4OZOf5rewvMtub3PscvsY7KhiTO8OVAeOTcbuJxqj9G+s2JQrH8/qZ8zD+EfiUxFM/1f6yfYZwFrDuHnqCWZnsPxwMVepXmJO2+BL1W6uu0NP8BXnsSdjyOxj6scDjBEjARMaAco62Q98NXqpAxncyzYWbeVtqFTJkxQy57Qv9AeAGyNWtsw64Rg+DODM7vBGux+DWnJ9ELVFg/Ys9GZc8wAvCutYuda7cMQpej+iTAr6Wgd9noOutiOvT06nBSM2krauiIA3OffSJ5Hw9N2HeC601MP0h14OI+XmrZP3arjVQh7NRSa6LVsnzcksZ5N+AL615ASsMOAp/Qh+SlLZaJD67FlN8cG+FtS4Z2jQMKLna7PwapQCFN4bZSNgX3pOkqEt3dYH9yPGpgOf/6Pt9U6ikFVVpXUDL7cooZ0qYn4ZFPWWUniqMJesoTxysUXiGQfYcYwv9lIMZC33z9dJZwHowwizMNDVvsP4pLg74upM1XzXl62tntrWzBuW05t0gycATxmBbJcR9J/ff5p/ll59OoCA/DyfuohEQaiTGSvYDEM8K3INFgduD4bM72CcaWY6thCYAJ1O8/YJN/dO1ekZFa7NWJRXLpOvfc/OzYlMRPyhpNXgXoY7xK50RKti7aVum9cclvRn+YJtWSdiLrZqKDb+gCkFA6MFU92B9O8f2WGTI1bfrL5yf2THyMrliqgaKG4Y1gfis0NBZ/Q/9T1Q7oa1I0Yz7XBwVioVWzc6XUr3lM5MbPRqBtYl7THHXne66pKPiVk+d8aw0MX3OY/Vb7PjqrqsGaku/AAg6OGWg1rYsKg3SUUwgwIXf/JBMPUp2hTSqn8QqvA8u5DU3JOiNU39e3eLQxjdYWwL1WAMYJ26Agpo7R22BAMsvOKmIh99y24/jy6WubzD5VMlfjv66+YJ0NnBy7bc9dDrk5Y0sN3P2BfakzTIDi48r6MsYvnO2aSWzm/RV5asCcCDuzU+LmGPFOI9NW/y3hUEIsQHEwyZvYmX1t7TIsBCxQbiUjvHfGi7fZTqx8D6r0cK7u357G1N/ngdG7uHP5r/R9Fag/2y1QEkfsbHv61AkvbdGGDWzcHmOSEEVaUSCWxDN8EK7JUxmcSAILDpZTRq8Wo+jDyc8yPx7xsWoZIFS8hvt7m+jTZ8kS/wkDEAZ9fQPdvLef0FkD03QO/uJu6v7oevU+ursgcMuiT7wlraBwbNkZz56KXSjhsdVctF0fhvVqQpFfOH5oMe5GBJiL5bzUJwaKRRrvtfK1QAg+owiHWwKNGrQ6QXjEL79zNfVpy+iRr4ENNn6+sUa4wR/vYMFz5ICtu6UWTy3JmFrVxnTWtLXAhYKMruksakSoXW0dW+0Lr5EJj6YIOLonrlxnWVx0CDNJb+w+/XNejcMs9RiIDpeiHcwV852ukRJQHqK4kRkLcbkxCPawLY9Sf7uN1NpxjGJWG7DH4YKf7gNHV+GtDoI0EeHr4AsAeenLZ98URiwEuCMaFsgI6Eka07D+IvlSkbhCFPNzO86MdDTRgo+DRxi76wvYtQQB6W8aRE3QlMyqD2LoUIjgqr3/vB64vGOogjAPt9gGaMgnVUJhj/BNTTsOEC79A8Imd/ATpISVEXj+IxL0Gk9bG2oMm8ozbDkuWhdAejh5bhKxaF7k3Er17xS3izfiElEwGzcfbX/uBvS7lKsDDX9aHaa7RlRC/ZJ5Rlnl+Wvyw2oeN5Hhh7dFghFlCZIfB9v3mf0C4LaX7Ee4U8esrFO/0FtHCiJVJaHRng74//ZkdK/FkRWv5ChNwFSoVIaNH/Zw8HRho4BIeWVVGGw0vlchA04UibyxWASgwfn4MwlJs4RBiL95DAr28ASP5KisPuGsrfzAt7uZAXBB8i8mpH2sjuGYHJguoe8SpnBWBa5GkcnFHpqTdivXdNR0vH7qnvOee0g2M/rHkWgWzFFlRnng/HV9Lk2NmuNDJfTfWYJsQoBi7XgzLhskGksq9tifcWV42UJKz0y2MBlxXPk+LJz+bGtVF4+EZb1xdJBYHlXKV8ZK1WfNWODDhp1wgpe3btDc0SHpNDa30c+JQZnFfkNY4lJeO3zfXhMYeFjzV88W4/KkyiPh6I5bmFPWEPF3j2q6eHI45qhpAssMGxBnpNOMLvZ8sCz0HzJBquaaaOb+SngqmNYxfZAkfC9z6zFWRou9SnZr+Z8ZGpCpo2qQGkSw1IMvm5B9AJqDO+pT9ZPCK06uOPRSRMiSBFIh7JAWoAs0DRq07Ur72Urd44N7yjDMFG+agOhku9wQnezgDsDc9b0lVFAWgsNkvwyusTUAVGAGM9XRs8PRubimwTzuHqBuxu+eyVKbWJ25Do9d+OIWkpU6z/8d4kErJ5HCzhH0+Wl5lwdMA6i30c59MhSoWwq1jY4jFSyA7SzBNytwifTI9unHFqCvHtFvnqiPWwErtuSJX94tfbrvcMyCwiHCSjmLrDppMRfvyXA4ca+FZm8JKIySTOVtE/JPRFSLyO8sJZVdyKYTcEykOnADTwkxsy7sU7gzQZFzDIM8iaV/zWnZD/976wxnFY1C+SebaRDIIGrscmc9w68pMkM8VQoSTZOyDMvKQyNUQB2VYY2AK9ckOmjbnoZuK1WYWkdfg6i0xdM/aT+ZUnjLC3rtd2Eeba6SvxqMiOT4dXYO9BgvdpkqKdOx8Otqy5QnWmeSFj7SHTW8VjZ6b2DynWFTr2xd/+wlCZ/Paeg5rTYR6GfPCi8yucK6vnxgAEqRwcoecR0jr4c1lu2G2Pg1/3tY+I3z8TTkvrlaHxEO6w/RUMFh83e7A7eMKWgOmrcZUH6Ywh4zYAzSEH86SyPaoL6X1jugvDOLELylAMJ9TKbhxskkry+nmaEOyb3Skw1q2UHPcHX3mjUtGOHYVs90gI5QXCqh1l7C7pqY/7XMyP+T4838rYrSTqhhF7BUiYPNJGdWLjuuNR8QvafTArf9fsSqbsFh4pzEnObGICLBLXdJIHv21ANdNhQPOyZ+qynSA399YkHucpocHYXYCkxai/0WigqX7Js0MwIdlXIPD+60OaxGUrK5Acm8KsVJa2klyyDvvJTWla6FrOymmDic/WP437UTVtg5rfxUEs1k/d9a7JZL0U7+/Xh4zXEjlz+ve/gikoN8mRhH1wm0kvTm0bbJDikR9/sD51pxcyvH0lR21bCSAhOgL3A6ADsrlmF06g06APbstJgHxcpfbofbHwXJrDpOxXIrBH0uFxb8mTY6yWyrT2yYPuYyLGmLveAHLYBTU8UPptRxQ1wN30Q80vnjVXRgfwkZ+TeCkc02N8dd42P1ZMohw05UqwVUlkCiQjjiZs019YbaNU7TptCVTeNgWkwiKXkgpF9wSL8AdIZADD39wVKJETOOmAR60b0C8CyAvmrSSisIB+MOIOvwFkQmx8/V99rW6DJCq6Tshj/vnXi8aGU0lbFvDE2j/JeiHaZZngjyQUB38AADH/0MF+6ee+EgAE6n56ItsyObTrxtF88HMb3vLssFi72VDvzdujX6P1oV3hsrlapcdX6IN6CiqmaLm1yVtoLh/azClPpdXMb6qJHAmNnf7tgGlDVjAZuF+sGnI/SYx0WB4EbkMyM5cRSJvs2q7jzGeNDu9Tha8tPVeQRpr2mHwfjawImd4S78xmsVeHj93RRInN5ySTjf0+H//O5F2peSf0BC5Nj6BQtCTbCYOwYo/n3tSrxUwljsFWkAjm0kdPit7Y8hjNJ8jEeDbXk47iAO4ZxmY1PXaOquEHiFe5g3uoh0JsQ3J1swpBLF/91wqLewJvZX55avEdbHxGn6kkwTEUHPCTn/60yEiqHDqRK67516Ezc6Dpzt4Sd9VjgO9WvI41BHWptDf6YQSnEUOgN62Kl2xQmzUjQn2vzcwBZmEyLCIcbZc38rd2gc6vPF1bnlwFW989zqXkrVg6KvkCQnoR8EZarWWYSqPK4Lm0/FXV1qiMWAMNVz3Udp6O5zptv54DwVuikEK2gX4U61d5IdQOXIqY55OBuzXyke12gIuP5mK102u3nWCwDLRlLBYqTXZSZVGCmE/6M/hov1K02Xor6Ipfic6UCVPLbz5sp+V/kSBnGhEx0l3sW1hGzQODSSg5rNtphJ7uiksJJA9WUx4teEoeR2khBTRuajzFaDWPOdnZ2cZAvuJNpnU7Iv31z5RGLnHih/eXIEFZXt32LShPtfv2N/scNCHGjxz7SXptDqS1R4z0pEL2T3zwf3OiRWDetsZQHkGeDvh5E+3V9muaPcBxAGmIrHj6I+hHdgRlwaXHyGXP3heyjO1GSNGyzDTv+g889gKKMCCfacxz/9ae8HzM3ni+cFTOKjPZGlZDnflcgOXFjVHCuK8NuZblfodQdwECJBCPEjo4lYLHCeshsmNsq1F0uGj69dyLsVMVYrnobljHT0HdCT3x14jdA2tPMdHM2prtMID9+CbkYkrVI++yeRkRq3fbWtlhP0nxKI9buZP9QkGEvkKdnRtnIdyMoHil63z1nVE9vQthsxPgw+9bJWVa5G7IKpVv4Qj4vCXUU3dGYTrS2ejTLl4+3tmhM9l6wNPfx813Fz8s4ZWXmBVFD+O6TbI7YM/GVT/UtpFLrZSgPlOl0aQqXJeeM9XFz47Yr5DyaeiFBTu8Z7vM66CypXI/oO2W34mOEY6+9nyYofODo/z1KiFFv9UPEY4+65d+i6hP7Z1fv1Kok6XjYiF/7ptrxU4iGgn0fMqOkW6Hwmuq8HKhz7J1UV3FFifPovWwWEH6A7lDHs4HYMYw02GuoFZU8h1HC5tcHSx5ZpkuHDnZo6dgf18ueCYWp6opAvhWg52BlClxU14EdlAp00r8qcWOKDS+zynHXZTiR/HIMSdUbutcXfJ8WN9mploXxGpwkztjGG/5BSbpPcGHjXikyB16eLJj6rT5XdgpaFuMJhjhrOvz7oh9rxJHJhk/apCQhYIWlAEfp0S9FE5+xDzXBKbrKab9Zi3HIYiR9mijjBWyNQrANnRFEHxa4+vluV9zFewFjkHY8DeUwB/YCrJlrRs3jYD+MRdfB/q0aBbaDZKlR3poBM9pTeIjQeJGhj3AXqcVeHxYfB+WkT1iOegJZo/YF5VmNw4X2vsnYae/tgsSp+Op2PtDvb/HKA6YfVAvFT8N0syiUEN6eRm7+pDanrYxDYkxz5xuwleay9iaR3vMn9enSNMjDGLSm7oGYoughI5OKNwDQfRjbBoShsX0/iIPCHZwA+Ek3VSEkDBTqy5h8U4kmnC+U7vg11Do6dx+ZjGsnWa5k/bhV1Fn9tDEuo1X3vL9cuaUJzmz6AyEd2oRyED+fAhxd5/jBzYVGvVs5XLh/etdgb46J8zyLr4biuZZvBQLUCy14OUMJz8YbuxqywIerdv/KP2qEE/MG0j5DWG73yhEqwELXzI3l9iOjFnjWo5r7GFpfEUZddSJ0XhQ1u2UROkepCZW1Pk6j4uVo23jAR3x/5a7YR5gvzUfRHxGq0jDS7ryXLdTZdvunjbXMJvpUBXLAC0P551n4GxuGmwL+MhiiuXb9OVJrX7imSNGamjeIR40Cq4qaaSp5wVptJ8x9lq4pgR6AUfxG6SRjhNzpk0njAKlmPiupR7BOH2fQV6PYbQ95yLmLs6NgoDhcrgdd2UZg0h1dmwcHTKPVxbIoIgorXmTyuNLz2pbuEJMxssXw87orPaPcYRX7qgNuBufZAZeGG1KRgOZ7lYY3VzsSWfyh9HWm8sgDQeRkKFNt++FaN1vDktoHEMH2WZw0qbh0qTLzpi8ROR7kSbMzJJq5T68cjutSrOHXMpRf/3hdRsbiJ7tjYY0tRjdM7PMPZbXsqVe914cbdhGDuSvvEeNIGBv/gS88rmy3tmgZHO3uTfuTYLM7TZMhhli66ZX4M5eHqVKREQz6rGepKaJn4gJKdwDgFzzYzSf/pIrT5xG2FBzPVNORJDGW2QBHIN+65XVhfHmAD0MUdnl7ZaayCeBXhyqpn9/KZmsZY9Q7/6oibLg7ghzZ2rhf4mtP62+68UgrfUugUTNjszdb6oj2NbTmoWHtsYBxN/4uNA57xhbu5BXenzEWQ/5k5mMePN/F/hzDAP+Ltp45dLtWwOQ/3tWBnuwL4vZzwhPsQzJnJgscR2WjzHhSIcIic8/wS8tP7zdZmF785qIffOkKL+oof8ZyLdaUKK1BepY14JGm2ee5Z4y9rwa9ZmQz/TtKpwDgcRUGF3VLh0g1e0Yr3lMNTIimPQPjb8s4iDlXv00glVR/pLQU0UHP6hhaMupC2sONZ/ydJ/qYTl7o2/3K9T2QN94jgbrhNef7xYwFGrPQGdcQu/IA0nJJLvzIXQxecy/VMvupo8jz+DFR5Q/jirMMIgobUFTzym0zBAbVCSbrZBuWQtMbynk85qOQwWC2S3wyeqxqrckO7N9bfZnNVEESi5SSlaWjMvvWk76TB4UjJSQuuMWg/JBH+TFomoQye9LFhCJlaTbC8udWT+l3uNq3fEDT5svxXUz+hhNrvlBJNEJzXb3XyDCSsHWx4dUSWj6bZfERTPeyCR/xNIcbm+b59fxIjLjN5IMFfkInKUhqFrbTrdGY5BZwZJSfzHu8FUYBub38Tru8KPOq/6etuxd5BnyQzVsenta942/+QaMEWAc+mb1YjFaNzp9EbIieVLMuc0IiLu6zUdVOl0lhdTZLZVWXDQudfmKZJddC9nVcYanF8EHN/5LELbmIGzLS0Yc6R5sEUFfak6zxVu5TrmDakcNLsugmvOMoV5mdmkLC8xAcak63iOyMorOR0HuoaAd/WaT/g+R9ceSpUd/+ZEKNA6qvDk3UBiD7gnDjMxmCzdPRBRpgKwIEF6EaUdX/T5kli7rUr4VnUf4sa9DmbTJ4Chp8A2XGQO+Kh1aORUrEjasvrZ+XOgvHCRBsQd7nFDXszMzk+4Bd2dxoaKlJQX8TzDivkkjmuvu4/3NNWT4B+nujTI8On6XBIy3y/3ezu/ThS7CEaD4plw0HHDeUsjG8qmlihOek3Ddt3KQolBHAXzjNyNBDmPMJGkp7vfGfscAzqsVoBWZQhHcO6P3MwMBrOFeyc3E0sLGWq1X/77JIKC05zevgegqaWzLV1g0ymfmFa/QpeF/GRCJ2xAjSub6DJ9s42JumbJ7d+X80hSTljlGjsqkMSG9BJ5So0eNeUQC7lvmklxFLGO8Mv4gr165rSw3nuzECDDSh8gLdaKgA1rOyM+IIMpdZaqooLetZNWoqJbpDirRSVQJmoCQj3nGP1wWTtR/Xf9NpoQiHwPJExFFcHA3JXrXB0t0g1HB8I4ALfQbJkl8mqYZT3QN6d48ExjY5cYXcBkRz8kEnz4Xk7jQROiXkKFo4gfSR+OMq8Bj+1sJhfpB+MY1QVrWYmEQXm9yyxmn/qJxvfhxNUFyagM2MPTvyQKHjyQHXtwDgngm5UoljfT1SznueqxYZlB422mp30eq0XdPT4keKeGaTh9Cn2Fuv0K4h9GHLB6X6C1hACe6NfQ4ii+rvsTJLeQIqphBu1Qkgq4YJlPXrRt60orOxJjVnKgs5g/zTThHbXOKGB4X3/jyy794E3TgJCPJpdaklEyxdFea9+I72hdccVzy8YIEOY9shYycigwIkvdf8QPPqmiF1U4B0HfErlS928pkZGgH9Aya147sNlULD+CLHLGm6A7qmf9XmQPNIZnJEZeGMDtOhSBmPjrOX0NkZs1j7HLg842US9FOgip5/8x9kFZcvnwiJg9hgDeC+909mmDJpb9FP3nYozRzYLQnrKpFgKsHsm2hoohsCHZ3BkGk56ahGCrrRt9fgsGSLB5PI5towNgp8FK4TIYu0HmLUVMI6KdzOLWXDbf2JOOdGFDB+PIeY5N7dxfOCneb1sup6HA1CV1R8ZX7RJ0p+Xd4Xs1usrNCH13cahANd+3WPXY2EeBRwpGEETdiJtvCqIExQdoSZ+xUuSltLyEgynK2zPbMx+mg/mdyli0oq7M4p+6qkzfydPCa91I14yUM218fFgbAM+PaYGJ6hUN1HeNHqqXfdaqVe8WadmLZksR4R8O/q422S8qgfNHouElrOpxEBB2G/vx9F3S+IimWgk/9ugClS/WsfpThi8FxEfSH5hW7iCJ/qO1q6MzPQRbphUZ7DaAZcODHfRMLHUIZmUX/riuhKWwXyh/fBWlQlO8zgN8PE0qPr/7BR47E/fxoIucfIFpDRS0YdeVhk5q/ZFYIaXyX9chT2KAdcT5G1dpilJtQuUuI4z1alAnlTictCrNBu2GUXpshQyiv5Nig06UHZ3zOKTAjClfZ/q0NMkWdAcyCTD4OW0+zVgzyY/GsZt6yy2yKbvK3Cs1iXSrTgQFfWou/QxViUI7A455H76b4BZpjw04uvQlhx3B/MQzTumA1d4oUohS9tsgyMP2CIbZmC4fynxk3qX/4tCNupfEqwOprBZETyywJ2sITZ5Nzi+fkTnMQZWktBpABgTQcNeh11ix9d6zRFiZQICyS8xw==
`pragma protect end_data_block
`pragma protect digest_block
39a966c2f2da2f7bbdcd709df033a6873ea7af51ac1dbf701f511a08e69d20bc
`pragma protect end_digest_block
`pragma protect end_protected
