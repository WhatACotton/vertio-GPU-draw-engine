`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
Lc1Ync/yKy0655vz4Gi+FE7JrxIpM4DHJ4RDLqfde5MrCM2cCThY23EhoQy1fFt0kNtPGACBtKakpyJAVsR/JhGlRvWlW9cveqtM/qPqi+3TfGiK1rWU2smPU19OA06Cr3G1xQG0PLIiMu3+TmJnlTJqhd2+WkeMk/bdi3yiewWmiFHPfzGhmiStOXP2H4sWiEJHfU6lV8Uzy5oMCMj33vfGSAfXKWL6lTkAPvhhIgheYgezh3v8WZVEdCZ8KjGZnsPeKWRGvKNeLxeRIzW4IkPhUoj0bOkQhSEdRH0ge8xA2QUycpL5VweRiT8eyVa0inwdY6yfw4OIHpM1j7nsgjVMAWDMCZ1VFEfCeFEbxOQqBJhElE6zyVHXoSk1Ced9at0RZS/2b4u77tNE2A4MmivR+08SdYrTYOyksGt6k3Guh6K1b9BUsRjr7o4Xip/ADSV16LBHaYXYFVDjlIlQGRIM4O5KveBYIWxkvvO3WhsI5RM5KXjfP9yRTSCYcT2c2QGCM6XOhIRDHtXTYgvbTOb8m5y/s8TbX54XpUqH2nCLcrIGknD5K9cva14VncY6SmZPp41X80Pq+9s4C5wpEsLtYi/7BHYP5IPhLGULQYo543uwsFHd+6BXAA6T0lVa6IvdMDtcFEsQtuPpPFMPHyNMG/u7Fx3gkGs8BckHYz7c/O3pevM3iA/qMd6XI0CA2KKFJh0aXJcB8Tuh4qELttZqyHDnciNKaoyz7tbG5YRl7+Xy9R5u2nNEOOjZVp8q8JlFH6MtB9xlAGYWcxbqrpg6WYURHNq4YlO/xq49kJ58DwW+KuFuLblm0m/L5PlSQkRrVf0BxO8q/wS1hllnwLsxNXUe46VHcwLcpkcyTRkioK85ZP4jdjIULYF5IiSSYDOvW7QqiOTDA3wjW/sBOdXdTnnPqeW62qWsLdFxu/0UKmA9z4xSm+zTk/qkoChjdq/HXqss4UENwgoYmKlxFibPrXECdYzg/DC1JWr0g5a8wbH4w0GMgWGxhwsgt9yXV8LYxJDucJ4UYdvw0+MqOqb4RFrTBFEQRbDl4RNEO6ozFC8s5czOaYofcLtC/70vOc8BGzI6T7cPzqFUuOuUTDpq8HOhDPpot9IZffwsuOLovWUyTsSes/7rEm0DrYKlNBt0i3AyfwYK8WQAL9Ejzl5BoDUDE1X4A2tCmKBPuGx70Co6JnyzwcOfE7zC0EoUGu2I5StxoRrEzUwZkGU+egb2pLQ/1uCLNMrtfZq1lO4/Tkcbp3kauZNMN75k1H3+V8XH6yVj+nyAdPkh1wR/E3h3oj7VVBUwBpoob0bYBid/XthrPHwy1VhNg/r9cjuKaps+FROUyBfgwg8h4Ji16Z3diWN9OoAl+u0vy3OZp5ktc7l80Kqe7A/VGcmbaiPYHsWsTu98zS192cq3skejCbsaz0drdr5oVJOgEw537ang213l+N/NSdwwq6pcPjsmY6T2fYrPGwFTAWceWq/ZlDkQCnoZ1ZX1MLEb2/ENaDkohC/Ca2YjQrW9XX0EMugM9rlm6GYI/rTobeaDdy5UIF1Diyqi0mJwcxLq3YWnmtiCAf2QiSPW0vJkVEP6/SP7YBC+D1XrSEXl1FTI7gW8wm2GAnNaZji8FnYnr4R47oldvCGoVG2QpukAruW/3i4Vdpde76P04Gnt9vB6VIoKlhNQKpFz+8rR3/s5ovVVvSTan7vu2xyftVa7MUs5JVt8cI2V0gSCe2hv++jtmql25VTF3svED9TQtV6oniJsnbgWM4NineqbYSGN2y1hTzXd6EQbcmqa4efDttsUc//ibA==
`pragma protect end_data_block
`pragma protect digest_block
8282e7451b07dcaaeb072e57fcb74ecdeb2c19eb8d6f38f040c5a6dad4e4fff9
`pragma protect end_digest_block
`pragma protect end_protected
