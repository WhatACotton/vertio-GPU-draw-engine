`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
U4SpM/waeaj9EahED/Ksrg/DOym2MeiQLBdmv2+nYOivGd50K4ddEJIqO8rDKBLX4sRNXsJYDc6SuZ+rcb1aG6I+6wr0ACnWHDdF5Y2xwmX/QtpVkNTzVlsE3/Rk1+c3SQDQFRkdAvWLEQy82C8qMSg8DVJfqLwFprvbVUJP9mRmknpMv3dM5Hq5Z0g6/gBKNG/UhnHa9YZELM7TaaqNn7B7irtn9MgvLx41JtpV2RHXOx0f8KvV7rmPzbWht05CiqvkSCONW5iF7V6bYP47w4DudF1HAngcZuBlbOmN4D4yG/UpveFoxpALgjjXVMmRqcZ4eGeTqqHT8xS8tNVeFxS8ZwcaAjhQlcs+mTLQ5ZSkFWs56N0mbNCstOlMWgzHyno1ofl8EW+Ig2dzFEVMmLCFVJZeyxS4aXzhqY3Bujp6JmzXf0mhq4jG9NmouoFwXRLwGl6cS0tFjFcWExxMOahmasUqmunR4ZeOuK+w6n/bwsC2Lc5U33kgQc+6LkOFk6HQ5127SdDBWt8gOcuCgXygYR9wbgKAk7wCqOmjBAW+c99vLfqDKlPqMHaIZfdzgvyGEFf52vvditFL2BPxCO7suyISqm296QYWRm28W0SIEBwXpgBX62y82WEIasQ7lTe3Nm29hCzleHZGtX5P2lRawCwe9uNG1gTm2+9S4nMEqO3sUS5EhsLVXVfJAX/xrwIYOY51EJqrqwCeLLSNUdcXiKPdsAkl+f8xUBz69+zD+vxlsWuV9BLmOwJvPo5PxJ2ubPnRlreajAegOw68VOuTMo6rS+hF2LAc7YaNTYN4nMLEnDXcZ+UmF+KGzNz3k+H+hQnhY9oAdDYZe8ds5p47O3xJKFwF+G3FQpUDPUFgcrezybuIPJMj5n6RhAt0U7/4jQ54dhvBTXjo1GDvle3Fjnr1Q2h35dDJ8rjszbnoGq3cKn/3zRtDjgQhlXU0/fY1ZBohs4NkeOdiZPm6Qlya59MPfQxnFjN2t/xVERb6Etvsti/Mogenfej8hHqSFMh1b6fMh9wIFOJc4DR22UYy7ll7EFZhtJapmDwHxG2BHaUy/gm2JEIixWqvJFnC/MAmlRpyB129zefkVNNo7uWg14pUKX1R4aG5Ip24UlJJjWZkOoa94wZ64kpmW8VeBN3W0ghwgvVQw+7QmzmI+R4IozAvtOOJ5CBydD+cGqfg9t7ONBwzDQmniWWbpYeHsv5hAnV4NlY1XPuMwoBl99yp+FW4EBIZEOjmgW/aupJGnibX6Uo7OhwNmjj7YbuS/r7tBRJ5Cy6YLAhluGxrvr6LcwuE/0oKGRvP+rZirf/j4auYlZAVhMv/MzjlNafHB+n0hNIOD3DlK4UPUT4oFcTcAUQ7nt9KEc5vkCL/bj+Jg3J4igIx1rqQQwuXkJS0+6n7NbmJGgU4O4LZmJsPghdD3+qKbH+BOzHEkiInYaA8w0214QwNLgFUElwk1EBzzc+oDBbU00OVychMFWpdLcjGpuzMiPB+A5QGdj//1yJznj2TAxFUtZ7A9+xJD7vwAwzAV7gyeKamY5YXmD5fdQvMs+mWR8yEnaiVB0ya9l10fk9pXN1oTqDvlqM9iXzpVS+xzLqDLpeKJCXwEauV1zoJI2HjVaK5UE6iZh+o094/40qXMMPtVDtGfkyWH1VH35yuheGUIxGzAu1G28snT/PMbpdPSbFw8HuQdsPL2Csd4cKPf8LpEvFvlNKqlEIlOObuilXcHfN9yw77JHzIRREs7CCaSF0hZBf2H5NX0qbhHO0C1yeDhs6jwDc8EZjiNsk4vxtbNOHBa3V0EympKiOe2nXyOonpF0Izh8u7DSGytyr9pjeoUQzK0H/Cv7uXvZ/vOFnMxvrkRk+VQvn6JIZxvsXblhm7RixMe6YrNNw9kwZAq11DcqInxVXeabkoyozNBEIcx/+Nr5OWm32fWV/O/M7H3H+MHAtJzKQgYgKTP9ukBJU2uukJ1eImPlNjjPULcg/EAmsN+GARy2kuc+BT8RwmFlbUQOEcq6VA628CrYR7uuOqIBvWkty3aQfpCGDWYdzaLP7TFYOYSXbuEbVzKt/uESmtigESbTEvIW+g66/Lcf/8mmuvMvAHjiVmlesLy4RGnNrdamaV2Par9oebO7skY7ZUTsmkYJPJJcMWNF1/gCRsPKSFq/t4ZDWhZciJOoVlpMWii/dTgxDacfhNyaBtli0ikgviqexlTQzTWdilh4s/v2yQLLXiFqee3Bh6e7Kouo+ctHVXQubQFSnFtJfFwpACCa6HwvWDLp9zlmY9/jzb4CN/bCnM12BWccNxV6/HPIrXHSCZxuG++Cu8WeqRA3mCjFJXPC0KAjGQKPle3aVWgZldumEppRB55T6DpmRam9+oV0esvblHGlTVBIBI8u5P4wqq6ki4ErUDYq6YKjqju+Ehv04PDFzl255Q/nkv4Wk9H76ugpnZJBD40XA7T5CoVY2Z8ocCZrE+pMJpthdpmv+mLvBaX2rVGddHdKAHK33DykrLGJslpH1QJ4ow8+LrOGYZwIu3+gXMHQxbYswjbGMx+5UKmI2wYyThAoTWnCQEnxYvGc077IDnVHv6M2m8hRoY9Qc0eN737SzrF9NI6liEkLN5AM1UtgQ/Tys93Y+xkEbWDl7cMKv0iX0DwKbkUUgCaaGIhPrh3kUj93qjcLxn/T6LclAZpIk7uSngbHLwyxn8yp45WQCvMpK55QanLlWknL0uJvnUfJDRFj6HtQuBUx2cOI9XRUOzEFyiL9q61Bhlk3QnhYgII0Hi2zb471kpSiVeuXzhfiBeyFUU1j+CUlfbpycIlZGExraL9ewy+D8TPOFg4SNz48LcfzmHZJX5golDO3c/maEYzGtdApC+VYRo4lPZqj2ZhCB6ymWnBuOiQZXikBpK+eGvR3yrEtS2ySZO7gxnOfz4AcAT24cfOb+3+p6PJWtw5NS27ZGurTwsaoIqKZRLwJYF3Q9CW6aom4vynYzxydxvh5S4Sd0f318zLYf1RP13jilQOzUz2RUoHSwL50aR/4AxvKFXTdlGEK8fitiTtKu8c8zgN90FbUO7fil5GDHe5f5U9DPA79rjAlxK+oGtDE4BydbBUiLNO3y9MZDh9somOQjGLU89r+MeunMwjhLui8Bxii0gBawLNcD4jS28rOK3LW5aeheHTxfKtyaMd4vP48Bz+OQdnaV02rEzykaFrz20phKoEjB6yhLtiaOLui5sCqbKNMEQAmaStQJmSW1LyEHtFEzAc7ZpkuGRn3aazmXBqEUVIBhxtAVdHCvF5NdHr0Je11RLpdQz99oMYOk4Er14UC2lywylSJsLOY9s1LRYVsFNgujInDKJ0fWK9es/gUPIsQgdW/OIglv++A0cgA034ZFf/bn0SJ1OX3xvHnmjRwyZtp63kFaQV4WL3Y3O4qV6RXxvN9ZFfT8lhdAllzQVthbO4UcmmmCFopicuPBOYDPcSMvgCSfyl+cR7OEZag/aY+aKLda+yCw=
`pragma protect end_data_block
`pragma protect digest_block
742ae127746a65fec31da464c73943113dcb42e2381469f904e243e9a2ca6515
`pragma protect end_digest_block
`pragma protect end_protected
