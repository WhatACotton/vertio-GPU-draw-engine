`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
he13dvGjpOJ9XgLaxbnfqyZ/blFTmiJBnZFth/W06diTzH2ihMewh3Zkf2Maq2sSWpBXASBc+ZnteKQWu9OpN7UIQVoWXAvIjKmJVVcXp8QmajTeu6GFsY1z504ZwgNGejLomFnxU+YUaw4J83Wdme/BQe3qA+UNU1Flqxx99mB75GE/XYvIcHTBZ467HE7wNCtwrBbcqlVbaOLELcnsh6nPQZRCutSEd0Do1dGPQPmoOVRBDE/2MOzpq5zaWYSo3nHNrwlbx7ZzyzWRW8Oj2ScAWkjg7GhHYh4p+NKbxgZTAIzBryQiVEw6F25wIDoXiBiiAAUQSaTWD/0y3djVNfUxKvN9kQW7KKfoSvum64zxx+Zy7ZYtqnUFZJBt6dDxCbFgm5XTcVe1LLwDrirRCuHBUYOHi32iAO5AZch9jK5RZTTMAA+JF1p0l8zv29dfDnvWnMgmeSaZKRCsS9PhYpm7HQM0753xe81Oxn4/nDW13CKNVzp6JK5OqhxvYInDdMHCl/2YwFQhlK5f8MlDaegK3M1ORJD8x3jx9FfPen81cdDM8+EAhr/T5H9BGfVCkLOieszvblbQgw0A8Hwbwit5yCMecAbE3YPTDPtmyHJCIBqA0O3SAC0mAL76uu1A3MI4ZY1nhrMKI7eAbvFTEtzAcc7hjF2k7gQ7O/s9pRxHECnIjd09JAz8RGL5z/sjcNlwydcU+FQI/i6VhMerjFGBumqEwl1M/9HE8HEHL0Z6r7UqvuNP78MvpqEK62IMtFPo/Q+lH9aWo8x4QUewQl9F1XTRMal9jtT2pe2kR4zMPaKpxhnJ4h9aCT0BNyG/EXaHR+kY0x8jd6FwGBLcwLp2gPzYygGrpJC6GCAPFZPnZRxEQL5bHMsu+ZYg3/Dync0xD225XZI4F4CzZGIR5wb2Q7CGXFCmZ3VdqCieP9vbVluXOcL7DBnnDqTp2YEyVl59bkI7kI0YucVYVeVQdaV1j+OZ3lv/ll9T+Glh0+z8SvyqMHGSRm1Yy6HsmPtpIdz/OAF10TskroSPK2y7R7eTwEY6jS0FQSOY9eYf1TjY2C2ty2GH5Ba5Y3Y4dJ5CvEN9PXoUfFTT6Dw/DvZB+GXF4YfAPM4tc80hpHvSoja9Dse3ELR3f/1Y7fEYwbDC97ZvSrytaj5tDZZfgZMNenphjDLNJt+Bvf7RK2mxTI9iOlDQYtoRRE+AjVko/EmFsUSR21wZ260Q5niEefpj4MA1mBsoG66gM55qArY4qnAE6z7l2AXFJwZiNe2TstoDyad2RSxkLqiDtu+ccaCrN5Dp/egSQ59Pc46fX6s1khxn8JGCIpymwGP2wzC4/rYCurU8xkE6sVMx+6Gks9XZxxZxaf3sypq2W+2gW0NEH7Ss7ZtQWMtIhgAWVkgLCtulcF1JJqOWNmlSUyK1VP2FP+kNW6FU6zmRVjFskW5hkmEl9TISb58ZZr1jGyUlWxehlvu0HX9LFrYPLJKFIOrfGWC6J/MMZOHyXER0YAtrMKqDGwOdK8F99RjZ86KXZOL/RXfkQRV9QOiaNUPE4BfM3lpFCOlgIC2/i0zuqBUklQqzqNmagnduFtbKCvWHWcyPAy/j0r/3Q75vppwPmAeh8hpD1NvO/gbT0wmly8wC0X1l7mTc5NzgJ4qYYFI6MHxjdtFCsBDbqG7jvp4a4mXpAoGW0ghIoXQCTLiYFSimA9Lp0p/YYQnOaSKrCzVXX+gMbqvBuGmBgJ2ZDzdqtTYDy10kOS+EWOXTvzpO1Ea4JhB3SBY+dccjUYdrNpjaOBcK8yZkSV4jtQYfqLMF4AASid4cne9vG9agpAVkGNL4ApKI+h3qrPeqOfdyfVAjtGoiY7yimFofdYWWkPefuFPxJt6fCst84mi9aWZF252mfo10owwfeDjyKzgLc4XFa844Xpk3yk3ZbaQtcTSX8rHXiMzLz3INtNWQe8WWOIUu6n1aDFBqbzei1eEFhUDKNUsdI3/jeOn/5Iw0kLT3uCLETa7o9Z+9b/b+82f7nB9lRYHSpZyUDILG8i9818JZSTZTK5ALaVIMJ+Pu2yw86q9rlYBb+a2ca1OKzcaYlDo3SqSCYXQXanntlzo0ZtPV+VNC8Yb0OP/FWpqq8X/VrioubKc0ro3zQyDnPDC28wnucsry37ED7s190L3nNrG4Z/VbAbqdufw9PjuhBR++6pWOh3kp0wCGNcOaQg2Hs+0pVGYccENdOtM5rHcU8hn8bij4KY3h2sP7vmX5kVhDy+jiIwXr5AWW5igyf5ZfLKujpWgt8yJiC8xl/X2GL9JyBzH1yBpk1DWi2BLgq3AT20ZHgmfoiSRpbF72i+w1q22xpnUSXCL93KCak3k95qJ6oJwVuJJz61XXYhq0/T/0o0A6rZboZaM1nz2RewdzoPDwsvOK9xEUioyrhPV+FShqgKqntqLkUXbBjY3+KwFyJjsb0I/sY1f9/YfW7NogPORL9RdwRTMR5qRsRC9FhgR4IB/AUz2zKwUSzS8Nd1vidTLp6Fgg92AnX9a0FEkBuH8h3Xf7gFfl5sVs9ObhjptiTW0DByONQUfe1owQn4Tl02w/oFehO3mB3RYPrPJvOpBiHTiTjeY1WpHO+wW0XT0kjG4CuWNVIVD469+J5o7WpN7fu1ZuUrNEOopDZCtfJLyoD/gLWMPuamzdQ0qV/m/HSUGT9PgO4OnDOI/vt/gz+84N4LWaierzjuxJfzjLKyuPJLJom7vhcNqr1+YeBNuXBBwz9UwJ7/cu3qR29ul3s1fY8/sjKjynTRS4bkbDXH6guUIDwLOBvGMvctbdaTwfJXAAJXBgntR8E4uMVVH1tr4OWgcXqfpA/VZMGtvGcFzHmcYFq557W26NGSestTEXYwsEggRssl5j/Hzb33N5M7qvfzdg32NPfVgxjB9S7ZsLgB+Gv/HSUy4Fni3wbLpEm9+VkvfbMb3GYHPom8u7GO+scrukgXatUtCWlhWKawEPYD4N9uTNJazF8WpbsGcN0Q4e+X2Re/IRqhfr/6nGXtjI/VnBk0FOKgCkH4SV4KxUr0OZsGRLlnaLQKoz6YO9slbDBhLZKd0dXOX3zCltspV0Xw3Gi8PKF4u7ScBmvrv/E/vU7a6xXMIRoOlamYaDEwG9qBoQH4lj4XFz1Staqcx6Cqdyams652aUXBf1vyGdtXppAXSn6r2WeSlspuOIPcl2KmUtXeWQzyuDUx2KjWHAojen9lu31HkM27O7JtezYB8GeonmAQ9TDDUd04de596IyRxV2hDG85WbJizEbwdJl3inQbJDREyzdRb/4V651zpreVCO6S9AKO6iE4iJBPXbaythFX+pKRZ+12yYHu58hfVo3KMfFqw5S7Oiq6B828gZxoXDULYEZPqKcAXrDcq+0RJPEyu6Zp3Bu+1vXQ4lBl1lTb1JE1QlrbZpUKke0cwH6qRPQJoSRprTHfDnZOgA3AXn7bGlfr5EeNAiz8zNtAGuXv2HcSFMUlW+vcaqiTkv21hconU0Ao5MenwYdDRACQyOUVn2ZsBIDIC6gXca8qJ+ho6yP203MNXIEmXylL/Ml22pj6R0g7llZXG1R45laqc+aLTO0A89AxMPAWGZ8a2Q14TxHzh46/aSQAztv3//C/ap6BPPoaHN67V3NYZS5fQ0WPxkhAl9uq1vn+vrYkxrGqBzu9NZLxsic20TzkKMQIjFks59TVmbhlxNovoD2uZGIQ6Y4dQuqTLjpllUXGN3C8ckrT0JZI9TngL9iEK1bW1Wz3NTZQz4bwWY8JoreL/m3OCnEDfvrprURY+M+10/Y+l/SZNoaUlZNurqjU/cfKn9Q0nGBnxhbOouFwxEi1DJS5HUkCADVUaO2vPMSQr0SumZShS3+FczvxtWHHYhoE2shalmYWSd3R4pccf9BgPDc2kjiq0bVnfxXZxAPgslKvZEOlmD7eUcitm1jsyc2Gyxpl7z5VIgwPsnOJipOMO7XTvLATkzp3T/7Z+GrCv2EdZRHL4mLP48LCq1ocUpmQlCCrnpK2JTMO1XUW2KRW2r2xu1ZbNjWppDIALszZdE1/twdk9TBygZgmuWxjQb7758eBrRICNENxHkF0klUxUYLvG721fhk8NhX5X3XOhIb1ln05KO6ahSRCJk/beKZaeNIcYnCcMh8rSpM3aIsjcFUXdANGqC1k2DXXg6G9TlUzzvrh0fA20Wvnim4lnQthGKt9k5HGooUkettVm2uAVDPD8Mb+DFU+l2KLlhC6ZdvLiYTvId8vMOC/dC4WQ88OkW4VVfin2cBgQ9Gu3gbOyvBS38iQA7nKzcsUjG8XQJABm80cKgUrsxtYlUyzQ0dDBpjC8sUiXvQUOUqfGjV6ZQIFZLHBkVvdGED3skR52f7epeaO57nvZsBseNiNPgbL90+sT9Wba7TYedlh2vRBBqf9VvRY3hzpaaRbGHwtUVlzcso10GOQnk4a/Mq+WQg9LutgxWE0IikOmmrmiGfNgmmbR1PAp5/HWC40weP6AHAIo6hYQA6kPMXRAiKddmipsCn+QzPWa7sl5viCP2jW1BWtpuS9Tb2ACei/Ru890eCf3gO4Jzj6N+SmxWaVtOr/ow7zXNT2Td4kLWCLAMgDVD3EGlxMWAwU95rc/R7Ojmg4GFa8mM65MKhN8BVh92bLtef/0mS1lihBkIDgdi71LXWjoWQiUqnq32ATAyPxEio9WKlsfx8nBo9fPtWKuiYYlNAxaI7S1aYAL7AlTKyabWSvl6i6T4ayo+ZRKIBmUG1fJaJoMX0zj3HoYp/WIqjIbGY5+V95AJ8mzObmeSBdiukgNo85bSG/GGMWFSZvpFQyZasvu0UgpklNshvzb/yLSuCLJy7+JJnT43fCSaXpTauwjszkDx6R0CEvCQul35Yv3QW73QlOP6Nbjpr2x/xtbWYCX26IaeeSV2+M6DP3WwRcHDKihVdSw/U/pB2JjaFQdkQF0XTt0W0puw1kUlzELnA92ni0fiW4ASEwtJjb8Yjjzud+GB5G204TN7K/T2jfkJfZfK418wZvJ98W16b88P67B1nd0t8KnibuGC45WC+FbztcPzX3+piYkanhjmV54mUzp/nbURM9WazcMpdHUeiYIJWI8S2Y+625lKkeEfGXSjz7BsGBUp1s36kO670Chrz734e0/QzNlk4MIa+A52Z/fvMA6N9QPawUil/d4ZTcBfKgkWaAMtjld0mDvz4lcolseMXA8jL35cplBzvTg+5AIhd5zUZe9V67GNU4GhHU7+jaYHfhJcmeH4qvWdvS9mYP16IsExhiHUt23Urf2f5Ujm1NlFhF7HaqsHUYaBsIQezTaT5NHkJIRZV1eGs39o7OcMchyy9mhYdrqARDzUDy7SeqaP42eyv/CQadHZJkYuZKegGlb06BXQ9RW38QVqEd0qMFDlkRE0c+9CyvKo0zWL+MUVbHUC/D93cKoGNZaiTxUkzTzLo3Kcqb5vUoGro357f20k8LdFBWbdyqZWkwV9va+pDb2VJYHfYOvA+YDV4EC6uo02YqpGxcwLdE2P177aHgpBgyAlAbtNr/7+l3pJowiu5/Z5PswnOilvq7Wta0n1fDxQK/ybYhMd0n6FHtrlUDmKWEPuSor2e4lgOw98sn/sCJapdC6M0pw5iGl80MLkWFTxUdiWBniZNOBT0kYEiMF8+698xptB65nPQyky2Eaz+R3riqTVHm01uAWnFBsnG2OHw314xyWLpOtRzDcxGEvE5rnk1PvbkDICuxIsS337q6dMCMd4VqWpuMvSRlyo5ppvAFiCE/TL6MhHaYrcHR0q1yqnTd3LlijmWYNLbPTjy3iCl8WDtW4RgfTSKuHfgQN1d12gaD82booBi/7pTeaCAspFDTpiOmcI3QutveH1AbOhQtBB9ZX/QFd+b7fb6Y7qBNSem+rpLyINY5A7I0CdUO7IENBHUA+ePNeGNQklsWWdYhUx4knYScYngArEtpVcGYDBxiIXbyrkz9je6UJ3l0bB3dImMBa2IABUTWW1hvM8N1qwraVoLKKsDpZa6SRRrfKbcWJo+m0lQyu8MHtZiAy+BdBcCzXcjf3X0gz2dJ3kVuPNgM1mfl97b6Qw95SFIiegfaZ+bnOKVQMilv+7oUcYo7T3zJ3rcVlyST+DAST68QgcY93BIOshXbrIF8mWosJkpWMkPmiNE/w/wn2cFumqa81O5++VMSmCTWNQpoGFOhyQVKAcRm1MRVu29Qa6KAvStVHTsua0jw6WkAaSIvtQiRnZHNYEQUm8aBrFNMcX67m6TBScThQjctjkkv/vk9H0eV9l41QTW21M5tabkArJwycl/6ZITsaPHgRSvffD6RfG2Y3hrg9WtSYTj3nBH5L9iyNwr5ckTmpUSODIX3PoXKvKiLN33lkUOzdLHbeU12R6yoAk0F3E6iRcw94cSZmZjZxI6baJ7a97lIzIg35YOKqBwjAeGMdauTeu9ZSo0RP9ZP6H+EdrjFYg6WHns2A8Tpb+42U0pROyDtlw1DofkRtIyWoxRYKqpamBX16EuYMccEt9fcwzVFcAyPwZBOtr7pP2d077PcD2aNp8xdHA8Lhtcf3P1YJExcwin+42JYP8eJ/jLxXU7c+i0VyaHMpMllyqR8Y78CL8CuJlMUjBxpfmr7jUGQcowp39tP6jGirTUQfA0HirckoK9xin+kFwnlfhH1znfuAIjmv6thnWP0o8cA3kKVb1cm1Y9BIFtLxutocyObtJsWpjXVpAdH1P2w==
`pragma protect end_data_block
`pragma protect digest_block
bcdc12a6b627fb375f7fbc0e0f9d5c032a45ab5096a5adbf89796771f535aaa6
`pragma protect end_digest_block
`pragma protect end_protected
