`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
XHKcD4cNqtpb7hmtYMnY5nrWS63kkAAzRxPqaJiDzz3iVB5CgcUFWaUuxr/550bIxTfFBCj8mXgTH7rGkuwH/n5L2mtNspFQmg1dX+ABNX7VOW/XRgGiViZvSpN3M+SmveeAGn/HHW344lLJxmUKWAfX1d93mkJVV8ZttBXJxoUfE/ORh79TztLdXhabn1tSFApNiM80DzVhEQJ5phkojLciFf+uwo6bbIZqPUeqJFSJ1+asvJjStGofb6XvdvOfDEqNXknJ7/vOXHY6bxomGVbcaeMrOO7SuzmRzKp9NEaBAyVyeU7IUcrN6dygoPTVS9T80Lv090/a4E2IeENfhf4VLSe7wO+LLt6xzEZ33RNZcFVqoNSzmOs4DD9B27nRgqUAH6qSri2PXhHopcDJEBFDvvhYX75vdLvcTTUX6pRRqXRTBM5ZwVv0OUiPNZ60LzOfm1PaWI8C6DvNEjHWShR9kIYt0XYZ+E9EiASbrCF7uTIfZTCly+CieviTnOC9k7IZ85TR77t5aMEZ3di6IOcOQYIvgoYedkeyiGUYgvQ5cirZMnL20KbCVw9BvrTJ4H+zmtFIgw2wTuEnGpk47vPUTd+eAaQ4EBOAVFhjK6xa+Bky/M0yYvV4e3CjEJw9NJzMnrG1y8nMnWmTorOpjaQTDKz233kLkeGxnu8PkXVZGcIS2CvWycQMKBecORYIGZVc8mKarj7rtc79/20kSFUGnA2+XuP1QnWkPioLDOgrkhi5gr7/KHpbaYSQD8rUSFn4pgcACd04RtMp5SHQjFUcng4VYkctaf/Z4EiTeLn+GwGiMFKu6Ch3h59q66hr9qZUYeE4VSgCgaE6cA4dYOUlBBDgZc+uvOVHgpRxTyQEP4Rz7U8Y7dH7GRi9srD/E+d6VU5X9F7Rnde9waacRR1NdLScgOMeivkjJ14bk6VKUGwqlRBIhR3lPRDXdfUtW8MnYF204a6FdpJcQw3puXfydoSEIG4Ib/qTUvayPoZfDndWnFnztR1Ql9GQph/XYvKocH32t/QZCBT9XtUkffdZsKO6W/U7HKZprlk8JAhm4HSF/TtM1/xQynrVDiGBcMj8RnzxqseggVlsJemrR25O75KgTQCye9/68LTqeKjqH0DGEiQf51Xg/a+7rcMpJTMg2ZP1ySk1j2daSyGWA9pvGv0numWzVQU87AQmlylO8iTejdAmU+QxlLpczE8FuW24/N+wrWSZuN20YIRvEG0JJw8wlbUCqIAJ77IcAf5JC3W9qzm68pRCpZvHWoHKtWBQp43VwWsBYJFnwudg17UFyHyr77WkKxIBwBLJhf2m1MxINseeWO0t+Do9go8TaNeRpXUK7f6uVa/Gralmi0BBBbLE1+xdjY6Xw5zF15x+VkYh8v7vCruR6J9FQRyx/9nZZPi441uqY2xoxma0JHgZcrgifB+1DaQ80U6jIpfxYQQi8NpRxy4708ohtnOqkkzYzNuNTr148XBxDFJkBSlrPceFvYyZQdtwZQsdrdXHQJxFQXMQls4OdYApjEBNThfif2hZ3RlJshuKsWBwQeu1nQOp/hAXtqG/VcJ4576ysaBXPMjeIhi6Kw2e2dM3uVu3f29o77y2DA4eMFCnYnt8+YldTceHbb6mXyQ+a4L+S7j+EV4bmjk6P+xNpj+i9OjhEgsc2Up0GfFO9jxqLtDIsgvjgMRDb26ATtEfL213fShmf9xC7SC8CYxDVvufA20k5jVq2PIr/slP0vVAwwpFj8Kya6Fd1HJ0KLH6HxFci0OA8EikZLIHqaC59D+h4soNqEo1+8J6MawVPXkOyKXglGg1S10gKtDe1/dNZ94xGsza7e/g3FczsodwgyK+f3d12CUvwBBt9K/yqpYfTioLlLl/uEEzL0vL/t9QK3wn0zsWbIYVOTO7GHRSny+mNyHFfCuSIHh8qyOUdCQySm9UbFNHJP/tuBtcrMDrs7d0Zy/amqRen6Qe6SpwgEzwmx6cyqANcfFW8pKhkcMKQY6lDucDOBXRvPtaYJDtTWTRaj8wC1hIZ0ODPUaFSJoMjMvtheCRXkWIeSJaBVXZhhKU2VYq/j06QS81TPhTVr4nQHnNTwmqycdoqNdFCTpOE0JdOVbfiUE0o1k/731CSs7L9yNGVoE1WET4DVBoGSVDlVGas/Huei7k2fACUs6b8Ut9JdFor55SeOedOpHeQYP5RUrmxTfjt/gaYf5YNqZZQvnVhVCk9J3XoSMIy0t+nmzxdbs9M9OyALpDmU/sHeUiGR+W0aGQ7r2YoeHYYCFGM93OOz8knsJjhjD0fO1HEZXN47wircRa9rYQ6mpFCYbQdv9Efn3ovocCbvDzvpGxefNwdiC3rkdMiNhdAeWtWFsODnkNcwl/LUS1IBjjiABf8/CWu0qDrdVuJkkKDMu8QxmZirxqJbWDpJgY96n3zj4389AQGFdBGve+Gi+wSrdSjE0GzBNjzIt5pVtofucywDDECmQEbnbjB2An3DosCYOlIA6JI72V2NTStaEcJcgeTFK83rI/rprQja8K0D5+1CQM8VGieNz61EjcCwZqe4ijt3P5goDuJ2UGxlYiHPA3Ktv68VJPerfVRa38SL00lbaP7VafqAKutDGuCCeJxfEtQ+ZvynQ6R/yJzmI/djKtGZq/ZEZasCbtB0fbE4kZMrXHM2J1erLQkncQ0f+j4SQDgbW020Ir1t6rGrqARv3TFq5B6v3/zDHyAiZaFGUfFbVNFLqDuNlyhHz1+HGtsx81yfDGViBJ5Fax7eLSPoGeT123WlJ/AH7OXgMzf1o6UPjnziTA7bH4qhAz8pL6E/scv1uBbiNDRBECNb5/Hsx5T/p00tpOeFMZhw56TNX+KrpFWrrz2DkIkAe5KD7sHI8w9xEp8vf6c2TZFIGq3YkKmrewqU6Mi2MbkAmA6LaC4vAJosnfU/BGTSFJ+c0WRYsHKqiQN8pso7S/6txGYfN+RjFaVF6w5gw5Vtzqt+iLyufPWBhn1DFu/f67bel2SjHw4KeKf2bLVc12bnPWH5DFsUNve9TjOpKm13VeLE0KtTlmawyCe3nyIg3sZlWie/G+e9SrPxzDR/C+GZxziKD/YPMpMBuizLs0/lEQ41ybSlu6jJ3Tac/xGe023pee0+RZlOKef2wf3fmYUHecIhrbzBTe1BDn9XODhMoY7HhfUEGw3VmI8RZXFk0DAOcnZAhrLJztIhHXEk8ZtdXSfE6Ruxye+bNZSojagPKrVQRH2vqHSCD6WlsBZ2nGpUTzfHAP2MAB+4vN8p36OMkmEoMfgrotB4QxMYtLxlC02/220uWXyvyQooYp+rWWSznv+1cgDDb88IxGyYuBrD0+sHgTygIm5j/hiLUShoWc8ORyALlDOlHgQ6PCEhXsGCGfS1vkcyHCVxP+ea0XsA/wZNOnAdenwuWroLpdVV6/5hnngDDx1to8MAl8FI1I1JriIe0IzLOLXnwmBe8FS6nM5I99cn3dz3irK10AbkkPrhNFP/BUY5bSL++KTyULiAwlDtK5J+qp8n0eSCuZO5UKoyueZ76z3Ry+2zuEEPdfwfUIN/PP2CcAPrHczj1+MMLoJ7zuMANJ6Ajkb/1kOSojrDO7Q6dYRpibx1lITEmnchg+TLmFaUItAEla8Buc6PilLfvt/oofdvJiaavYvGXbpEcPY7VsZN7F5lMp0skos0nD+x6hzbNiXvaONEeJLkRfJtituIWKKyYVD6mXHj07S/SVujiNpoIdAuZM/BvSOA0DwUe1hn9SZm0hCwtiqaUOQwhJnDO0hwIvzcH7AAWJu3M4wcgVjGEcc5xbnzc4HXT/5LCyGvW5Emb7kIczacZEb7zDMgSOyZpILbP4nqasHLbbHl8FXf4sMaj0SISNRJxQkW3c8pz5pTAusVkzwUhoDqcERd5xR/FKvqv5+CCJi/qxlFu2CpS24i2u4l4MwUS2MIYxOBrMq3olaJGCpPPnVwIWRl6Yth4Six5vW4dk93ffnxnM+rl1XJ7suZuwOfW8RiEa3TVUI40uwrcnoeviilQ9e6VJJqOSky6CLhUP8ZeyMCbBGgdWwPx0MgSnIQshnCh80xpLYtO3rIETgeQcMoRXZwvSCrTxNir2Yt0IQiQdKIPmRjPz5xPlZPxL24cIApx+fwFtVh78jxRRn4TRwInwxm0H5j5fLoDF1r5oEdpEmvyKCBRr6hzKBwYVngWduKKT1C0plqAo+Adl//LkeOhLHhfbMEv+qSJn8yeqnnMJPCRPfPXeaDch5LRmamJ2Gh/4CUZ1qyrYXpxda6vLHmnvE+WmbN8Gf3DLAvLRYXkGYno9BtjrdBt/fUx1/wlcU/pVw8UhpNwUNb9Xol9Z+YKOGdlSjP+SdVhEZixWdfoKnmlmCwYa4Jp6vbHiLpeHKGT2+oFIFno7matslBUPBLG1lOnpOkq26n0tENnyuvOM+fIF+2guvMti/w8LRCobkxtdW8m05ZGpk9Y2oS2Rexxg8Abp/2Yafj6RfMPnLtS0JW89HgyIqeREsDaGX8ygeTwdluL38elw04qW69AtKCVigl9EPwMANi5IzwuioQPly5XqdKY0Bf2VUgUtg7gwZLd1fg9QbaKIdxX+iY1k3D5TF0Z8N8rDwe6eF2coaUYfpLDnGAIFfCQ2VtxzblP6P5VqfTZHETI7AOijWnyaVZXtmhImpYjD4RtUjTB0x4qdQQr/4zwQWMJbJ4GCwo9tbgI9XYCtryeAfM4fcTJymQfljOoL/2j7xAUKzrf4fvcNuN6bo2xYwVcnce7t+G8L5Vq2SrK+UakC8+Tsjva2rfQYTPQ9LjPpFNn1qjumUNGKwRzu814WMg/mZ81Aet1H8UdiRAhFIhONpcuhB9oSDHHp7fc87sRybDY6vg++WDpgYHYR+7qT+nCDs9KlLeRZIYYR0kgp3YmiYQWSZGxMK4jLp3JmOd8iRd8AshhfOWguYocXKIKhZUfNU8ajc7lpOY21WJVokGz+88mw7mFyBTK/IasfLtLdvDXfRoNo8MpB/kTfhfc+ep6hWDt+4JLFcWXaCQTqnWmjeKHXNHmCzmTV+xbv2Zw80rKH+WQs806F5JK9gtVf5F5pn74DV11lLuyHrer95YYsuvq327ge+9Dpq24Q+8z5bK3roblURAGH2fJp6egwRr1EIeGxTWEjf7BQm6ImDy56/gV/qXK3CZtSqIx1jgAhae77pB8I7wHz9WLTZlUg+igd3A9PpbIhFSU/1b/2xfL0Gww1hd72H3WYj+nQeqSWwoJwPEBWXyySD7EyMldIO2s9VlfB/XkNUYIfdXAoCjX92UhS3c2VSpM6VrTTgDOwKNIP2TFzVvDR1R+HrHzIv2BZWzJGCicR3htDV1T7mDKW4JaStVthjb6NE9GkEp1+LQ4xOoym0MgrlQxoOP1AVLLc7qz37/WJEgKFGc9idFCjYz7oS3ylzycLqUs5FP/RfCn+K/pDHZD6Jy+5rICk2iV7XHAQFZq+D/kS+GLulXX/GiZaAo38Bc9FXYf1eWkMx6jqLQrQcNDXIdNWcGxFrmRYq4Rq6hoLN/l2vZqCTcCy4NpYO2U//5oR6YpHtkcWufC6Y8VQ6VFF0sfw7PN+PClDakpkEN+1wKztCJKajlnyZZdCW5TQSuPEAT4GfPZyBQEwZ2f665DetAcGneo8kSNvdoHHcVT4gnVxb4Zp9XZIiQosrX2agzlVEF3Tf22tY7DRqFX7SdapR7qu73wSZB0N8/1yaxEJaf3C0Cd2NM2AW0nlHQQsKDSIHA0xqPJmZdTqkfIPL6/nTNRpO7rh+AZAC/YEgNNIQofwfrXqEXzWdTpH5FuF3i6UWKaZsP/BBRTMQ/3DOw0DZw8LooRRnFAlgg0XJGj6cdHl849Q/PFvJ4Dw8f3fUt9aNbMltResTiQkcOEwK291aiNx3cNapJuqyp9ViLczAK4dAf5N5MNrtzpOqme0Stz+NZkDg6y8x0rCUu8KfsQQK3zsjKFNnaMatwYizA2FAi2kQ2zmLXb8mvnpCVIhRvdd7BGXLTDYb9T2yzfrdcFicL60Mpc25Jr2GFzL10LLNmAX3IMoLEyDALGQEMqwcmgDT54sCKxfPPY94gbnof1mX4IaMACr3ldqHLzHo22lmfev4/z5qt9SqKf+seLs8RumiZuNzXqUVViJd9qz6OHVjXyPiNb+uZjiXHpwbwn43MR12ecvJVPVIqk6tA1j3NjE/Xirxe2E+PN1jwaYKuEozpf5BApy7OuNpmP98Oqt6XNa3jIqTkD03o3LN4nz9fg/W0CV5zn1Q6NcmKHJdSLe3ezjL/NR0HyYklx+NKG1Iu1OJ5Ne97t6zBwza+qtqvO0/s8RjQt0G9RlbOY74/C7mlMcuJUjfxksB2nleXh7LzkYD/Z+1PTCZAIzmHqad0seVyZjsxpdficDxdVxDpZFajCjR9Tx7DikFeXW1G3ml5CmKNqPiYf/3hddFSsXZE38AkNreRQLdbcvjhFH16Fgb9pMo45ABmvEfPyIzfq8uGzIeunm9wYpY0RDsP2W67w07s0FhH3zWpuektsxscU0kTrN1KWGisLE7FDtLQ5b0bY8ezOWHWYJyOWJZ0NHr9Hy2VPXwkTbxJlA5QJAwZAzDn7Fxm80smPpX2yE+cHG+Yehsqlwa44q2coqU9WNUuRMxnWY6zhwkOsmacJLwiA0eNKPOYT7L7kb6qJlH4ZGAXpL9LAGze4EmTwu5LMnDDpRzwnnIq/kp7GtuiE1zi2MG0XICb5AI2cRzHAMM1A8Dlj1CklMSxPAkVcyZSouxa0JhvdBbV/i76pGGNSb9htLEwB9rdf8kanPW5GWoR5khL1md+urfnaoJ8ZK/aE7YB4aeWwW+jgPq5Jc96JQ0a2f5mRHq89ZiW9bbA5Gsux5lJNNTNapIdVJDL5naNYKxgGtm9uheKf0BnXR6a7juQ5q/YDD0CWoyR5ruTPzGNYH23/oUREdDc+FzFj3wUi5kjrBDyZAQgsvoIqRgvdqxinJmaZRKU+TKvmpLeQG4exuyhQg8MlRRLhMffimVTcw0SEryyZ+0FWj5Bya9gkXJ8XE1OO9v/svDPDis6iCqjENHNs/T4KoraFA13047bt3y/ecxgiFBEmZwco0Vj4AG6nr1Bl2zIbwzQZd9G/qXvmCzWuECUgLy+lLpNpt+fe0BWlgfzlT9w9NRipOrSiXsy084Kx7CRt0Rs2QCQsOUVv0pTMKvvWo4FoJ9sgPNt1tcD2EE4HjM1GonCi141EFXl2tuU1b6C1u2FlSRhi45SAmgxrK7JyjGg4qyFdKP5IN2PuGxkgRBC8/RVtWXpzDutUOO0fAZjvzzFfZiW6/f/OzBXOqb+3LlrTygcR/j9HpmbskODP7hw9Y/WSxZC8de4d4YcIQTnTa8JA3m+gubooK0Jq42PsX+V9qOSCYYBF/KP8nX+YCDcT4S75I6kSX14wE1j9DwbyAT1rBKi9ibnDrOHTbIzKkH0soufC3lmrnwLOE1i/0l17it1XSmN/5j8el7uoNXcVtbLeSXe65DizS/ZQQCr9P7kszRrskjma5wrixLiRF/+bR9N8acqW4eFvqHkIXF3shes++UIVYHK/SWn8X7c03cyB9cZpu487uBAESIB6hczq2KSOGavH6ohWw2J837zdY6NfUuyF+VA4kbli8V56ZsQhDazLm4wAhjbBEVccVR0FBIW4pXrhoOA5MOToumMtsw4YkpJmSKGUdhpi1K/Og8kGJEwC4aoQAvJ/HBNJUdvIDsmzMbb5g4ucQpWq9qwKhVhErRCGT+leFM2sf99f9vSXXVJGaH9JmSY3l4NgfjwtZrGzE1/1gIkCmfBMgndrRZQ6h13v63qeE7wFihn+YvSQFt3T0uFgQnqjAgOhycOuBRzlV9FWwTL7dxQOaMVR36N5f+mFQ06pqWlsTyTXvot5/Y2d3h95JI4EV8GAWkp0XlAPq4QCHDhgdmrcq3B0eAI3Drw3uPC2WvBQDRsTvNaK46BmvgATaX2JvdnKINl88XrxUjFo9JA5b8AcAxpWsVL7Dk/hcldsMXsaaMm1KgsFDZgKOxelskZFRXD4d6OtRixmZriiZAWCtMUkl+tHEOp0x0WTtwHhapPtSlkyBpH0hF76BPDepI0oUQwDvlo1YZbUA9W3KpZQXmJXCHkzB24GXdtATMSDWFiqZBIiSt7l9plExBvn0TvnFt9+86d4g/swBf4jAi1IIQ84vt9i9iZ1rd8lSLms8RIrD33mbJmtLBSCe/G5L1fJMAGDS5BA9DqJ11apOHv1IsZoL5ytONIsVaBRMcIBCn5NA6bMG2SYfgy513Y0iFcJj51o/ee8DzyzginSJKVygDuU1FMnSfpsSOP13A5yFCvIj2A1/UZ9AIyZq2ujUZKZiWLUaNMTKtaJbCda64gkIUHxcGIQdftPIQEr0hQBWpSVIoxnJBc9NRTWjHHDtEijKUdP2v/+n496FIY70BYoLikEjcOhd4qYIyjffmrsTOakZKmjtHu7ngbjFY1eBH5VFuXcXy782aLWCgqcevN7c4RRXGE56TXk1cEi8dACDXhXw4w/n0LgoYx+n5PaYAfvtN9RT1U+i/9iLf+Wh2nPHOwa7WdaIwslzfwaGbAwG+JCInCkjF24sPzMJO8I/xhwLB8tSZ8W0OrdLibrkNXRJ693QxGNoDZnVLKMQdBx88+RCmQsZZSJTYHUZH+LCHTgBdw7pp/IklAb33eNhR3eWEg+c5xwy10FsN7lenIKgBWAjRMJmdOyfGO0ZGvSzmHlLCzyKJ3CLBzIsfQgB6Bva3qpkRqmYBmfRKLyAW8VxwraApjmCUFvysUe8G6KMdT7a8Sf24AfC3wWiZj6XFj2HRE3bt1ha2BP7EI+rk3ArE/MZotvCxH5wXYKomXbLAcdJOYgEgpFXm3+paUp2vPoiCTRnjUQzTneLZoxcPV8SFu5YKCZTIoarIqiqzIUADoy1P6Tk4MKAmIjmdAtYvgvoP2GBzJ+5SMtb7tzIf12H1vyryKervu+Kz9D3lZlhikaVm6VZ/MK8nh8Jcs6v0hkKKByXzmuQGmOe00Lu+JHGf36ahwUTHJfpB2u+wSvEENIrMpMsGuVsCE55ah6ogfcC7cY6p48mjQTLGkhkmaISIBta6C49U6PRRxN7TesJraL+C92hGJKndV1/Ia7hoMFM7ESnyYtKN4c80V+EQhqCJ6QXg9PE95twtekSfsMEy58fkJjtAV/a82XECh3Rw7wz2tDYbcuZuPU9Nr4ycAzdvnIeI8dWC/mQQnGTF2wZvnYYBK/AQFCGaGVbdkxNAjFwa3+7/zRltiquSa9OQRsp+DjbV+rRwW8icTSPKO+iR2T79dplHZhzMzyoqz3CTKHAOmJwOGAbcyT+56abtjnATbQ+MzBE3p3KofNW28Xh9jkXeglDcrK7g8/fE3LNcp9h8y86kw/SjRtsVJQ2XZuAnD2BmplSBEn3FUTwKgQBBvStmEFY9bET8G5U+yIwpx/Q5tY/Rca0xKZU6KsbJBiCNyFGeF1+VzDrIZGeyqLI9FAvt2FnpS7iJYL1JCEqQEENxUzQgwlZBUcMWAWU6ftDYIizlxv2OvVui45vojTzkQpND9kfDs3YVLqAUulTKkG1CKFWIBvZN4Uo+VPRAYqx3Qz/kmTinjFFVykrKusf+lOaVUrMDkr4dLcRis50CuxvYt5EMF+1SjbrVxxUJ4pu5rgJMXOP47LTpdWej1Ljg9tSNesIQsTFBiQr196RsXVASCvu+KS91Xrtr7zrvVBgFxSz/VGRlKalq6I1vUjCar2QmkFdaRsw08rkeVCckZrGZC3GnKxF75jEhphkIyxWVYN6/bcyhR6aTo/PLe55R7CcCqmxdf541dHWtzrpZRCOAInjmw6EBChldaPhXYNkozw3ktCM6k4JpNMBhXL5KLY4eZ0By1OBFT2iYyHfgjrdqOFQVMpmd4uqECJitGs5TOLp9DznjkAIHSdy6CH+XDNnDgJm4K+ypeBqAg5tMLS0D0fD0byaJyu1MVv8hGHupLad+OA8GcGJqYTjwo4BOUbTxN3BdSyYe3SGl4FLWcCU+l2/qUDsOTOWwwuZxziP5qzopFDZ2bq6RsVvtX7u5HOsl6g89tEvHqwS2Kofip1FS+bGzfojArom5l5zV0ekXMc0rIIW+Iqx5P3DtgWSSV9mk59BAsUERi+RgNy95kgyqPaRHSYI4jHJOzvPHKs1fKxcf7CGNZ3HPooQ91pSIWjhsT5U9jdDRMo8h1bETJ3/O0Rs5hZp0I8ovr0sOqYfug06pNt7kfJFzdR5dMXYJZq/0G2n/SdybpgM3CX+cZErrdKbXF2+AJc9LnwYBco4m8HnZLxFc4EoT8qC7UsizvQq8tsQMSuKP3mOLc8fkC4G8XErC2qH4U9UJ2Tu6DxPZk1wyUB7/EMPVfAekI5k0FQDjbarAlgnEvIb/4eY/b2omhQuIKaAgtMf2OyffRI1LRQF+gj10KyyD5HlplLWb1L31/Yx9XcghJ4r5m5qgAd+uCsXrlQK2RGZ8HGVspZOhKnzlcsWPU2qRLIG4X2W9ju0jV14SdcM1RZbZmXMVS4fuu6zaR9KFDDKR1WGC+dF9Ztw8YbhEgOfGMVHMN460mXopHtDBP/jcMVZof0dQoyLCoAaLCf+NVLqoy10DLWFz32zwPGJKgjZPfJwAG/rzkVSvFEHy91/04gS5qugD/RHNnRCqsx5/LiKjXiIsD/KL0SoG0xny+d3KJdgoykulb/SrDcrPKhqkStgb4nepcq8aLyiPghXd0Ww06FBQKsCNjeqf+VZq0BOtENkZvwxH9oA0eNYipeac4hVOyELBuPOab3MHWAPYarQRUhk1B51Gyo+ekKIyg1I1OGEtQbXzGas2H1kP8sVdSQANUCVCu1y8So2A6X1w95ygIqK1ULTIdgOTMANoFt8qD6GNMIuCT81ZNgjIfh8oFUvwJwyZ2P4kZf1JEaZFOdcckQRQuKna1lML8HalX9byKRr8zli8DyBrREcBBTltFLg3mXXzBh3QRzmbq8Nk3QujlMEnMx1E0gKI9tPJWKiMaBflA4wIO397nzp+FEnYb78tHfOo79vncNMXEH/Zd5IvlruQ8oSnJO4wjtmQZOOqYRgImw9mDsZhgtqkMyAB3Z8AWYq14/BA5wNa1Z4lbDvwBvPez8hTfE1Eou+bPLEMAd0lg2whARBf4cg+uyDpEgAAAH5pvlj1PaaPaf3/uDiRYgZI+YKlLmqoNJvLHb0J3z+ZFT0hcPn2SLc3j3RHUhT+MH1jSY1/F4Q1qvoV6lfxHDrz+XudwY2pc1kInS6c3PLHakXDRRiU7Gf5oRX0TKZXHym3JdnBrvR23820AoD1lUuZICvMEFNZd/JD4RdXk8G9t5l/MrDVLRtp/rGV+d99Q3yXXcrpjHdjHuDft/5ViTjem60bcgLzWIk8AGNnOPw6Ww5ShVbjSEopvfqmcKswGjuBeqxEYHMuUEWINWmDRBuTVDVJGgFpuxP5aLagITpyekY/YOzW0CTQALsXw4Sdf8Wr1KS6cdSZVAIPrdF/uipXE9yJIUUGVct8Ve6bmSpRnOGfQFt0LHRLW5MaiYt0K1Bh1KsM9HbkbICigSDe9qMhR3ETNufTNPUCcy1rs3vvRs9eqUg26vJIpiWBNBXFgt/dWajGf3pfzqLvUqY8cXJiz1oZQs4k/h4dVKVsmIqybGw8ofjrs4mxICr7dLztRcj0mqOFBF5v33Fb881tuYFSKs2dhjw2rh1yFBp5sqGiSzwWbZ5sYAwZmfBIt58MqQNJgy6lB2DUN+KlrNNUCpahX7BtiSF+9toTf8I3CLEkv0OIYn8lQXtHfleT6yn3HyyFHx9V0uzuRYGA1Ci74Te3K60tBLJx/ypIOlgy8hm1QMidzi6phSnP4j8/ACHzLfSFn76+yUYZwqqMo2yt3GJWR922TyOzEocY8+361fPRyqH4Txu8SgVhey74mMtrVtiTrxJl82jg1fUK+02iTccX+MFl+3ZrU4eBj9GIjLvzay1P9ksdzUlxu+IDenBr70gBGgDgIHGOtHbCkpLHUjxWqr+fuNit15FjTR4fNpcZ9cEFd/4itVB1rjR47MNytZRJqzKFxGXNeZ+se+nTR44QhH7bv6MdpaJRXyteWsqijvEBTF/nc/lP8VvAtZVoC+uUYG4MTJ/Zafs4UypXW0NUWkjNSytMVJi0Cj74GvJQAL72ZKgTs8CT7h1PF4G1mdWdKBswVrZxjM6ie12+eu356F0Wv2SCDxDMjVjWP3rrUrMDSq7G/EnKzvKKt1ktgPXTWxkDqJHP0TOh7XeF09ipkStrxe4CANxyMd/IRu1GLhv0zkVZw0gkt9JRs915rUsJmHGA6yJqtrGJu70fqUzsWiBEwHNJ0q6jnF+n3wr4nw7oXQwY7gPQ5hT0FdSyLxEOngIPnVIFrjfi3yw7oSDA6dw178BlyVJLKffXN/IYr5c55tcPnv7/BIncHZ4Agw1tcKpEa5+jp1PYREBtYWGWSoAwDdBLx0n1QmuBcQabx2IULXDG3TC0HBPjoaBkVwkBJgakO5FQ5XJClBuJaEJ3HrFQfOXQ8m4I51vBEA13AQujzpY/XUTjVYG3dradX72SU/gQsAQJrULtYRmRYNPLgBhgYNCY3fyUQFQdhyi2EiNhxhabBOCRkwdj/q88TKqwmueJmQ80GY4Z6HrBsRUhPlySKFvZXEOcLI+comfiy6zzygaLjwQz0ps1FhAFJhYqQSnYVrcH05PZ51V5eKKQauC/S96bzOjD0O5seGZvEt3++1ysEd4hfMHDo1/aZQ74+CaYEEQR7vlwquYng571S6ahwhBK2CC5tiDCSGxvDa9kkYBmVV+8ccPAl6kkUD/OZhnDB9dAEjPFXI2LaLEho7bvoPm8/S2EWYR/7+HT3Mrw8Sc6mkabMJkp838Y3JLV4IzGUSVzYTh2mmFMrNY1O9bzjHdHH2I15iqCIfIQrQIrShT5D8QOWW0qequWUlURyAO7PCfk+CMUcCm1Nok43h3496VWK0gKKiNhs+Y+ynWTWLVG1UrY1j0G4bXLvYFs9IZvvU71UnJO8aDhxf4tQH6dJuyy4tfNfLTCqlTJfg6df/zsHmn0TMqnxBp/rY3hrM5zRtixFJBk8pVQRiRWv57+Skqpp9sJqQB8rdBQyZhowBbxWM3XUccwd48TG7jHbhWTDLg4SkIN4+kpZ87kf4D+t6+FhHQlCE3HyZSWzhNKzCDhO1RgC4kIXB61gWhktxul39D3a0u48SIq3wq7kBwldBb6EuZwhia1y0+evvNU9PKFsd2QyzyhAhcUvsOe4/A2zaBnu3KFVbe6fuFrLCLzIxtOd/d/R1evYwgzut5VOqlAIio4R+OsuZCcNYkVwybTbn+h+DqkREfMS4MUzq0eOAaDsQn8uCCMTz0DkYnzQoUNQWIbTa+W4lYHa3Ag81/cC0OC2F5SgBMKjGA/yPd2nNumk8Nm/nobFsHunNtupcwjx515Vezi0uMdH5icHae2J2APqFcg39vs3f60QN8rdRFozOlOQ/brPTMvpI/6znb0yJScSL7xPI/4Kz4rWjf7PbnbtMX04xtLkuB1pulZGAJ4kGCjYlDVOoO/GPmXLYxmeyv63AtZ+2Y8OLm62CJHtj9SidtJ/2tbZlX1ghq0ghKer60I98VhK/jLYovGVlr/1GMDXdMkelaijk8KlDX36tGy0gTx/Xf6qE35/Ng+tlYLXSucIxBO7SsJMxm3EsXlI/VzfIi55kkNYbTt4iOMNN6HAKtQ6RtDk+QAsoxrZBT+h34PicMLTGB4TQRd+HYfUdZVZovpP1KL9vJafRGwC/N/J9zAX0peNuVTLlWKORZ0JGXVVJ1YGdbTFFiIlu2SJ72OxZYvCINxZrYnP/5sswglX3DiTE64Fo1rGLj5IlXrky4acM2qnzY74spYOLEpLYSuYqZl9Vz9rhOmRSx4Ue4tI30VVKf7N6lHEmaacBjYhXxdge5UupJV9es6Qwkz4ktR8sIby/x+xXf0U2qmqvIVKEh0iVEV1N3VWXZPtIS5GHlkP5NGNHUuEiazZ3kz/hQLK0j+Cuz4qqqr/7BMiXhqKwZ2wNWntXOsOsKA30ejJz8BXI86annhvhUQyyD79DWGA5R6JIGwiJWev8bRtlFykyuJ/7/RCyMAuZIaDFoc8+lofAMmDmd2XkqLDZ2wZpzovE2nVUFUv/7MqPcTX1TN3BcXVoeUMAy/zZUb00AyHHR8In22C4cdwurcIMNUUOWyfCkpHjNqVnyTu4Q9w7/Lqo0Mvh6yy1haMeT/3AXoS/9hvXf8rSva1XMDD6p6/hOT89IQSL6eOYrQ9ghmxIGbEVbb/lM4iAHM1H8B6Puz0C+zJqec9VRHj/U8sxjHZbAMI9Xfk2QVBfYuOJk0HwdSPYx1fEnXPb+ViwdVI+U9/t5IlrAuxY270vlUVo9Mwdi9RkYFCNFt5pEUsYVxLHI5NypI+Z6xPHmVpLO2lq59hQKpwmnKaJLfavL+APrgxB4QRy4gOX1LYQG0AFCCZonrbW4HsgSKXZ+ohHugvmPtrjUvXttloL6uhc4XZ/3Pa5Vlhr/afMLdWlmCmDJuqsHJLkuO5vnPeVpI3IU072P5e9a7/6DQzoBicFaZB/2Lzf8luSALrjt4OQKBwNAawH1TF0e6wY5ZgdNDFI+8zeN1xsU82HJ45wKGnV8q5KP7ZP3x9euUr3MwJvOlPRjp5hMy0uAQ5Zz2XjIUViZz8bwX9ifJloCPo1rwTQ4xCmqRXboJHO6iHPti2Fm8eNxv0zL28JVPVUPVqmKd5XayyCqJpYkzcbS7Jj5XaW24cCE60kWuPcKlB5gIdP4GQRVZA6z3t7p6JrDPv6YKIBMTEnoJ+3NMyUQZO+RN3q+umzNfxh7Ox7YITAI14Xsaaw85iXXvVyC5nf9SAzGDaCK6Bdyhne5RAlX4vRqWsjn+Tf4ZzLv0AsZN4IeYY9mMOZ3/n9ObnThCqjrPi6UwJrsnD6JgOMEUsHYkkBlC3pzhGezYXm3hT3x1tgC1yOaYH94cmix7DyLIZOWromUXMBGIGBkjjHhbzPMySY+dFIzfBzij08kwJuMPqb/trOp9EIVDsPy4qnqSELYNSJLnZstl21vbX5UssRSltumnoFYM7NtMN0okddLL54tteMtakXbEIuw1FMuY6EkPpEeLFBhAUmmcTkljfm5O0mfYu7JIKeobMKkFdVKGNRVYtfuUWChD6R/CDYwlBPcnxuRqtVp3Cpl79KMZfty4ZY7tC5kmJVEdtwffQmOw/1BEp6IpgooOiIO/H0XszMCDRa14uANzdWLJRRhZ+TO96pAKZkkyQq1rP3tRgsz9a7rScAoi5kBec/eZ7nAqnxE/Jlc8ALfKgN5Dc2iEFA0wpm+Cazsnp3G4z2CQ1MyEavHe7RYBE/JFdFhWea6mAuc747gxcK0eu3LOK6c1ZbmtSFG0qbnt/oyOMW1dps/gjykfpPD69ux5/4bZ2TVQn5TSFo+aSgKwEmGvCb17EaEPMrB6KDUGLMkQWnb58YfrE6SIdZntwzANRGNl4ia9yFAUtIn3LnECLNTghoTjLFxHA31yMoBrogolD3Id8ZrxmhRzBIf/JDtDTDGzFRmKaAH179fpt+rRWtB8miYjV6EQS6r2Jq/2ijYRZ/W9ADVL7P3Acn8L7oZEPZAZW+cP7ndmNx8ZprPfGX+s9Dq4D5BLBsd9ruu/gMymEpTrJJWgL/cik1V1MDyNInI7Zb8/onBCzqebzn6PCqB2SpFHrT061VVRoIWj4BictqcO3fiXJ0t83zMpDQcws9dcALFkO9vVnToLd4hVaoPBtXvDtQrnlBz6pM2p7zVn2EHtw3Nb4scgUqFIYvU+b9jrmNYoONyzsmH880=
`pragma protect end_data_block
`pragma protect digest_block
a72f0eb363e36de06f8724b357e731a66b1d63ffd8d18db203f61af81fa315df
`pragma protect end_digest_block
`pragma protect end_protected
