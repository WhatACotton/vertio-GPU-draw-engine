`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
lsJSOLRoJRj/k/PhMgfsfmHPuFX1/zrJizox4HGSA0mABLTI26D2lyS1r3JFyYKxrlAfd+MW3e6uob0v7kKT+NP311A/vm4+o1fdNwcNHiW5SRZ23vG2GDK4+Dtw4UtnVWf0x9nyCPsmzfJIpufEQtIwYXqf5+ePb3/pkwkLFzyU48EXXPIsguTCEkGPKGxDLOu6JlZCKzsEW1BBt0eumHnTfmIi7fRqKldqcppvpbKPge9Q+ZoftXjPtOvptizYR7loeNjZMwiHbDWzGebXtgGEYm1ODTPDl5jLv5E4uGH2Rjk+Cg0+doX/VDG+dYLTJEBAx8MTe4opUhikyS2ikrp9SeDZQmZ/WYR0Kk3cyQwGXYwbE84xJfhPEvya/BOe7opeZ8j0ooTYiD3Tu6brOIlgcDBesbsrYVKGrDDoxf8a22fE3K5ZFMtm+RcMfldc4HIF5r+v0LxoIXevNWhz7IBGIIpvBB3509LZC64tjAxGXVmxAo2ofcj4sS8TkveApf1iLnJZQ21dHRQ3mbnQ7dx6K+Kzsx2jgYbgdyAFph2m2N6VzEA0cYeYBXk6J55xHRw7raH8ASNujtc2UG9Zg7bnXbYyKKTBdMqfMd4TiVIkCpKy/gaoPtKR7E05JUohuDo/UwyRyZmJ9CaP1XXOJuytZG1CHVnhsf5ZhGr7zXHOvnh0Us3Fh1FWo1QWId+1BOm8kyCp8n5bcddrV5ppt9VACPOBfyF8cfu3Fs+EIwB9FNGtf7qinxkieiX04nBLcT+c+XU1tOMqCPy81UXaNFwxd+yzRE1gwuZ0FyRG5gl4DCqfahpsnxNe+AxTpZUOqqZFZP2lD2AmpsEIGxbY4Zrzg0/xzBZRC0pJrYzCt5bCH4nz7ysJTVQ9r3P9fFJYFjuMcHdQzv6azmoDe9W/OM746SMFEyLxTerp/DQaEMDeZOQNWzRNWYoWSYUQXDwCkr2Fj31MqxDafNtR18OvQ1+yuf0UJPC2GUEZa+4v9flubxOzH1lETZi6f/NhAoov301ZUy/6m3PWK2clonnUvVFwcbPDqBhsV5V8Alh8MAHgegXKidbRDL2J1bZxyVqOLFPpY0SOUi1PYQYBEvRJsaEEhm8QrShDSKZzygoNd1z73wsL0is8wIA5rE/Ub7XhdfWuVkwYTIHZ9k9lI8u9fLDXB2In0F4cUwsIHca76bQ/DBmvuc0mCNYFDdKc1wGurKqrAYj45vvAUhSNZQX21Jm20SG8uyhAcQ/2NnsZAIO7mCOnesewYBhUo2xtF1kKkjtgURWKiXhEqvuPWelMA04W2B+dGNonTS8UXFrPRDmK60xBffcZfvSzpl++5l4tLGbzF0hYJQwg/3KcSFzz2DlGlMQhzgUMnjCjH0yHVGTajaPNlN2wwQpAhR21Vv2U0j9ga++QhP07xQ+grmDv7mOfQ13596hWmAfyijgImJ0UQaw25xnPCR3f+CEeCpKZpbnlGPullZq6OWPp2CGiH9rPTBITC8K5l2v/AnSlMC1NJBk1bMA/uZE4fkA9h5z+f/zeIVmSyD/FlqVQ2gxnLouRwiknE9DQb9eSZnAXTf49FkOaWR0iE4JOrcF5EPECHBabFbwxEcEsveAdKvH0SKw+bk0aIMYOSZuV03BwEkVvVpkzXYr21WCj5iP3k9ko2/8WtWmVwvIGwfCvdAjB5Rn2xBvdU576rLV9V2d+Xznti2UFZqAUvJzBaT88rYQW0mYqTamAyfhWfbblDzNemqZKpJQLA/53FCOhsIH5qSKhYXiz1i4haVy6bxxYbcv1Uh2ZGf++PBweYk28rLygqh61+Uc/4qPlrTTbsEBLBsc0A18bIl1ZYBoMNPct1EnmxyXMHq6s1z6ufiTZ3KGI2ilWMO3kKKs3s/4Et5tHrXQRXe0kXIG8xGb4gsBNz89DIqWpk7VACiigq0cU8RomnphiD/Q9uycC7hSLrwToCahss74AojLhV6AJBrz8KOCXvDwglFtTDeHd3WvhTu6HTSTvLqXFn4qK5lh+byBUKpCRW7AiaFfDYTZ5teWJxcvMEUDBb8roo6iunclgMgxKS98bzYG7XLGxfAnGi+j0pFuL0l6pN33FwkyJ+Wms6NjLJj4crOcehJiNx+y99HELXn67kEN6PcKQpBIq/aj2LF+Io46Sc+O5q4Ae4a+th19F3eTsiRRYR+Ofu2kOK3X50y2LzMZozqUz1vh5OL+dzni1/NOxKt/xxMh1Fi7VNmGhQV73JVZT5SpzqjbJyooVjWNV8FWCeGBv+sfvYsYJrLMSkGHwDLshr8ptto5unVgp6boxVKsaRZ9xjzoU3cQ1Conq/sTBrqyFgagAyk1z+o21zvj1pK091Vy68YRIkpDiFCA12KsbJl760HSFm9LwSa6rv5NGSF6XqjMPSASybA6NMohL6lbjnpG2ii3orMgDuBZLtOhHZO7akAy3BW7iELKDbpXElw61SzvceAuLgKD6Rw7jlLfAH6MnRUDYAwLk7ghHLum2eySSuXAuUq4E6t0gUqYo8MjuZ8BNCzXUPVFhI0tyW7rW4gS9BRF/T8DqmKs/Yl3mA8AFVOJC1f1/1bljBjuaaK0jKemzoiHah7ortibagj3YmT2AE+X+qOMEtwSCv+7OCqSU/rlA1Wu6oNtZMvEwSFV3fWtb1SWXpafzdQOqDqwBw1njwugQ19QFDMDfwW+XNBod3xNLnQaB0FFRsWL4nVLaZQmZEB2O3l8vBQ8Fi7YCUhJLMnhko6IvTIQImwkPi9KoZhIcp2X2CcZLtlEInt9L4XQD9B/WRd4Cx9HBZY5gQhdIWXTTTEFa72HcTz6xzKrE25X9BEqg+hWnvRoKrMfQlDukJCkdYX/uzNfVpJNeN/5HTmNA94J3kEClnG12Ee5qXSy8qTRSMd/88nK4k4UwZsPyQ/dFCUDvtTQgb82ZGYEpGW2Fy5PAgBfkw0vupQswpCBB2exOEZrTR59MNAemZg+0I4g4wLp6SB+O27mECC9fUq6mYodh3iP4IEsYTqmJzBKWZ2VTE9wsCymkRiKChma/uUJClHR67OQiN2ip1hAXeNvVJEYwudf9LPoL9RRBGXyp3Njt5LVU+Apf7ipzTOcAd08GHaKM2xJ75RPw2fmn4jF59heONb2FqBn0NEW9tEiTdQquthHy4p4Ysg7JTomy9Vg+LjIHUiHYG2kFQl2Zj4cE064wBlfBw8x6KIZGoVBs+lchUZmZSWGYELfnG9mamp2kB63YsSaPlfhN7eFnuKugNv5WhT8+/0VV55nmFtDnxfv2e/nqm3M5g8Rv3CioHpXh3x1Gk9nruB3eE77ZZexI4tYgiHHoi0Ana0rLTJji2GkGJ3ZXQV+XyOZEJ/bntrIPic3mc/36HIhK6bkbihAou4TghFkO2OC/ipsA5mUZ16FA/qWm6wVV1/NRgmpsyC9v8Zw0QcARRt1lDqC3GSFeSS7Y+orC4Xy4EjbbmSmHNRYiAsXVxPIyGrEobAw1GL/ynEOS2gCIg8PVReIyBu7yhkSntkp9T9+yDrgSDXiGi6w/o/ATxaBVVVaY3x9yoakmO7LiH7Im30lM+9tL28NOviclJJTSfMjqnvOk7kXvJK/Ovx9w6TFBTHcHvBkys+GWOGp2ACJ6nqpSfnuunZXdm7k3GRtGtO57CgC9apwYPiVKw9Yqp84hEemMTy7RtckzZsRihb79jg2izG2diPN+ZNVV9KFmpN8EOJ1iCrjQShvCbstb18AKvsxFXXgCxfWmmfkrMvxEnwSqiKeaPz9VG7LM6BCpQk+xZTrzx3bQYK7/9687ze3ebi6cGSTTZsENCGyTux9ISNru3QRWnLuXRjUM9baVwKhgrwpKC9hE5bkuaURDVbhFmZXSIn0azO0OS+vmehexwBNhwlAo0bQmsYuxMfO6uUpqtjt385HtwUFZxTS8XfKgAIjbqjPc3FTRep/v+nH/FPYdyDkTl+xqajGCvozXAs7bvhqiaClb2M9ivhZZjqxhYe/yOgIN2bTOxG33Bz1MU/L1PeufWsNSb9Cb25Xj3vTBoRm8o4iVDMc2gpc/kTHCjy0ERoXINSCibEDuEoOM988c99pPCJcSAwgTg8YKiybnPeaiGgKsaaAMj6TNAY75R15BbiySFqYCU583dfhw1nN+R3iVGQChZApMTQDC9j95G5sqv6vOhLpXPT2+qgVDlQ90nOzcCkqw9W0pQ/btrD9KBRKdMjyk9w7wZX32vn9W+XP6sSB9vXsWaKtXxMpM3tf4WW2vDBEzx9AlOwnDnLsaYHqJjZGfyI4pfCqITE5a6Sk5dC3ZLRMgkF35FBziHh9BVuWsvpqdWyVjWs62eS5301I0PAw1RHp2mnINcMAMYz2UaKgjGAY/LBzaLpQRY9LCu7RG7h8gpMFgeXonxr1PQbucg5o8j9LEHLlyuJKUHWuEOXZA4JW9OB1dr/jrvxVlObK6wfEvfXHGFZzkJNiyMnrg7zIhjV4KmDlIvtmzus9bVwRzOvSlSkHpFkM+FLtm9mUEXv5tRzreXzmkRKOkk6/46MNa8IdOFuq8+GO63UaVd/g4bdjF3gZmUMY0pD4XCHVEHfLSegQnmYMHwUBSZDZyxLCh3aEyKpx25iGJ78S6Gpb11K4hrE7zZdAevWJatwr8+bsidLJCfYv49LSgZk7RSyuehVhY6Fnt6wjQxQaDlVgemxtRp1ZjQ/sm/Ejq8ia+X/l26GcPDCd59T/Q0YuvmUfhJtpO/xwYJVwFv0O8zSKmIqdz0sW9k8EOnqzUpvNl74svb8tNlnXS9FT3rdGY18uLFLOl+VkwDQ1Lb8JUz8AD7VQR2Md+06rsKUejxtU46hrGH2Zbccw4mUwF2WbMZJrNhdPqHLDaKrwPLZbJ4Wr69beEb77Zq3mzpf1Ck4C0MN5QVaop0CqsUszWa9uQgl8musIvLx7JKDDNv7pZelb9yXMm2CG9KUlTYqJkWUUdFXAQxcfgTvwxg0rS7eQVxhkdvDhLJ9UiBH/DEnVWOu+5sE2ljewoPp3LpfYPxJE3j/gFqn/D8t/6BSoVziEOIcb+aT/Y+hdtyaYPNI6D6YskpvmyiaVuxLmFP72tjEvZzLTB0ZEun60/cWJ6q4RVK+zxxLKzwu34MfKnA3xVL+K6MRWCv1w/8XfOnFpfgX8JkvWshSEeemdmGeFkSs3bSG5A5YRh5sFhJSQB6CejzapmxwAhA96Tf9VGtBugOCfwQbaJbqkUQSb/5H8zPFgv7FUbXDtIQFVwQxKbB6oFXTvr0Wgq8trZnk58YvCZ9wLHVm9ecMEBCQH7Rvk2hXT+3axz/2nK9OV/dZaq0PfxM/GxRWBIKqhK36qQp33BeYMxWwiia2qU4X37NC/loFBoGtV9ps9Bv0FFrFD+7pKvEyqWdwG0uqUOpupCIqoGeGTNPHI+TW0e7aPeVD6i5ZX+PMA8uPuSwI6OVuUoyLt2sjAxlL62XE18D2LdA1bwnZ02ywMMTCpTt+ZrRliLUZCsedmoKd2yoIGBq8egZnU8nhqWMVi9rNhGuckFicwpS/fT85zgEEwlo3Puh3KhjFrZ6+2znF98KsAJjlHu1KQ40QIB+RP9zUwXXHgJSHP2XRnshfJEe9MBos5p5CfFHCNYR/2pCcRlIHbKX3gVRCDNSSHgPSsp4anlWfoqCUumJ/yRgxLupgoV8wn2Z67lyqFmHV0aujZVnWSQezei89lRw2Dxs+VVx96IzCa1PoRBn/ghiLzaVKnxUDmDZfBo9N7vSdDXZ6SVIw1RoAXWlZVh/4Fn4joXZ69wb37VzTJD6T2lxLY1QnJ0xLs4Ys1+N7BiKiK9kUqWCxUePf93Fp56B4JFBnUIbEaI0IpqwlbUTa7UZsRsn36fz6tGN132tQsEvA2sDeIkQWjcbOUNL+vRD2sDjjELot+Mdc8j0q5kmOQr3zbcpz/kLYkinojWOA7AwURClV88I/WGorVzd2DZGwsisxBm0tdISMQGZ+ySqdVMrAce/rW4jwI3Kl2KO7YJ67jGFzHFFeqhVtAfR6t4x5p4u77onSrFWS0CuGQFe9Uta6HZsnSeq87uHN2utGlwSrurUnxb6Fvznsgsj/6IxCcyzNMe3T4sDUzBlO6evwOImmsQzFBekxCt5IoqmPVFHEOjbLiCz39bdas7b1VKh6ZsXaKJBkhPYUOwdaCbj77I7c9bTwBa6v0MJNEw45smmNahqueY4wIbskHDzHGBhLfJsBRo5vwSRVOMrkhecRHOFMkdyTz5fnX5BgpCVXX6JO9SapkVtx9DjLj+QPZ36/IrFPDX3oTXll745ZGqHKV0ns1T5snirdQy7HtlWcol1hNeplODXhLF9zwSJ7kd/omn8sMBfHnjsVlRX9IF431BXk2LNqSoWB1aJlf0ZdByQkmaHl4xtd9QM8fOtFANgz4PokHkEa59QpJz9/nlxLoiWEGDBDyX1siAUVbDG+Eu+BeUxuFUyDuqZXZ4xxOQsO+7NWXT8BUltVEISiHISRXpvUkL5Bg54Oln0930nqhIJvmyH8QmE4nvlVIMiWy9pTiAREMu1t630ONxgjOzf3DyT8+A2wt1ArEV5nJXWBP60b2+iZ7nfCyCsRqBdGT+u79AqqRbN6u42ZPL7ri5slQ86QIV3hUBolY1GZz68/Q25sQZah95Upxt6VPjZOIqF8M4TnPPnRjuyieTSseyvaClu3f9orDiCgwHWQldX+PNe7WTVxZ32NMc39+3SsuyhF5wABnlQVngBE8KwQh/VN6blKfJ9q9j5rhwZ8XOgWafio0UE8gKbYCvRcJGnx3Swutd7WskqG0B59pSO1zz8p3G1Ox3N7cwywKdlzNjsiXWPK3VnQkSK0O6MrnrlQ/to1qAcRwiOh7ObFBAuBsRHwqTXfnbKXdcrFDmvRZGd2qrzdpF+u+LhfqiYfx18x2Xqt0tUtfW0mg9rMPWrtf8KUOyA/kS+I/2BbLumxoN1lRLw57DHNYjluBmRD+y6ppMMZp1FfB6EV0pSfrHKEnlCregK9i7VX85t5WXSEAAsryUpBDOFla6M3k30FeXZhSocrGeU8SsWsrtlZTgbgyovECMrpB496JL+JBhhNTLdFota48LMmMzg/tTc10NHZT2gZnHM+/Iutb69YarFREfS9qm541ZenD0hhQzrJRBhd44uhCsSwddRI/GdJbpA6p9A8Zk1h5SZ08FSI1sesl4mZVjC5KZ4Y4Jbdoh8B1JzWe8XhhzK/elMVfv4qWnKbvgxeoQW2cXftsqn3fHoheFdsS5Qo9CW8xCRxGt0xpfyS4j6n4V2kxORo2XCTOYzX0ITW8XxO6tfCOqP/PcIIuPyUXYnby15mk1GUe2oa/Ja7w2axMElsER5S2lN6HzetTMeJsoFo67IktOt0sSs0e2k9UrOK1ePrSS367flK6r4rHJhQZaPqTrIZ8CDxqNgM3yWLWvhbizfu+HwJolxYm06GZPpowcngK38b1FqRqZIzXEP6U8d0bMZfpCen4V+HVxIxkXiYGIYRzCKEoy2tOD/OUHaFbVIWH7tzpZPO4vk5UE6W/imFja4/CKVfUqonXjDNpMy+mCuFrqko3DtYryd1T/zVVNJk0ZFveK4l646O6MfEyhx9L7BrGJ61uy07qbKASh3wsgjAOSxN1CG6Umcamy337c7yXhsEBbdQF/SzI77ETNqEUmXDAj2q5vt5b5qFzNKJI1FBxj9jkcBgE4R/R4fyL89Z7blkGpZw26/ZJmfbPYkv+bfiEv2t4NhY+bOOG4ulFKJDQC+jRj86NcYHLv/HKHDasUS0UZem9kjBsiiL0eCNCjzxn5BmRuuagnVpFkGqkUBO2xvx6TZUSaDj1iOjNydOlSD+uRQ6DwBcLIlwxuGGNvLGsyYkmf+8sjiv49Oy7yKvRddJeGewUpvRCyyCFP/O1BYnSGMEgO07yf4ESh+wpcquBMFsEHbMxdDjJT3M22P88E4uSM9sjJxfB2s9X/USpytMJwa2fejdAyHdeGGqkp+v9YzlarSTStSVfcwiAlR6/P9d8+mQ7JztJYp+UAyza8yDPL6pNKpJzCWTvwt9sKXTtkU0cSHutB01m3W+ilujoptOz359NB4vsmWPal1uNHCvIvPVtHWjNK2+f5jGNcCLXDkjcqWGWiMFVtDjXviJjI/USO2PoIfwkyD3IylV1BuJCGi6vBPIz/hOMFuUuN93SB+Ws7BUPQrgdlj5cPa3Wuq25Gd6LCl6gQ+sINchzVaK3b9NLEFDfecx5JF4ZE/omSEHK9FddNjbRvgAp6vh1SEfG3kbFlY0qP7eg/yV/kchPSfGQ0u5OMOcBWFaKrClf75axzbgMbE1qe/P5s32GyOcsWepFNZmu/W2JkqqyWUM/0CkfqPm2ThnfB67jUQRRkmJuGtbwguGNCxPjwyT7rzeFtk39Tt+FB05qsTrZJE1fRn1Z3+3i9UuenRxT8DJ1v97X+l/uMBB9xPYdUUAPCuYQZrj6PTt2z2Xh/Pqrtcv8io0HuHkto35R5uJVMov1xBgzJJdKWTzYg0M+kRqkErkEUtTCMkmjuQr4ZG8vyRJlolyqTJfgF1XwDyhOkYovyJMbEv0TMByLj9EdIVnFgbmXOWHYsOB5a5HGuCYspYCLSdqcXlfsFLQJQwoiQlLCOJDwgCP+pFUpjWxOTr05y46WpFUd3sqFhDLW1e5AFzGE8WbXFHH4FrPYixV/OSOydU9A8bhZ35Dody9pawLU47fU50U+E26v3DpX77MqQGZ8mZ/aaP586nMjGATK9nrljoOeJYsJGEQnT5nIg4O4a6I5IVtl35TcBj2HP66A6jBzZuNk5PDinFf9TOycxQAyMYYVj9KOutEVpFyQVxXr+B5e+HpMpxBvuZLZTXOV1888sSjwARepMka16jDXIsFA+hLUTPv/1C5gw9VU0FFDzczAh4WkGzeLGAf2PxMEwj1px/b9ipRPyJOiNcamrYlLIUC9QwGjZj4JFz2gHTpS+5h0HVJ+epqB1PWabMQ5eR+TiFIetbBffFsceFynZhjdm/6Ac7XxLbplm3oFZ/ztXom8xkL+cgiGszokucdydyC8ROzRGzqqTv5Xf0XEjCcnjcRvl8fTkKFiQ0hMwgTg1DJmZpUGDwIl/q8xnk1DZRMzJbD21LaIeUZsjZd1almKYP+CCxufn6Bs9Eb3c2RHxx+G+XaVHOxK/j2sIxdylBkDD93bEOcqE3ywCZeOAzgFql42+jpixf2ohhRl4eZMlC4gtPipwu5PJxY4IrNuwPKaOSwlv4h5SQJ274sOGiH+tnR+CUXf0ihPuEl08SaPcNP3JJhO5VbR6ExkuxH0VhjWpCYO8y74py/RXom9QYdxxjADJLaGAjsOc9hpV/n5pBpUoP6D0XmL0LUePvjFBZy2NlivZVg7KZ07gahtcLyHWmgY46H3NW9oOfOnhNe3neFWSBzt8ha/0g+kO23o6J/15ojIdyPGrKOwzD3klZEKS5vJStkNFwpuMlsyMvyyNWnDMrxYuISc7z6uL8t024gCMM4/zK4RiH26io7twUm/eV2VOsCVUXpkahQ87q07HsQMgZH5BJ5IrtQ73fOUh9BJVtxJFe2U6RW30j9rLoGQd2lkmTXtOMmJUEuGw+S7QPP3KZyzApThSaNRtw+HcAOXxlnL2HGCcX7p4rTgSe/7TBkxCtTpwuDPLyoAgPMfwTtoIDWGqzhOchdmKIbkuiPqAa1x5xC+4XKhkBZInfrAOUHhkuD8SlBRdW0y2KmaXjZEQgTbY4f6l8YW529lKRoABdySN4csnqk03GjJlcjDrpS2uOrosf4F9PVaYKMUTxHX+adgUQOuSLaXU8thieLkqZ0JEjv4Yi082uoDQf3mI981XsDl9nJ2wjPC6ClILC1ZQCYDHo49lgU8AQuDVGUcmyiCWtKqyyyaS2igUKFx2vYWrarFcYnYBUZv68fIeJnLAuwO2GRhoqHyZaYnxLNB0KWd+2fKhh8iO/+qwmUByiTsT8YU4nRY2pxYyu1fad/qTtfgCs8IW1OMofeoUUuAhdX99AhzdE8UHPSOGCTEiIk6ZcjnGKqLahGP4NlfrlG2uYGyGurbMkflvn+YYZjsJeGcgtjKh9rkjcWusNBoWJ/a8TZOtG1LITi1a85rxXBX9yVuxIdMxBqDHl1NFvLPNyJ5Witp9D2utYl5Cf46VUusUZe9HxpWgO9IJPGEszNnsAoyg3LQ4c32mfRbWUP8mlsZZZxvt17hvG+3/b5aqE1ENSc6PqjfotgKKFSuMThXdK674paycR0ukUMJncZ6UyJAxeG3zmH9cCear7VWEDlcSL0OCqZ5Ml4A4YvhWjfhXdi4mARKl1lZU2y+8iTlMnitdcc+3zbCJ//TMBYnz+9U0V+xihFteYIqP6pm8y9xWQTcYyPoHMmivskprRqsONtKKJ4bhnY42pBdVwGdYopx+c+hPirehiAo3evjPLLk2HCfk+D2qR8teSk4xOV4pa++wHiG7DBsfaRbqs2FT56QDB8pLH/J39YUqHHERU/mMEWis6v5gB+yxgk83IpPrttpRNFRRdEcAhbJhv3AvA3rHUtfzi2gut5D8BsPPzVZzmLAFU4Xmh6RsjjOYwFWQYZgUfvCVLAxeSF2A5wyGChv2I4ZhM9u52fWv9zr19jtMkUOuie8G0lcaKdSL35ybmV9vHCWqbF3gc6xCOmb0vY/u4mvSEkxBbPQCXTO16NdM6ykIGl0yJvF5I66jWhaorsYvO47otQwQHmbTnTyIb/Afys7sGBVweWNKko9oDM8P7hj77kSfqys8kJbUPe/XKDbF9ABfEZIeKgnQPPz/Wkh4FYBfz2wnnP4Cp7JwJIrF7ii6rfo7q4+UjQR5hSARAVvtr5cGL8EGy/HhaX+VQubGRG4AhrlXf006V06gEWoDc/XchaM4mJzgCEmtOcZv9PQrzBgB2e82VbaeOtrntCRrC8P8toYZSheUs2i+kneo1FQMl2G0g3yCEhpn9F6pZd3q+cfqIBQVVKx4o7Di0EeIdePbAdKAXjGtx3NzBNC1Mg6BxDlL3qE+n9Rs1Ts5jABhEtNPhIFtWBNdu2IpKqmz+z4xsdBEIFKl1JD3vyebajQ96tINsxfeRLrRA9WaTtrhY2WwM003eoGXwxtZ5CuuLUr3ABeyvJBXgaf4dAPg/TytkPaHEoCEI51CyDMV7Da9cnRspe/2RPWjV12/7XJQ5hmBkltyDBMf1ooCqEgY0yxJD/3gSwP7jkSlxuTsWq+fzv1X4OyaFJ6NOLTeqpOx4Qkkc8XwHxoWOyvn8oetPqtIzR5iLdsyugpUonx+0h1aet2PNa8dGJVYyEWPMp6QJYwMSFBrelnWX85f/cvxecm3lGXMvClJ107gMT/6dBtVq3WWZXTpNe6+IO7NSNepMW8EqMfRCG5UlXuy15Ry+qwBwAYoBrQv0IcFW2hcI9VZZP2x8SUAf3Y7vrUpvK1v6PW8YO2zf0dpn+N1K35p9NUPeW7gBTQFP4IV5wKkd9kUtVgUx5jSxEqYT4Fdwt7BWw1GzzKi5ymIA2nXuqXdmeNLqAEyGaK412yjAyOFdPPmqryG5SnL3Yskn8bUuHCJ8pmYWiUMXRTFoqj9+QgMjZFwzGfuSuZkeugcYTZflHWmNSbe7gtE6UabD1WlQQq3Tc/Zf991NeaIjfGcW+WDTHXzo9aGIKWWXfShk2ddp9kmwRLL0kJHjPawByI71uxtpZmNHMwQXOWwWI1I48DJQfbsvQhgEPtsJZohKFbj1lk+w+b08mtNEIFdj4GHpSLaCl1SXCN0jn5NNz337DsdrEGHILb/Ujy/Auc=
`pragma protect end_data_block
`pragma protect digest_block
257045df45a33930a4a1e0d8430ca2e35e65ef1f106e0ff027338df0de9a3bcf
`pragma protect end_digest_block
`pragma protect end_protected
