`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
Wz4hEU2JwSULsHhth4/DdAxgoxzfQ53k300KZ5Er8YrKc7VTV4xjDtOZhtxfk+/JCbixxZ3qEyylwbN3k9/dRl2SvnNn6HwLUyx1N2XwnAYDchyWepy/F60+qmhF/h36BsrjxpaFaJ2k+NET7cSUKteoJYldDSVwhuEOD5wK+hpx2m3EoQdf0mVOLPNuF1hZYAMgAphhV6c2iKDzRFFQkmRiKoQEb/IsZxkn63EdwnBsCK/2hJETTE6cZJUX7QyjTLX+gBIl8pAjVicX6FO2mQaGcUokmHrITylGB5klvXn39ZuixS5DGv8N8Mso0YFH8dgRXho705rW+UXcf6LhG7rqls6Hj//ANUHJ57TZtSN38edyGXg+N9CAnaa/WdaI3wXD9BssDBRs2AefL+ebBUQJvwWkWtJfJWUEFDGZ0VfHBniiAU96l014jfhR0cIUamUXzwUOUek/wvWB3fVu2kSypt7tw2YD/0J21TWcmOZyQGoWfjapmCzBKSK1t0o+t0PeRR87bSc+W1S7i3HCWqs7znK7FH0jbGkfizuSqCqKdeLofk9lGSzQaCjr1aAempSGc4KWeVCDFvjLoI+U+/RSTol7Dj/2nLSUTOKMl0RqfaNxd3pYBz2Qtld7NsM7dm/yKsjqo/fbzpEQ+iRfCiPPVpTWU4EyZfCRd0CHGRvydOI9EYUBN+oF/I6wl6/DkoeQi63mC60TqWpwcZZ8oJ85/ZEn0oVosqPJcRMDv3PeJ9n28IDNKgzsyJmopwgKtMD+yJFgAAr15MZW76QRfh/IFLwZF7p8b+hL5PveFnq6rSEzt3sjAwVzXJd/R6dkQxIkq1ttZ402xhDyKdLTZloy+R0T0kjklkkwK372rIpAieiflghCkacqhZ1m3uKAkZ8mvbXC9sk+SXRNU7VzIOCUp8ctdsxGHrgZW82R2MSSfr28PYv1k55nOy1ePCi7pO3hGvKvXSijDFm68hT4n+QZfbT+x7dEF52OQfJskz2Az56BRHNqret2/0K+okMSf5RtLkHvOLlAfBoe7pyAJmUMDSKNFk1m3OeUrF+87Us4Zo/Wgz1V0a9kX/1pWYmkWTYq8F8hEFK8j4jbAHxb/n13/W5uG2Q9cAYMbmTTB4lYcXhyIc5krPhlHgSDBb51XubRn9q+GZb6Aqr5GLRrIOm41crzsVOYZEk9Yjx7qm6f1J3oTcSQY74v2lCOy0JFGmtUga9iLMJGEjljAppxyS8JvYaj3xltkl5Om/cQCKbwguwiA+ovNKbEkixLsIpVFTP2y0cAKav+PffTfVh/4tkf2iVyA3QtZf/XPTP6BbpMbRx5nVhT/tW34U8ep2hKEU7tfjYsat5/qi6ifdmKjTDHiG/u8mpxKjnt1qTWCHCg1kGfXiErJTOx6Y10CyXJin+IMI7PdNPpdEg++wbA03JryvkTCyc9d7crh5hnYfS4QfF2chCwGcJZX0BIAAyc99CMfDpA4Ugwin2fu3WAZo3vygp5loOGkxRzrRyCiVFk8dRLShO5PQyxh9UrqOiMhY6adZDNnEWa86BqROABdzTxxHoKeT4OOOY4+wxQrNMZrcs19H8s5pjp89egzffK9xyS/gfiLO+km952YKChv6ysTPMHpBz97u7e/Zg/aokLWOySg5CRsqoV6xnqKRVbEFa4P8V4iKJs3cd5tlheGu0izeT3mK+zEBg2IYZ6kXPHJRAvcgXuxLn7XYyqZU5EvGrATexI4bZZiiJrxHpnS8EYz2FAakd5/l7AUfcK6S2FiLDBjgDtVgHs6MH17juXJbv7bZv4c7Yc4iOqmL0N8oiJd4K3R0nOxhcAEL06hoL3GpVLQjbpZZRm6/PPiqesuRsWLRtDhidfPmauDamJJaPAGSyjlYBvydRWyS3RCY12HjEjDHS+La/9krCJ0qYAVh8Wx8psJSECI7Ca2TlSCjSITpMRRTjUXABU+jaaSZ+6iXP5q1x9ypieHfFvbzS09xcihSWMeiSO1e7w0yVOSGyblSy5ZxrOMDOfeKXtEVqLhffydzW4x2qHXpvGdbKeoa+UuOkcaSJi8qyKUKRw+Dd3zphjBPQyoDX3uutrH+v9UcJIVgsjX7AulIr0JhAoV194FXMY2dpi2H+kqyZMjBsFq+NLTZb9hDrSjIFw9KNuCO45O1Orzps7F/NmJT5sFkSqDDiac6c3yzgOPXwXFq7MCqH8NdyuLydM2yWtkbfnqkg74ejszfnXSOhBzb1WUIs5/XjntDZ8SAtKQ6yAkEzmqfZMd+L9oPwYhQEcxc6uCx/aOTMEISs8lfey/TZrYoZLRzQliH1bQlT4PzmovGk79+ebws0shMj0RtKwYXlFmy71fUb6YWj1Gr49irrY/VnplO7h4X0VVE/Y7UfnGayHWxXVa+hXoxpGcJYNRMZv/gnZPykK7fZ/uMZe5OAG4ZTU87j6Ha1+qusgloiENuEMrmuIgslYVR20eUwJukoK71IgU+Bl0UEdPH74a1o23l47eSkYb/m9XUynWmnzKTqVMIZc693ryHDlbXk1Ku7vtbDAt+S+MpTF6+0D/OcELDVKcl/ryJDHxU1O/plfptHLjWauL7/UhTiwEeeHlm6yFX0Va6XYr/0ddgBQODoczXIsYnmoHuOnfOT9NDhkF0n6UH2pig9svmhQwoEM1AQ+2wahZrs1zRN8P9Wk/xqywroe9w1r5gArDqMW6bwULQPVnbxNpm1WZZIYiLfA6w47tAYngSx4mdiOIlWYxaJ9or3/MY92mDtUeHcyiV3rM+A+dPNrj6Lj5dmpjAW5kXLfitdXhO3i9IuLWElPbTL1qmKi1stausRw1iPDWaL+8NwqCEU03sVhKZ1+ZzI5f1eAgSRzkJGMUKrJz68rf8zjaeNHh5+Aw1PDZOQ2r2Kf+cm/DsYYX7NpxNkog1i/dbCkBReveOZ4VZny8Fuiac9SBv4Dtn22RRF1aUg9yVEzggLFlBPCv9WEtYFBEklk5YNtqNgnrLe23Sqq6se9yM3Sasqh7wZXLfp1cWcnDtHVtrdg9oFoxqu594tJ8KJbJbOJ2YmPG5UpRp0IzEgRvYyP/Z2xnyTp/OV6cDmugBKKFqvNW7QNaraKiyOCI3D2Gt41tKEVid00B/bg0lSiDsosYabYskqsFzd3w2mdqd8lw7YJ/YBXQzky25hfwCunh1/bfV7p5Zwt4ahPqWifsQ1OL/8OWytL5yH4TkSz5HvGZ+YMWL8oDAqMcefsvgvzRweZDuDUTPCRXmiygpWlrJV1P1ub+L0xWr7HIG8Y4U6UudibFDXAKvUa/+ivn0BMRpp+Yj8nNfbpHxfuvYwhI65l71eFTcQJENoN2pMvDttnot9QemBPDzdMgDsxy/oWuzOxPU/dxqSo2gXhK0U9ERtCPLx23sOSEyN+j08kInU+QuAyImsRZUjCcbmk6c/68PMuhyuZKU1W9o9xENe+ny3+o0/BM6vzsX4QAsGKsPHmEHAp36uEuwDrsEqqLVbVp3M+/A1cyuBeSnuprlTHLY1kYC5wKmsccjkSevggunkWJKPibnfBjDL7pS8NXPme0yFHxiIyoPTplkab89nHBXKybhulwxda+EgqM5WPMk8YiB09iVdd+b56/tYkYqOHBGdhBSdcHZWP5ZrQ5UaP6PrxZrP7h2DzPmGFw1t0BzwilUK+L9CF8367ZU9ipvDAi8cSH0fr8K8pfJ5JSy8AyB6f+AMbLxal84J2Sum2f5R2ieJSywBebq5U69IZGLJ6e3UhrKHBAoBfsDb6/TWUmaqMALpVo5qbO5RwkWHsAyjrK20Vwr+pDCZbZfvyQ9WCPUgtuDlZI0RVortdLyK54jzanLKv6AmA3JIqjd/TuGsXPtTNDYl1iZJaDyFS0+09WcGcsMKfHmnHEljtCpqFXHX4PMTQCxs3nte1LNMDTUO6LAj9NHL1M0cEwJfZmR/Mv7aNDl+jK4UJ3pTx6yTIi/1Dhr+tPScHfUTIYk9xGUrEBl2UxoaMQhWBP1iG3X1CXmzyLPGnvW6TNO3iMO0uuYEyWGgIyAapuOIDFtiU2rAa02LgnrjiCowi1jFLWdLRtPc4vzX+0FIRXAIAyRgSaIu2q97CyIWI7vQWt8v0bgA6QtlK8ZXEX6W1f5FVwwvx++Dm5EWVKE/AEbSMTuPe70d7Uris/exRiUPPCppNLzcM1nw/xZolqbQaVsz3YFtzljd1Tf6BxJk+JQT4YvaXPGkXMSu6G+AjyP3tfjH3Xqy38VNmj95VSgme8RNnyUv5KS1K6TUm5WOAla9zrANBGvEwalgLgel5fYSMRTsyGFCjcUUc1ZFDAx/7JggWo3kP5FG0oWw52cmTk9bvxDbRruO3LJzEwySw7ZZ1ZhzasbwI3KFDSSTi7FidFdirtf9Q8UBRPOGSQyJzmnMcE2m4JqCp21E2Kh/jmsjWz0n17V8t5a3EfoTCDWe1W+A/mXYKXeiKl27TzPxRrKltDXnY/ndsTulWbd+VL3IxQY2puPKno4y5/VEXcpsACc/6ezIEjhVoy/sukSIivqnVaJSBXPT28qijgyCb+00vJVspKBlT4wwZ0k8DEqY6Eb5KssDN6zI7HhC93a+bsHfnE7yS2BGisK/QNfsD06Yaaba4tSBjjnYumLDHJNJ8D64P+8dp7jJidJH/16bQ7D6gZcgALv3PceDNj2DxdThz6ocQWSGD8LtvBE+5RsQfG79be4j/rIUt9zYfOfpRnu9bGgJT4gbShT0VlQg6GbGfN59Vnwcv4Rb6NaZqPNfL87e0n352u9fGOKhiEYPJqEo4xspyYoEyzXUFkaN1VK2k1sPz+gCfPcmX7pbw3CmPZykxhE5KhncJYWLy/+UytAKW1wszD7/Ma9eHFA8eHOlMZQMm5y1OBLELXBDch4hkaJ+Sm/4iCKbkR6kcLnuzyOrsVKnlHR56UTKNHYerqrugnh5Ls/TTUGlvCF1dAo1v8zl47setBYYx6C0kITfCJ6x1o/BiAJ1unxSdhUGXlvikrQ+SVhg44F43pb+aSRXLD+yZTxiceddEGCU+aB0GMxPfVeXDwRTdGbiOpZXZTAdVaE01/0Z/mmX2cSZLJf/c3dxf5iig6TSR7sfV8yXfjM64va9hd6kr0VpQpgjlrswCjI4NOQOTNLXMUCIqoRUpTx9WTMv03sQq6pr5oQSCN5DTBfpeEBBzra494rsOxY3+6nRZth7RLxwUReUqxThabmYX9CMJ0Cu8n2csqfW68MxWL2PqPOC5vY0CxuNMsQy10Qtifqg8odRZnYkdd4CfQ26V3WCsJGYNQMt9WuEePmjml3fzhHVMoloveZs9jGvvUN6PSu6xK2yxfHzs1C4bmNXmuoNSD0Q4IPWr6qvTB8d8vL/9GeLEdzzrAhm/BjgnZmS/JwcZ+xKyc0PhQlq4PBhRy+TYtOpu3J8jcUSzLqZoHG4v+ixwZsy8jkz6FzDsPsICnU+mBPLej7YrUwIgglKBGPr5vhrTK70u54qCdmQpPd/0l6gTsc3Lx4Dwm+I5hD/RbEFX4dhhtoi1vs8e1UKfiJoRRwBmIFjdFzMZZyxPafNFhH5JQjm2ojw16RJhEoW7ITLPxpSi02vdpXDhNYEEPod3/JBvaZRbJzEkoAMj44dv/CQofaquPFgiqQJb5FCgeo0XWDteScvRFwPRSV4PsmSgbCvXBUoPWe1t4thPc6jVE7QD0dOulJj7WiKGI8D3Lohr9/KP1cgDf+vKZeI96p+3urgiVWQXxueBk5lFfy0aII2U2QBzR9bVjhUJjZ6tSF5I7GbJPw+FmF+l9Lzs1EDJFUr804S31MdpB6fOwfrc0IByMysHIe40MT77OxaSJAXvipr4CW61KLemu/4CwRKLHaRDJyF7n2EHV8R/kVP3/5VrQzFLwTMJxlH2//L8fk2rKeGvK5kpV0nqjedb9zqpW/23/8gxifv/E6WZL5ZxiLIAE73uIKiAjLsKMyEjdlMZ01UlVyfPg5kt7gBMln/ru9i+tmwv8d8pg5pfiwM0EPGfE/oyy7tuKksFaXobj5FBjVNMGXqa1BWt4y8/A15v/F7iz45HX5bXVlKKd2TcgiwrUGj4Go89CzxV4l/p4+/7EKRcU8nRrnYfCoZ48CBs0Fg9/FyKfthWT7TzpgppK1FUg/7K1zC1ykHTmGNg1GEBaLwyJ097pdg4dmdnaJ96Y9ZL825yyQYuuKCZTVrqM3F6Y86Oyswr5lcGBkRiCO0zM7xm2Whf9+TuxRe7WhZwvsqKEHTRROnm5rx43Txbx08ZoTGRn6sOwBPQdy07Do4Ordl3+W0JmfGJTOCjJGhcfmlnHXMwSvzkoA93w6R3hJRImvK+bQ72SD+2XmF2WE3gHtupI2fkjDD0Lm/4622iceIkOcdt83e3VVMavtj5JQ3hxI7DtKJfRfJ9CPHmRVVYGZD5PiUFx8e+ZNawcLmXQKZmYoIjwxbOYMqk6q1FB8172I0ObCCEc1o65K8CfPiyTh1g39Y/TxShiT1C3kvpjfgoOaj36YXadz3/pafisqwX/2gQDFa0yY6IcINj9tPj4piPjdlyRcV53DLH0M7X3yhpV+KBFEWZrHC+OlEogX56pK72XY0lFkjc95m81xroDj0aAdSf4JZCiLIjR/dm7ShRqW2aktJYhoysYK+cXrqQ4jBRVTvt+lRaMG1upjyWCwfKX+VKNesnY61HCHfwkCoQIrMVDoE9+xFbvvyz4VCmUqdV2sIClG0Ao3/ODj80ASnzPyUXD9u7lDc/vsbeFgpzlz5kiZ2Kw1aAeQ+ED6AtDJKmSPQY1anpbMHkIZv6OVlu8d3UE5PkQq39Bg9eC3oYSqU920hclTv6xpK22wIPbW5II86wsvi73cbAUerLk7SZTftRnHnmk4wLWrnfDy0ZTY/vjeQI3bOa9OI2Jt4hmcHV0Ece5PGPCvCYRMsoQF4hO5jsEtaCauY1sOj/TJeQvBJuJvHUR7haJwc2w4uLg7LyNfBbwJRxZNOA5fT5emAvPydFghhvr1ugYI9B5Yx8io7c2e5VOcsllZJbloC4HJ+ACxm5EPsbvq5TV5uy4sboEl3uQZHgrMFmXZfqyqD4PX9sLa8k6+jvihPuqSkdVIP+znKFrwSfmDMLvcPF5rcsCYheQK75ouw6QXd6+/EwfB85YWhK8oMb1t+P0wQmLJqVsZoPbyObdeLoJmjl6rLk0MusrUHNoQcuIxUekdnKTApGmwK7OIxMQfqMudqQXzisL7sNOZBhHWK8ymIQglhANsGiIrtSDzTzfyPgr0aWFissLcVo4e1f9yIsiv3l0JmitKuK1bOWRNXJjU+sioUL5Su/ZWBzGB8/8EnNQelcYl/ZKARH63QsMwtaKqX+ot8iwx6+M3fsz5mAhAtmeK/CdB6mM5PtohtVF7915vtd3wKCa4Mj7Ce0DWUVZjjMRfMxZxdiXZyY/N6+JQ8sz0QyUsBMLRR4MuGJNe/+w1YP78Yj4xEy5DUWK5R0DBpIZceAFM2h7sL+vDLJGgmjl8Ir9oj2+C9MX7J6e75ULvqjbZZnnL4NbNuB2fxtFo4hVWR7yH+kgr2nHe8f8JToUxq8ENvlqwBsajaArDCBN5cYff9j6ZLzd+BWP0yJ4niTlVHDWiQsQrckfnIavDimW2E0gtqDTtIJ3u+JmBVAu5sIT93KGI0ETo9q67b2Hm3w7G8COL77jS/YIzgKZZXFsJLzu7vYDoyM4CYwn2LwnxaI48JUX8l4Lgt4s2PyswXkRs1XsWoNaTZxldJq0Zw5WpuBg+pzmSt05eke1saUpR4IcqKqtzGkSmR6j6Dmh+tw70WwxJ2LuAXI4gWvH9KAjrnHmOebewNwbn074oogxyWCHJNd0PInqhzPjv6I+QtSzrvZMxJDtcPAPdvol8bZj6YXV5LezYVBs3bRPhU8LIuK7z+fgklN001guKyPlie5el/Zehc8AusrzszVt9jiig7M0nuJ9AeXHpUhLTYp2ZeBvoYModDoNgFiFR+pQk7vazOa5uIpJgRkpEsuz8LYOo9XA33cRv7fyPkoTth++gQSXj75B65tXTFP8Eoc5JOsgHp1qingRZlQLxKhEBOGI9ikFLEdZE8F2efyU5BF8UqjRecwi7Ez/HNwH1Ezfmq1QVzF+0PKrUXqH3RzFsR3ntLyoqeBrtuXdAr/uAzsYRtI0pOwknAcvB2oZQqEJMdl3Woa5J31k6HrI1eyGwZG/JrSoJkRu4CdoiNBYPSU6s+D/bCBtEuwnt7DQ6SR+6RnebaEsfexSRokf6XRtRJQ0aDuoQGwNA4TNkzQxMX/Y68ethAYnYqdV6NZRPRkTCdm32VqtOaSRJLP2qIJcYwGetCD/gqzQFAgJVrd2CAeAnsvKncdZzp/wbSQnZXGov5NZCLiUeEXvhDgZiF+7qH4S15eTGW8QPj3FXklZx3FsjmVWLXqD0nMrHMui8Q4FbVSJJ3+HfT4bD35jEw6Q2gr4JhUnPhDChnv89lOde8FYEgFLgy9ll8JX2S3RZqIEb4OWI0F4Q5KEkvbd7oGH0sTeaHJ63/Fl8asfGNS3BJzfAsuugiWZlsFbayNLUgXcGMYTVxQ2PW6OGyhkIXVXRQGv5hyjToozaO1IDjZ9lF+wx14IKb4X0rDPUuugDyvafRRMo0vi16SV7F9pofmr2Phw8tfQBsGe4bJ/RCuZ7dPUzQHCblWyxbrWpGWSdYL4H7xVqXy798bcjCgPJwURHNfzCGGpy0e7lWNjVF2Mq6aFX1nqdtjRceq2FXHaJKsGUGBZx6iEOObBuQ8QBJGxw7soTKlPhbFhdu8O4WO1u3mQalomBnSx30bgliWHJSk24XqLLQRuNpuDvek6lq+6fC4iLCLbveRQ+xbFKCYY1Ua55f6S4HDTqQPGZ/BX0+RXkDpOYS1e2GrtmpCLSABsXdUhiMb7E5uCPdlvSzdRVSJAiwPXMQi3g/cwGK1w7f3/Vg1SWz8nro764cc7+jJQC2c2Roknpybd8AwVV9ysNfwAoPOkjmgrUtdNqK6A1HUaaai80tc5P0RdfmAm86F34AzeRrffuAhiCwwbsZ/fyopnzTOO3ncA/S7wk63+g4liA47FHO1FO0/Zco0aQWoT1GJnFUNzXVUBJK+pqXOU5+EhtyHc66MdoopE0I1NKiI6sim/sNvK2ARDNUrZzrmCkC0Hk1d38OpEtgT6dNg7VHZc4VbkA2Qo7JZ+VV3mg+/jtLWDkfHsS7m0u4g0KJ/azpZ6MTytLvCMdQKxTHAAvSvBkjeLGfTr9ajt1d3wlgLLLpgKSUGpCypsBjfwjO2oTVWGepnk4V5lvcfl+Cv7ELxKjpzgCTxgfWUOUYeBiQtJPNqZQKYKChKZ6OOb98DRinjvskcNhes+GHuuOLcu4Da+E/xCdDKtgglu5d+AgcrSJsejLMKTpijERdzX+NbrvlAW451q1eWRd1xX56wsYYgVqtqkl2Hvy/AMRYYxH+i7vGCOdOLIkuTEBuyEOrfkqpiEWOiVSzXhus1/O3unXgmnrHV1JgqSlGvd1azweHfUl6wwiYc46vcl7dGaKN1yfjEI3mnmBRZF1skbCaOduOPwtG0W6/z5glm9wSvZggy8QwFHJJwPDE1/6S/Wbou95mdpXEPVVpw8hgyNVClGplLoqCUzf1TEBWCWzPzpQCEvjf1GMgX61XR8+TZf6nTRi8+qL/JAGePlhtFmuGPpYGTwuWKRAM1D+CGzhX803/wOd8oWcPhcdl0rjXhFoU0RP8Q0O4VHmZJsAsYdiLgtSXNb1RRFxzbfhLqPUeo/HfBsTRsJRNyhECzWEgzZhWr9CO8uVY7sI8f6OaQiccgG+jPSvRxvN50AlsbYIBwbvS1k/S7t9P9OMrDbCQtwmMMvoYGYXisuj0DDwYg7P32sGYh+N4kXS3EK0bjZpuIn9pX9cImSCw0MPnPC7marz6G34bpOauVhNUH1KQaBwxaDlZxBD/vSvkiPKS4LyI31QZo8CLKfeMJ1HVFZdgoNPHZM4edwqtoQfJhRgac3C/oqS3ycWQ0+k03W7+DgHyT7nicQCTus2tuQves8gvIgR0zhNFjQLKJN6Fzw9sKQJMCgGX2WMveewtxyAB2JP4bhgobXx/avP69EH049+mmUP0SU1Z2mk6Vvoz2GqoHs+8ouHn0vd0dUAaKzSGjOLpOULC/Erm0dSQSUMfkDGa5qME48MgJvJBVoyQBvPFgCaQDxfohCuSs9LM+Zhja3OPhQA7FtNDIPsZZQN9Q3xgOCKzchjvQ/YinGRAJpfayizfMITazDSnHeRISJKBs6YEW1p1HhRKA+yjtSoFBsQFTgFsPC3mZKY9Q30vdi4EBUKerm3H8dRasQi5xgf32AEDJm1TqRtkwULpw8SGMJqPNI1oZh40rdR2IwDz+ipaoTRuJsVrpyWFNN+lLdPoueZWQnDtSQRlguvxqmk0gXjLdzdfSeh9Heu+tmazA17yEqLFw1gLRuTWMt7jhXzlw6ECC/aZ1sxp8HEE7Nt+OJ59cmrovh0wEyATGFKKN+AmPw4plktIKwBXItbyFTn7Um6Z3B4tE/NrPb8PDJgoznK1H4sw7ah71dbRbIrw93fyJaM7YhtQ7QacqIGHTCRIR7OO4gYCkJE2GG4irQd8gopR36lHBzk88xAk1cHdB4GXijGL5Ah05bGaiYlmRRYZ0v2nuY57fsYrfK+h1GHctACnNgLgoRI5ZZNDMz2GudCOjzcRuW6lb6fNrBL1Zik+S0T4zqFnx2gDYNey4Lii0Jou1DCmSYzVxGUkgQ/El6eE30XAOH5GUpeGLOkZ6/BP5m/9YFG+xWOZymX7NBG+SLbRD3V0FIOfDek9hebG17wJqwVEdPXSRJJMFRgaHj9bFuFaH3gC4cJ94LHYvx8cyt4BDS1JRtxv9G7yPXDil8HZIka1t/ezrG+VGCyY6SdvAZVOQq/6lz1sUysHN+8qKYTXRz51aGQt6Z5IVDsQbzFrep3q6jeObhDQOth3A35/hbKmqi6G9mqWS+brV44lWQVHsuSxZ60NFbLCwRRbVHNkfHRMETUTC+AOVEgeLX0/XceridejCLMYowhc2RP0YFfdb1ykbGlDiy9ciQcFvXBhj9gCCh4FaAI9FmMpjEBklQfRhyFLpTl2pwEI39fvSWEargw4bOANG23c7VaXcLMpfpdX3D92FEdihQsGtxJp1rZcrIFyjs/xYKMc6Uu6bOnvQtQR1AcW8x2cZGqYeLNE3efQnAmzZrZs9wtpxGScqChPB8fUs31feCdV/JBP55os+UzAcryzzplveLn10LtDHqxDcmJWzodaalQd1WmwxJ6Wlbib1I9a++C27nHUC8mF65tWULMpZuooJU2ZBJwfvpCVgMlT+19qyl2V9lWGmRUGA+49IfjXtrg8P+J9wxK44D01xrNhMuGv4z8UTG01enMeIz2Ph53GnXGqP1L9eDiYgp76TzcLpsuSutvJs3M6SrdEBFFPf0sgzS9vmpo8BtC3RBB08GthaPJrplsNOugSlCyxxJKI2RqjB6HwJDbrvO32JUKcGlF4zCMSJ1trR9PB6dTSY24379EQ2B0ZbYy/NEJlSVhZ1StQXRK8gHC/dwnhreRKjVnX8maR2xb7gKOE5P8s1wF0gfUeldVDphFWAW6i8/Osuagi+gKlznMtiuS0JrtdU7oQNzt8fECT18h6BtvdsrYg7Eyc87h7E7g6dbKs7JyrVVEGRFEkznWoaPagIJD//rfvttjjV10e2Pa7ZpkJaPkPruW8P0WnehvDjeCGjs8lpNjsXgibktVMxu+cEWauz9YTCZQbP/p3Ia+Ts0MrXPjabVux2js5TQpQ47SlhBNvbO6BphqQ11z3pmZBW6WQb9axABW9NBNi9ntcuHVKTwFhJG6MhX+NtDCw+ysOBNR/9wUWW6xQuhApv1M0p/wo6KWPQ0wt4CrN1NLiZ6GDYNLCYgKPkJTdKYXDVBy6/GngrmGVmyN96i0dC0Puc+rX0w/V8mbztQw30pQoDgfjbluMXuefLwkRJzTP6IXwy0sGWvOdgz2aQq5Quejc0iEx7kuI/j0GrtFx4ABCVPriuq3BMv+ECXo3FY4JY69iwxhzzOr1TKdEQ+WNTUCtaMao0o8VUYzwAnjOXAvOsZPiirPjtkRrg9vfhiQgdXztnnhe+lN/MKck+buimwwGzayo9UO3PTiCdGmtd1kUzha7CFuXeg3yaIoKxT4pbRcNqBoQFfk+rPOsmwiPR1+UGIxEmYhNFL3IEm54e0b+MCApF27GovKuL7ygPZqqInmbvvTyeF72bivGq7/f2sqJTOQDyhz8W8lh2MqO1ZDtDhiRFya3cxnSg8I5TptMGIHI8vQDorLWnoE3Gwadq/E2n0Vs+c0+bS6bFvzMZGFTyePpLNhqNV6LTNUoDBiJTIWEaF7CXeOxaZrjXoQqrxxAHdU/FYiM1Vho3N1YKBLdcSrJJQv1/hjiO+fZ4vjc0HRK29A3dE9jvoO3zJ5jjY7TFECmUIPjTylV5A3InVW4NxhTYSJvz4jXJ2S+ufBDErzeWzTnSh76AmDryn4c79nyCVoIDttNd7x5MRRSaLqaQFtb/ZTXeDH9/Bwuklv3/MK0qGPSx9ApvZ+3rYFaZSwJXtkgrxi29ieyLdjWQydgEVGQ1LndQ9yXS7OUlEFiLv2zbTaIBH7YpP7CzkDrH4zvMW5rhomBttr8OuVAhDmLSfveNCxfBMWyBZCqM2Tf1p/oq6h3rY0kwWAONnwFBP0Vw5AGhgSWv+lYyBwjaoc6S+lWiSfpDvm+wPx94bLuAkaNVAm1oj5zUSu4F+e5fe1/z2dhqoDvGXL5KNS6bDYY0FIkF3jEa2+8ddER7A4zbtINjRF8f/PBdwvoV4qLw+oAVG/6eGaFWqxmsfwiDIniJVbm+snr0MNgNKV7cxEROT/jLGRXQLuGHAWoGIqRJnubB6DDx7fEmnGJtm/HyqNvvox2PBbsdDNHwJAhGcRZuVW7m+Oeb3Mr6lOouTKFK3dBPUM0rS9W+zOam1e+c+3LWl9yV0zT+zOp3/+FcSqpj5TUI3jvi2qqSCRy62J6SwTuFDzGmuuhN1puC+l3OjFlVdhUnx+EF7XYKnm/KxL41J7OCT5lT09ek3gOiVdXvzRwQZiTzzRFUa/fFKZn9iuSB4ncVV/VSR2lTp9S/Ua8Y1cowWHkJborXKZaF0C9NEYs2uCPQ41furtpHBR3HkHoGQh95wrdE8Ey2MzY51sM7IoMvKGWCRUfKMZP0HaArMN/MLJseS43TsAAPg8s7aGGLQdd13PUhwhrSS7bZ9cyNQg4S12ou0MMVtVsx6mmCC+O6ZzaG2eUbuaFxzR77mFa6UJe5P5O2uAHPvEfKLNqgsw3188yvN1PZX+zu4lX+YJikYALvBrpeyT6/m/szDm4vU55OP69wGvMRYTw/jW3/juHG5JfqH7OwMY5aTqV12mfMYXhHXW7+JAs1mgqsSQMvFkf8aqQ9qUqEbXsrbI6NJXZCjscd/mD8l9DK/Xvpn6sH+sCakJlKBwcDiQd0ssugHRgXEUehKQcXy7MBbbDCdtXUCWeJQm0pQSS7M2dGk2u0zYLpcy7LvjiDl6olvvsUlDxtZr9Vqx38GsE4AxNdbNgqRYjuiEJ3xk4BC9iK9YS45wvlCQpMnBTPLl5z6q07vbnvsp3NDCwJDt15C/9vDzRRu99U39MUGijkcA1pMj55RKF1QNRGmnPj1RJOILDptrK2mthE4Tg8LEam25OoaEvG5f8wBzAPKgszKiA5qk/02azh782T8DOCu/Y8u9UHpDBXFmgA66kPZkEdtHZzcw9Fwzkn6f4JAG3LmyQXkHGVmfTWXIeQiYBwK4NMlYWSl8+/wsFa633KeCep0huCYd29DngcZF4qq6SKlHsmBDraey+UQK8WJ4iMarUt5zOUO8/J7lzjfsEo/swhfzenE1AoNllkJKP6VrwvkEa5X9ehMYBxj8dstrZFkTvsf0xaNCdwN/RFjVnSIIbFVDx5bZ3K5KroW/tEj6Yj0vLnTx81/HKlJ1kq20gA/V1F1wsynnZ6fdZJSxwj6WJLRAn4zIJUKTp8a5v8hlKES2z9D1FqbdiXTMFpTv2ysVG4DqHNjRJ3at8UoH9BShRMq1neHpd4BtIAjSYUPXHjjyuuM8Gou7rhnvje5CidTkO4Md3Inuzj8xM=
`pragma protect end_data_block
`pragma protect digest_block
dfe76e4628b53b565660851fdde64c3b1d323109933eb0e72c91a3a35f7baa26
`pragma protect end_digest_block
`pragma protect end_protected
