`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
osDZ7wBG9H2JjQy6xDNijBVuErJHYl9ecBRTB6bR9ZpzjacCoigS4o65sflQvnx/HtC/nUkGxDKUdJUUc6A6eB3xoFANYQ/2vS/gsA431BY5S0Kzz17WtAopG4MkAdFcPCpSZRN4nmYBam4ANfQ7hzFj+Ex7LPCcE+wL+nTxHanCvFt0tV0DU9JRRT3ClibhI3W0dickvF2ku0gSPqf5XNVGe0E0h2J1wM2R42/siZ8kvO7S5+p71vwRcQDrwrOXfZ8RFtuT2jObDHzPRpF45Inrf+oQFWFh8c53gaBRrAOQkjr4Ate91YqIDggmicgiFaDoYyD6wdbGCg1E5K5QK5wHMo0VMo5P8CJDXu5oVv2Apd6Hw322bhrEZSB4czBXa9b7vj5HTADwN1yoy+V7ry7Q1MKV0u1vuZLrMcZZ+016ordxyt7n6RPbeD13XQHP0c6IgCtDgNPJqMVWNHeH+qoMlsFC/iCAOosn80pN0TcuqmKeazbBeaUqfSINoHdrvxYmlCR6dq1JuPWj+HSDa+w263I+oDlVvQX86cbgxcEQhishvMQJ/yeadJaYNJd/FFR1AdYtwP/5YSSHKOeEuKcDSgPWsw+ZbJqX0uSinz91Lz2sy/SQp4SfaG1bq1CGeXp8OqKYf9etBN69HYBaI1CScC/AvUsZUATQTTlARNvYYjnb/X6iKvrwHasIcnuJ+MjXXNx93xiv+lqh1uqckaT5gUIWATTZvwEoF5/vsKM1k2E070nbJxm3RpOr5vGUxT3bhkTE1nm4vKFjY2gjSqAtRxOdkMVlFxvU6hm7cNnquk9RWMDvpuRn9DU+qxuAyY10kIKzbpMXxrk1peaUlEGy/OJuZWEpy2i1whrcdAW9qk0kCSHlvr+3SCYwqspMlti+HLeeDBd/J4A5HTV9NI/NwtYzLfmkywIFqFJO3qIS7L0dt4LI70uhaRxlg13KnqixGXGjkuAQzRxLyKjajJ1UpAPxz2dyPegUEeEAFdr3cndKAt+7IOKxHnYwu+7qRdFXg39Xywh9AMxGJqWIbUul7vzyC6Ski5odCZQIWtBZ6wIa8RlcRzQshPgnEFfcpIrish2DYIF1TV3o3vcZrki+swligsKUkGHlEQ8zeHo7dChvfV4DWB6NbIeaIT3sjVEoSb4hlZFF4agAxJ/OKkkM0dcTeaeTyQJBMqg9hUAjDrny8/CbFpyxVRQZmNGvvE3BmcJCimEVgyi+smwg+1FwZi6fL5/ZeyVbj1BqR7ZHZ9Bt0dWD2nU4B77YLqr1yjEWrH3lmDHyLQ1YswxbKDT3zIEC8jnfpGeUFrI5JOpRGgWYqJE8Ny9aHSVUSiiQRtBEjYCHSi42Re7Df4Jwyl1KxvVU4/yOjM7Fx6k0IVsgBMdUhn5jt7/2IxhKJDhzqrmummbRYpYXJQ7nAZxVhFxj7vJAxa6NDR8yPSsJbRRx2yNWqDxSn0x+RTQXp0ani1nFrOLPRx/iHCB2xlB3C/b4kE++RCcLY79AxEvJnuW1WmlCApL8IkGFhz8bAw144yaa/xjENKkJkWjQbCcgb/NzV8AG4JSetJt9sX5HDJ530SpOavl5d18Y2hLDwta8XcBfNWAJIioD6ge1OOXWwbLIAMpxMcbG2HkkqPWj+YWQcMHsa7nhgyxkR0an+xmfspXPugOHeJJOe4svWsS8n2hC/gzdPRqDKGTvMpl72K/it/U6YaftrW6Tz1eWoyYKdhB4EIdpp+e2g0aB+4tqY/rBqlV8cDWdDWxBGXUCiZM1TjpyyLxth367QdBdx6rX6okwWMzRLkI8+jqcjXJ3lZNcSof43rncwnHmqBuCFb4unKLtVRcJ2YBFzi7+IchZYZ5U4qq44qPnOGE1ZIrKLOvfsYJ50EyCCF2+bdyn37qmTi0/UIItGUYi+08slFBLO1pKYWKx09g/2LjccnFnk3GhkbkdI/FFZ0NMpG9V9y3uXVLRyZfmZMoo7YqXarEWkBbbsUJ1RLaa14s6SnbZp2sJsF65xejg+bpnY5Y48p7C6X/fTnbQTPceGZZoPabwyhyFird8Zccn/NPOLnAkMF3j6JLblZ+ACPi6KVklTLxgQAOpNJ14/CFwQSU60X0dC9R/A7q5FRze8BvFYFYz34y4HWx4gUuf16gYSnRak5pQkanFz0rHUcHJXb5sqJNBhjF/G2KYpyFYfdWVnD10OOTvTqc8bm4GZE1w7VReDE98YgppKK+TaUl5MrZ+webQSSSwOaejB17Qzn4Ch+9sTf/tO83artU/qQWgBuBiRbAOifD6rP6UxOOO81W0CssMmw2OuJjfvzRxBoRSprJU6waUOw3nNUpHTO4uksOqLka79mFTIBdJ4jcRxMaoStcJj9RH1H1YifeaqMf/Z0Z/yb5NAoxsInMGPMUudbFyfS5gCKO3IEW8a+tRcc8gnpSJBnz9CywiBil3pMuYGadovtVeiat0XJx6EGDydC1pfnlvswmcI84Ysa0QX/UURkcJIfiGzPy/fGoNf2Wfa9kdRK/wWbDoRXFjccMKv36WaQE++Ksx1JQNph+WhHUpABscK6NTDujG0e90nSVomKoo1wCTFREDgLy1uhNAW+IebM8SdJ6bgsPRUunguPyxthBrMK+JVcUoL/uoOBA9Si/6Htt7q9+vndG4YeV+/xMDuM+LFKiP2GM74Hb6rHPCYfFXDya7+BFENsGsyGEelZXIFIeDK13ppXzg1NVvMBDQGXIW82BDThV6szUypdcpyXEdWTUiHoGtyJmZQmGCqNsubNbW69DNYeQdk4nt7YmVo+J5JiQ3d1FhC00nio3J0N2qqtPFIlN99SFtOZQEcAJHbq8xlXdt/qDey2n3zN5lUuBi0qSxMlElnD79AiA/VFL2tjpzih+SgSHzF1ofHE76W8qhaCJxwkLt/uPhHtOhRqq6qfMoZfu7oA6crEsahUSnhqy+qTK+9PSeKSglvhnyeQJXlJGdQSS+Pr+WzCKdheNuEI9Ke3ZLhqXSYKoWcwKwjG9kevi7g/CTvRbSMeHtHwNmx0IQfMQ499IPoAFdso0GuZuBnL9SdMHcObLhJa3NmoOs3wBUx91dLtj9MShGtbs7Cs3YUpR8u7k5lSgqQ4o43ApxA5/TnGufYp5VkndKNHZ4no4TctP39YcUgprv4oU2iNUDVZ0Wl3M0eEljuDguRyHYn9HbzezqEDZUFCBAR7X/W4V4aUIQesT3tV5kQJnv1nFZOeqFxUCK18hlw/Y3jugbg+Dszhmch20pA96XgOiTrnocdikS64h7r+ya4/xHNCxQCz5XFHHM7dxN+WMX1vcx4jY6fQaQ345jhQLlj3wjaITzpPzhdei8eDuCa94XPr51yjEfLxADUJ2WKNu+f9ltTHV0f3PEDPdiwC2x5vPLROlkMRA09hU2fondc8MHetMkptEC9Fm8ARX8ppSxH9BiNmAyK+nN+ZTvQPVRHe525za3oEf9VY6IoEaXhGJxklTGCE7eKQfLVwuRr0f3pEYYHX46WmoJr6kV/DLLr28Twp9UZWrx8TU+e7zF6/zdI5Y8EGQ2FCRcwVo465/B/oPlCypNyOFVa04puJpb+pwO+IZ5rW44tRZhDtksSmt3aTsBZRlKSXRXTPfbPa7ACxZVPQydhWkvm6W4hRbHwBaqsaPX6J0drSUe51fv97ZWYRtd+Na0ryAp6FUgWtzUrnYST/6u5cVVBDUFuI7TlrzG+hkf/LgNbpYdBFDnFZQ8LLKjOTN4O6EMTKPSFgHO52vgXIya9zJuioquoWvjL/G6DYiHlvxjxHEumdwq+JJMOGgfj3d4KOoMSEsV2Tx0mAPMGpL7vZNu0xWUo9S/f+tcocNFZSHg1AAUXVJoieG1tx+/bjHH64m/dSgmY23VED+IFxnz+lLWJ4OdQSWVLoNfAdJng8v0g9ZH1JgEbCVZrSMjelLEm5pAIw7TPNTc9k9Whq7QSCWAsPeNq4/ebLTQPVukopbqjV2IxCkBnlw+z+TCYrWRap4RoWoxN+DgZSi1yLcKLXnQnWd8tLjH3J9l9XLAyIWq5tobEwBtsbFMtMxtlHYC8dM9kEiunLhksttWXsxHxkJeuGd/f+vaxDN2ApM6cASlwES4NuwqJwLkEQ95JaVN6VK9J6LGp+hw4rNFMRhKKzUpJpLNgZl9CUMDjmsaiRcd8Jc2wjaBlRBivKKnIfB1gdeWemAsSU10iBeql18yOoeGMGSPu5Y0VUwLpN+Tey7ss5b1SFLwehuvR7dyIhPS3MEeOXiJp9MxPcVQNJMooMN8+vvD0V9L2ambgB+1AgEPQl9zAMPcZqIaazT4faqSpMJBRZ+qbFizmRu6ghgJfAwJCeP3QRmP3GqWxgQdcHRVvq5n4fO1ECAB/+gJ29gumxR9XnoGPHGKp92vpDIoupccyW/uWx65DLE0V27a5jw6V/dcqf0gq7VjrcYingkcosjLu94PuMLL6Z1ylw+V+oNzgToYg95KVmYuFAI5IkZpE2VFrJ0iTDpFZ4bK0nhKrnQNTl249nLNN01NhU7qaQwFqPQBLxycEKy7new7AQvQX0qb12SD0G/xyIirLvGYGjWwE9aIgo2Rinm9El8+98zI4gPQU2F0CnU9cb0UyGYXc65MU29K8XhGdWA02EWKeQDXMxUk5nCdqKDqHlprtIcCJGZCUbE3sc7X2+R8UZPQi+fqZ5NbnulxeXW3pJ4wIduYRGGxeYzV4IUxOLkXQCSFIWCusnbcYl46Z+CTHVBqS2CY24TLZx+/venJ2lSh6eOFcNlv03KcMDJzGQebx8EWWlQDrqVYGqh9Ze18zrPggSjfLtF7WlIwVxLqNvuAAbDGO7s2m9UTC3nDv8VGUyQ977p3QnrQjv5IQtH6mvwQbkUWr+nGbrGulKYULewsJnSe4qAic0//9/ufm3YkOcD0h5BaqenIKhLS+Ieusm1FeAlgfur/kMGF0UHr9E8HD/bEt2UpALHD1DpdUvXYYQHlcahFY39Y7cta88KAwwi3LK3TUMHLuBSy0dd3JUrzX9FTmxPdXwKzKNslwaavBGr2m8wwWzuiNN9DxDzdiTRiviCmlIm9gFfBldE+iGTSISjyb4/6lDGOwtN69lmdCtkX4mydSOTHCPG71t1Xu4Qw1seBDL6FdvpoOn6GRP3cHEuIa6jGrsWt/ACX5NmWhbXadm2veB+/XGjGGGspub4IIbuasj2RANIwrrG+FRGFuGei5+FitUuRhYXGIS1R3Em3TeaNK2hG00lmHOg9kefbEf86rL+/szt++Gtm7rle6lMKT0i5435wo5W7E8aepbavdEQB0o6hofUqY+gbPMZIXgJycrrqm/xUDb52PSzKmWHpeW+eXUEyuCsUTMkr/bNcafuRx9cMfLRXHXrqqiDkJOJm8fWrnPN97lff9bpPiVucKdImV1qVKX6SDTL49sTOih6X9/PZjTcDS4WsSNShlC0/SBZel9lQn3nJIPqFWtrmLbsjeVPpMwdaCZb9yiJt8j9qKX3otLQykTs6cN2s9IiVsFFHpxgnvKDHx5eEkO99kDkvjH+nAuiuU8SfeeQyF3C2vl+pqATQ7VFz4Ik+3B5kKoYeszitRojLGvvkWRj0V6E3xV03zXdeoiyJN2Nf9jjAnT61s6ZdMuPMlkgau4LWzb3Vew74FdOuI/y3I18XPxqrPF3AcOMZnixjpvwnuXQktlC8AO0dsA1klTWpO83t1aqHEsJyhlZ6JLXzGo3xzesiWbSWTbF0d6RRsK7KqTthfVadmYTzxGtZLdWHiz4EdtWjoJVX5fFWHzt6/hnp8qJELzZc4WAo0ss8WpjXuaSGxppe+qBFUsQRr/9QJVGy2Ps5UkpPAuZ/AhGg8Ae6Shd0ujAjC5EhMtW03LnqP3/NiDZ1xlxPmuZ7TnSk1UOY675Hu7iVRyGlt6UKVWdFs7cY0V5WWcZuTlxlv8koqR1Zz8C5z++wVs8hS6M5Kfotzq6+tZCfVbu9WKOJwMlXudPqZQgx1l0liN8elagI0ObJrtepn00fVxoUkbHOJG+Mv0o/KTTbPF0RBAn74iJ0BARSzjlDXILXcXXUeF0gI+oubEjZJthM3yMqcAOaRHx5FD5S8cFF52uCVqqu8yLGR176GSjBCkAcCsw+9naL924bjkM1c1dUFTsKaVQrSaBdemalmPKI8JepEsuZEP2mvSmXNbAfnROXwH014r9WY8wpU/fdKbx+bsTysiSjuzSydpENhgEUKYwoFIJdksfNKZDskX0C0mY1gr7WOoQzHI1EeVV5/hIj2b1Se7dl3/NIQRVlSyNZBpiEq+C92AZC5x3xcSUiNHYhXG2q+0z9rvT4F2rIkcIa6AiQNgfH2GDCwratMNxEZbVruOZMpEcfPr6mbH3I3C8Ume7/gdlXDBABp6pU7SrQfcNbKOxMuH1XDHZrpjP1tE8dhq8MXWkfX90F9aKOa4g4vWigrZTkw8AAtupw0ULyph/Upuna4REXaFlSIlxrx5PvF86Zu6v4oXmipgpxFgo5zm/d1NJTQl6E/BT+eMNn+3mrMA/Fn7D0RfelVDAPHfSfHgJzCgzh0D5AJpYSEew1NfRofbkYxzdDf4s97EVlaI1qpD526aNy7bYAAFIsE2Z6ZU/bk3frtlcOn477vG8QizyhKc6Q+akDrE9nKEBT1ZAsU+eUcJm0KE1Ghc1xi85ZtehiajbLy+lWk+NN2gqrJCrB5lsZfVebaDW0n0GjHQE2ZDpqqIh/6Ypxlof3sLPQnr5PQ1Zu5jfJfFlw6sHcX8Pcw05hOWnl8d+tYRULUEKEYhR8pOkAXE6ijf6Bta5qVWSfy8YQVYn66caRvjNACJ3HwB9bYGDqeWI1hX/m6Vbt+EQeUyK83GIi/yXnCyf9342hKj0jtV4fhLSdZAKyb3+9LQ9TY1BYRHNtWJ5nzip6oFdU8q4uZ8YayIHMCDo4emiMNMW+qbazgOB4hAdk2hwa0abedDSyST99FQIme0rcOxuKp3ES9tyVzhYW8crXL/Bitkc84/hly4BnhJiAExaI6NZ7LY95zv0XmjfjKkQ1FDjoB17q5+RdhsuX1xvG58+e6G9obcqJvskCe8/hmPjmSgeO315ineJ8u7IcnBjysW0dupWIx6SJ91KYqwDeq5ZWY7MY5FM3h1toIQQHfQ9DoGyKMHgRZ2nlMUmECCT1eKydSuD51b3sasOt4jR5j0NqQRGpem6wRGlDnjOoOR69XxAsVEGolAji+fUrI8b6TGEhOeWxXLKgvuo+7z7ujXwYCom9jguj/wGIGz1pbqcYHXiUjruSoKCJjvPJFz8Uzrf75LGfdNZffQncUDA4UsqPbCRpC06lg4zYDUbfkzvLtWFJVIWfHjKYlFB1awblDGY0pmHZiPQuL1EW7AyIObcxXiee7lN9AHAgs9ZCyBhh7bKinzrGOOmP4WVtP7Os0Kbin4969Km0eVlGkedDVTwiIBwKC2XNOo0C7zD2tYqWtBALILYRp9TDweuqbwGqDsRZB1eGD8Tz9HgtdGzorgu/Hlv3flzw+a82NT6kgGEsgdyg+w9bh+OTLMFNitLNZBI3I3op8Y41EEdbss4G5+07VW3OOu3SjefOK+tBUyVl/c5BA/X0gvEnrTJj0tuUhlPzRBTQX/vedSw2RTKFgoaCFCERdqQ361yFpGofwMhXMjxM4SVhWckipY3B3EZXferJPqA8EfUpP1D8s+KmKIkvwgn7PcHCffXqzVDndHywUUPtdYb2038SxANnwaNFwNe6aH7Y6r9Go0RAcxLsyFt8vWxkgkpWai/mVfWpHnh6AO4t5bCT0hqIE69SCrMO+aNepbxrw4x/0YLWnmV1khawlg18D+ZfU3djCRbfhbjzngr0VOll6ONqT7dtne10Fz5nGBv4g2PiyWMgDJ6nBuF/mMDVwYa50qwpgUV2/U5NurbGxzkf/aOl+IZZmLscnvd18rmWF+PXwRYd/lH1U9wJM56eXWR2hRxI/fPaq9xpxzihbFTPJmKH86QoNXUYFyBXTg+S+wo1wdIIV/yLoF8G9sJd7vm4V5zJso6JPLVJINXSPOoGuKZY29jAXz+f3I7Qgxi6JnVZ5QjeCb+Gu7LEsBy9os5XtbM8wqOO44KnyzTnw/M3gBPyYiUqXhjBlxFjp5hxGcF1qZ6zqXiVEFKV46pBzUmBURx6FJO6Ytfi/mhzIL13tB9A8z3yVzLJW2R+6UR9wtm+7PObvEMWQe6UitpWTamoY+GihTfmi46nDgG6tB+mINZq5c40xyFODEUu158hAcY5xNZx6w55tmfZK0q4jfnCSwtLJMgYlKmV+3z46nFILYbXiYVHLvRVndq+7EoagWOYsQz66qNrivNZ8DXR+bmMm/Tc0Qz4yEsh6XosTB0+LIe7IMfNB3D4m2cUzBlMvIwHhdkEM0bJ7zZsdqI4zreMq7MdI+n3L0S8FODE9LKpZSFm4BzyA44fixO68lwWuLmrNLFMpYZYIqx07zWaXmQkGuQwA8R5CaMu58sP8CDmu7tKxDu333QKwafTo7Cvf2ZcVkS/u4FCaZLpzb2GyIsEWyBoKKbIQf6d3RNOVNFnSucO5oHt3ZXrcv9HL5hDU3jqZ1brf+fCRBlnGxMW57Fz0XD5GytPl9Hx8xd/p2ve6AWzJqBkVSv7pF/eG+mPdgsG7cx729b1B54fK8mylw1vAmAaxjmzkZae7XVKVXRnSnT9Y6auY8NshX7caNPq+6qUpWmRyLx6bWxlAh/eQR9bajBfIbbUmvaGndkMNbKKPSHC7Vq7G3wnju95xX52Xb7r6SSqdbK7BSsChjEYpoMvQjZSmhHhnC5cmAYJIUstTEgtAB73dMvCizQJnmy3Ef9HFsp2Y3mAwt5y91baE4GLHSrrghRiI918KMJBak37y8HnHI8sm5Pnq5oU+oDmp08fWZ8KFwM+C7PZWE/xrNZcg2ob4bkZ1GCFm2bOvS5o0jIHKuAnIAVGUke07xExVEU46aU1wuJ4+x9ggzRya680ftKF6SSS3bJa4WdtTjcePaYeCiv794ALApfT6PoTnRTPmrx8XUTAR/iLnUJz/0/r1iSK2nnDjiHLvr1AvvDg3frXw8HrKNXLX2TGVz0D475b+VGtFPV7l+yOOhZo2vPMu3TThvv8BG7TJb+TABK16zXFwgQfJhOSMqTFH3iH8QqVcQ4zDdvcRo5zdbPbdyfPTIwrXGdthpNe6tKQh3vgqVwggIY3VmzjyQXl14kEOhXyTF+0oBxIR12B0KJkkULxHEq+MfV3647suITmjA9F+yh5BmYGx9udld20myf8ps2CT7884/JHcAimUxrzritWpRKr0K6oiWLTy1vquOmCEAAznzMzshNJuLiOd7Rj07mWl5SdKppRoU3YJU6M0TvFpGsQv4bfW9yCgJljCq1cshBU8YHC0Z4e9K/ie09MkngVyh1YiL23fOclTYK0U8oD9k43l1FIYwqb1UIMPuxaIaucWqA0r6D0IEydbMMuhioC9td22aJtS+itA/FP0l8IKemiZIp/v1b9dAWA0IWZOSIRxb726x70emnGinhN9HEMXztfCLTq4w1xm0G3RwR+QV7DolLylpN7G+XMHHmLVNMRT4ZfGc2AEVer3DtPgMSc9M+vVURrduUgRNodTQCs8X216o5O5ZIYPNupy90ucrYLDg08Nom7eOmHB0CKEL0rMjh7yEHbiapWqYLRwWBjliS0DzQC10e/VuW/eznf3SDcF11isF3SkyOzPzlw9dwURCyq7aynB8hYBFBEkG1bMsA2h52NZVsGRbtc5E272QEBANT1H5PGvfHfxkdC9JStSYS1RD19dN5YW6dgN/2H4uqflzDczn6H0NAg5zRc/6/5JnQJTbAwHb6Sj6JUS8+hCOl+w+a8SuDAWrAkRBknKYBHmwi5qmOjFw1IxC4TOnM0xYGEJ4HbPfpaTH8QSq8PHa708m5OqQDrccOY6+DNTxKmLaW4EOSkVwb76xIFyjkZZKDJilrTOFyrtMWTiWfNwJi8f5+ExlbKeNUATZGSwWWEG9tq4cHD5fsSZxHd/kgSQHmqnLVvRVmAs65POkfv/pwpg9pVlLsWw5BumnQFO7K1ecrt0AX/yX4Tt+OVPnZOfdz4IpU4Bf9j8HCifwtePflM/5vW7NASScKlJIRF2fHLH8fQtyZ+7cAGhHKtI23NMFjiXDdArjenC5MO5kyEZNAClC9e3OgZdTID7vPd3C3k1c/pkb8a6zbOBxzFQhIF5np5HD1wZp10bBSscW+bWyT38wiYG/pXvNSp3LJ01UeYx+xX/JHe63311Y7PAnQPyeVAFBvQd+gt9CEG5CfoRD3tJkxVDdFRTEaDQpWoGq2XtvmkQ5fDRfBPDAV3rw2/BeQKtGZ9mwWp9YFFKulr+bx43RernbjLvqiMi+3M38qtZijQJRuKHxIyGxkegaDsEbN+IX4z8oYRD8jmaHGRE37gJ4QmT/HZbQ05qf7t6oB0gBNQ1gynZpegNkSAhfkPW61jPAxWgTTrN6uDY9Si9al6jmV4AIuY4wVXZxGstmVTwf78Qd/ee36N7ZwLwWSWmjKQ+iKGT6lSmJA7RIvbzT25OjefvWRFtedebWn5+iSOC5UxgvfdmvgPcfrABXcFB2opZDZHkDkeP9MNCaQbnNkw2EMOFp25jL5M1OOnZqDSZCjoqaivwATdECQKRkbNDgNFp0U7p4n3V3yIBqkNeeV9xPa5r0L9SKvyP9i0i7ZPE+ZKnW1aggjoPhlJxGivE25Z8CbpZefhQsP6an7WIarEBQ9mgOXO76hPDDvdCJx5t9WIdSgy91vEJAS3yYvAMaQJtnFwdxPSWC2JLtu9tkzk6ypppsDRT5gTD3FGG7xa0t734+MlvyH2xLIOcByjTb2GyXtOqS5s1RmZyz8ZmU4zHlvUtrCmIiw9trO8g43kg+Zpr7uTN/VQ5mcEgwL/s275fSbDbibNj8dqU8cAG0z5SYRHo4sTt1J294SxpFfSeSuKEgtXa1ywn66JK+K+nYfLX0q+J6WXec5Wk77sfORqCvidmLCdzSeFF31S0rTMiFJS/47sykFf4XGDkslgldKyAekXr56cd6HL3feInjD/80uEe+hB8K85whLPFU3H6mWC7cmommQ0WG9HSOJ4rRh3KUQAA7kGaGG6hv86FmWwIu6hN9VbMDL7QKq1mZYRw2x7IH3Zj/8IF0xrLNGASjhPUv77VBT+uFizdB1mqPy4c3/d1Ma6AjX/S325fO7AL0luFvymUz2SUIAa66ktKPfervP3XCsk4IG7zQ2j4kI4zR1ZDnJalnRKr+KAgK/ohAQNfEHl6KJmXkfOsLeQuwOqO1Aue/qPkT+yLaph36Qqy2UQAeWys64CFK0+QKmByD0WIsLz+CoHIYR0L3oCjFQnuieZbYUaxWd9EqXKpn8+nmbVYNOXMVjBmAdbKodWrWejkJYeZ0u2j0mUpYE9JuyjSvKUrc84FI8D2qxeNCzhDSmRwBt3hkGPI1+i5QHBAMXv6eH8kq0zU91qi3PI+Kzg3lWvmnD6w3kJcksalSsndzPzjfMvxVnSUeAeK7vn0b0N/NwaljPVFMAVzrrixWJ8XIHOaDmatWvCT00fD/1WGQlNjPUEcneiuxqTHZjMX0eBAuRXRQOZZOh2fSMlhk3LfmMCVqAkmNwyyoolKRcevz70v01NrKvns6F8r12MlWx7S5Ar3gEVi0fp8R3JpmPisMG7baeK3MjmLA2s8J7aL43wjszTAmTVFOG2hdVpIU5sgm2vfub/Ct6kOxhy9REvp9bVEnI3W65L4TGFaRJUPhP6gnv65LHYbExFKpGlXFoyEL+OsGxpU5SridjWCeFahh9OZGdfs5PtKyHg/sfbb4hQpIiAskANoCqoXYK5OiDUegBj6zQ0ZS8/uEXmm0YJ//4dxfNFWkRn2GMUie1DNTzoRboAUwnXo1l6Z3GG/zxYoKQz/uApCTHokIo37BSUBjgcD0QNCHX6bEabosF4KYM9C7AIy7ZNavR6JGlYCy3PdhRaVl3i1oolX+57YHvXv1dVDSjyCHEkPZhScfiS/LGbmHSjAspcrB7ywn7gfZhfDuuxm1sZDHh5XmLEaKGzO6ANzdanAaXyXOocbd+7sImzMQwsWGRds4vi9xQ0UqYwDYGkzVHjo8jRRugcu/uCUwlsmve4YYvtfvbSxPQBOScCpCZAPUwWzZ4p6rZm8WF8S2p+lZuVYIEQLDQuHv7Wdqhkdk8yWN9MPqlnX4eWtbWwJbqnN8NETsHz2KfDBRmbAOJzxDwZqhgbPIHu1PhPna35/1XCWcS6RYrNuugBrBvjkzRheb8KJKc/8E6sPCq2zw5p3XWyP33jUB3H5zujSRcXX4bImWqflBRZaUqBMqIzqccdrM5Zb6i7nMxbPlupmdtaQvrFf2K6K2ccYL6S6/98G5BsHaPZB8ig44MdS6ozQQQgs6v9MCQv2al6/4gFfTWo6DqJ6FxRo1fe9x8YZ9fTPPUU9RTSC41VYS6D5kOQW1WEKAvuMyveOGX2e/N+AA+3f+K0EPrdzZFq6Zw4FaDKfneIbyzYJ1pybTmFbIXOWjs1fEprVnij9MGbeylZDh+Up9+nIMT3T8OXoxo2XWFjVk9LETVXtK12s+aAhi+OH3v8ONm3/+KkodEk8BvDR+UfgGU+ohtTCOKr8aiLc6TnFW8MqHp7qqRj5UTdXYfWtBtVCdE7ZV22B08rcDs/XerJXkdsXGHmqp5ojK9m3PU5Jcll4nBb9MY3uzEDXRd+fjH1HAHL/F3fqlj9hiFPeMQMZY/6q64sWD9h6OPMxs3i1h5VWhq0GwJjda9/cxjop/I2N7ylsPfo8VxJ2kiT2XgoiJooa5pUeFlqVvvgLOjNphbkuv6y3A8nXfj3Z0KsTxXAIJGptkd3YTosYVN+0z+a70LPMerhUpMqMcy4XoeUQvhHMLVzjlYft/eD//3E5odOaphv3y2cG9fo6x68/L4IN1q5ayU9mrUGQ6Nf6K6W9FoF3Llkc7AXPRto95ly+EVMEsskxR+xJvv/+02SajQTEc4NG1kvck+Vn2S/Q3KkRkawk9noq70ohYUTXtYwMaz4jEqN9cAR5yuJHVEB+xrYH8AevAgzM6McbL9jT/OzHhvt2gbUVRD0GGpI4vRu60W5utjAAeZe4FYFnBRm1JmGSuAcWF+Z2BuEQF6Zl6JWEAT2ARlmuiZuh4ENAMU7EIlRMAG2nuCBqfMrhkeUK3xLP8Z9hwziS/j06TygO11K6dz7MtHMhfxMd0Ms3lTphuhG8/9f9ZVRLwHcL/ANNl6FM6i8GFmMvBrOA7PwzHIlm4U44MZyA5bVZATLR/KW0TYlntOrT3hxdm7xXMgKIHu3oOOoJYM8XBVRcppyLlHMT0PacVIjgYl/WXrS/YXcopgv+MkxVFDz0HS8H8vBPjhg7+Ois+pHILCShXql1OA6zdSjlNZATLG8ZQR2rvvmXmZhwRj7XUtuwQFDOdMO1b6ah8CG7LEEi9ujhT1uf4L0X2usXFDO3Vb9f8/6PEeemilv6xcnS8o6Voqecxv9sAAUuw15LquEi34hfTvYj+Ocl9lQEapBBOOOBQABDvt5Ib9GQGqrVWQEFtIUaSVUW6h9Zg8Xxangh53f2slweBGKS3AN3fOgPgXS+ykBAzeR464x6S9RbjFAtDmtXX9SvtH4jcLl+LLgElC8VD/EDs2UHigbT3lAqTi4k+mg3jWZmxgXZ8VfCNRFYUQWFIEXWHgy7i6psLq6rlFsPjHRY5N92GNYsCDV5zidrvvSjfXyGd3Yqy1wngJT1Xn1koNJ2kaGJZKCl0toifN9WJDgz9drH3LYE/MbGiDyI1URg8jp2ARrJ1g5D5zbCQGfUomDLZ8qah1aLF2aqmcXbvpEUmFvHYdKYOr3zD7JfkLS+g3u/KnQ5jBEADTofmOfKN9KIYmfarYyX3zRlkSfiFoKLlsxcwz76RFYLQdUyYO+XZD7SYv+MSLSo08Y8IJ9rFwnGqqanFk0y+f1QDKhGG1EGbXvf2WC6/se7DKDYSP64iyS+NYgtmTlyzvDupiseY/HlUu7j5OmvLXtvVuY7KU4RUEGMOsweKSQgsQwB+Y+8BkozE+7aGjz52P9nFmD23EKQElr0/Wyd3PbE4i9COoKhUgXrPyXhH0Vvml16OzaZJTd9tmlh0OUSJs5v55SBxOG/TusBP+mYSXxvsosvljH5Tahe1Aa48dfoxXn25IeWZk07r53DLlNZ0ljyu/vRBxdj0OLXYsn/hhbFr/zWQj2CSdqX3LZOoVRqkFqP1FEXkMUsz8u/r1D30yWMfu4K0FsLFz+6SmTVEjxwq8JKkFig1/1NmdcEoTP5+D1AOAVApp+8FBQZPk3nd2YOSwgoXAfVkWfJicMO1jZxPDRF5FFuT8PiRASUM4g0X0/42F7/rEZ1TX8kyjIf/X5iF2QmgFYWMuFmO8ELJzIQ3rQ1IHcJI+6D/VHZi5mWpltOOZoRdTLkS0xNc9cwL6B8D4cM4O0OPP1WANdPRvpqWw5CjqHMLBQhZAkyCc1Mt0JZnKbpuCOT+4fjwVFMVjlpWAPqb0fk/tUlPHUZmBJlzdHR09RH4KLoVfTN2g4pw+GkO+qJi0PjG8hCB1Wg+bcpe8BRDssYrO9GpbAS1OPtJBIOa5gzA1dUskUquf7AitSaSk1Eb7QCg23Mr3dZhkUJvi1pPXIK60ztL5hDCjD6jKyoQPv/YUsCKmQdKqZ3B6F4dpqA7k6OyfFv0U4DrszxSYMnEqOe9okcxFh/IglcXSza3FcItZ1ZB6bSsumxBoRDYmPAABzZQU2OvMKj2apotEMnCuiZkVym589g9lMJLK/U8FAmqlHGBxgXrAGVNYhZTuIYj9lCgwwnkR+RKLaiQYNCIVoinoryKuNsp81EcisbRq293uaareTm5NC1ew8KAWvtwcdegNNrXbDYUp/Np/NU8k9VSk871noYcDtu9HDmlZ7RHK0NUDIhtCztoy/Lu5S3vOe8x5FBlD0L07gInqGl7gZggV4dRxrVaMbuJbbYTzcJ3QoxHLoyyr0JC0AHzoZXcdGy5XuTx0O6gLWDb/jmUYSomW/hqUKXN/YsNGnwdb5d0L87+LTAumDBPgTsJM9axqsJu7jk5aeGKmBxGT4SbMx1ROZy0Q5A3OwAKXFlRQ6JDOIb0EWDNZYGFk7R0XnmWOykf3O/foe3Q0Ee11KxNLkxGyzdPGzD0moOl+g9pekCalVi5XJ8QqSnQ8buzoJ3y1j2MSPgKjwdU8eUC3p6y9XvL0vVDf5ej5cAG7Q
`pragma protect end_data_block
`pragma protect digest_block
c8843736817070778dca1601bfe43645369d0922269ae32a6ea52037e360afe4
`pragma protect end_digest_block
`pragma protect end_protected
