`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
nCDzuUzCQesTtYNAC9ymJvWsaKnS+DBVwasM99q6hSPOK5AYAdLusE/+1lDs+n2tDjunbt2RxRYkxN5LFKSLXIdITEDxmEavn37JZPdluFetls14Tfn3nxG9P2IdSeZQZmouNwxjmnXBCn+bBORoUQfHX29JGQDDpWH5n54a5inm31tRZbvLKZ4C+PLPWFPSxnsMJLuFsQChgEyGMV/2/CrdHF6AbqfOzg/4jFXZPpBh4iYoqq3iPwvaBcEzOu1fSA9oBfCiYDnYOiA2BOdWRa1sJmzeRHKkFciVtWpwAQU7EsS9GzyOUVjo4LThIg4TY9pTmUVbnGO6SULCP2YiIezBXdHSLhjVURU0R+ZS6IqE1OZmUGHUYZo0Bntimyd3lV+bxl932CcpoHmEs9hKyz936G+R3Bz/Pb+Fl4m7mu5EH3bEr2wJls79c2ChJYkrQ+F1Qc0LoAq1dExBz/4GKj9LFmmPE5qpCzylc/yz/YwCm97/j5FYzt0WZG4LJM+TVe3wf3MJj9kLV/1SwRl27X3Fbp+IH90q6Jav5hArCYEybPaVsGYItyWZwr1ePdmzESU5yTZJFOwftYqmq+ROxNcQd57skBtEyRkhf6jG6mO9WVgOr9j3huJk/p+AM5WOXN67lLu36njhFF3DUQ84uv/qfDxVh2i4BbmQRdwEhpEwoTDP8giG3TC52Wn1NQyxhlZx1RMBXyNTETuOZHpDDbbijsEruczzLJknmgs74yRCTuO1Jx75YZMEGVgCd3RYNqsWtM54zJgn6XNdostFYacyP/6n0U3XRsb5Pg+SO+D0FIwE99jo6sJjGxkBs8stELGaJV73+OKLMkV5z4nNZdCasWjuvkaTge2zuF3RSmmFWVxZsbsetmiPEkD2j3D9RRJKRCxEURO5iG4jZrbTpEOzoDk/++d/n2DfsuMFRWgqfE32dBENsc/efhtr3amvZviJh5sRNyZLtg3E4WAcjgyzC0Ffu12zZJWrLeIRSRaH8gvPeYZk5Insm3OyBe+6ejcVZwD+8sO+0CJnXGFLzRly5sNxFYO3j77yEXChJTqwhgVILbwHwxXuvM0swDZD21LndOMdVavNuv1tfyUBeWFEnJioGliukg9H6DZry0Erxwb2yyCuDRxVOrAUExlvOv3GOpsfPrsKSqbfgDmnwo9Vvxq8NdOewJcA2IE9e+aBOG66GwXvsINYyiTpdV2m8EvIevVN5A0NTvW1gMdkMwymmlpf8cg8th7ocPYO20cokxme0cNsQHFy6xFOJefk5v3g7qh3l1RQdTiPVgvzPr6Poh7AQslFwkJ6fZEjTqVu5Gz1KnzM2yuT9/slhmqEgpszyayktXwMJdQPqHAdmA2U4eHGI6bitwg+MKQM8cNTnMsOedJU6LIdUCGWm3x8oSqbwAKcXHusVdH5sh8gLVqTSdkLQVjo3L8VsmKTCug4zRKqw011AgoJUr97Y/qJX0SCMYzr7WtvrQnOQjz/nfCA3PUS6VLD+NvJpT7lVJGwSzUgTUlg4ToWGnG01CY/lPa3RiHmxf6J40my244VVKwyXrUfzXdl4JlenHkH2Le4XO37G37OTK+gbd7P5lGGC43qr/J3U06C1KBPiFwQ9/et2JkId+DKAmrGnngdIEns6PG4STgul+8sdF2KZnnYog8xv0qD1ljPhv7vKcOguG9Dbtt3A8tgHWbHAOSgOaKio9FrIT8O3KgfxBOlBNsTT6SBoPm76Sn3Fmoacrk6SKynh9wYD/d7hwHfMPeVIM8ouhCRFN19YCd+lusFgsSFpYP3N4onpz6mMpJgaWTvHqzw3GxtaOk7p9SqfNsoB9b/ANmxKM3CYB0CoyYk3aF/5MDXXzx2CX9JBxjGHLQhHhdIEbk+T5bALFTiIvgnrR9N/jVBLFE8bqHX40IyISffc0zuzf3dv4Mqi4l84lZuUH9hkAzlHn/XRgd7z11ahTNQmQa0SZl4qgPauBJtby3fXxFCl74mcB+etXGOW2J5VmnEO7J4YFMYzZ+zgEXP419qossyGQJA5JOWKLm9hfnKryaKz4ZG1S6ibK+ngP7P57mB/L6XY0zIELQPThrBktlpgqnQ/Q9OXGV7FZCM3CsrrfLvBevGWIZeQ6MyFAI+MKTkMElmKwFizBOVGPXkvbdS67pun8kb1epoN/HzKvW0X5/V/KatEcI0eJkn0uo6GuiYOzxi0YQGOaTqcxmhySiP0WLpVVNXlOWoTwjGcNMsEYdObjGWre8/Kpq8AJcBB1bjgSAu0SkyIxcYBHcwPlpSryfOYl81gb6KDQxrEejqXkRYC1Ooe+zrFw5EpjVxmR98qJxn4dYSN34Hg071xWgwSyr6joN/S3Vr4Py7c9RifHKvZdxoGpaPrWowReb3XsW+8rtx5hL/XOG2L0Fg3cGjT/gf0vCpiCHpBWLYQf+7KNr1IgKwie3dJmmIxP+wiYwsBCEyG37Q1ra+LV/KQbOfplltAvAG+PS3M9hyCH3JKT4Qa7UBFg0ZGeFLEkVtJn5WybsS9ehr520ui2clYKCmTs4L/lld5IpXFb3/G8Gw6gv1STUmkn+CvO9cMkRDS5gqqvBmoNIeEHdjJXBa2U4k9fWHTTQJprv3TWr3cDYC1Zx/ztbh9Zx/WlCThB8tAcSSbMhI1BQPHGBwEAjelo7XbJmjJUmC98ljdPvdkqdX85xp27ZkQGlV3/R3CVCsxEalHebzwzfVQMopCXUvZRx41ivpeRL3Gp8zPLvnbJt0f7b49KhMM4vrA8Y2PuP4f+U/OTsYuz7OIMPBa5cQNnqO1IIPaXVPCkzpMLrWVeQx5TzF3I1Y8WLVzYrqkNhRpT+2Hvi7wF50ID/zc5r6siA1hSgxZMLet44RsphN9ygaPZxcuUDwVJ+ssvSFB2QQnXZySdhXw1Cagotu4qofmJanfgxUC4M8/aPoE0FDLUGccHMfweJR2+z/Rh2hMEYVpS3Ky5ibTksIyQwti1Fd/+Ta2AETt4NYSorsOQDMo96hsK19uBYMDVLnuJ84h4sgfg3J47NVtN/PsrJZGCBucxTC8kmqrfrmMGAe0JtIH5nkY40o8qY+ktvnit+AW5txDBYNSaHx0QQuI8AIhR97zR2y7/8UM15TmIyQwAEJv/aEZEP/f7XbeAFTgCRJZferNicUMPqaGYpQpbQJeOifWeZCX/Y7fU2yMh08TOUgF3PAlNdBRIGYbOjeZE5QhzhomLjnQCYDuyS1gJBzmGeig4jqht13jT2YaasCr1d/58IcxLykulgdif1Pq0F9biDVAqCFMWZPK3ZM5AChMkW8n5TSIywXxlf8pCc7fTs3qK/CNF8HcUhPge5W64hNCtKuRq/Ib8gwJY1HPdrOxW0IWaFwtNKAIqMZIvKog+oxpdVPrngZik0ZEZYHvxjguNGYQMZKB/WPHXeXvxt4GGmXkwjYnofHW3ipdk6fB6kd2PuZC3gcuRXrEYNhJk1SJJP4l0hZw7P7V5EGKSEJUTleXDZmIS9vR0MecvyhQJP3qRzJ3LjpI4pOXN8Dcmf+XubBC0LVi2tGN/uw1vR22aAEBmFxCx1xnKlTrXtZNBXr7otjk2RhTzTEOZ/KJwQppskjpqhcnRlbR7UAgDtKGpGSBgJ6VhzCIlbY1X4FdkjjAhVw8+dPZCl5+v1OUz0sW0aTjEkVoZq+ktxfyMcfJjP2Pfkt26wquOYelFO6jmEf0MYO/YRYQbe5bFBVo/trlz2xVVX8LZH1aAmeavdNI2Phox8wvtISHHqJPQ+Qz1GwC+Etqj9AZzim20bwlrJJQZ2hldbnBsH0URLkvxDEhpsESSiYDgNTqR1LCTtIpaU6u4YVWmYSoDbeYYb58K1qE7XhG8CZBqysv/dW2Z45dqbsr0UGjMbU3moBfpje3WqUr+h6AouxnPwchp0lrgxxJkZRi0bYpj8cboqDe34e3sRBStlqztKqcKLSErKuBq2zmvBN//Qehl9YHr5TUK1pVFdsXoeMqbTwMQUkEZfu8peTfrUXiF+zbXcDK75FxNF0nefzQ3m6kOIf2RVf5A9arSMpxCv2ZxHdSU6wZXKdmkDXSrzCMOMz//xJmI+pzVYga6T7siW6wMajU/lO/KyDZuvrynhTTbdNT1NqOAsgyc66ltMCToDm/UKb2GgyaFBBWLL2BnSU74f3Jl1OJ6RvfahFzrJsZpnyOTjBBCm4wB6VM6OQNLYJeIZyT0egarzBOlVKMIWCxrwGMtIMqz6EdvCAsT6qEUhCrWKZpy2hgKUdmTolg0dRNdi82xl4pvUA8ZG8IixoTpGxcl9hR6hD46AFIrPhEHN52PIo3KrRrBvgWG+TeYrJh9TVIGOuVSLc5ZGBrxZx/Zhwr8VeTjy5lk7jmGoDkHCHVKJqs/orzHLfNrIFtcfjoGPVELGQUqw4xH7x37qwSWX5wWQWGX6iyiem8bnF88BPTg0BJrU5VbVFAU6ik80zStSgTxY+Sn578Oj5BMl0vrm96D2FeR0Kda0FyT8h/mBddmywYWdKpjnNn7lGvzVKbF2Baqu7Qyyhra32xTtH6FuXumNUGDbVR1kUD5oGa3TFJgwujDpWxGEIsFR2H8wMGFoeCwFTxkRY/0CFzrjc8/bZRLgQAArow6dpdXPFRz0YdGxpdaRuQSe+iH3SFNFdUY7Im9lgqiYBwhjjxKd1RfCjbwVEDDRTIbpmkZx87E1VxoEn3cHjQDO/DRhe0uhNEjU0zGoQRMGUkj1QJPPbH8BFP3u94mLGnkhzHo/sqryhKBrNLO9NNRGpzPlkVluQBLg4LcOc4+EQ1yjC+pDJav2o7Y8ZxUgO29hhLrBd2djWJlh+4yCp+wl9fPOw8Yd5dMqP6YBH3UnWTQ4JDv5UGWgq0CkRcTI43AQ4nqN4huTk0Us04L1fINBQPYJIBoql5QHVs2RnmMEykdfOgdhyLkDa9yIe8NYkSdzHkpE+LlLlDIpHzRoMBYqEshBOS9pINTf1wD9eEWUKdMR+xD8ciF83jgQrSTC1jBM/kqEiNckgArpmCrPqBz/Yws6BvDY2JzisvXmzetz70fOJzNwiRseY8jwK2Q9zBfuxKhRrGjT1cGEJKTni8FjSDTGHwRftoj1TyXiQ9kTuUXa9BnBDLUALxcF4MQ9Juiz7hOwJutbKGcfDwmQxvz0pM1RBgAw+hBdiyaqR1pIvlCqFQKrrwovI/7+KD0f2vqUhU3MtXlhATrNFNuPmIvFjFNvWrFC8ZGQi42IDG2RRY2m5MsTafnYU86/uRw86X0ixwOsKLVN+ljXtjeC/aWeCGycF0okWloETd8jOI+qDLkDR5kK2QajsvI8VOI+4OPixLCxKDPPDRj8BXvjh132j+4DVjV73uOZ7Dr7gcvQVH7QeeANkiboGzQSfDBwx9h3R1g+dq9r24K+CCGVkuTJBnQBtPlYzLRTTgXJ8x01IqdJxzeL/AMriemLv2HTHffFPRmWOCc84YhZHov6vx6b5D+m77M2r7ScjLC0+1kzhNLO8f1pHADhQCXHWqt7L3Ku4B+d65in0zl3I0qtl8ZkHlJeRiVLrfp9IMx1XShvgQ4A1AxwfC+DVYJP99xsz2LOJFg1ijG9YD/eQha16YfFEyXAyEFHRAmY26zsb2mIwxRUHxZfEnUOJv6KbIuMOK5fsgxXNxjjo33QeW4TO7M5whi/tLE9GDaxlP+4V2jfsKQQw/jQ9xShhLX6Fc819HEgzvJ8ZcI6/tM7mncW+QQqAEEiJCyV0+MAeu0ZOPj8ff8M6fAYZXLYUgPn92uk41RYPo+GSqWgc1PZhAx7V3ndoHCjUd5vzFZJsM1blniERUpC6i1vFySetSjoICUpjEiNHMaJGtVWHQ+t4J6T2D2ChasJkB94yQUhSXzcEgCimsMqwT0iq2zO9B2H56oJj6jfA0YmPrAkEuB39p/SDO1oNdxisGy4Bd2bU3CDuY3d+8brUd/stq+VKww8gToYdSuYkIzLN58YG6jbrbwG9ze1uzc4yOS0AUe30gODWshu3fLgqWGi+bsYFcfcQqPK8hMQk6HYXEvxNAOUW5GuN2t8q6+8/+QQyMjrPqW434hCnU8Vg/1/n8pWnFNJEOHet0ReCQbY2YVwsydNFlr4XBguF9VFm0OJMTxLoB3Z/sTPj0/9zkz3rz0hRU1G9IlVjrLnlZBSFFOja45c7fG9F57I7TM/sVWN9wJYHmRRUt4epduIpYP3A7QKxoYPhDqI+cqxS2W7IDwHu3Fp6SP3MawvE7ABuZAG9qNs3WRMc3B6ZFe96Im3W5ibAqbz3zT8ZkKrXEUhy+SPYKFucFh5aYz+m6hoq4r80vE+drV72hCEaPhmKVrqg/Hz64dbfjftDJWvUZb5XSbPv8fUgt/qcF6SUzbmGXue3UA7s4Qzjzo4X21aq40GeXtp9HME/6O1JFotxWo5IuUdkbaovfcNUR/aAEQ9eRv2ZWkM/fgSl/DZcpKoSHtg4Q8F7QdnzgR9sUf9RKwDR61S+/7YNcq8MUa9oqFH+qiR++8/oCFiMc6l9BPrFA+i9a1M6tJoGb18IIhHHU7ZImskTo9vsn0GYHCERVpITtr2vOjgrWqB3pKe4YDD3k6o5s/P1TVixmE2I63sTNMpKBZ1+CJ5i5hwdCka7sHDMgjxeQi2j+W5zPz8INLrx8lzFQlZYFs+p1k4YLTniGljXq7CVeclBM/kdd0Lj5Bzgwpxag09NkZY6SGP56nJqqpVW2SIoF4e4WAr1qlaZhRnp6zNk7OvfKnO3iVCZHg4tu3ZrV8qEfXyLFFPS1EoovP8632Qh6REy+kkN0P6EJuCFj72V8aDHkQ+Q8zMyBw9D3b6cbq9c7RS4T86UGx/+7lv7tIExnJgJaJx88hEQHWoXhhBe0iwxkcMYZ+5C/VUZgUD5lzwo4pk62LGtUM8CM5DyC6uXFuXyq+pw3adQxTD/I0RZS6N2R1GSDt7WtW3N5OVQeoBbXfwYe+uWBhlemEHWhdIcSJEdO1a/jg3+WlB/sh8OVNsbKwDUEyDLtR8dQALcK42sO/wks409YFsxAjTZE29nSp/XIoc/FJT3EIfobQ1kOU6h0mAXWAznrgULYMiVJp8neXVx5Id2JEwD/ax2vNFanDhghNbcXKgPg0+lK0K6D/gNKi47BvdVJwW4sRzD1jfQS5LFp3lV42ZgqzUyHnpV40T0/aXKdOCKDQ4WJaT/Q8sNleWw7VR4+vsfW1TAuZ822HozrMMGcN/WnLRsCcIKARmchb9Q3zQAAAAefRv3eKX8nCgMHPXXKpB78kBHjO7CgP5RY8zO2ssvxzD0Iq2YQ9r3ixp9Q3jMujj+1YgbYMys4wH+TlzliYfRmsfZFDPBAYjjfowsCbMDBhsFiPX1uBme635eFfIhnlReQ1NztwhPkpybb/Slmkjm4pZ7fXPpnl/DyeXzUoxAasUvLIxDJ82+y9TgDR4FPgaxqpxJk8jl4OvuDdXqZAf9I5NyWI1fQuTPvMWllh8m6wxx8Sw+Od+nN5Mr7K2NRFJOqSRyqWOP4QQ7gUlyF9b2KxY2W7lm+UxlEsRWFVTOqrx8ZCuchnCYtpRHBagoh160qWVFt1rL+dzJj1AUTZU748Psx7IKZcDbPX1z/jIDyoRySh5HBlkMcdNCMFXP1Ycgtzs36SKme5HZDBZEKZLCz1c8i4YfqG4RiG4LSIa3tjHdiYpuBYfzGCnYnPMCjz7IEeg0gxmz/rkxwfYUXjEVxl8Ipfz2s/3pQgvBpHZcWZjtgF1lcpOy4AOTSj9Qbncvb5UeebANCuGh2IF9nIyY/8vj9TcSD3TlETDWgJvvdfUqVrTULZhK3ECyBVcydzUEu5xlVLbHjtVvjFoeFZ9l8m93YhZPiXfvw2zSsMB6o7Rsf315dVempBHnAtXePp6HF9/nkBqQsbghFiy3Zl5v3vhuKCq6VYr2V1e7rucutJFTaDHOgmi/UZoL6wY/akGFopSP58aOsgdDfCYCDkOjE0aN66/1nfKR05DsjRhjJlswuL0uKNnQhOgsvBTqR5KlCs5pl4YRXyut272wHuBQ+QJKwhNWqEkm1o3GcWdmAt0f7ZAXHHhG9ZKfH+46L4LWyJfqxhCtvwTam2a6Q0Uicgvj/q4R4ejjkMN7AyB1CoyHo0OJDE9FBYll/CbtBBpPwoZnK8wDlG3mIvZiZ5xuFkrQE6poi8ADzipao6TI8Z8UY3l8GbHX53UneIVPjmHSaTnuZC5apzQ4QqWRH0T4U9aAJ8bXtBjggHIC2wZ3RC1WlIFRPeIEY0/ci9N8QKt3n2xvcQDXr6XqOR5J062MyEtndnyQikuSrEwoSth9FoV8DfXtBOsBRbKFWsPt6JkhAG/MRc2qVOUSaLn3LjSp2I6NM5W37CaSFQd5wjjcMqn2yvoq2rtVJspzYmjAtkA8jZ/CEIkIawKE7+YmyZBSnXHFnSh6ZuGaQkL1baIJ1oe1CE60FaP/naBAWhtgE6y30hEIpV35OvgawHANxIsktUTb6LXIE8qbgHj3qS4ip7ptPDnFH6w7Zga5kcqlv+t1Qc1sg5o+PxsAAA0oDvNuSQH6I95Z1CGwXc/m0cGumBhQAvkguHjiKjw16WkfZOcnF3Yuz2Hrd+X81hk/7bZfL6TBXkZl363MbAJM2GoaNVNVoztDvxgMflURVUJzPIbL8FWwB37VfgkB0/eYEuH0Jt4gKLmCr4zAVVT3kYirF9DH2XKwHfFnEbX40oxfF54/QnlmH8sXVrZ9qRkdMvhTuPOf6KwWwVW6JyNpwpsbsWvzuwnsKdoiU2hKwxTxMAqPI97B/WSoeL3f+SVJ7B1WYd2NM+8huSa+vvRydH1AfJEnDkFTVvRLNtrpvouC1tRorND11okM6+qH0oQ42hWsFUTEYMB3E/OXbWq/8Ze4fh2JXYRAMbhdKXj2VjdhkH6H3v6wUKNEQJKGKEXMEtiZ8mdvTh8r9TUC4VNGGzfZhkFB/K7kWeHpd2ClysgXK/gQQIzdIRgc5KD2dreOkMe/+TRJsv5+hLZJaIaWfsAax64aLhq7JTG1LM8yGcOEwf1buNQIDTSFSTbpOlE7FwReX3D5JYqmEWwqHZIi/XpFkI8Ue/Y3l0fN/SJVycdVR0B7raS98xOFpBtB3JePwNInHk7avwqqgi3T4BQKpBUNZ2fYWxAUFimRwqeCgyKhsUWXoKarT45BNb3Kz02d4wDJYVfB1nPXCco4wAnIlyx8+B4rcIqobbxGVWpnUBkB5P7MtxT35dg+nQa5QaPOENE792x/bgI7U5NDw08q1CAnEU/BVmx/3lf3mqDrNTyKWdmAXSRp8MhzHnSFCcXpxCWDL3XeFlV48aANbbv0aQgXqsUNTrfwjjaOLGhS20yLRjGaUF2n+tAY1ocln9esOGoMix544+Um86sKNbPNwnoKBbjWAg9pGvmf8ki/SeC+wZPyaxL5k+3UbdUSTIm2N8PEWdYb5jobupLn5i2ALVvCc0oOWgqBn+ZQ03XBIef6PuNvSGCwVhyMrtHMdTVCZXPaCIBtYyshvSGIrE4e7dkQir5MYEQM7Ukfhb+igtm2s7jTQa9WQtDW8n6LloJc8AC6eEc4EyCfrl6RIwbW0PkjkLpB/4VKskNyqzjxfuA6yYw+y6qSL+2uB/pSqJ1jC1UbB/6JjGWjg9MbbTlfkTd6/Jygyaah8zfnoc6v0WD1LC8rk7Ov+ztZPHNS6EQwAIe6ZXCOEJEyJQEo+YZAJ8UgSOwLVTrfEM1K+AykSOLyKebAx9b25Ve0guJgAMcqz7E2aJEwsJ3tfZ46LKpR2VQoQnPRtnXdmr/JtLwEgPrVr5IoPookBKWh1Tnw6AEwkG2w1cx2EE20HrWyYvvCiK11PfW21t2F100uP8pMXw5IpI82u0HtpBgOwn27y7oCwez2NAZMGpFG+Uwc7BzjHWq5u8M8Ek26G8H3vX9PbXHHy0w2EZJXyNDa8Y/8HsHzCNTZW0E4V/ej5ieVkwyojTjrwVOH/HiC8aXliLTuW4zedJNjkpPVIu0IwoNUvlH56+VCyl4vIZmyV38cq5J8wCBshA548fFlF0CeihJA27Gwy5vMW4TiDAg9SbsiUvhkhh6F6bbBTQK7Jy0qU53BAcRgDc7chUNspuK9+9hOjYJ6FwXVZqJa8D5pm7+KbfSV3Z8WIHmR1n4xnRubeIhxmKEDdUDyA0wbL6ql0mcoGQlOFVotXDSAiBWR7L4L38X5VQzuM/s8wB4lzLI5mCmb7uyM4Byf2powlodwO1NXZiL/CYVTziDfCdtT7pW3/tA3v953K8GgCklCJD5DoWKhF17h8fbeANCPUT10CXaz7yJLfBRT1PxsBOQvncWy5RdJF8WYwpGItG5uoEBQl9WdPdyuoEPZkjvqDNr9TLD5N4NGeF1QL3Mm5owwyv/qHQTEsgwe6xylyzKARxiGKT2gfEIxGQj1nbpXiRpQF3kri/frB+/xcoEmrVO/Yn1MNGNSqIdWF0Oz0F/LLrTzsaOojnpql2veqD1cZv10/bFguODE1V4Z8oRFsVErZfli8s8I+1Gph3H7oH0nXr8aVSirZr49WKw1bMA9pSPaKLhNYYyh/YoTdTLRJCuhJdm9VLW+83D2ZvZkF273MfCp6okF/j6cXXHE/sVW4+SPfFP0huJbCPnl+nuxBVl6sfmHbkAuNexVRg5NcGHnCDrnXzV+Y2uqUOw/Fp0CXuHjbI5KAe7ZDYAK+4v4OYE3pBoah5D0r4WdI+P+Abb3ZLwpvQz8NUa+Sb6eNwKjmMKzG6Gyzy+wDCc4mkOHpNdER1vkQMMrODHqru99OjJZJg5YQuW4u5wgmrQ9EekZMnNfo1ysVn61lUS/h0VTbWZyr2SWxsu93AjLtzGKpI6m+eFvaMZI4LzEI90RHihnvXG4rf7sWYbscAtnwHmzQbLxfvaDmvFcJoE/4MrFPAkhlH8iB6ac3TRVqjr3kzld0b1YfN5zxFMAnKupqvYqkzlVHy8RzcKzX5o7kT9IXnhEHYl7vu2OCVE7lq66VqHEDwfNw9X5X7DztvaGkpTGCUjpPmGX6lpiy8tWDxpaF3xWY2bwMC/Zjmbt1HV7NxjdtQ4TMEUQr3o+wg2t2Imu4HyYAAfyxyscw2M7jT7btsOfA8zfRP6AFAuOIBDoDdAndzYTCZifST3PE1B+Pt/Ije+vKxTD/R+2RmDUKx2MQvDj31P2S3/d5Lg0ZwuHw7viNOReh9FJ7epjUnrk3hFFd8VuXs0XsidT8TDJfWbwHl5MVlK1a1+TIaH5EWk7trDqUTdWQyUeK5j2o3ZcWs3lf3b/PKYPyTSIZ+ldyf023jrrB5oQplM5nQBP8QWI9jvmUdy2Z+xj4XYztaZVMtXTeFX3+o662bhM2SvjMp3FniAg035gxOK0TC4Dp8LtZWyuZ0D82/4O3vik+Fd5Q9k7IcsvN+3DVwXFDcwq+ADCd9DR/aOsE9cgNvRlzMvPfMAy4dYn2P6yjSJUz9URp8hf9U8QYa+M4Cesd7NMutxLOAwrwztmCIzzWx2MWUYuYXS1QRu9iX7xSM3BYmgS9cNI0ZcbFDwLv4zG7YJxk5alNKG5AHtBY5qmXiJVS4Mo3ujmFUDQon+yNVVEdz+fXY6rFmXAmV7Jfn4152YPEWBUY36td+3RlWGnmJwjx0DX3orWXWKVeUOEKsKfw6gGTUpexLtDoKY+1Q5+Qzz3Vvf1u4RBYPhG4dP3I7KNBiDjha3AStPPtlsqJVou70zg7n1BkyOMZtfsYCPLIl4PZprmwpW+OykwNBkBt/YGYXvGbKI2KOz+7xxhGFLL7EKVUNfbYwOKrCqcR7+35nYmEvxSpdtCG8yErJBi6jU08ZbQqNHLu+BM/CoOg+BAo41k4HpAnJyNkLv9MaF4IPzEdVin1Jfq2ORcZvTi9CL8cPH3s8IthbqfqNiXu92ZT81/oGcvoZqaUeR09H37+xbTQVI3dM7ophkUCGn3kfOKouobYzdT9DutnYkG8c6gl3NYNHPgnx0p75HZx0nyzU3/R7lTZHTA5EOAO/nk7/V0EKbtOuFvovFuYHFLAm6+rZyqzRoGqJFAXVylbQw3y9iGksVyxJD8matEYOIeIcjZB3kgWhxY39bjtlBVKHDNoDTwbBKQOb55mYZAxkAsa6U3eOIRtWl1B0JHUZuWKbCO8gJpP8cNZk7OIbpCIIVcbcVZq4YoI6vvt98mBgAwU+DIAFV5UIUiMunxToPmG1jdn4pFUJxPWAWI7XeOkoXj3m7B0hHSsvkEXwIoH5e32yRDjwM25f1S5iacOFzVQohf9U6kFScpe9emrRK+8shRoKqjWeaiYixR534KXXxHzANTvJWr+RxI8iyiHEVm9Ogx55c8aUpNNX+/MQG4P9zYKvHvH+vyViPozj/q08DZt5c86CCi3lWFYTtpOki9FNTYl8XQdHyrOfrLCmjCkJ8s9oClTQLAgSysehzZ3PigJEJm5GVnUa1UKHZqClTQ+0I81V1Y0POluNRMHYIwmtDrTzx6gYv0bH92LSeudngFjFscyTOiINfp+vt2JaeOsWOoSBy4AWEGrt9cWS4HfEV/qEM4vTrH0v2QfoywuPdRCLFBECgtcsF3BYNW15JdJyvaeugGzZqgWKxnMLV+Pl3DJ8hfYr7HfWza3pdEhA5Peq7tEh5XMptCu/RBbQomhbYJjYtrYbKuDUalJ+qIQIdn0nhOBqNnI8R08A6VcgWxWwSQ4VyAP+IsO4gOaj4z8ee9405xKZFFObWvHTeGRKc3undrTEQFE/yEEC1XPhpUBuGX/kv83Mz8b5c7oIxM8e8NYZk3kVeTqQGt/1S9Ehhz9+5F7Pol8b1+lMtUS3B6A2LqHQIZTvdYPejgj5mrYAbz5fRQm33cGZjEiZDGmHKva3/YNxAbqECeF4HLfCkRIZmbv9SRVar6RZ9uo8b6ocjkln7gLVlOLLK7cb1fw5BKbwEz6l5u3/tbVpZrYGtniE/Sw+swd5XvVHLU05Z1QD6YXUC5j4xmxqS4KMFhG6elTJLKa50wEllUVg4C9WVfYUaR3uQ+C+YEi5HgoYMgq24xWS4vC719+DWKHcD3MUKGUrarkMbIHeZUpb7w55S5gMxlHgRI37nrO/h83/zBkpv0Zplns9+y7TTdPo4Jh96XvhqGpfWiDVcyFw8Qvj3wRRX+INq7Zp/z0QX9CimZmWWzQFIMyJpA5batOMkUqFfTRuxiDotlRyb61T9UVIXzFrHQiLDmExDE0gzuY17hBrehDxg2VMtvrE7tneuoRKb8dDQ8wDYJrUf0TPa816n1LIL9Q0yVOdCQfYC5TsGlL+5gAL1spd6tAzNj2fxt9xfe4XFjYe8x8Ml+vfWrHzz11zfVQ3HOoR7ziYIu/59wa+y9QM3ZI/QtNEDPaXVfvhPthiWnq0V+VAsBKGpcGKa9J/VHQbap79PdLQ9EWxi2dEgmXQzynnd6ZI9VNtjJQwJSKJ04yLmPL43zUOdKxlgFJzvJJxCHaQhp9XyGXiV6LYmlzyzgd4XZISGs2qRjOEXTFIjazsYZuFyZs4MZ9oYPcwsdXysY6DRXzkBh653ISJwzLbfio4Hi6IHuunVQQoOjdF9HtdtPawZLx5YYh2XErpfDyCf0iwqSZ/3YJSe79aOd2cXYUIlXP5dToHPtBo/yBT9fRJoLxCXLlqI8USg1Cendirys8qIpLItuL1qn49+NV/6Dfmt4fQPHR6KfprQDF/oEdKXNOTeHR+Xu7SI/6JqlsZU8talyFpRyaoPkJKBBEwusmGzifM6oqXUhTs132Fi7a8LaPETgRtSlHDku+7EeSeucE2rQ80SPbiv3Tki8bJep0Ka/rpTyH2twTMgOXrFvrNxANLLZxwDHfq7oEKXfX6UC21hSiA3jS733a2kVy1Ni0I2QiDN3bauaFhGEVGwnmjc6qU7MeXTwrKPY4cZKjXLsx2jFLpjqmjRMV6QiTMsQKZHFhJiPz0u5SHvmrp+1e3hgYZ3pNS5fTswUQNsPQR2ToK8d9c2VJTVyxcTGE1zgedkb/y7fkU3g2jjYuLA2Yg0+Zc6Zzg+0dwj/L2y9txF+IhBt1KUa4inETCNdKoVAnT97pJbTJKqP84sQ+GO8jUZBTZVtKjvCGagXEqEUKU5W4keaR80y1AshjBiXM7/N6lhh94gyKZlZECuAx5YXQI+KJ72hkwy1Xe/RwAvVHbGwTOsOu6v5KhCY+xSqTQeqvaa+AmGh6Y88iXVQOYO6A/I78YsFTcQ5avPA2Brj0d9DKWqKYrbnTHJw8GNf9gbqe1GR4Ox27/8nkb8t6eEzg20pBGKmkx9zfYARL2OojEkRqcP4XGTr49v8dw/tCgArzgBPz+Iv7rhCd9ffkN554PfAAbRFv51ofXF8jGvR4SL6Ru04rxFy3XOfmfDw/3YMbL7eFZ4WFSmxgQp2YJJSecLzat5saGNadi5CYgqBTm/bMFUWExDBVsoKC5Xyyl7IttOfdqCzDBiXZeJD/jIjiV/rUw+8r10bMOkZBlsCKL410ZM3m4MC5NN5JEDAinidY/lrmayM0wqOguZjB/c7THcY15SJwJHnImgZ7LDCkSsdlxHmZ+6tgU3kzCWPm6nfwAmokjXy1L9iBuuwMlpuHnMSE5vTEtJTJgOm/R4mmYTxF7G57ThDExzDhuPp2w1s+92o32IV3dQPhcrGCWb6YmdPbaVORUQJ0ikR8OlwunlR9VnlxkmhJvUlI6TNIueKuoUJqDEX2C/cEPdB5DcNVFb5pLYgM4iP9mlbKQQGFKd9a4BJrot+z0Q+ZX8kjVNIzzBuVSNfsGMTeLauyDUQKkefujEwvY1Ti74VQxciQ6X11XHsTSTEqYav9zRLaQS5edg23VpFF/XfLbRz3MXPHo/P1rGBAbHlvwYResSm9t4fiILBDEKBV8zmYFtsXbmkdcnVNdOdjT1Q87+JAyD5XLMX1aNfaSyZWjWmcsGdUq2OHxxVfOH88r7v8+OCmZdkRpLf+qrg068tfuy1uGPbDtfovgh28sCDdr9Dl0MvWCOaasLXBtjpR+7MCBvwTgIjTjZ5ZIbj++d0adZmiowJcya17DOTb6Qq9WgI/Z12G6l/ndwiLxmUwrOfLjafT8aYUGRqMiPtJHzPOkUyCEpdWnHaqWvBP1wHPeoJX35+8TkiKeBPTOjPfgOFCM3glyPdtSknzR4b0XW+NtrIjcIebig9fy1MLKYgJtbgiTGCYcz8w/9+BK53dFI0tAT1Oaa1oonKHhBMWppgWHii22PtgT6wrmi5EuIZbr9tBEbTevFfCv3IhNwOpDyOmBeVAnOqwZ2MizM7BtMzK8jhlmdZfewcat5nAcQq22W7EWZ0MzvC7t33SK6r5sHtlodHYReWBiOC0lLza3la8hyYlffAly+Okj+musWloUKOBC+ZbrKERNwvQ8gX7k3sxmG0WdduLRdZ1KiL90fwXwAEWb7H4Eb8imbcAloDwI512zEhNr7zI++VZUcXk2yqsq/9AvoCHOKKNKx9EjDfu68qg3t85FqIwywiK585+U6PnabwCElhXLXab8vno/Po8mZ/In0Tw7aG9fRL36GkWUS8mzijd/kzAoCg4/AaG/MGDYVgDwtcOe9BBZAupfHVi0kTwSNqC2HetAdmUV2MXDMrynKk6uZqjhrC1bZvotpz3pMjsmVRwDHYRvNbNKhbKOk2FJQJA1p859GcG6LirgGKl71kGz3csXMUYRswfZ1yCfXBOEL2z28Ra3X/RKwGQfUo4fxDzlIyyq63uMiZ3g/A99KKrLFwAmOIAkEhuBD7QuRPsb9I6yw+9h7QqS1IGZQLTZPYwmoH1iE7/eXUUE3xYK0lXzGoVWxEjRv2c4B5R7RWdLW54dEB/IYQGVDFMiVXJQVBYU8rFnXG3krTCea9ZEgK3Bz008/DT1z1wVisGk2pgqMVeqre0SE9uDuN4ke/i+X/Q1ItMQGPUPEHzQ0133qNIZ0+Eu0wqhmYBaiejwhUTA+7bVNsxklTCnMjsglq/wE/LYhFZzPaYpgmkvlKxZBuRvXMh+ZyMBVy3spYjZmmAg5K1btxJGfbY9BHCXtwvyggyklG0P+Z/e6RIvs6RU33aIm91h1iX+/N3g1uYlr2CYhZkXKJYWABBfG4CLtgeHqEgbqh8csAMOXw4Z8q8DR00sBUPWUUgUu7qnwZsx1RVxGPqFo3qmFixKTCgRv/aIVozzDqa3SSmBO3F9VjRWbLiowAydNM7e+UggB9R3Vym+4LdMqXcHCVnY/8uCQsSZekrkma9Vi68VSIGPWxRa2ICszmpcAgDVscIyvz2WeRDRdBrHwb5O/t171nRRsKcUSvprPzQGyaLHAHUzEcv9rnt3Biz4E/tMF6iNHEcfry1ubxPr1qbX06nUMWdmHretOFA66b1hwF+I1ux4zZId3foHeR4n9X88o9EM9b7ThR5b9YYhqHXco4q/32Zqch+sknJOUi+r3cxeYFKlb8a0ufDNmytbbDFSEmZ7saLr9bWtotvC09XmSKQJrHpeGpjpXIabs5tddHWMxnVc592gZFEtmrFBP2yLxKI4RBBjD80PonXWpYoiR8JEXGFGnBCiNRVBOYNvVBZv7ZmLzpIt4k2mV81GbUwQPt83H3S6HZ6k1BC9vc5xvy2+bXGKTobh+kqEMeIScEx4mLHjVbq8p7VRqdbBR9XoDJKEQQjW+VEMfkMkMPd1XhRh9BNvR50yzCehdyVAsLQqL0qMdwYPy77lA05axLox/tg6h0Yv4Vx+/7+1rynwRmreb8mgASz9000ooAM63L3jQQhhPDs+nS7sYsOXB9u2lptIV9dmUxK/L1HLruSjG4puwC3nTZxb2j0S9bbED+gzFzoTKDtpeuOA8wFL5tC/WS4UG2z9HRSE/5pC6QGIFkq+wjonxQvNHcTRfrOxXdX8SeMck1wocRbYfyrV7aq40MkzVySOkyzh8IYf8squeHpB4bxQl+pHaop3Hr1/PAmTHUXURoGPREzoYHjm0ETyzDHHOQ1WIsXxpqsi5XOjST5VPPp53yNRYN7pAE/eyWsCqewD4Rjh/cwW7/VX/v/v1q/wdSdJ+pKvdFzoYGjSXQ+uCw869NhPmImlzDkL50c4rfqEdQ4BMazwO2SNsi+n6rf8nhNzRvf4S1sp9XyyeTyIOGq+glAGm6ykvPS9MFkjLzAQJeHY37e1ZUBsYtr3QF4cdBJTkHbhHPf3d9gawaTueUfbRDEiwuC8XnDIO5OHLvgq84kdIoUwjVwkjpKGlC7McA86JClOPJZNg6oet0k7jg/c4N6ms4Z7V9DdQ4mv+YqX+CNiR6u46sgoDmarG98Hma70yIh0z0ZgRTKFeKGHlFmJZW8IyE470elo0ggZomw22KGrmbwgm2YvG0HDulj8I/wYCgB6YCkZMYMqr2mRqoGxuqoGsKJpvMwAM9QH8d2RjfOYl37sLeHeCfUkvAmjqrcrZSf0iATP614VHkWPJlGiWNoOx3V78Z3zLWNOymZVUZIItECwjPy9t/tsQjQOjDcQzXQRWX6y6WW0n8fGWJwPPGYjoqO/hQXTdY3xK8ckTcjQfXW1nsVR+ix4LAkAHgem2ZjMrCNzvE4YfSL5gRPCHXCl39QFN1YBdhT2qXIlA3Fild49Pogb/6mzLw39nMoDSYvFPNxv/0YalC54x/yRKArXHtOPiIYRWQCTH7/HCYkDcC/K5iQrNLjPTDs0/pAwI6qfKSrcDom3rUWBUlA3rMt1f2mgxXVwMhq8QJGywNkEMv4ULK66n7o0S/0RbC97pDsb1SBDY+C2rNepJQ5LoTeMH2zW4Skg2JrsYIBo6Da4+n1uO0IcODLNW33two+mYLL6d0VtMz1I7ftZls/L2S84jR+b2HVAJJ2knh7/4Rtakz2eCWIqBOS1F9XDfLcp3S01FHvAmxgBr1dUiTdqHxc8qPu/2/1cx4J82sVqZDKJErSNlHUT+7qKXsfoIX10AzJe5SdsMxofzcAL34FUXdrh2ZPt++n98oXADo07/IBN5jefm5LnHm3qzBfumXNx6eIcfiHMQHIC9PZnZNx0PGYFNyV3gG/1rRn2O69ieSOngc5NUxtegWuXtgXgWwDZNDg43rP3LqCZRrMd7IphSOJ/U128XDE6VuShMH0znjAHbrTt61EfIe1e4AC+9QUQP6hFGSG8I/nbFRtWx+rpQlck/2n1ykaRPntaN8MJAMN2zW+U8K4ufcx33Y+bXa+JD821vu36Om7sSqmHb9/N3h9oYp7THyza+XB7K7mAHQJS+WCH2u4UZjLeN9QiRh2+vNzXV9CorKLuRKKi1bjUjLPrqoPlDnVQzK+wnT/PSf4zbC6AWctK+odx7naHBqDfBE1kBTytpiUozkTVh3hh424d7nGBoRnRqiOfkaHbDmkzMMxpElIp5CjUXBjviNdWGsHuAPElxzA+Q6IHx0RGcQntkl9S8EwZuVCX1CFZGb72Bd/vSN1hfBQ/mrBhloAtf/MspzwMJVS3B5C7OiMNv445k2bTfKwTqiQow6ssPST6x8nVKDZrVlFp3ygGBk3iZBZP1F2GTs1rbMJ8/MNxi0kw4wuVshl6mmX22S63+vhs58Z4djw6g4utQg+6lCKmxL9u+nEzyOuwGpxgT98E08jdtl1aCbcaB8Fe2Hk6MWT6AyiQX0GMZcQGcHlUlQj0YI3XQXFd2vu0OfJyd45iGLiOSgYyq8w2P+DvXr+fNZc+NBtaZwL3C/r55VYG+rLEW6cWAKwtg8vPDujbxZPTQQKFTBIos2ahbYXmYQtZ/juQVAuE2xptQ8Yb8Vxmw+8m0tCd3etttPLEBg+Ar0ZmsagYqU82rl2AsZhaX2DxD4l5tFJ2eJUqZwUDN5ewAuT6utai4Oc2EfyCBPg9Xya+gplQz1Mb1e7Zmtx9qwLQ3Ms7Nng5tHBwFpXKehVUxVywlcN35s8aICwTVJ822LgldWsNomhFpskYDl61OLRd99ngDCbyw9A3Uo+TQwl6U1n9CNfCXJpwKSm+Lbc1f16prRBMRwQglvXtKA8SnetEkAPT6dmHHHRlG8LjBqyR+KB63co5cHdeA4oa0spckiExy4QBxV5aJ/EA51NcMkkOEj3MpKAAGt4zCvIQ06LXTfsh5MPARvcvl8pAj/vBmu7auvxAilCSWtSHOW903imgTmmeegEQf38uPg/TiSzBGPfS7ao2Cfb+TPTUgNOBlhlbbBu6sXJxnZZWISbgQk1u4Ihx8mvIlys9N46x/lQsQP2rL2wmpw5MOus0A3kew0Jemj1PFAC7fxW8KkLAzLXbBZN7TixDBbuy+WV3wZ/QpkfAw//hHWhm23TvsHe53l0HVedpmvvus19yLxEruR+taIrrjBSaqzwMShx3C1oVUt2zkkvUOFcpuP5+ASi2y/x23sAPvFJf+OqMDopOXj6kUQi2Tr/rpy97BY7ZQxhnmrrV9YGbRI6CLhNNZ1NC72mMUYDflXC72sWsCy8t3e6BsRkwYbBA57Sz1YewgTaQwlR02OCsWmieo/VE0zARGsSRyfGj31OKttatRzdD7sWVSNONcc+0cjy1TXmP5XE+M8R+LxIUbMR0u8jBHXynlpJDUfX+H/7oYb67+o2HKa5myl5NytjdDt7vdmUP+5xnOAiBOUpxYCpxsiflJ5Xy+RP5ycLX+q4CfcFVMjGFqzi7PJDqlG4kaEmfqOltIlDD6jQteV9YQ4w2pSwNpuCUXUNm209M6zwz5HON729/rCECb3M9bs8t37Pgcfy8ISYRBqewmzD6NTohGOmsfQqAJ3A610tscAiG9CKGfXm8uWCtMSrG1BwzUUUrmMkySOejhiV7ounQARssP8PXEfrUHWyD+1b38P7Sy0/WcFb1C3JdyQ6YuPejt0t/qB0K9a7lsAV3hOuG+xHofE/VYccGZta0xIPh+keuKebbOAi95IfQdOMFVAfdup3T/yLuEfZEm+68NQO4lRdzppAs6RlfM+g2LGVm06/ny5TDHBE9B6dV14CtT1ROGhHiCN+yLvhD4p/h5F02PzWsKq59GKpDHIht4RFG9dguVO7E+GXAGcS6iMEMW29FwAvjt265sd/EpEXucUCTRhZmBT0GcFKFheMN2bZrqkAfiEYCoI93b3XRGVwrLHqOc9/dWYpVnZPy4rB+CLPe5DyYicvMybsK8jmxxM/dbdHhgrcKC4hLK8zDkOCadfH9SIEuGNwbTAjOqXH0Z8j/qpecebDnnW/RqtCaQxvKWhRtNIasp1wIXxLAsLZsFGzDVn2jJliA9L3nlgu6eJV3Db1ivN7DzsXAOVfVlDDnlkW3etpmrOSnpS192uHoU4cfW5pE4r/cNFqDMTPRna8r6OBwsgpsgFj8FFlS9mz1VuugZR8roAz+mvSUiImb/1DulDq9eHtjKajSSHxURdOURTur2bfFCrQRYq8z7/YR11O1PIYQfNu8NBvhewENH2iHKPIfd4FEJ5SqhGwwBJ0jrqlI2IaD1k/w37pgL2h8t1Bva+BULsnyukWV2gG/Ot1r2XpVyh0a00ESlE5eabhILNHP7WgMlA4/VOevSlbeC355+9I3oDRTin/xBaLO/hHkKPVnN8c8ZC++SiAEXjJhzcpssC7oOV4k4YvPEE6By6t4FnsEPSY/f4KM4bNLkcNlsgWHpnSZEVZHs4sY+2vk07WL5XhXxeFLkXR1ZleLmpD1pHLo7gZclqthOdMXpYo3qgeo17fKn+jrfxTXA4BN1hCc4PkUeGOXZPJDXh6rHHFOQRvWdecQUY0n8aDVLDn2iFhiUJCiAKsri8q4Knh/5S4jp0S+GTNHGOBO95d/BfsPvYK7mAnifEK2+aty+RflQJlBvBkErutG70HQZv+5yoEcWctg5ntxupcYMYcqkpRJ5nwZFpB6e7EJGYx8ZhP9iLnNPOLjk6Ntc4lk+y9RwtdelewQPrJDBSWVx/li+O0bZ6mxrvI3v27Z6BhtQ2XchEbY4QX2ztTpu71DBzqvg3Yz65G2rTbks+OMbG1gRz0mqxPmPsjlpd+3kOFKZ9YAR3AWf9SvFp6rEwkqOXWh+7wmL9b2HxqSfc7lJ56YB4IPoHZTG5qmK5LBNKgefNLnVEbHfUt0MfctH1dkmLrC6lLHT8drgg/n74Ygs/yhxcX0EXoH8rsPjxmBBshURhLZYNq71fBWkkoPaL4m8119ksZlSo6gMRv10PBcwiqkpBBhp8d7bBB+/EnE5CrEW0koYwjYJTQNys9J19DBa4YrIbnqLWcfAmbt7VNUCPauEFjM9So1dq57JyZi40HwYUGdpeDRqONLPSxnfDXiEGNiBNKi+XIQ1Xx9eRgg/GD7X51urWMoywcN1Jsw+J7Z3TKQI4h44QrdSZTPF946C4r01og4FFauEs4yjMmuErPFyimQn5YzNQsHX1TROkqGFraL8kHlWAmL/FVeaqioHDZgyXLuPo3GBEVDUqCup8jhEVCrQsFQ5Q5zUozZlh/heQek/cpak7x32ljwKO3o2SSigDnK4jV6eFgKI865gly1PRstJLygsup5vwBgtwfiWCCK2dlj6fFUSqWyeZlk+wV9syrvILZDXx9CbXcoHK9MfTwsZQSpq6UV/KQL6FTcXANJSTpEaU5qq3EUh9kgfHI4GJ0WOOvSiyTovbOHxusa+fFlJ/UjoGFHmNFkkHSiMQxiseddDRhW05WNFGMFV9Wa+DYNcyzNtFCfOj1gjR/CBOKFUOgkpofI/cApw0vPde8hILk/pfs1OzJGjx2j57vrol0szrainossUp1HNMKPvgZGnxvWNjnL1RpfHWcDypbBLRlZVV2Xma1IA/MmPu+pimkZEVeUfB0dHUNC6oXfISQpfEBZGx7A0cJy9vowQkyeyTBCIbakMKMJOARVwhxiAetwqK6LZeSg+A9vo27b2o3jyUyAbT4Tkr5u+2R85d+22F56iuobBBsEQE+Eh/+pM+fQZZ8UeKEV+dig9IkVV8z6czm/eW1lPhZ89yoLUUryoViIsqrSSUIXU/kFW7GvHNbMG3XLrG/BTounlArPr0cOkMLqEGSj6FbkV8GSvjGW5U4V+FZG4KXsMc57vg4Efbp8pZXBVdoa1eqKS0Upy+ns6/tDJaxSBJaMYbck+9tRkSUl8pvJRhr3hURJZSzER7fVKGiLBSC//NxEZBYjNCOiLk1LToX2C21DWTY7x5Vq7A8PZiDo4f8QNTvGCoO7WAjC/TEhGEsMnLPgcOnEF9b6i4Bva+PGhZ8csr6zMtnInFwoB2oF0Eu+nJ3Fpw4ex5/aDDylhGCLozQWCzhwqoGvf6EvkUAHc5uY3ndXqHCDE5w4RZ/q0NIi9aNc5VhCN5G0Yy/mBeXuXV12PrS5fTrggEltB3H4bGkkMT2Cmf2Nn7D7TbdlbaWOv5Dn0HxVBYMdUioH40JS3nZUFFkO1WnUcY1UQL/GmWbZ2iOu/piHoxNcxt09kt3jPP5F/ks1TbwzMBmFDrgBvz8B9sHIwQ+dG5hAT4YezOIux7t6trceht3ZAGQdh8h2b7GZcrmOD40yOCSr7UpVJKlG7Z3tU4Q8rrx1fae3wxKXpg5E3DamT8QmQtqg4A0V7qi5295BkNUKjhQisn9iHmKy9hVMNzwECT/LKiX2edgd3mMB+JPQOzrQnttflAu64Tpub9OiCegv+S4CDIxIQvrGP1ku759lXVvjRH2L5U3ywdGIvJPtpD37m4JwUWK0j8n/FP2tuOB3bFm+Sw+2RQ2LZAj/C/gSnKrI7YsTLnsZY5oYXgpWJt1YHWctzWiNLHUVLFVZErTnM2S4SHkv7134+cpTFq8tMmmhYWycXYNJJLqVwiLO128B3soBC+b4EqIJ9bVjQg1FTpY1/nNYI78UCrTJDVz8P6YxpBWkVfWRnlMqh3oSxCSJr8A0BtRQmC2NZxcsAgLFeJJG4EktIOgTCyhFCgRhpVP9j14t3lx9epu6FtG7KA4NrvUiDLIGMtLjgXEm+OTPeGDQVQdEUry93LcwI9u/bmtBwsQvWtvOH5lOUc/I2LCyDhn3uvLzjO+kjhnAOlp0sg3rC6vM+Y3/SzvNVBzFV/WVIWV4cmTqxFocbDfML5yXUlMnDAwNRq6Q+fdP4KBWaPO/QndbYNsDalv9NB8KePmzNwn6vRKikRaC6ZDC6WO18w3ZvGAIXIuHYQoiReOoEWKQSWrwrD7244QHm1IdVZ2IuzgB+UYpbZbRAqzih014c/mbLn6pS5BXi5vI6enMaAkGsDzuOfYDgvzQTpdoOCO98j2yhEq1/KDrExHveVmLpowvs2O1dYfFDl+PSHzV1yODNUKdnK+pYE2wz1Vbp26iDa4+EXROx0p4WM+CamDCFWur/Yppwb4o9MrcO3d/VRvWS1Gle/eDFajrDu51mgDxaRBcq2PexyeB/uJWy78EXnzuCsC/VCMXNT54RHzELn5bKBUSZIy0Qp7Ndz9AKSmBqP6xMLUw3EV87hSCQoLjJTY7mC9yy0Houlcf4kqPBGfApPhI4iTTa8+O91QRMLodnse3PT6roCFYiX1/2S4CCRYNGLyKiI0rbpR9fIcpnabvZuhOikW4PvS74joesNqYy/eNd3SbZzgWIbYoMqmia/woVhIb/4Mcz3ydGI+/Zy8Rp6tFC8ubgkKv9mTTfRqFpGiJk7p6KBozWpSdR4TlharLa6I1SrqWd0eVDWBoezotK8n8oFo7H1tc32aAq3i8Rcders0xvQ61uI93hWnxJwBW5SQgMgA6UOHb7ehzw6PP6fT3zgGxCCXKcSLc568uwfV+ChgIz9tfP6QyydbNUOoLk9udgswQuIejzFNA351CqHfOrZZiCRQ1oNwxtSFHysnlRg/d2zLg6Qey/N4jKLXuL+yJ8mmiwD7eTLrskDIN9C9qWh0f+Ui/6BkJzyp2ffH3/EoR0nnsYFFahWOIgnZq/t22mQEbGLgAsGqyfvg7byiz8vCsjw68vFzu+LPxN9tyuRds5FoPcII5x76vpyhqmJCwhB2rnZuU4xzI4CGCZnfMPA5IvvmUWm22jBCPH4B5CnJ0RpSyfslqQKENHc7wnOeOpKfQiSQNt7wKiPQcB8HvI/R2yfvdHggr27AxX2wLrPVfVFZJONLUHle2gpnUhS3LySbdQNxCeBUj4TOCfTkCve9UbmQ3ORtq1KpyWa2P6u/rOXvN/1ueutppPW0oA2d6183Xen0PRWA/4MLred0Abgp6X3lpSr5KZMbnxMk1Ljzb+NdH23w3S8VsMzpEl7MXVkIQTr3FObL3Yewtcq2t6RZOBJBRXqYEMFbB60MG21MTQjhiny06p7rvuAwSCEH6X21ecx3yirPd92rPHO0L1jkcFltfi/z6FKnZj0s8Id2LHqBUwE0CUsHowzHSEGmczVUkobLHLLOkg5aqiKjYB9w8SoXNwfvDuiUDoh9F1yL+QfTx4XG22GSOY+ijKlX9zbaSHuCCV6o9wXoqBvMEMUZQ+kiD0c62jEfE+CpPiStvzdjajjsi56ZtpK+jIRCcVgu7x60zQ2hBHn5Vf/CktqhT2Vxxwk0b5owZWCDPYlM6gVYuPsFPmP3LDGU/fOuAJ3LL6Y3IKSdbpjEg5slP/nBT1Qevzb6vpQJwGg0hX4YUhvCo6LR1qTv1Cg0k4n3PetyE0ZxnFbC+YniLETAMrYEjB+Np6B9mzDgndPYjCAaXfbICOoiFufIt8TUrkQVXh2UwdHDGAuo7nztuFDFZb+o2a51F6U4rItmfm6T8/SgPZ/saHkwPH1Xdp7YVsAuKqKFP9vDccSz6sfpf5/JeOjRegPORmSHQ9Emx/XU5qdKap7NCpRdJof/01a/LDF6o/nHGVuLUVOefg/uwc1yC96+7ra4j/OtDYVoWksVtL7ttHf2MAVCHwirduBKgB9rpOCI+YbnUCzmD1kEhuFTdmfM/knu6GfKIHv2zghct/FAqc9ADYioWC0pKFb+O3obmL465DX46hR2COLqZZlPJhsk7uXPerI/zbdUWyN8jmF7Qc8jWpNWpV2U7KQ1DpCxqIDehEg49+pvyUTRRMo5T2PHwQmFQXtNSrqBAN7eATE1v4xm8A2YpATTPydgQxSat1QFm2FZ0r/ELPs70WxLDMtPqyvaxZucJO+8VHEnkaFi9lAnmN/+9awpCrHloyONAZyygDJUwgy/+mL2QWQV+D1x1ZDLG7cEHEVBel+aEQhlMeAwuuX+zZUH3M0GTX7/6A81q63QT2vmJqJtJt5zgKEn4/3+0Zik0wtfXOQZd3M1LiJSZoYwpbNRBH17qSeVeTA9sFoBjHZmAQNZ9nwRzKFHlnIEg9qUx4jasiRWsjza2dWAZ4QVS9GFEiCFMrE6FjcoyTz3Q5Kv0QYsTG+6/KBaNuBaONFHnjIaJRQamf5Ia8KhR1ZOYKww2N3GQj7c003mnHH1fzTQ3uZ6YT7D2NYm36gNPwX8O4P3kCWddr8PJ7Kwpq2gsfMsRHRY6aPw7gIHgO55CKIrEmOKfbKNan9KzSFodLjg2PwgtM+ifsgLxuRRoUaL7FbZmHriwPinWRFseRomEg08dYZxiTzyfgYFwTjBwKkDD/m6oHg3PQYibPfbof9jiM7AbLtUrsZlmkaA+WxINucVHT4obl2ffWnYkjSxuaYEHwYZSHysxs7TtcQ6owplmJBXQA7TxIyX0KbLCY+wMQzwTFQBumrKhbGvn8JUSf4r5xw7GVWnrYnnV4+sLdfG0rUs7/CKz9fUB9AluiexaWlKhlLPWet51yT/woVxPZmMm/62pysrAQYBg09MFwM1w4lcthTqLwpDyIvzcZNzFn9XlVIolvkCb8xviJXlo0FBxrkboY8HtplXen65mUd+Ag06U3wAuicmm50ocd7kybuMt1ct/cBFZmtrlJ20brrPY7Eoamd7xOb0fT/zcFRwAjI7V6dZmh8E/iDJFf+I/BeGLUN3QLbjtIZAum4vFBQG12/DLIft8w9odKVwiEOP3u56WNVD+yWA9xl3iowz3wXuBLtPk4Ydw7hHVnLBF7485CXijIAjY/1bAvBYcqFKks7DBq1rzd3/jzOlVJDB1loFF/+ig7gRxiBd6S5s/bOGHcKcPI5QZoGnbXzHalqZWXFn6eGiGWXvAFjbOWKU9MiVkmijEVG1/f+DrnkPeYlUO2N9wJU9kVTnsMjQ9DTLuZbeXGB3GJgc2160kJZbJeqvoGxii/xAv3tr+pVdEt7ebar3khhvUbBrX+y52NNOELb+98Umw0zCFIxBgddcig2HSX95+yiIsUQt38Cd0QSqZszM5jNt/hR4cksH+c65FQYeExUrjyuO2IO4YaP/5be2eU2s7+RQuFeSrkJLhvFlWFSds5V1cxo7sDEsN7WXuNQ1P5ZvfcdQ6LbBkDVPBgGJYlq2ESwXFKCMW8WgGZKF0MKvgfTrLR/tbe0CjcF23XMPp6j9ARWFhaHeanX+IvjZOBhcQoDqjq+B8zoJPLrn6qvIKojEHMb4+yGxPGWin/HHCxdKY5blCd36NHhOAeWPWIk7b8vitvv548huVDRD3D2w4ebcFQ8LRubtEc+EakL/qLnXfVjQ8DOxwXFbTezH6byVyi/kDdfk0P5jnsYAY9dlNfUFszRSutnY3kv8lf4HCIAQw4E6w6clMbB6F7hxMp3qb7rfTr0d0wTntPecFFwsLiQYbbFUrGzpOkLEcy2Z/ylqgDExBi8SuZ4iRthw/dyrmPdQrAQ/8tmeyevEpivwhFXt4LViP0znGqcBZJ+E/LVlWYPXRWK+HLc1NeQzAHTpVnvJZB4NvIT71q8rUuAoVC9y2XJ16ZENT7uZS8oeLKkQEVP8OeGvX0PmnnT1WpyhWNEghxVsgex/eFx3hZnhwHJV/ZA7z7REobduQIkgwsXU0z7/z/lKADNphu4Ms+39NHowfbAelkNX1+xN3RVXcxHSR6iQKJWw8xgVSTmbmI9NxAJsvEGj4kRaxnW8Xgf0Pl2pMRGfHKrxPzFDxy56SyynjPFhFuhQOMBy8P9Dgy8HfC9sPDToQz3uag9CLYdXIhH5cZ5ZZAKJBhyxr6pyoia6ttWq6ZppRCDUlaBTcjCogZFbqlKf0UmNm9c5dJmcsqJENR0zbUjDVc0tkOgvmHBOXU4CkRzJDSFucUd/wXhBM9t8wSnwORScp0D3/98CUbG59CdDIC7RzqjqjLP4uLn/990RGqVH6ic9C0Qwy3N/wMVrl4usl9UJESQPOk8SYljeMb1nNF8KLG01NlvXgWPD1hxknPG4kE+G/pe3Lbdyn/RPreqk9NcZkMk8IaUYJStVKG8FTBYt5CLxzN343ar0ZpR9nfVJIzrhcLl31gz8mITKDA1neXajKcrmKSAa3tk/69lfczZqeQh8rLIAOKQRJSY6c9PavO+xb58hBpDZNy3XfbY47l7UBHfKK7W0+OU/SCPK8BHu0Sid5nxH72xzr1E+7ERaZ+YrhTTr46Rb6qBljsmRyW1cSdLBQmb0azhzsf9qvXxOUYJOAjJkf5m800Q6rLR8cCBzB+/x/Kv+h1NRiejiH2XXXY/rwkgr3TvdwlqdXtSzv0a76xJSlTxfWzt7m4/NgsI6UjdPAKrSodBubiUPfMptUSnkAuDEbGvmXsWE28GZzXTM9gSB5nt7HriKGFaCXm/IqZGDvG/rdS6rLEX9JCXov29jEIJ3acZNvGhz/ijjwRQ4ZKWoqruvCAj087gSbT9sWurY0ta8JG9dWje5g3kBtGAsnubH2D1nGqomaBCj6JXLef2KYMFecmI2coKuoS0shrHR/CO0eS/cqEqyLqKeVzKDqBCKr+SisWNMKicqUXEvHQrmYOYzSis+wA8HTCy7fjadxnzkF1yqcQIsb9vGt4sAUp7QN3fOIOlOTuhrZxfhMq/SbEbVyrYeuf3FZRpmKkSyEXsyVc7SOlD6nOemi0PwEsO/6eeUJSp0vTjzQgsPNvKedB778rL94xYp3T+tWJhEywknA06EH/6kCPB8LKGT2t9ouwNzH1aIo7xlClD1FZvG7E6vRcGCUq5tae+hDujXetCPLAS6dtXtRhJqA+wpfxSjnolJQ5aQ8MHfnJE11rpwi3NrX7nxzu6Xdedu4BGy58r5Bbsv8uwSaban7MgQq9/Zi1FbzkJdJeh9Ar8nY2CbY8koc/a1cCXl8n6Iu4OIop2LKhof+w9tKjiGWTxF/EubC4xSWLtysw213msGDYnOmAnMc3npQQXqD8t7VCkv/dIBor89E9ZCDGD8ERNjWkvWKK2ZDVUR8tgwBvpmFa4fRE/UW9qSxh0toEyFdou127x7jdMLiZdw84xd7JW357Xs2roFIR5xFCV1VA0vTQTegWwncu5KYto8xeAMr8kOEO+AfpmFM5d8DvzHONkJTTA/JlcuvMsWHBL2N7y2ivTzYtKn9bYWKvtAxWxgB1X5hY3nTcL21PpXudoT2IEoGSEItey+A2DXwrFxrtYpVF0h09tA/2pS2F9e3Kk+24zP7Ty48eZ+/HLeF+VB5oE5e+sXMF/nIZZg4aC24fZk+hG3qTHcbvaV9AlN0OjjD2Zmd2/1/wNsGXvRxhFIagAaqp5yUabG5quwIRD6V/dM8he9cMFMY+qP/BZ6h52g4Q8Z68iknDfA/HLO60UEXMwk+E8mSxQ79wxF3O3K95jxuPfssWXp/fqHcPVyg4ensJdZWuumI3id5Xm/UwY0bCaVKDelk/EZuMxmYv5mmuGWtOCivoX/DYmi4+zTSg8KbQPMrmGBjQq5noCIQ24DraszJTmEysK/b44BuT0pm94jAoB1+4Z4oF9C5iIvVHOWYoG+XOxrzJmNhDFphJZQ2LveK2NEDpOGppYvTAGT7uXP39pqBgh8kE5nqQaT/p6iIxhCepXbGTplSkLYkBVBam2I9gEoKs05J4ts2QcCRXh5rSpCZk8GVOJquNvqnO0kwiTgMK9DIwnJk23iTmWAU5DdLRcOA6kkavQADb/Ik7kqQzl+/uygROXtuL/mT1SDRzgTPjyRcG3xpHasK0R1Ws1XAEeharGzs5slakWw9DSdX2sGYEqhvv1uODLfAmvKFCxx4UasvPtSS40UGQKEEnA/19M5EbFkkdzo8e7rXpOLPrf6Bhir65K9TPxV08c2BOKqJRxz9lN8XOo6VKH//h5mPa0LIQtszqlGas6PRbpT/l7fB0iycBr8cCsg32/9GyQlcGzEEGbkq7aHDxu2hbtrQgJvTkZVU9w4q3stDgC8r30h3U1pIAjyZOAdRv6FRp43GAVKultfQdvw9YiUbZbcNdPMyjhUIWjGwWeBBnkf8OiYGXTcvxDrXaW2+KmafV6EKBWKxESxZpDUpGsw2a/4qvmc084L2TbRyeMQL8Tz9P75+9BmmNMW42him6ZU6/zGKLcFZNbKz2cITvYC43xOD7pZWrxfKJpXIieojV/Mxqb40pz4NtjI2EqiJyve09Pcg6xymCreWlzsfGgrkywMyD+jZ1/Lor4TByro+9cg3LJvZNe6HcUSVIoAajGulWSMfAHLKUEfJpAerie9UugQ7GmPN3SIUEMU8bbOtXqp3S5iaf8ZpCESC01I0ABpiy1HuvAaruITu0+HBN1vPskZIco4rHDOubDsATECECtCKM3Qaxfxi4U0xOkiGhNDoCgD7fVlqbO+YVA6wg6xzCwaz5hgy1LA2svok9kLooz1RrxHlwtXuG7cGBFF18GnCM/mtbCEN8mUn5J7YDSz6GsOCz+HxDBd9elgvDi5hsUEInULhSdDmwxqwLWsFriyHK6GSpciQTdTJYJy2iLtSJa07f4eUaT5nXEwqav/J/p2aMvfPcGU+a8UvGz8/PVqu26ls+0K1o10UcOzoAJSYrxDAnQhSccomfmdoB2KpSdEpIIr/UGVWJ2AiRFyUFBM6EeLBaN0i6maR2D0VKxx6Tpye59dq0y89qcp11E5uuR8I1mwIIBRRwbL3jTJr/1QE/6UGxGNXooGJzP+jtRcFHYpG3DEGsjHcm7hlLfqE60j+1NYSF1qehaADJ/5EH/b/lIKCJY9XRNE1xa2amI9RiBhTD7Yr5UwpC3+UivcxenxoxhIzfXedYDFyFKgIr4VZLW56TpshwYe+F3S7Dsdv3kXytTpTQPkjKFfpp7kgnUoYpTSt52s2n04Agez20a6pFcZaVXhhK1xgWJ7R2TcL6vWfSUfRjT3gCVmRg/f74yFnI892pSBKnAdNFQ2DPRWJHXPFnpGbUvNuoET1JybaRXRmhhS9xBUwPCIxl3BOiZGDOwPd9mwuhktanMc/JqXEzwa1IyBKzY78OdNtcBQlIqmTrpre3rHv/iWWCcSl1c92i8HbSMTFQCZvbuKE6FcYg1wtLIiyfM9S7wp43uleCslJ7r/TXgwBEP89/yTVrmCMbAMYpc+LfaxRXLPEHYYcoOwqEZDpq4KmbljvV5ggqYHI9qmpY01Oa0+ztfqTfCPnaeGPKvQ94Zpxz/fhangf5zoRwh2dplhlDGZAdVT53OMAk4+Q0DZwLiz/F3VKfv+s81WuRqKljuODDGTjqQdw6SE1Zf+aXuapvcFInP7MjHRnXMK9N8OST+KfZpHrd+Q6K7cMLaPpDVD2UfYA7EO/fJjaxdNZrQFPrY7HWMdMaKHe6b0odtX3xEgpzSA7nc3Dx7ID/ZJ1kxCDD/Gf1HzpEapPm56qF/pMlcnQf1D0m6Xga4/GEsFSBcsO9gAzE5o4beerbCMHxyv4V1GocwnKc/BlT7UEf8jWyPo6Uof73YsStOM8GJecQKzos8pu0zRY5r9e8mgv3Z/CITQ5ywn526rnliQTVVcFeGnKIdPH0otBJ1AIc+llfUwOwX73Wkm9VS7NKxJAy0jBGaD/nLRbKIYUpauXsoC5Yn0HwQps7UtacpQe+ErMMBwdr4JiskAtGjnXfKq4VUNz8E0FM6BTqhUI7oleaZ+k+0k2y7r+BFmP0tj9+yVOMB6EGxPNr9z/JNHPScRvFqf8Qzu5vmM8IBMLLDPlvGDQANmb02xzP99K73QdzAJiR9R5Cig/KFUf+H5e0AvrfSofAtIflEOhRRYBA6tgHP6e4yP5DJtCOvMHc1W7FGlrls4aVOHQ40qB9o41MUvMBKU7P0iGlTvGP3V3PyrjwCKQQ/YgTNdGaiW4InYKp+7nrPJw/mueFAhoN4yAAb1Ujxs154BG90xaR1v068f6bIvxRO2jrxZ2qzkfKKxjiNcoYoFk8g3+Cik9a080434PnCEjuzw82gHORNrbF/wVcRiPaW6PsK9TII8cyYPR6X6AZIWT572NE/xA5FQI2nMWqSIELp9PAFTncFtg+P3DRxS0CzP1nLMYrLpe2s6WwvKtvvKtRznNrmICo37pecbjSu4wHPW9kTaMtQi92997y+TjQuWLuoTHdzcbGzoRwPecaDh8ViV7mUxXQ62WsAhhTLJRBqtnBUZI8j0g8/Pm9Ev6TvnxMDpVh8caoR8fLBu6Wee2AtgiQpzt2VV6sED5LEIjQQU9N2BAp3s6ZADlDoe9lKmFK00JUY53TcMbXsS9iGYMeIKTy0HPRDv7quBUwUG1oPwqbtpeRP/oeGpdDOelonQmQ2EV0BmqzWoyAzBpieSFH4obUfzAMhVLkB1MOtUJeIXtlOgMkOjeKOYCytUmBnszGG09pu65jLfl5UaaYIrKzAm9wqfqzLpxDDtkgtmgm5MGNo/MQrx676tHg2uuyx/seek9yfiyI2uTr/VxYnPULsg++O4a5mCxsQKtNw3MZZG77lw5LHhvlY2qNgLzsXJyxOhneTtslonljSDqM7/7JUlc23waZ2ooZUiR0MUYSlkcvID5GE4mQ7O4BIZU6AP7WSXOChVzo274cNX3yXTdqoUDAhdwyqcPsNRK1jXCPZpeaMFSXY97Jx84gUdgJOSZmu3cUIvXxFt3rSStZci8rtMppcLALFJA3JVlEVmwMMeNFDuFE6/5sJg/BObubgMr9SuzVo8Mju+vi+NnGaGOV9pveu7w5R7doFArdFbqTYCDtVcWNitHP1xNhXWkfOzK6i/mUs3GNy9yvYTrSNpaxt64p4IpBa0lfGqTw/2y73GeAWNFg5MVYsOSWEcFVpOWBGsNy3cpK0wJr9GYcn9Io1OKL45A2/xTs04Dfq5MwBGJl+82hxvXsy9tEzGVZtXsGVAoIUihuj5gt1/gRJ4ydu5jpR6Cn/Yqm1LaPmmr+u92LRU9Zpejh5N4r2hBAATvzXB9vpeVqdn68eDNqWLE1UrFp43ZO+fgAjy4ESIF4AmHuT+H/vvLRwms6QkbbfGFSfyyamlUO3jsBMLHt0pzvIaF7ApBMU/vIhNEISC2KHIgOcf+R50h9rBdRj/o5i5twXuXWivYMjXWTNnw67q6WbNJvun2KL2jIjLBghxZPZWxDYJUxlQ2PqJRo5VuVUkjVHMxS7/lXI2GKBPbFlqZU7NJuxpL/dARN+W+YYAYFjdPTOg/5b3kPkktzBMZzwi4GPCe2WrehPT7Lp9T/O4GGx4ArHGLpXsw5pD8E5GvFiamfuztkDNEODaNQaK6I1kSjtU3sewzvEPu3iXArbozRfRW6FpPoxqmWQaQ8Cqu4CgQ70MGEL7rL24fSCZp8qznGQbYmbRKv0Iq5ewWuZDevoyBwniazPqeMKvaK06P7MyksQWjIQasZT+UwGydpEsGTukIjw4wTiDC5H85giZ8o0Cdn9QYt38deAsEdrOPfrf2HKNokwbWvY6kUDWlvW6dwxiWKZyI3TvzkVV47/cAeNureFbT6M5ocxVdMHxFSKSLgXowRY4Li8RS5NZyir3w/E4FKHNXcZ7owacXdORJUSSXo7xNnXo0bEbTuTwMKIKTi3Usm7f4k9h2xaXGpOXl4Bcye7BXlcEGL6IiiwIdAPZOZYTw3/OGIdJn5g0Nrt4LNWyjy1Nb/oHgoc4bku6wHMkqjgMNknWMReyVqoGmxl8NAr+6dbeV6+1wbPd2UEf4NO4ZyKthj9F6Cm94z8ZuKLWdo5e2SjkXlbb7sNWNeXYRpJwfS0RY8PgvSmlHtegfGYawMeROlQie6tH4dmUJIkHe4JBi6udmPxrDlt47zyASXj8D6UoLeJqZT1sKtSO1lcM9/QsjQZu1QzajQBoa8BhOTndqGL5rsBqQuUSF9e6gOofvAH+GYKy+wZF3dNDbqZHzlpWKFsz4QNL035egEcP4lR2xiTe+CpdWu3Ju90wuNfLbVSReFiZQwlU/6BB70vfLX2SZ0kNCu2LtqT0NaGemJXVRyFaZVvWdA4ud76a9s0FEyIDks0c41Oxvrt589pKbbcE9ZsDEpUuhzJDZ+FuiqVy4Nn0JhoJzzaCPUCbZe+viGpytRASIibh2crKGaqgBNdtuV0v15+Pnk5u3VdH06kJwPnzKAYw/TMGIY4SjsUO07wRB6C8uRdVxTVNhA9wEsL1IYMfp8wm3oxyL5LI3aru8DLe7OaefusQSNfHqPJ90m8EssykCmHnqVOL9aPmCZv33I8EiuX3xBwkz4S5Q3c0BiZD2wHxvi1HQ8v2J+BPraLMVg4kny2AMaprnyaw96tftHnp8Eh9fOYtUmKk47T3QjZtF9r3LNxc6Wk0YSZ3h9yqF1EbNEkIWonJD7Npui2NwEKTuh0M1LY0tWJvLN4Gngl3xUXDL4N/VpbI+vNPISiFMD9or2HRmstiLlsCf/OH1UAOQhqSxW9DM3WU18jMfu/SvIKw3vwSNVNkeq//pFEK4dWxX4K6ZqENfJaSzeHgv8kC4eIr7IBeRukwznEXsPh197ePcqxgb+Ydt9dcOETViwgZqRKPESHie+sEA22pB99ZlqWGWxY9pcXlxMYtVVQuRVUNMGOXh8mVJD1dRO5EXkJwZkxLYuX6ESTpJ9bdH38KmJEeTCfNSnSwv4S7AXEho0YuTd3HQ59ffotNOIQuJfMoIprNuhxRS56eEsdAei2rReD15VXvk75kogPNZHUOwK/sYjmmzk2FKAo8dRgprHAnoHZZNlG7VtUWd9A2A8at2TgfgOPMPcNHs7WPo93KCgh8MJzU4XSEPu+mxBXa+iMvxqRVTJgmM2xpbAjkvpgpVtQp7BoDHHokN4gmSl6VOWZnbsc7UvdjOezB4Go9GANUXbqg5Idjs2cuF+u4Q4o5wzhllgOGHSLjny4MEqxkghq6zmuS9rODow90RPsh7oM/D7u1y1sK0IShfzWrqTxBIsv9+8XLxVtxtxo7YP8dJtkBAfDNuAEimW4w0y+JfplR3XAfSiVPcT7TxaASvBoLaauqINkWxAngpQkSxGEPTbEq50/PKrULhz09Wg3faK2F8F8Zq/F7MB64cw00TgxNuZXyxudIXqvWFVi8UHKcE0sVAtdsw8XBDtJa5GMlvcZVtFoejL9mdzkER/hsEJzFVYFt0bUH+7EZDO2vJdlgyN0+VPJPHzhXvC1Ny0uxDLvbQ1jodFzoQJEb94xLttAMWQKEEXohfNtGAWn9aIGfvA4npZPMMXR/g/wpmj1ka9Kw4qT5vool3VZpfbb+yE5VRAsaXNdxQPL07ZRiNS62aI/ahFYTN0WtpaeePw4tMwII8YO4FxrOdr/P2CLCKbgDrmTDOxjbWzpXC1lggd7XB+usPxC0huBME4EDnWgBffgxlqu0Y5NpL99IjpDtALZuV583JszUyOB74oPjyNSxdIahWoJxe1Z9TbfeAFGaU6t+yEt3AfO2Cn1l/14jWmco9CH5c7Lx/vDm2P3+Ws6yAVLh8SlJyt+ScXG+pAc8UVll3ga5g1Fak5nGXyeokX2hDY0oh2W4jZ07dq0rvWhQ1xoztZB1MvuKtzDYbvA/e2OW+kTgeZj8wo0eJTSxCuQVKa9tqrdCk76J5mZLCqhbztf7FkultcELZuKS+slKt9kMgUZ2+waubHwTa8YJqUtsZ8lZuunYNGn2b07/Qp37WqEl4q5bnHDlfp4cpwa8DDl5M1RBrILXflGc4OkVnmaVoTiuMSNBE2oMCN42zQeoxeJ5CTvJ+BA4ypkvZZJMj2SEhl43a6yWQgS68dsjszrCHTGG6RKRzjFrNpwxTsqwrM9NrGMrpsvCTGBJq9MJK6gF4oLHl8k9jG6QJkYHyEL9Sh6OnDx1RQTnHZOgV9mzz2zytAK0fSsGNQzPScL61mmRoidRKEZuqltmWWdZcw7kPpmxSNaJzNHvjiwBpWPG93e/jTAlQLwxKEMHItRN2PV3TGO/YvGOzlebqWsWtLxmbvZNQkQj0Crs462Y2YFQIWd39eP3K+5jvWbfNdXt1jSci1qpdhLrHT3VCe3tHCEy/0calbpISs8I9jQiuBJT3kdb6Xq0Nrp1HJVhyfKGd+yNA1UOMYsWCo8LLyFm7ihSrr+1th9FFTUpt3qZjeBRGZD5CHWAZhGlvSEucIQdsWiYgOwuduJ7Cab9zfCo70wkOXnccL8nJwjGtqPTdSYAzyWs8QHu3vpleZW6kw0Fpn1AGI/2rlXpfSQbixhvqeh9vxe8An2gIc3+gbsdy9icKHlIUYkrDvm5sS4nj3HIAgKgZ3GTR3ZzyFbTlHLdwZN3g0Xx533KKB3FsGloXYtjergb61KyrNlrTdFE2BH5hYXRX0j0A/eWB8HH3uPnYulGMpjmgmzfIZj5pltCI/IGyOBgcgw5YbPwQT9vpwct3XA0xY0tZS4RvT5RZyu/KuqVE0H+iuOmEFxx577K7gNXMTSCO+Pb3tjNGjz36vclu3ChcMn/Dpgxu7lM1i0WuQMp370vQ+IPw/ctGRjaewkvOwAm8iS0UqghFOLviOThXmwKqaKYEUGmsvuKkum9+ACqkpxXsGIokRbCxbyeEFAqfGJrJk0f9hWebo2Z6X0tijDPeFNNn7aB1SogAH/hNA3DvBqIx+icAM0JlFyNVbbZKwU1e/kYeuX5RJBBYsoBliLaOTQIj89tz44rCXTLFpIpOMAcreRLRn9isT6FVXcv8w5AfbR+b9ensfg6HhE18g8TPy84TCGq8GVxduubrThm1d2f+ramyxczqLct8Pos2iCRXVnxTcUyTx6VKIV/LpQzWLTjw5h10cykbSbFuTrjKP7fL2nLSGHIW4I8Bt4R4hWYXqNRydYZnYdqhgq68au8MrG/8QSMTRPfEQnX+LPLG1nOQ1ZHtLYEZcC788Txp5B8TGg+T+TMnmtgSxeCS7AqTBBbAkYkoenfiCR79Jlg2KcRcB84Lfmkxvp6B+ARmEhNVuDY6U4SKuFGFpKEfPSlI1DO+U1RgmJdEVUhNwHvIW3vgC2rZ3esTt2BpphTDJ14dU+NJhoXqoZoNpLexClrb/+fLFyXUmZrMreWg1tvHlAymB8D8v/ZE4EUjIRLfoNVvNlYF+4iMQctR8MP6MmFwYJ0YD6502qEqZQzuNuSc2bw+dC4OCEcK+ZCmkey1ayCzGySB25/hEXgUAqesX73UGLfRVy92KKsIxp/DW9fxhjVhJ+7j9Q6Lzp40uqLANAljFRVynQkgBfkoARLBmCQVKNjet1TVfTxO2P3/UBJ5aRq5PwFr4QFvydR3m668hSgd2O6TDv9PByMRB4m3VYHKc1mLxGGDoS3HByQZ4+Tgjm8NGL38lLatzSSNccBFV3bTNRdgIkkTybOnr86BPniViGuVFcAV0nwXp/fWXJRUNPj2bEXsdUB83OQbY3WDCrEPLhEQmuNRkfEGUQ5mpABBQ+hqCtWgszIaVWiVWB40u8L+3LC4TNOxxD3nfWvr3Y+HVNjnplet4iItW7VD7OGnBcSxxdd6Qvz8wpml9fysLErguvRf5wwVuYPpN72A/ybnl7SZeRj6YGM0P61LGYH9uZTMzx4Pa1veRUMnYVPy7Ml7gt1VyMfhnSaU/uTh0H1zpHvS2MLGcu/+ObQkOReL94tSnrvwvxwVUcY4gMl99XnrPpKtA5d3ts6NLo+14ddfT1NlIICAOcqSDl9LEiJAn1Iqwt2X2DFIGp8zOpAv5gh3ruL1HEFz8d145mKkbLBwo0Q3QHWVcRFM0vSszzOSg7JYV3w7Gb2F/7RbzRUfCMQ3rKMiDgGY2PLS8g+A3vzXrKjRtOaD8NKtJp+5vYilpKfZcpCsSfim9z41dpNCXfMxJt9fXVot7zYDrrfIf+9wLECApNT50r2Clh7S9ivLUckHYs60gXsuUElFvQozP5oLfF9PbYCY97WMWZQHw9opWDU9RYaq1qofn121rG90gjrweHmAH1LpZ74PbvE8cMqgyXv8P4Pe1L2WjUHinhxYATJUaQyEyfoKP3IouZDVVS6ndUTOZGtspD4/JGg6cHIU5q9oGeIOJtOTfKNEvL26MH5t942tAILYAGYd6gaqOUXBLGokvXtSF+QrbUc8tiMvESL7WnjyoamAOCaiyM30IFrhHs8Sv+8IZhzcoNHAAnhLj2/1x6kCt1FPi27CQsvJ5pmk0+H6XVnqhZyAbMkaSL3k66eAzIjSRmC2lJOdSvkRj2p3PuV91lTX9ul7HCja6o5OaPt30kEo3bOYav9mC5qVrJk654mdizGzyiysQCVYGkDKPryUeOXp5p7q/1X7sabx5opFS9IEFwNi9vg/mYHmgf0SxndWcLdqdozwihxvDqfI1v8TEiteXmOn9HrBoiLjRa3fl+r8W8hglRKquortRnLVr2AEtuEsQnhPGYX9GfGPXmWyoEml/0fTISlpHHvNyq14USnkRvDrYjXP2lPzaaty+2RBzTP/4XoBSMJXUS2HnUmzV9d2Wh3Hbf+OcldOGMQZFk7CHAdMrNIb34IjZyXGGIScoiw4n/VAYx2ZpM2nXYTq9tPEIt7Tmp0r1mdH4bhqmK9ZQXCSFeIi5vKk5QsdytciSK4kJsByr0gxt2LbK/Ht9BQZuXmfsh0GtuB63SGp5hO+/hU8KrGBlbZsZZ+0hnufrkPah/4ES5b7qK2IIIk2cE+Y/imGbQyxWUmPCvAuix/JYQc87QzEQhj5xOr0NYjoTmwaTP+Q+hSknDlo66v1p2W1gtsv0RjRtio7DsHs/i9cQ44+lk4WQkCUilG3Qim/feWsnAs0XlAox+KQbbGYrzLNTEcM+MnEYQBYcNRyHaIKM3X3ERnZUWKaXaSbKnhprB87w+hcI3hAN3dcVf4nLvzLqZK+27i0DGHUG76YTUCaByZXGCFajh5hiM6gPLb89ChJycdtbz/s4HrXabmIp5/zR/4TZvhF0JzD3IQ5LcbFTHO/KufaqtnhhACqdFgxR4etbqLefHPRCJJI9mjPyjCzabTVC87YRAZiBxtMTg1SLFQ/15HzjxurYLuI/TvfHoVcw2jpYdQrajncj7YThduOGpCqs0l19mczMEKv6lAHpwZonj9kYewbcwoNnj/srOs03jKUEgqoAh3GpBNwwn3PlqHmNZSf6wXvV7u4w7LjTRVV76ePlouvG3mg6KOQMnPEX2wr1cmO1bincxN6v0NJ1vYmbfPB0poZJXrMd9lKIhvOKsJZPPSd12OW7CUQeCm60HQQVg4WG0RpwL0w2npwhA8E1rgO0g5KEzw9iExDKbTQlKTdCAnfCfwuDmOJ11Z5FkFzo7PJm/hwA635efO4rL9oGg5TAC7Rk55ukrDYImpkqcUlPlF5ZbBXd5wyMfLUKKbOxwua7Jo2RKZ4izwRhU7FMNZmBXiQWEP0wWEfkdUGobcIQUhujsACV4yDe81ib7Gg5p48WcrQsIm12Ui1eLfG9aC6qqJs8f6Mjol0bdpM58C7kTFNVPSTgAxQOs4oWvl9HnLQl7vk6SSa5o20jR6e4pcA9PwG0lZF7yOErZ4tDMXxXVEsS4FRpInOqbmeUv7DdMi8J/HwiEGo1qphksDYwmChwJIduc0ohgX8dCOpduzBc1fMU9pkhG1h8QyU/dNUJHdTdTYGPAbnskYHgZTUK/z0zfmTLZgBQaEc46a6k/AoXzo1IfR8w/2vJpAqb3s6X1kln9BQjL+tSO6NnlNHqmkM/DEhLp5YoxrUbn36wny222u2FgCTRULeHPnzYipP/lbEPAxs4Utdbry05wFn2VtOuMtJd8pDjBXM0zbNhb7I1/SQov3O+p1klPWTPQBOQJH4nwxIJGqctPzoJmvTJ7CoZXv0/iBU1Dedrv416OO3zBWykUT+spJMTUj4PV9HB6EQflsdXTdacMPybDE06RMAOOvIwZemKy3Y6NVrFO53I9Xpi/zWASC/497T/S9zAabsEIlKyK02pKPz4eTNh3Iiu5W2f98VC7TdBt7Q5jsWUxEpzLPA2s5bR47OUY0mfdCXAHKwDPcV8qf8mCWOlHE3vdbE2lSAuFz0L1qduwee5CR+EW5iV1953SwZGpI6mtOyXKIniHsdIiTsQhFC9IBDLyw7CvaccAApzTVLZvGsTK/5QcMODXp7Zvz0ZjBN8ehUe+CNCzeDLsty4FKHNvlROIcESJJpz/30JhCSrWKTbojjWDX/QVhm0inUIjI2X1EeWUvkFMn5EQeO2nGT3cTekDUQ3moRKdlUxMcsu5Q4v0KRYlAcOwsp96vYx4b8D/1q2t5cT7P9ESqgFsKR+Oh56wRL2N64ztb5YeN7QIJqVTKJ9pPFkFeTqgNYXt7IGZ1o6j67xx1Pfwnxe4DjO3GbZfvaNaADF56TyMuikPpnrRWbwZPkblu8UaAg+E6WdnD9UfH8JfqdHgC52gRTLtGNURojxMsbXl/GpymCELrSayMCtMycDmHW3PQPAnYPNSr5kaNjUWR8EQqD5t1OU6BDfNhXKs5kfR7k8ZvVij9msepSKtyAUBGxVGgXOVx24humGiNRzHbhKSSry7vsRhVSI444PrkeMtF3tv5vvVvFRyVmMR4PF6OxUn8Sho+qBoH7WpfYgpJfSUUQmK+gGXmc8hQ2bCvcBc1Dja1Su925jj1wcbP1l5Hw0bjTpwcnHr9NzMdwjj04v7iGhWnigKecG5JeeYJNcuf44bsZPP8XngkS7Z1LRUVDZPdTvqkrPpAIZ1rYhyWS/XzHgbxz+NSau8r9Erv9V0CwjbpSbxmYYKYjE4hkUqXibw+sW6Bt66xBkykbzfMOna27caLbDVGFcg+0ADa8OUn56X5kO+Geo8at+VHQFE2d3q4UaRacYaLjGPkEuBzDrrZm1oCcs5d3sAdhtByDFODQ3y2UeHYTvn+vt2fBNA1KglruTGPqoO7akN53rkQGqviVz7CHr8jSixhMdQRo2LjhWaW2HUUtMWcXYr/QfAHblWqBDRU5i70SBDdEEEjckeualSa3jhfnuJbQaBHZ/zQov1cxzkZ5lwzU6N
`pragma protect end_data_block
`pragma protect digest_block
d82f9e2a9141e31e2bd3fa918abd0cc76104733da2fac96821b0352f6cb8d3ce
`pragma protect end_digest_block
`pragma protect end_protected
