`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
sKiSYU54OQVczWRNRfwEjyxNQHgdmIp0iZiBkbMf9r6pP/KympX5ZocfSpu5ttTKPuMQ+NvofGgiUFipmVmqb29AI67xXxO3362M6VKtkerpIqCc737/YXbdJaID5jHFCK7lH7DNAi3URBBzS4jXSG0T8ofzF0INhybJrVtldX+dRh8bsox9FS+Kb//J7A8iRaHtuV5VjYnQRGZj4jw7gDWxkmZIcnQ4pTAIJsNRtDbdzPphu+oLcXtgMfPy8sQk//ys6IFardcoJf4OiPHoEmmQFEcIpwt+w5z1e22BeCneyOc48dyA3CeajIOfMRgMVkQ7aTsuXtKho02WPNtURI+EkmWxEY5ZOApSLAyW9h1g4KvZU0Ky52KX0jkc9A2bs2AD+Zq9+6AMxdYM6ErjMKzGbtN4VaOnwGmWdOGqyJJ5OLkMvK/RpmapletQlbWrEfbREHO98qnik00JBLaOOWlRJtFKqQJMNK8sw+0OYcHbzEaGryjyUaV0pOUxLZK5ypJonlwSPzQJabsVo+Ap20usL3y8r5YFo0ZM9r2MJ5RuXDg6zS8IY2l7i+6FLIR6Tfqo+0yIXefzXnaASxqrniKJv2CD/YEMnxesKxULSDW6bNZlJlvUQGVoT/44cq44d1L9baVFDCj1PbOcWwGQTS0cgTloosJ+tgxBTs8tpqC/D6iWqlDmmKZ/0PqfGeRM+W2vnGmEj21OOpDIFA0QStdDa53U7hsO42PnXxJAQhjtEaVEFVX3IuuYPo6JlgKdD9N0Fd1tL8vJ6SQbmORieJpU1DET3A+LMKw0A6E8GbCdzGWY0SuyuMdTstwkvhlKc2wBcayu/ZkxfiGZO2qGwlLA2z0uFGlT+KUGY3PDYauFLtqR/nPL7Fo9C2tlowmXh5vyzZUhH49cqXy/KKM7zgaokV3tMmq1c5bZlXeaEHiCR29tHw9TghY0ITy8k+4zOtz6z/yqPzfM2sfynFkBkKsS9JjVCE1306d9lZu/Vo1BsjsJumS8suKXJ7WY774o9AY4VUO5Wo9GpJR7O+KqDvE5aEiXw0nf8/bw/uOnSeVMJpOeA4QWq9P4L92q1jGUWtKzp17zQxUKXi3hebbqyH1TMSiUxpvXEWC0k3TbQlOXFv/nPUzHQVNOTtpsfMwjKIWdP+f9LvGCLzfda9I2k+5u9dona6abXKcUfp9azcFCXIdXb2wuUMdPuiGxYmP0wy9KhSpCcNO/wsv9JTj14GRvYMNN2ufSj7P0/RD7kKo16Myej1VJq5cfwcmX9/VPTdbvj12vVCg+6mdY8TeLQYL1QyzcE80sJ1qIEwwhICLoy1kALw2hWAqOZhiJ9fx80VoR9i54p3jJV/2L14fnt4VJTQcsrgsbSVZk0NiiaUcfxVinsAbNG+k5C66TiMrLP+pMIBJSBoVR3a6cBr0jJ9Zg1V5SdK/7SWu9OOgNROVGzIMkvq4ZfVtxCxD1BTchk3aAgQW1nFJPxsQyaohU7ip/wGBN9CBtCU+DbYA5FtpKRx9YhM69XmbYlrwHU5bfaKwIcNzQ0S4vKM12JyrWYM+4Cpk7Y8KDzd+Tpo3Gbxf79oSVvBjaH9ha2bJWOX3M8Gmdi4KF4HHAvDCCcRrs74aa1xbteUguJIZeYBfdXjNRVQYQRRfWpkoK+R89ImHo79oTleuTQ+hWuzygCqBWcLnAjupIcADroU9Uw8ufhi0zWtWHVFNMwLgZaht6UxbC6YLxU9QE9U6bM4OzVBmFadx6FVujMUVCIIo4H6n7uiKC4ssa1XWy+RhaFNcI2Qu4Vd94Se7RKi1TBje2xs4U1tgXWkNLTzIPSDLUTSWkBurxTju4q8j+ubhEiMxKjCT/+/k8mqX1mGijuNrs1V3qblkTrSS157569WUoKKG7rKjvrkxNlw8OmOYVYi2dHZWShBZ3wZdEZxD2pYa0COPihK/LmNgQMkJEWP/W+4/cIW1PyUMPzRLSrf83RsQcZ2IZsmwxfuRN5nK5sZeliOgmngIXmByCiQe9WqmCRXOptyXgWQ8FDB09jgASsJx36bThBjqp4N7TYAB/xcyisiPS+Ry5bHQZ9H2CAGFAYnU+QyTzYB0ZogQsINYO+uIX0Vchs1AHQRzLhN0qaXQN4K9OG5TzjUNuHNE8cm4hUR32E0YGaXiG3vVa4a7k3ycoUo3mNaI8d2WrDoGDAMaDRzugjPkhG3MN5ZSJAO/2hdcfhhAwSKF36vGw7pWJJGMVM+xHDhX1aOVNSp+dbuL47Cw/c/lomBeFXjf1OHCOKKjB9OTM7hWBHTETphf5ElcxEddZ6ItI256iMsr6aCUMdlL/NTa1XofB/adqQPBlAKZcCJJ/yjt4BL9ht9jrdojfPB9TPyq/8EPoXjhIQzUrddg+dbzQXt0YpCW/jsd9gSFcTnWONpVWQtX/L0Gj6bsnU0pcgAzcegxwMfwC1ArzHmTAXzOgZnLA0g0smLP628o7zCUmvJ5FxPD12HVxT6qZ61UeXCGY5HVo6Ky/FS/aJVjw2x0O6ugSuHo3KwQmOXEFbZN1tUx2dYf6xC12dUaedDQDM6qAtuGem/29JxoK8+i9BFO3w9eDC6I2JHrzNdeb0duvd+VkWErkspJV18Ht/cVQRSRAGWgll3rGeD2hHGn6tbHFzQxjxDW5wz8RBDQYVILvVT+esTb1F/BYByCSX3HSxM/VT2evd1m5RhJy1dym1LskfNkHS4V3zEzcop5DvYvAisHFFOz6DUHo16rRrhtmpUx7f8CdG6o48zPwIQ1KZE/JvbLTsn4w9HMHNLJG46UfW5ORxt0WGihnvMkttEFqyHHB0JxuG+HBwgSTNEVuvq2FTiQSF5AZvWU6tL4SOYrR96mldXjQ2m0tFcWOVxrzYi5g9iCIySUt4Pq12HRg0f0skSCeRtxbM+WByS5RNRCgAb/767ScURbPsfkItf6kUWsaQrbg6R8uLaPhEMctoakVXL5TRzW0w5DbpNFTydjfVRm2VrL2E8BxbbUEjGGXhse6aSXkjH/vwxQgZXiYRh5cODzE2EnGpyGdyVgDWewTGndr03S2e1ow+eNCApl5HUoafWyYwv6WkCrBrMMXxISEWx6T9WEU4z2XIcteLt5pHZM7x1ikMR6lN2xjhKyMjCXSlXgO3Avoad+cRUGZ8yA3zJ1XxA65hVu49qlLyzxGH8vR4TJEmko6f+QP3xdkq4Govo9B0nFin/EKZ7RuAgI60p2/VdyVPKN0QnLuqJk6YFlsKjKgZ8xNg9AZ88a9hkCz3IKMIlzJyEjWjGyEOuhqnFDviFiGtW9+D8lxnJL9VsrdRk6Oud+dEKXzpqTJFklfFRo581RC4nrjebqPVmEO9wyAWMoA3bLB1IEqyUZCVuwlY+CWMTaPIAWSJkCj5gdx2QrrMGDedQ1+l82mfWe8kvxUDodOawflfvo8v5HGLQeZHT7b1tL0v/cdTLFtEtQSJHExyySfR+v4Gwp4Z28yxPxARn74yNdBAUbQe33LwOJXasKbEk+5DsvtmtmjNvOrj9Qb27rDWrJEKLpMNUHmnv/RWyRhMEDXUwHgNrJlGSyM+UlYlHHXIn5OJUG4DIM7b7wxIRUAwYvfslokzAVv7M/XSA2ACuOqmjlI52COstQ8/g9h79zIJDTqODzeeBT7CX515y7JSqz5ue8aTVQiK3apZiUJ62R3qerDXXK6qDrI3yi2KhjxffWZjEZ+8aUaavisHlOBmZWhot7ylIpbhxaIBi47nY3hHEZnvARrF+bCc0MIAZajhUB7E2OiEJ2SNh29Ii0vAp0LsEHKxBKBx/pV7sMYAMb5q9rFHGZ+aSYvPdGbYzQ81CTft3wX0JPVxkXZ1qMxQDw5AFhmKFJxmmOpeVfOJ+7t6zD03w3zM5e9XZTMQJY7emg76kzanz1B1kB1iuFAZnIN/Nk34e37qLT8j+zWngpvNa6R2+J89ZvX9AEuCPnSnZeNt0NuWkJ1vyMODYhkkHEzKZMWUuYYax0ooRlwuIQbV7aUnVknGNBzVlVQ4QDxC4qNS/P/glLoHVbNIkDIz7W/mff5S66GhH/jAgZbJniB1hnxLZtqum3Izo09Wnlvh8KuIe2cO3ufl5aSVWAYdIcaMOIGCQmkV9bjNN5Gcb2v84RZGQVJS1gI/emwMsrBleFZeCJ0HfK0MKIbFqsH16W6tWcvMgG7amKhh3Mya/HnpPULVfHMWhM+0gPKDPexdrKK243kp1xiYZU+iNi3z7dLBAjz3wZD8Ldk6rxbayARdd4UTWk9WW8glxvK/t7X2bEarioam4KZ/yxtYnzvL0YtA8kWgo7lkrZJvweu0AgNFaPvYt6y5XgvUZHhdTfa00lqGdm9YGYK+rBlkIxwH4w2AUOz3gi2M3EoCfnsBE/QCHchsOlJwA4ktPAxbYwoTPpJWncPlUECcehKm8k8S6vRgna7MB3Yxt/yN958Hoo3gATKasy7MW3JNqGUIgEAuV0jjYhiHXN3FutqXp3HdKxvTt+np+EOtavSvl8Bp08baVDVX73FsG3Kn5UJxJ1z5DRMYeRhLODv2OT1Zfg639ZNgYYvDBrIVKOeQlqqOLzBI+xl1Jw7ZqEU0Kt5jpStB+c0Y/4eaMvS2JZX7VJBeqGTWTDxPVC8XCutyZYyqkbLI6mlkNU79KRNJ7nTI44aSdrE2o8Kvso9s00AtXaC5UZ6jaWRbDZVQv2wdMUe8j5iJmdugiH6NtEMOLaDR6MD6VB7wnjS2zy715wzcC5UcGqVTJeSo4ICAX/1ciq/M4yH+tlHW5GnSJTWx9M28bJslItnqIdcMvbLMS+L2J4EC63GAHxneyKha2J2UchWbfdP0xpG6zD9nQMXy21eBmQaYkMfci0+/O4G6FAnzwzdBCekAvE/k8XNsVcZK+NEQcabkmp/JCtKm9QcYW8cIGIaqf0+k7+PwUudztU6Xh7yXxmRXj8bty2IZWz/hfvMLF7s8V1kJE16rLC9zhPCb03m6ZAwSSUgE1FgQKs5mmS82lFSKXJEQYyLMaLn5XimoVKm9lyceEjaB8gI+gG4Lo15nTcKVYnVikEENjl+cTL5s7x6SYTbFsqG2mFRW/M2uKdyEPo0l+aCUqnjOTMnGL7vLwWIsws8xXJ8rrhZGSd0Cr+6cfSlXxlMKJUpNfP0DhvBZSDxGW5NrbK/p5Zyz2e6qPQwpXFDNxiza/fv3zxHMhMh7cmYZQIOHlktMnERw3Z3vS1NFU2kSkbsCSXI2RbnlkE/ReTycroE/OhxVKbZJ9q2WjsyCy9d/I11/rKdAoS8q172bj4Ea3u8jGb55ItlSxp31nomO1Al+DXF75McqCXBEUxxrJL0giKU2GepjFrg2SDfiv4dB/FFHnDmrQkWrqYIDqAJMxYgbgDr1jdBdJ/fpT9nUsL+TEt3k75CmzyPRmPcVD0BqIavz64gBq+/1f/iHIQPH41BQuAjUIERfcVbKcBpJmhAeKNrDIbSsxeRmBWo1E70zkpOkVl5/6slk+KIXIZo2VsEVmG03h3t96EAeQkj+ll2MqMUgBqbSt5aEWzSK2QZaeBCunr3KuVoNFni7sYlbRRY2Aw55mY3BZ9BwhW/zuKXk3Z1ik08Rb5nU3j/yWCZdei7CQwRyJJLpxvoKJwLxtA1f635lrrdSKY5ql7/jDzDuO81nhIIJue5L3p3eVwpPWcDdDlionISUPD1UJbUrl46RM6+AalDrj6iin5SOGwaq4j25eU25MgRORBgrWZVcigaKefTF3QjgBnZ3ALLaqyb4ZaBT1B2HYJ2COr5Sa3nei44zAMgPmbUpTvbaO5oOBDwjQqt+wufYNBh6fvbiJX2jXSxCN7q4aaE9OmlQezN60q2mwKw4WOMHkGjPK3tt/iMQwzaMRSy4yKfOIHDgDm2Y1/uZJ6WoHCHzEooQ9OPyzuP0Sx1a563CM7AX9a79e4AsnAwl07IWCuMuAKS87gl76BLdoLOK8pJ42B3XXBJIlytMbA5iARhXq0MVaCg+Qudhe15wmMSP54q4ClmhRAOF42unkZdEAVPNPFeB/O34y8hCPXBB7b/ClfidJCbUuoxdNEfd289a0MRxchgbqCTQAE++ZisYIwtFpsJu9wRnK/4+pwKqNlvYgb4YDQOB0jfzomU8Gx3tLxVWjT9Rfv5mxrdud0xOACasFobIXaVTPuS0Az1N5GbAMXJ3X5S2H+XKQC9ij4fUh+yYvnuxbMh8KBPrvQF1n/dtOnwzzW+E7S0N5SYi0rBl4nlSAsbuk8fjeDULogjgrbXT16b+Z63emSHOdaQ92rJJxE3QSAQ+pIRI1zzxnKNFl3q6/+TVHZUtHcJApsVNa5zMKFc+bcZIT5tc9oGFF27FllIoU7WAFLbzW08mAf5Z36e93oIC5EhpV3H3wj8FTBdaRndzeJlHkOdfRQsZKIerejubnmsL/XdoQf9zdS5qztlpvfAXbWnmD43kiEDzbUBzNcMiCetJNkVj5gALzP19YW7b0X/gGvDt41wVLHFIQldW6HlsXQzoZ1yTCIhM2HexgdUwb7TJpDII/0t2jRHCMngcrKyFB9IlfrNsxt4wGi1S1XKSCY9/Cr2QU8weM5Et2gd+5ErUu7uexl0kiP9lfGn+QM6ywHZM7xR8rNnTB8yGYt4DTtk64bpqd9HVCCVa7oKEUURBqznEcBvXbTIX0q3iE87ml8Y0T5n2ozp/kPnOmQ7swW+hbALwmUr6HG/54yv+AsN3Kyp/aYkAg2bj/mdL+pyId8NL2M6vxCvX7uO9Z++6AenFpUpL4Re2B7Egq/TPFvwEKEg1vjSOGx4l4taxUmjGISmeUzm62g3Zx2FroGlV4/jOgurKEfNK/yb0ZQXLEu6tNBLHsrDBruEifUNgdtQPiV8l3F/hYDICnroSxxi9pWlIfACMJSxv8Jy/SJRCSZXR7jPSwxwUCqYXo7avrbiaV9KH/vSKxgUpbsILhzTeTQMSUtHRDTPxLd4gHP+8kgV2QfghrmI6nGG2NidaYuM7MDX9ziA9C+veJ+lAU78yi7OYGFUu1CQ5JV2MLV16BhSDtuv4uyhzeDu6APyS14vGE6iv7A0xKgi5Bov6ML8LqoDIWH9DfWq2+L4vZkbHUUvBxInu5B8LH92xw8u9x0WR/ntySVLK8TBeYYZ3JI5rC+EV0sYRqaUQCNE2yYb7sz42R0z+xmAUpmRHUmvrm8uCEX+h6SniIRkFZzlE1ncmUPRP9S7C3S5SFL1+Z45kYYhyuOSHoh7Mtzpfk1PtjfnJP6OBMJVR5E1BlSGjccvmfbTfhSoIilTXQDPpOXb5B0M56OUC5CM+yfiub83VVnTu9pdG5shq51Hg9yzbTIFavK4yCZFW0ZmzSdztOUIrjkcGqhquUYN8yQ0OWIZyUSWiJzEk1qkrLknSASoPjsOwdl5mlxc7E5xl25OqmxC/D4AbYw7vGVZ7fnZJcz4q9Dpu20xX6PzSBKdu16+LGi99ymgWu7XbNHHY4ES9qS2SaSqrg/Eb3VMfuCMzZODUZYykySwcBpynBjguSVy0+YXAO+RAokBvXKicuXSyeFep1XnS93mCoPQ/s1cFL6tksL5PiC+P8riWgBQZWpJvvwqdXBYIo7Rp7oLYe/mnEfkiYM+ydgwibuk3+kgjpGicvIz0Nm5eZwasDFPNvpU6dHXzWzjCBK1P9nkn+QVszaOkpT9v5YM9wpdMAjRaQ2D8U+qMtHdyvi822A3fsfgDJ2AcuK8rSsuwVEBw81+4aXMBR+hh8g433ToVPmDlunZ7lRV4uPrUFx+ys4xEw+o6yWZwxyeDmdpF9RmpAeNzVaq2lWgkOASfpVYbh12EfRnL4oJSOKph6oODCGXEDJxB3OSGg5SDC/WJoaNPNL6NMZYXOl5g7Fv8ZnCCpQsXeHskC1Dpthle6UA43yKE/5YSSzd6qn/B7755L7NGOjigSG7syO1BxLauaE7sQyP7PG3fFeIYBYE39FALrL41aOVJhp824UIxe3QtaluEYOt6QefIYfL/S4+1mPIFSSAS27Pbb9q6HaBOW5+rD9WEUcG1AXK4jZGB79yb6K+DyDQsoC2ovjOIQCfJ5aWD5GF+AN8PrRycvSyQz+0er2A+yeowCrzmVv9TilbVNZBqX54q9Of8QnWxBtQJLUFexdqOl6IhTqFILOH0olu2jD8Fyx9rFFsqs2inRrfZyqnUnxHCOqkW15aNqmLxk0u1mgPSBoDNmI54ZkxNTF0/0Hqxv6CqBuxFArGkSZP5noqtB/rRPufyTDXOjPOElcgiYLtMxEzg59nbylCk8u3nq4i/VrmDkVyuqGnb162GvwBrL0jfD33FCMCysFGJY4ZFcPy3rNh2lTLEqhb4Rsg0Esh13oEluuYVY5kM/nFVQzbk2IuANlW/q5HVG1oi91zwVtIQeYLcnCAXJBU6+xZX6SWMGPoYeJaS+zkvhpYPMKqmNM4N4i0WotNYy5MoQqVYUZ/u8a2lUzO3LLmetfWRZKSn2xqKiMFCqiVJeZHJuZ8HDGyQa/pM6qIgpB22lMiGkctD14dO/BqPnyZ1p+MjTzqSCRmGdvoICQ8p9vmJQdyJ7QUHGSMVuUOUalO+FCSWifVyrSlONYe1mDMZegoM2SFPQRM9Erc8Ksbrl1hEEmIXV4cbRxx4YU1V819JTOYoiJwMtQnhGd8dIDPuocjULYHFp/9/mQJZuvHUBaE4363PGw2MkzM1hLsnO9Ur7ZIYc1vjE2bVreH0e+v+9ZQi0LkSJyltXjSpzahdiIL8MGaLgm6y8GS/kyAChSIdSEdCOsFDX0BAE4ZaLyW3ZghCZ8oQ9UveuzytHaCojoX131D7pAI0U1o9zFAs5JHnyJzpoGh6rEBDOYgHcZp42/0c0HnVGX+4tSok+C6L5QIxYqk9PCdGDQ0kWn20RPZhG5r+gKnCqAWc/1iladQ5Sxn1hbUVqvFlglWgCHzTzLqKRqRRN2uOGpC8kYx8ZM9//dC6sy5daYWKcszTVwxGGw1MlpEevWAxw+cTencXc8lZROvCubVBLpUhYjYX6RhOwB6Ho4gZUkQL1vBMm9RsJU8Ty58u32imGzZXymaZYc0VsXzJx2SitEQF2VBhLujYsnSKZZvbv6reviGg9K3B9uL/4yIPovFGGcfm4khoI6tXECAbi6R6OrAbeuiX7gAQukTqtuTghchFxPuM+hp+w5CKZX21i8yJ7XMRb5Pp8AokXkq78QMUlf9nPGF+bdXDuyfB3ge+GpMXTe9Mw7jIl8tb2COOunXlnUKgB+JC6LaLJ12itBkMMqcVkEPWN8DXhv55LHVgcA1VEP631KSK0koo+99CGsQOuKrZgdLkxZSaHF0WTZa2yIsLgBKVM4Z5s7vos2P8be6KTy8/9ulGsapN4ecpOdPLf0qTuNUIOS6SPyJ3ALo2fCPuJomvdnUTLE8I26bmQsFfLb4kQ46RDH9+ba1Ya7exb7M1HkuLJ8vx51RpykH1+829rfuFLG49GRY//GlBPgDevBebh4Udz/nDZuviQDlM5HGl44P99y43wGvDm/u/8pvNOiiX/a/T0qEJb7LJllbI391t1h1CHKrC8SvUIx6074V+ApHskwh4vhv9YnQQzFlCfAIWRkoLaFsrxLUklqJ9Q2Syq7JHOjzOshlEqq4V7MY68vxTEpKqWwPAfEDcLtp3LbQH5fPoOTHfzSJpuPm6ja3HA9GQhWhkTpx+wX3OHDPpZ9NE52IsItaxgsZJ9EbiWkRgE1EbsLornsMHVnAEr52m+J49aKGEDFDawJYttPrTBnataoaps6T8/vhZY5UtHE3udcTnCJJixgRTUCKi+3G4lKYBtf3TE+12hNwCTG5wReE4Ht1JPfAJu0gn1MzJv2qXzUWOdDB8o2epZeWcEzxDxDwjtVtWkaNaNsxOIW8DMgd4KUYnIBIS14Ce3ax31rQYzPgny2291JQThPC5oibOooGFiaIrwcwgoEP/5gXBUdMY6+8MHJj3I0VjcVDy5rDeoXHwJI744cBabrrdmYs54qhuLeLYMQVhQH5MykCtOU+V3Kq4q+SlhZjvQAHq9YqLePbLOWYY+w3KeYXjDhnzgzfGuCP6gRZpdXDEe6Q90PUi8fjV/bR8iRtm0KVywZy1CrXJQITmMXm5wv7H6HLGDJ00Xbl0F4m87mf4EhO47sVySIYE3O4PgzYHjkNSx/OCKzIopSyVT/A/fF08n4ONhsrI+wq4TAOoekhge53QJ5qXSfjPxWS96UHrlDexgKAeCS/YbMxSTBXrbLb+eNaL8TOwWbFGzbYttraN8nIV7GQ/vYIVT9aq0ZKrZ8NOgvY3KZ2B5IA3iaPBi4WOQTNkx8AFVFBQgqa8f2+X4mgGgo+Agl9d/wd//RXqbxBZGepG47ZP25x1k8G69YWq6zeQi6eC3mb9lRSiTiePW/jbQMlYBThCdpLJBPV2fGvliaa896BRsgQE1WjG883BFT5cGj7ZhntqXoTP774NfjJ7efrxnNq0K2mbMHF8l6kfxigLbYMX3rWVOkSXeIKf811yrpW2goRClHXeYyUxvFrjZoTle3EYf4BnyTAQFclqYR7sJOvfQIwZ5H8a4DcXARSeJDI5F+Y2zUEw1GrlusQ/jb/k21PkPcini8wPbHpKloPqwtOb3+BYav7GkeOHxsstlwhR/RFDFcr7QoiDHPvMeIA1867qn81QFg61IFtrnzCwoMq/DbLa2HEAzXQNcdQQ3vo8UWKkiMq78AkEc7ooLKiQKotGxPdf9M9+7zVUMJvalR1+ihDyXF8XJS/5urGKH/VR+LGbJEY8nj65g6Zaxgeutb/gZ8OZKjhi3jlAMjnGlPDKgzoUf2qKtfIddzusGgAgmlGNyt2w9LNWXzGrT4LtscrvYGr/zGBKMm9lwaPUpSyNfl+ht0AzBVd+AaiCF/dveGUEmguOkbuBS+PpbkLbDQ7GGZsOXuOdLG6Bg7Abtt5yZK4+p+JhY8qNhxmQIor3ztLQ4PzgHN1hLi2cHRiRURoxXuNd4SkR7sklrxDMryOk/gs18fDJv0hVeWaaXWYmqRDgIRno71W4vCLQXNloU1Y+IPfWcwBWWlNCOyluGXqhbCcI7eb73UDumTOO9IvmLxvZ70e2HHV6YbpbBCQi5hU9Acl1E2/6TWhoVBeUv8PmDxipIVWl11XqpjhOHCd6Ea15YGePLfMiSo60714wRFi4oT5jShzSlMkpKJdAR6fxP6VT3nnx7pqhuQqFn3TJJmzoibREypJifYYu4k5JvvqvhQoC2MqidIrhkJsgEfiOS6fadI2TcUGAkarv/Hsgk5/0V8IHmddEp9VrNXc9XLVUrbTNN7WeMsmHt687brm1XqH++zShjMlQF4U80wYYbX12YIWRCj3OXyqLBnN12aRgaRhB5oFHIZUbZrJ57fymSTFgWswhV2SoZS6Pn6UdDQ3/XPKo6cpt0FJay6jgxOpuNZYWRzjZ4Yp/SkM1MCqqUcYGpIxkhJi6SjCZUvy0VIcHQwmAy3BKjIPZpvsN0j/wUUDj63S/rqxU+mzb6loF1RndAFUOSmV2qyyPbzvw7NQTl6nfTuM0PF8TL4uTqeRIcjfKWrhdZqwjwW89f4QmVTR9dEju2O80SbY8WXrWhwr11ttuYsP1sihF2NdoeIyKFYppEXFhmAznpfF0RFZeKFOFCs/f0oBPtOIr8mlTsc0APwitbjPIrtwPawXGE5F0M0XHANTIIyUtsPDKvhu6tBU9j/YHNnjfkwUmJLDy3pXRlRgwyUOX/zXToQjrza86raVqYp1Iin/uaeB2S07bFPgJTHVJYg54/PeKlAgl2pERY/xIH0P628=
`pragma protect end_data_block
`pragma protect digest_block
a65266627f16477090c592cbda09ffca5695f1dd5abaaefa1076098556d77bb3
`pragma protect end_digest_block
`pragma protect end_protected
