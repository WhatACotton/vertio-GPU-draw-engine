`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
+ym95JLKe3QWaFdiir2mvKcYvq1ylZUSVsk7l6NSgd/pHi5/dVKh+l1yK9JE+tO7NMTkmrfvXp4PGJBKc8eBoId1gndxfGvDfRjOa4ggo4z1ErDU6RLdgEvLKVd32r9xdMKuBmwL4wYNb81WwWMuWlZKsdHh5C7WNEdOAZRL/XA5ReR6Gv9T1LJhbtCjdJvCjwCUY2wZRkDs70SaFN4HruPnx7ylRhrGmCPMAEVyWWgQ4AepGIcos/dB3MKdKrlS0DqhDoDVjHPOY+M6oe7+ZL+mQj6tR2ahdmZw/SJQUd136F/2PZSpTxoYuIgoqKj5TSr5HTJnuRhuJPsfpGtecZ8vuJUGG6GJnKXpQXxccBgHcsEERFY/Ni+WwNHGWG6cBSSkC4nDreIALMmKgI3iNf6jyDezC//VhFmaymHzHlLI3JlGKPCOjbZP091coFgwG+sy+o1TRIbu08mG/hcafYT6YRi7V6rymA+Vpzflh3A4ddtTUxNlTyqZ4VFEOsNY2X7sCPLWsINghcGjOkWdjbDH/wtKF/x8IW0nxiaw/rB+hb0QAiam3Taam9ePnyqz39PyvfA9yBLuwQgrC27loOWSKhVb+yaMXIRLOy3RdjWdQ+HZyM0sZOvs0Llafq0h0Rtxv40XSxLo1+D+EdhBlMZkG5G69EVAQSJQLQKZ5VSugzpIb05eGp9o7W8EL62j3k+hAuVcGjpB+e1PsFVJbXWnyBXgIkM/EWr7Dviha7ZeRcpZzZ82SNFn9KDaP5cWGRgCkZzgvMxVs/56I67Mm6veKr+CH56rfyJfI08HX4orYBRo+5UDSpOVmvex98xfHpxxuZXHahasYlEpGe+Z/ZlKxp2mmQgWy2cCsWvRBsHeih9xS+wvcvtUJ1cc83QQZgYKBmdte8gzK6IIWOUfM75g9yo84bfy7ags4N/9IBVCjw1TRD/hJ3jah79zmhDPxlvt02ULp9HkW+JqkJehNNDjME/sI8+z4MU9D5rsTTj1qxgoYFpmsHvPkxOJ9oE1iSb92fpFf3I1bX76ftVYCOTGP7s/s1K/NabXxGyKVk8HtcZIRr1RSgRWVz4QegvQGt7FRzLE5GVCCNm4zr/MF5nXN2yiVvwzKrrYRoBsAgFxkgU0mDa7Jm8OrBU6cQswQ7Ag7hnfthoHFWbeVsBC1QYrRHciWYfHLJy+eszIuEDESnJpDkZfXwK7RqfoMZB725xWVEb19dR5wRHUjo/fB/eOL+6ZgwZepqNVi6oVOY1AGAUt0/QKfWwBfZHdtV6vTMc1IG4bE0MVVdBPYZOO+2/KYmHbgFbc2udPp8r0GQjktofxGYqbUJ4siYZrnxN//FXvJ8jmD5jBRyBQQeD5O4yO+YkZ5BNbSyrFveRB4S1uNcNyM/J+R4ARqkuzrQ2FgbCjgSTXeQ4mUW/IvLM29v/QmrWK9vK05PfdPAtCONS4/LJnNUanBCH5xWpyRLVOkJNWYw/pquTnrPpoAKDs21Z3g9ulqlmz2XIsyMzjgrXntc7OfYpWLRL+LQ30MyEnhjC2eCwb/gcD/jdSRxgalN4yU3LjEpjPTevaRZ4nZKU27RiHDBsq191Hdmxv0B48rt+2bMtwz594Hc8WVYpRTK96aJG0/voTCGYY5P2smdJil+Ca8gylj554uo8wdlLYfJO4dAVnwUD7aizgLj5R1IseyBr5Zrs4yM2PrU2JlxaOdIsfJlDiA+h745N3jGdjZXH33bo+ETcJKdUXrCD6d+Q6429BcPcCvltiaQT6dqTEC0n08KtXV5tr/zXt9IAMC4G+9FqTcdztFaAGrt+aqV/U/7/LhwSEW+A/5CR+DXoYT757h/s+7lYjMAtFCVXXes0rQcytpqxmn5OLKnIqJBR6Tvv+eZy8C//B15GkcauMq2svb2KNRtRSk1aH+abNnqskffMAhLpW8SPjHsNI7bAt4gitEW65Bp06o5cH8k7UMOxyeOPeFS1BJTEBBFWUqXwLuZsgeiwfubJcTWxlTa0lMaejOUMLEPpTQ5uWUk2vkD+ZAvsJ5RSqdlFIgfF9GqID7eYyCTk8abYOYLcVeu5R1HdwB8nuOGTjtDbpNmx8Uc7HTKHzorW0/nvcCz73ezvIF2CvmvU1y8CaPFGxjnTkjnYiPQVr7CuQ1reMXerDfFCoWer+sIM9hqDc9tGfHdOR6WiRCkBaH1g8jTKp5sT9xkuGr+LjjyK6D239v7B9yJnyT16EMmLlk2OFOLk3WfL4O5N2KIDc8/a/ulNpw2gRQTnu0j9hp+4uSeXs083x+3NCBGGDAsaOyPGAJYp0IUvzEtF7fXH3muEbNYKr0kGWv77CbjhvdzR49GlSWycXKhloalz8iErTML2YaY0HBv3ofebwK2RAKx025euQ9x3z9hc7ErBXUPZ+KTWtC4aXoTG1jKrtlBX3EveF62QU4TeZyvBvFmNdC1tXrwUZpxEgumsqLrbmPFXUyjFdBBIgw20yaH4a3Cpjp4ZjG7QycPUXYZ3v7alH7XecpkoTFhHEZY/hWISmcjW/JXbtbjHaEozuuP5EvTvy0xQ8/hA1P2U5Q3vI89QUXBMBF6hfzERupqy+ekB7Yfw3tMulnyYHn8gq5vvSReU88Frklhy6tpdJtE64Rrfw745cxvQawxrOT/JXGHJruU8oCdZyA3CE9AF+Bvz+2I8idxnAHnxPG+cgTI4datnWCvb8SN8jSxNeF5lzqE51hMRkMBzsGMcSV1jMXRU10MOpkChjnP7OHWiC3iQXYv/8tPttdi9TG5GIs+AHnSIAIdHwCunV+7RTOqHAM0Bj4EWpjbSBxjNSp7fxROLU5npN5T+hkbzpvnwAGR7rNde/iXFdvAfvTJWSGr4R/0vzpvnyWyUVhKDfZzdCoRh6CRGR3cWQIu4cwPY5/taGu3myjFwgyuRy9DqGo+9ocGl1LkoI1y7iCRjFzUqaOJ7YnTR8dxn3kDiQpFpdP0UvG2qwPeA9MrolneofxI5L5TBT/He5FzyeMEEHAIasvy9oTrD1nTMZwRh47uq5ciXZmCrNPsr9Vxhliok4uqmAAZy44HtoHMdjz9CLugqyBcXJz2aFX/vz8+awAtnia8bqtQ7uE87Fcwt1FE4UNGQumu4hszjDCWOpB3v4ls8yKXrPDvYCJhPvJXawI1sg8EEfR8DJ5EWJXSvdfgvYCrljlL+DEtaU8l9HKfZqDO8Kn6QrAME4zxzfFKO/kmlKr/8Vj25WzDMfY723gAFaNbtOUdxAMxDDVIVNeJPQPs0d0sCLSQQ7HQxayeGLz0GJvTLjv0lOqMPOiRQoyP/cq5cTJRZg51J5zdjB+aysdnhRXil3GOmzVAXKeS19hUkne/ePaNTV7poSdfLmhHRqKo9JsW1lyXn7UTonBk3cQfkzC/DxlO5qUp+OZFXofGyQ4Hdqkf5a+DgcyBAuZDLfkw5zdXDuYDL4zbziepvHWInxknoxmsjmQDJivbHxNeDlLHuBkY2h9xe+g7r6vu+hOxhif61SA+CI53/+ZiagpPD4rA3N5mPWIcXKA/qHmcetWhykjWWfRkrNd65I5V5uHzpG9qeRp31NNOhjCUapWF8edihvr6D4xLHXt/Q1VCjUtGunUmGt6TZwUIMOTBwA+h67fqhSDDgOsataeM3/JTxb0pitNvtV/IfRmBNQE2ozYIJ9Ks7D1uWM+krZMSBf97PymtKq0OdE5HR2mN/Uf5vCUnThaUQgNVBBctjO+X6Lhc7EGPhR0dErCF9p0CCxppZMw7rYuR3lrvI0pJZZuTzgM45yoPi7P+1IVkKV+WQ3a/vGchFZRweigYNCjt1pgzFgPx4xe5qs7bhcOXVEeiraYn8ong6Q0QiCKdeFAaS05eK5/gqaTt+00BSjE30YhWoirX9d+NW3n043ySeh6z0gFVEiVH4MsCyIYZqIZRrO3vElWb3UBujyaOnn0fJmLkdCh4t2xzHdFGTAmYy9STDF8yUeuJu0y5vwlWmqYEvCI/J6/zyEEI1xRzJ/rQbY8MQOZ9cdPcokVezfnXkDWgs730TG2d3wxuLOyIGWcfe6PXL3lOMfOvmeJsP9jqKulqV1+RwMohDfH6oIcNvKUamFXIwDRjPTME/92sMoc4/YLwtvPYGcLo4pP0GseWMUVbNjXgTZ8rR08QHz7T6ncA0cWvSegmRcnXDYVLCeS9DuhI3ULKUrz7TvM+wCKhcLOM16y3FT8iBDqnHzzOH8VIdlhdJuGK+ZrmvSklPFg8WKYvBC+uhcW8lXp1zkmxiwfuw+JPrK4fOSVmjkYTokP24Xaw+rfydyhJYAxheDoN26NLJBDOTLayPz+r55LWI96Bud3QczvjbvJoh/XToYk0wcGt+QjaqwKUl7wBfmWvcYYNU4OD4liDhv1K+e80N3/X6/UKN4Swkzojuf4ILHsvmTmQU2WG2j2ZnIp3DkWZ71xtNJdv0duF5BkE9DpmZrY/X7+Eca4szref83G/tWpuPbekzqCLa1L80fd3cuPHfrvwlXacXKP1KHnkprc8a+Nfz6P+9vgBJAcDVPLHPR9UKn2EKow8kN8jVALfjTl3zm9IYeqRfsm4RLjUu0u9xNeCVkmlTSX8cw6tJv5X80D9OPdHN8Hpam0XP51uiqte3gKYx6UlHxenUpX9kPHl4zSxs2w/5MByXu3+gEfXUxaSrNrbXSrJ/zEczE0BkvXad9jhf0qkDUMotIRxjSSg3+FA6HwkxH7mO8A5fQKuSVkh4GYYy4jg0B94ClsOKRRvvl8rwbejp/+2eOcPC0yJRKbs84dvm8iSid/MhcQF2dz+w6kYkPihh9Cpw2BnRBK5wjwp0qavsRkZxDrp84pPJ2L1p9RbhXqRWrfUik7Yo9q/PF7Q81slWbJmk13CVatiW9qhN4GURUPqRxsg6DoORCunEcp6CiwDbx1M5mWmVCfQ/SL7MNIJ070Cv47mmaZ89mx31V6qxWkxtGHoKEiR/blIEp9udvKzjlotRd9hzWyUTr0DwzLu0LqxOTITAtMzi5XVrU8n9bdEXSiw6G9afg0nhb80Xqd5yqnT225bAlckh8yoYH1Acx9oO+IB2SiikxqQavQUyBicMxkQnRSLQoNbgA1SqZPMGd+z7o6AtHgIw7e0zqLg5rpq+vfJ8pbnhX5Sq2QRLB0MOCBrn3tQL+D/5ChFpMDzrQzlMJpnSrv37EULK8BGNMMyq8jBm7T3mA3BriL4s25igj0gU89LdW+4WNn6MPQQPoVgJs0ZoXR/eyhOn33Xu4jZG6P+i7xuTN8maMDHbegNmvNAMt6yP7N80ttyjoArWBnMCAjapyYBKNwFcxzGRY9VXT662YgJi0Ey4i45YVrwZdxpA2hpOFl9blsV/w3f212jcqXXl6iNgqAAc6qzLEIk4w5L7ds+v9YtgwsNj8QLlM2KwhalRDf4351N6YaX8L7Q1sNBbPHZM8rXMqn8AmP0ahcQpJCjm2rbsyw3UR25yXVa4j2kkh1Z41XREhE9gFN4P79Y/oZAdrP0b1x1vqR9VYX6OSGpj/IBWXr81bCZSsmAxKvy6V0vHLy8C5fnrdyzMpDDVPItP1EoVi+VOcKoyW4ZtDWriSF0TQ6w6MlbBxszkD1esxcAZAEdoKl9fTyVTl3pJ1fllwSNLuEhD4Tv0AxdKlhNMeyTLIBd3BjVGAaNfik+EgXWO5SdwWlQXm5u3w0IbS9FA7TjpbNIX+xwJg/f56lC7ikOImZX8qkVBKhu3vYUukP7K1MQFrleEqhSRWniSomYs5SwobXkAy9F3wccnHVVOiH4aQ+pFKAN6H3E6B0NZ/rfpvrxa8OJqNCr+naf7vf+eQHKtulqUOfn+daYJqS+rimoLxdeuiQvRqYitrbKOVVJ9TOD0jPoCOiad4Z10vUo5d0YqNTkI0MG3zPWMT2pxpkVmP06MoUjrwVytsd5VDzx9uiu/H/xPG9ScHMA8TGwDCS5vUEr+LfKrQnhW7xXChJr7tfpq6m7VskT8jxTHTGKSdW2Ye0bUSQkNybUec+InHC2LkPmDaCFtOSP5+tyQI5gB5dnjgOjhmDBuOtldLVfivnmuYLdXG+of2iDx3J3X6DzVNivizuLvEeVEMRv8m5mleMqyHVWovLBkYlb/tCUnmMbYXmSaLR2hTdXZ/HlJ6qa0rKS69Z4j8RLKvhkG4JHso26IC1c2gFlEgaGxSKD7dq+qPR5sljU8bdYqVv3DU4ZpgU20+pOdcrU/UBPkuKifGo0XOhkbQcmXNJFXvPU7sHqGBW3rSh1oGlVIXfjpiZU59bQA0kHtAS/+9FbhnjSEQ1nZXHXlgPsAxGxtXgXVyTnVKeG0kWzV/a7eGFc2iYZ8+R232S1PS5N8Ra+0J2pA2oIG+H/odtxcob3Wwl/DCGVzaysVWtcORE/A2v6zbXWMCk6qxKvE+oNzdfC3NJQThzd5NjEtPNdgYg9LANBNayYUuq+x5nScPEyYhF78jniMJZAETmrHXLuROTVKxLHb48ErUQVKOKXKIUe3+WfPhnVDgvSr3EoPanf/4vtBE32AObT8G2Q2VTsNDYPTigQNX3seErHogtjomWyaPKmsOw6pbd4TWYfxVw1q2deoD6DJTOQGrBO34BRqGDBSk68Zq/aLG/sC3p/Lw/7lqBtq78LusICw7byxrAZrRidjSmkDLigwEm9tmaz+VuxJc3TdRmLtoW6unU57MzwRdeG5IO4V88H9zWZ91rNzoXzoaZqXa9MRHJWEOfC+xPw==
`pragma protect end_data_block
`pragma protect digest_block
d65cdcd27b095e09ee28d72e6095aeedf40475e1f2ebe89aade8d339724b9a48
`pragma protect end_digest_block
`pragma protect end_protected
