`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
xQ4Osx5Y5TjWsCbtCtO3FfeX9M5MT4i1V1bhChqatZSR1eqDRNk02HNTFhn7OoX626PhzlweXhINTVmpAJkyyxr7ELFnqBBIfUz43JjSqnt9sspAewbH1QAWYLK9FMWDcxE0dIlVfZywlkSAmKdVDfrJhpHxKvHLVYub4FzuOzeK2nLZ16XSicXDFIwyr1DfyX5cyHaWMeFJgtMcfcy8Lwuoj1jkQp66CpXtRBt60IR6VwsYnP+Wxc0IGw22rHvVJDLlcOqMp0ASzBDuGV5a7fRGYm2ttBxIsNaL/KRWvectX7cIiJl3eP5YXddYBapsqrnRKCOGEIw/wFW087660Y6N1uIlR39zrOByigsZrkJz8hSNNh5bz1ebonmjBMqVkN1HWfUk+21g6Q7gsDJtPX0Z0phOIKijI+CgXM6VzJNyxNrAexnR9tTmdSAXpyRfg2dZ7dB29fGCzW3El/Z9fX6qW1vuaDXno4N2cZwO4GLpPBj7T/fkHWM2VL9Yc5+lss8J+etHhgED557ucR/aGhaOMmCjyhUuYS+6arVIcfuM6cU+QewnNovuTO1zRZA5DR6QwfIHQxOscknWXwlcetkdwoxRMAmjtfHdzEgQOB3TV7BnmMoz9XhtQyFrJXkzQMKyFTJUatjOr4xyi6yM2ZTPE+Xh5cMCdx0m/XRzsa4u5QdUnSboMu1loY0V7SsTN/AvPAHbRnvADBXTENTAauLHf4KMVYtrTxOBX/dWeD+Uq340sle7X2EMlZCTUa+SOoLxPQJ3jDkDYb159/aByPq8Lg++YocNiI1WQRmCD7O42CH7Zbx4o97J0iHqgdpZRUgIdrhmFv7gklOtxU8930gjALI/S+l3FqkkXD9vJyypxnGYQfllNGS+UkaVVz62vZtkfJoTGDf+5ywLMmgq5q7bM6M+uMwRNBhEkIWsJWIdpPJA8Wgqt8Jv6DwKh8RnwZpNyGWa7mvRw8jqwRYSnqn6k4vdX/1LeLmZNupZfAkBNRAWIw3BNbuZ9sbtIcZNtDIcndwyBuU6oF0FQ1s5Lo+5pyhzi+UG0nWL0jy4vC7Q0mi0DXQYTr5ZpEy7WO/1k6QGxVHAs7UOzxae32TQE6miZ55eyNCdtS/PzTUtVXiD0peWfn0GqEqmDwf12BcjRNU/Q5R6avxvjadyGFr2C1mzdHbF0BbJYoFeVptdkKnu3n3mJjlOwqlPR3LxSXEgQ89DgvrqPiJhVj5NKXEKXDs4Bz3iGG4vk5IAtI1z1Lq29jlyoiNwH2hH4yTsvHxx/tBXcxZXavptsS0S5ks5l7P1ovgyXwOgoJ8PoabhCztlrTfRvokyISUch6OVuwzOz1OEw+6iRyvJ36UvpnbLsunL4ROHTrQeOtYWF81sw50AVLFzcLB1ulI5P4x5X45hcy//IM72BfuFl3Q0/yYULI5QnblvVcX3RIghvi7JxO0wdzlsIKoznipynbTyRb93kb35n23R8fa1ydET4W/6X4Fzhm9NRata3opphTkGBmjhXQM0RUy3wJeVdcwE+80+pxPx+C3lXOEbhuRym6Hmne8jdaVmZfnfPdNYHy+0gLgL24ZmilaJoHwWq2mOH4dTc3JcYcNz7vZJWryF8uy0c3mH43Hvfs4EfTA6XMxNosFtyKtUdVVoEDu887pMy4/ORqUDClZV41yXzH4Jf1PlMX8qxxjnOC7W+a1yMmqt/kXEbBzK3npLNcEBIsjxChgP2s8RHDPHyUvvincPkVYgdR/sWQlxp42SlN/pHtVhL+orggzBxcchreUooGyMEi1Y86z70XQc+cNpbvnUGXDgEmv5c3PoqeBmSKOK+kUQPHjQEQ7hwo1pbc6UUSJzStUlyZl3ji9ayQmfxGbJ0oj3W0P2SKUgJFGysmmU19fTn/NMUXUJrvJ0Q8kL/f40a4JxTGczCOo1X5XfkmK5POyCsvIBj/KV9a+YDLfVzLUBY78NdvK+2LLXiISURaJoz4KQGMqGFByqUMD9UjXs0GhnmJTVg4OJlYTrAoHAz3YT9jpP5Oq5BoZo2eyWxMUGXH99DKPN7WufdMPT4VcYGB0P/jaoFzIh2MjZNGpdtflhZRCHheWcvs/DhYyhvxTfk2QXSD+PpvtgLvY8mnqeGdvZYKcUImQKu/HWlzsBVqNam9oYTmai+4gs3Uowzka2L30r17gys+oqiVcnaTr83QuRxe3rSW0drmBZ7K9eG062G+of+JxNXkS7U+HETrlxRRwLEuLQ4JfiGwRjQJh5AUxlTF3i+c/ZE4IOYJecfBj0Vu83Lg9+JTIodU3xlYnSR9urRWGg5KPMlK3Mf0lvIXpCZ2xHSKLnhn4G2HyQqwk6VVml4KkMzzf9QvVqSas3iNFtMywfJ3u9zfOutDItyB+9UnwTm5UjWjlsBo6D6K+ZXxeEgzqSHj/ZBjizJeqBBAK1RR8LCTJR2bsZgc8wAqp9vx7GfbfJcofHWIYmkIURz0Le8REoZCyipNVuI+FDwPgGb+EQiHtEHKBgZj0mQCcKfxnHv0yvCy2js104qb37PkBQFcIZX+8XnNypVvt61NKIOXWzFnJ2snJvVq5mEJd4IojnqHFktj57Unc52iPwCl80PcywLlDIwWKcTXApRkWaYh3CDYZub/ENWenm5qmYNRx3UNMirEnfPllWb/bA5MxYc18XGZxUvNyV9wT2Y1N7I1CdYlh4UP+V9GXOe1/+eVg3/+LLRGaRO27DfIUjS/eoaOpbauZHWbn+nAvynG1GTa/hL0oQ2aH0BF50r/pOfxONGS27pu6K6/zbDwJCMd42A6y2wiuFauXUSTw3MRP0fozD3Z7UxRku8RXMwxcs8IrPiWRLFwTQ/XqD4V9+BCPrLWkTmt3xnlvwZYsIPloC9GiONQt5sIL4liSMSFtiMSNdsnz/Ci8tMWO7ICQbqQ70bV+jTs+hgbJV7Jevn7r2LyTUK9NGptq+XQ7H4RcUa1CB0CG7xTWTlZ0UtYD9VC4zDdGfmjKrNDpDq4fU/vC/TipJ9iVXSvmLlwxzexzyvk9ljhIQEQnx6aqqQZuhoenSrSrmg7BVxkvdfFnFiud1Lo2moCqIbP/Nc2HOj1ibJPsnEKqG1VjU1712xoZBTBDTw9Q9SGHLCDslIA6qK0fuVbAo7YL1szjfxbxqhqaR2rMiRzFy3hKOBGvVIVD+H0i7F2iAPTNbMfUpvJAZto35VU0zv/zLWkLDdY55VUW53qgZ0Zqy3zDB8EcdoYi7Kk2MTz0d6dUpWKiXzk8jLgmEj6/BRePFzSwnQ1tah6GTbUiLHWDuD1mNaG+NABxqAdOeDGqDPO96MQhdiuljwBg9KAt+W0Ixqgc4xyS07rK/Cl81GQpFSXPcH2/mgEQYvNFgnbJbwcC+9bG0EPGrfWe7YyaPZXKFZ2LBoHvr9tyLZeNKysK/lhQEYjErMwjjeiU56u3jykCd6RC/P1eHNCz0RR56zMrMkBSCGXKgMrrXT04iLSthjzx7gCq85wgE6e8NhBOxL3hQKIGv1e1W7YpP1c0QzYO6vEYzbRfAEX4UKOb9EkQGIzE8sX6Zl8fppRbnnw/F5MS0cdclSaYAEDU0PLY1ZbIR3KKNdjMoMxnft9RcvpMipBcPpTwNBo7KFTLNvfgm3tFVwH2HCT1VpwBn80hrn2b2mC8rSjwi9fy66C6TTMLWPR9y3/niMm1Acaw5WXxcfQ7+dA4TlyHRv7pq8jNt9dPBn3ynfWmTqQRHxxqUw6sm7B1BwSHy6tQyPOgnkmuwOUxIKjUCO9yglFHmGbY1nNDlFjmMk7q99mjBDk9kf/S/Vt3Aq0Xt10SwnOt5ZMSZVNwPV4/JuYQqDBDVlhpz18rU/Op7KBvCLxEBMz96PYCEYPGMBvNxv8fBW5iMot5xmGTUiAx7qD4p6lD6a3hdbAhxv71t2d5sytlDh/orGE/8nBcpTpNUlgY8942S/osMELdBWw6famEPvkU0xI3VjstS9Q5kLrvm6KSJddz7csYrpgXouPpTsawJ/0VUL8iHepjeroLBHu45ASByjq5RsuLP7TGcMKHgYLrIvJ7OpEOaMjMOjtvSj6dPzFjaqdegxSGWl4hxKqO2fEFCjmoPaO9H9vIYQNgp2iTs6N+MPoI+bA7moe7iLjTfRngg4d5J7tUlH6jtW2epmrZtKPE8g+Rb8Q6+gqqPrdQjVg+DX8u8dl7o/C0nV6eiE0vwvaTDX+S/BI+Rz2RUXBYaRXocV5r93trludTSvNirYvd+ob94m5YFfw1DKOx0LR1U3HTZKxndY/ImNg4wXAiCcLCb+S2zDR3iPhoK0FnewL3k7wS4Kt+lORAqfYGLWa8fCF6JOq5XK1DWz8be84DiYlxFfgagOdH9FSz2LE+rB8pWln4iBM0IE0kuwBUKDNlLUU6fM1c+/ku5BKyzftOWPnRksZp3pMcPeL6v3xMpYGsLIamrnB50+vvJc/LJ2MEUIOlJPz/ERWdItmvaHjLSkMqOtb5uhMHOEMN4KgVLPdK7lnSgTRaNuO8oh9xR6YYV2vHybNGC5c3UxKX217bZtjF1Ccb/ZKJTq6+vw+IKuHNcLGdRGo6cFvCnNYZ4tylSpvc0j82uZtapPh9R8MVTICg+6QfWBQqkKyDhzb8m3JCPNAmwo1zFp+xTIM8guOXXUcqEWuMp2gkngOWHearm7AAlNpa0oTQMaPpHWN5Lg2hg0RdglwKzv+rUO3s/TPPshAjgK185AcJNfLkJJVmJ2mbjJEGPkSSiRRwFd9B0PRSu5YeABhtWZHBx6P6BsvbHPov5a8X96hDRMBCr/Vr5l/0Vy4Jz4+4U5mcoBIeRE8JB6Nyw+RQ+YLAyHZkdDEqiqhLkSFPaa34iKyIX5Ve3tNSTGcBYh58E88YeBa6QTi8Dq0zy2fCy/qlW3LCj/Wdv7wCegllZjVpPoMOiq9GD0VNTwxxVhrjDz7Kl89BnWSH7LYQAoEUKTfM+ZGph5hRR+OJnP/BzeWALRxrnJVqocaiopT0bHXEsvnGfW9WyZknnwbpEBj2nLHfjgRXGYltYBvja552ltoRR+IjAGUZuHG8HsM42QArZ7X6WonSALVBQUNUn7sEMzcZH/9WjFnsTAmL/xLr9R6YX5X0XoiGhR74E0bUnEzcEQTB96Fcoyqlu7QSwA7dPIouBhkhcaOV9sF4twxuss/4A+e7NfqsqiM/HrhRfbHprQSfiQlriM5zr9MikBi9wFPfR6h+jcmsMWTWp2nnBg2wJs+lbG7/eoCpnEWCWBwj9WJnBWpK5MRatEHFdbwF/EScCqMAYmwtTtCUuM8ln4fYLwdB/hcUofgXta7wDRdI7FJGGklRyHCRak2tx5ZwzfOpb7qp7ZSC0Equqg2nREv5xVAmOapVnggsWEbvkBDS2WiAdSWsUGABey1hmDc93Sgr+XgJ9RwtGaIr5Lc87n4rREvOjOo1Zfh1tpHKley0INNYDqad1jhNzM49v1JCkQr3Ez/A+g6F0z2IdzBDebrMF5+ALdGi3l21s3eVtd97PmkU9fFctB+KsCZRoam1SMocCtbA04UP52UsJ9Zt6gW73jd6TVNhQKAc0kkBNh6eiZpA8g5bYCEaQKdhB2BfBS7FgOOSqWVbphwGqGmtqAKo5F+FbKkF/FbxncgoNRaXTc3+46RJDTn+mMLPBZiQHubEaTjfr1P940cFoMlZYJTFBdlaijKi7L7tBH8N7xpi38niFQyy+IzMylbWq//uYRF5630FRiu10gzQn6P3owEKrFu+d+KX22rfUaSO26sNT51fNIgqwvX6dbF6//DRTdQqhJK7y634k+JHtD5GP32I0LSheNAUrSHmVZhVUi1Jt8kiFzW4Rzj321Ta7NLr8kDfJ0QLUPXPzgFT2awx8IbE3nhvg2OIeYje3AF+gMKy90D3TeoLwSlYy6ygbDeWHdaGBTuI+/Fni1R2YxNiKhQFMk9cwTh/ESulMQUnICLtFlk+nFRcmk31Fs2Mu+KMKyf1mHdwG4jElYqpxQlpuK9tT1r2DI+MTFnu9pR9z3aBr8Wbw824/nC/Ac5wqxT+0jAdLJ2hpP9TSjcgz1ZHFFLBxORBXGXEsMqQNOOPp14CPvIOyt12GyO2Fq3RUXPjWkBIljrs94GTOTqJv9W5DMnjTwOJ3CpuJHWrgNaPdRHxGlz2l6AigYXtqMX5D6rrp3lmKxlIYySsh81vh0kNDhc25zJM0pgevDtR7AbALDppilXSQvtqfwk0VkjPLSoUIDiRvgpy3VBBz40VSGwtl+5lw+vvt53YerFA+Ymua0RCpGAbxdwW3RDKupk9KEEc+2lcZea/06oxLthparcsWjNo7oStmna9VHsB6xYhcxkXFUypJx6lcjWVW45KP3FKTMNyZz2nPXslS0BHnoT277FgoShBX0kDvYCG6Hf2Jxjd2XNTkNcsP5me26enIod4cFYAicM6FV/tR6eERvkRgOknPrmViUVyIc5Zf74MZIFHwrH+ZwOmlOJB96IH6bIzHjx8UhX3BMG3n+mM/nxAa9FoqnK5ihyBkqowfPQVUFQ9Rw2N0ofaS7ftdd2F6Tv/HznooVuiwEHi33QyQBg15OGti/N38iDbk6tyRtdIZNYWf9yyT8XKghKvRNnMusP60Sm4fMALvHZiAPfj62sT25kiQl+2Yj/jlkVSKlSfxGIQinIytAWgyrEl2sfHIJeTlC1Z5Z9Vc7pnPErZm3G3KNUGPofD5VwsBp3Skoaqr0rM5GWx9UYEQ4Cx6k2OVQ4ZloZe10sAu3Fsrwf8olkPihfj77F09iY6WmW0nMKRtBBXWF0aIu/SIzgX5Whl95bz0Kj3vJaAQStsyobuwOOt27LJgAC1KDLk6SXwgx080BvfmJlEasy+Q2Gf7i9Y8xo8w7FZaZeQHfC3I4LzLjYTKNFiijurJGDm/ZOcNIezd4oQ5QAUuKhfJoS9ANrip4gS877BLoX2FyC5030lSbPM0dXKNdaIRahIau4v8ggnI8wNtTNAOhZmQxYG2lCQ6M0w/NqVNomsXzLZghr3Zt7nWkE+NTy96IMISo3ppftY9sXBtg6d7lOM+SP1fHonZjTJ+uIry2PGNPzQ9F+M2yxj83BUsVNjnwjks7fqqnkVM9gIyOsQDfZcVLFloknItYUnRhBFod1vusEqyUIwqQMxtxFJjUoo96qoushGmn9bydw64MFCRseMYEEeUHWAD2TJ2raXYtHlhm7N8A+2NWiqSeTllbYzk+FDBCX8MJkiepeuaONvuHl24IDEAkVxntYUVn5zg793OdWCjI7OFkCL3DN3mrOFiq1fSrPvSaj5FKgwbutkYAKILOi3QPEtcNeeJKGGEq1sIZ0Fbmizdmc4gY0nm3+EQHYUgcHcp5c7hzJOapCZCUMNuXmS8rMtQiKIrYyNZ1rqN4+kh74RwyWFOsOoBQfMCuqFAjUJO+MXFOdcaTgRsnImOSxefxsyHbeTyjp7DG10gpWgou5GfTDvuw8dgg541z79tnScijbexQmCnMZfP8XbDtdzDiYvWLshV0AJ9LebFJleqrYehicyyaftiwuPH9rUeiFOUoV21+u9hK59SEso1PAwEfHu6LL9c8USBTFtABkA6g00+HOpm1B1Nbk4kgY5T0gJcdDeFDs1I9A2MZlHhgbjOWhw2R5WD0ixR9EfzXqijYwzx/vlu9Y2dKW31094y6Ao7kwr5nMhFrTZDD9BojMnsHokCt6Id8+p2VddkEt3ko2AiIbPH67yKwuRkDDVq4Ag8/4PP8ipkq5od9jdVPGrTLgmyC9ZWgN7QrA0Yrw5t8c7h3TJfhTnxYx5DXrhohqQSD0T260kp2qQXFwb+qonkdNwE+FEWREpZryYLuiQzB5mp4VhxcqYvl8JfmJhQcj7Z/ojQ5lqJ60XQpKgbyOpt323jU2SK8TVRRO46ijLKUMiT3ax1bKWcmMgNZ2Hmu6cR2A7whIfK1xfvLzla/wB9252gDiHD0btvRbk6CH0IvpHPNEx9OLm4iMS8o19UMvsGral9vfkV6Opq2vvGAUkFZyakwL/M+WOEojE/UCFF9GbtlIuFy5jT22FWRUyAH292py9ZlN4JX2YMmuD2P7rQP62tykqiX/AD2d41qlguy0qadi8cAo9/ToGSronAQcGd0h4nBETcu8Kep4rsRdT4cOAwaYX9C7R++74uENfuiGfcntrBhoO2GI6vxBX3p2N1RqCbtpBQtxeZZfYULteaJZMaHRRka2W9iQUzOLmy5IF9rxkpXrLYdB9LESDyOOLxuG/HIOSkz+VnJeG6TdrVx7GWhgiktGyfJAbpu9O3bas5ukRVaAN3MtXKu7wnMNItGWlLaFi7eVl/D6xTQpgrPlChC7K4kHgaHNoB4B97LR2VF8nax+CD/Uos4JSgdbww7Cf/QHWGyqQGhxRUE4C1dYERbhcRjilVS7hNW8fC29i2cf+X2IdpPRoNldquYYXiERPkfIbbcN78euUAlHQsAmlPEO1vHkMY+EL1a2jBeVAQ3EOJKv0DeMmbYebtcXnRcXnYBbfPPDeGD9XPsEqLwIbPGsHPCsvEiwr2bYdO8o0IAZnHlP38xl0JCmZE763hJSbW5D46btXuxMhDahCFNKAkmI/Ho+iDMNJR6f9+EcbuHcbxCd+1aDPiHqM+IuYqXzuaCqmFa0cVgXa2SuWOwe0Te4AAEz911LH2M24I/ce/LbEYSZHlhkv0x9hJyeUuh2mJ7Y86fVi1ZdoFOXWW2kQtd7uFkEqb1TjSHnYLDM+57V9oixkNFTTFxXFLA5YJ96O47NEco4njlHfnS74WycgBaraLnlV71GE5hfmQP3gZU9CeKWdXSu7LpftyuVuTPb+2w4/NPZnRGRiqlIfNaEs2d1adYUGp6CiEu2uiyZ8GVg0H54PFAL3GqZMOgiwko2QmpkW6VEgzWKov4fTYFGLEmvm9fcZt8mfQXWA/uyYR5MdWvG8fclrIbBoU/SSE7+4pr2HSIQjsR6BzRTkz6KfaamiYDnr8XjYwL8IDFQUxUTD7G+FRoZyD+XKhKQ2eEMKzfdYxblEFYiKcrxcTxRpLo2QRsoRK4ZnjAxr2PlfKK771Nx7hf+2APaAX2T5tvkiwC9zMKePAf/OKepI+z/pv88EHTd11rf/Nw+sdomlE+nWcaqgz3lcgc46QIQvEpVwFnZofTkdXqZcBkUp+luS6n0Lx5zTolrFP2rggJ0aRuO9AkuOFkaKGG5GjSE8hBcoX0z3n0Zv9Q4Y0HarRjYyiS+EPrg+GIIhwj6eDyFJr7hA3BqNl5uwZo0WP5SEsyKgZ1u5mZ7ZOpMoKyIUqO1VSaIKxwdqWHxyyLUkdv+bQB1LD0lxSHitw6rvbTy0zlJ9mPqwFSuveazISzExufspAaaSpg7s07D7vCwG0AJWaiZJ/DO8D+XkkXvudYSxIWOqnsx3uTwN8NBxg/Ro5MsQWLEUJiTDTPGYtTZoIYCTpXDxpQpDWUdHTxWXMXbOu9iYMHKoYyY/66uSpA4Nnd4+cJPer5sucvgYo4wdLOKEHUIqu94pOizjaZa8e9BINJF69jLgTJh06m4KbEz2pSxqXBhMRpGwkI/c/wF/dX5uAqmFoXmcyy654wSTfhVuAf/F1OB1hRTowso3Lk5XRUwpTRcwnd4hvQN17qdvg2tvgk8QXz211SUZV4kES56Vsa3RTzdvfrfciuXl78Cs9/MpqhNkYkJV+1EaPq8jBnnN+MgF71zvkiFs+YegC1SfDLef2l0PV8MxKe4NOTcKS8qIv8xlQ9iTBl/yxfe+UwUBIHlMrFD7LWgNrASQAgOsSyt0AqDoxEW9mFAcTTxm/6iL9dFghMyhmr/6j/dJRn20bPknZ/6/4Aut0ZwwC6WZYE9V8TWDN46nfhPs5cpV+xuQgcgLscljmxxR0esCqP1nrQRb3aRlKAr1x2BtR5Jr8IJVc4o0UeSTTfi6o6m2adCJU5+QDSeyoUUUN0EE6IZke4NMhBID4Llo5oGDvFtME79qk446HtgyhCoFd2TwFIRwCxKGdqwc6Mw1feIa6RlNESlMYoqjtxYwEwS8ztB05M5X4+OuDuI3BeHNg0fbE6F++gWTbT07yoIvGU7opa+eKqhe3XQ6O8HL4trpRrMYQ5Yhc2zPiJca2QcgXOnKBtwQqemSKD8hSAF/Bur0p1TeuV3YtAnow+OmQufn60IF0PK3sDFqKd6VDBWTU65c4Wkvde2EMx/A0wO4Qpt6CcRU9+uJQD1xB86Rkv3W7gqZoivQSEVFmCXuyqtrYDYBdmMNpRBLmJS25PYHklg0pNIdJx/VVXdXalzjK3p5UlElcORYlxSpPvWXcQ/fm9gfJVErqIUqmijuCqZSqLVIMx4qad50a3FloJGAIIbzXpS2NBtlVshWG8ynWwgB8xZyNoOrvek3jd+XRhRTWX3SsjZi2H6ENfdI0yJjoFMUMFQt1Aanvp9YLLNNWyX1pKOLHXXXdhkl1aO8GuV7UJuf9qstFWeA4pXVNnLoZGgEo2IxxyglZy5JYffcEAavS/vN11kIXiB54i4kjsEg7ylblxkFrxWfzlanRqhdI18gGbM46EdP+Sts8pfh8b6NYepFx6F02UyuA3Wma5/ISczZVmNeygl0AZCnEvVlJCNzjaLRknNGh4CtLqBj/4ZHTEZ8CG+gblE03g/N0MbFJDr+xX1VxDDnrl1wzaWyCY04lexwgb4XnPB4Rd6HZ4M4rQDJs4Tvqo99N+txFqvdc/1qSmNohlU8AlUyz5/RH05SzmYRG7lZmA1PSP1Zl5ljHrdXJp01Q9g9mInrb9b6oeSsPza2dFGntt9PQGMxPbAudHwO30AJMEWtfY+oDEynQb4Jp6oN089urNCEYSP7HCXwnSv8uTY2B5kLN3N33LMqW1CYrNNVpMbGlLekgsrWOMtKebrzSg+6myCTYyn+tcM2aaGpqDh3CbnvZvPI8Bmyo6Pz3dpEHgnfvGHTLtJCOx2KH9Psd4JDmbNS+KW4l+j+nCMR8PFuk8JZmeYMdDyR3U47UW9STyBpSCko8osRskjhKN+/M61MsvxBwXMUDKeBnGcG15E9saoVNTZXtWnjCU6HluNMOzfWmGnCFPuNGZIOxwF+EHIU+Y78HN7i4gT6zdplBXLwr2Hfwtf8WtQkGLdMn0xoEsUQUxYYp1ZwucecJcZ7Mqb8RH3dZplQNE/udAly8ohp19WMn8+X9dekuN9udIa7PQCQtV53G6XnVamGhbeLrZfDRWyIsOx2cx4KkhpJZ9ZEcoobYbP1d0eXNTqcZmWBPcF1NMGMZd1Pnw42+a5IVz7cOfb9tZrneHmU/GA4DHKKHlcUPI09r5iy8Zqk++wBNCeIftuJbe+HmN4Ct88/KhR4w0ZJIlCbcd9icV6B0fzqDYKg3Ri8tMkv47V7J78cX7z8mJJ+cGs+MJHOD9A95fJiZiFiodbkRR7VjIooRZs6985XYETOa4KXH6CuCNen4sJSqbvQWSPlOfkl36QbrWf/z0hMFwHvc7Fnwq25AlRYKBucC/Jfd6IfS+M3gFFX5BlySY+HlkMaBeHC7ClqXFdwhQDDvwLHeB88M42kpDN6W+ztPKMrI5FZreswiKMekMeV0ZuAfDAMTsJW6PVKMCkdY2tXV74vESgFjXh2qNynWEYf0Mi2FS6ffW0YAnshRO/IK35Q2pdTQFUDD7/mcvyRrxCE5KU9u/I+lxmzfN0ZydJmLEur1CgrDzkU0fQ7TCWX8UUkHGTehxl1080yudoJYCoRwmWRSwqx/EMayNc+479NVrdDqoSGX8qQTwf6z+uvjn+QHJtJiKJqXRVukaBp3JgV/ry0WyVVE5UoBd+VbqCcOuBSn0Dec9oPIs6/ffhWmKh0dPsfMhgpvF3fHH9TTkgb842omtp3646HicC5JcOc28wOXbNum3imNLUaYCyjmU6Zni6Wsku+tf0puX+ZwZcsdCLiWE75GxuMZeo+L9nmlqAWHwClWzs6rNIyNPXEpW4xMYKUACaTnMiAO+5PDWUSIRpnIe07j9qfGSuTEHFBP092PlGY/GWxmjw8AAEI0gMf685IaQktO+DYl9MDK1Ep9uZKHEu8Q+hmyWz7DOLgmezoHmjnc9Tolun1WTITyubLJt7YxnBfoQL9+528I2TqYFG+4yZ034tuY2Z0aSn3mn6XA9y5a0wtK2nAMb4A2UTqowrc8Ct0YHkhRNqBlDu6DKiOMezkqPKYS8uyWg97zXhdexHpanRGCDONaQRDakUD4H7hzIwJsu9Y1/cx6Cxfz4CNhI5l0rUfuw6tnlMiuclHCqvaecTUdWwVyv9ELimtJMUXVfkoqN/rf1BI6biFaui67aQsQJE/4RUsWGu/C64MU8pB2xIKtixGyaL8yxv4fRHbx82a+dqlzDAPdYcJCd5eBSKgc2kwmVQW4HMd+kVG+N6ixWBCAYNguFODpypcm6D9QIyIeh/mzg/do55t5TWkcHXqTlhY8cDAsUE8PG6vXlUhK944FtbRTA73JAulr1a8JXNmh7wAWyUdkbguErzkgOJcyCHrCQ0fYzZTscpr1hOQU32vz0jfoEES7ma9glVkT9beeJ0PYsFjrs3lr5kwIxgaqu1P/WUznSGNC7rKUv/oLV8IgJMfMT28ZZ/3qqArQgMXb6V9PW38LGCdJ4tQwJkTLzhkI7CEGf5GKOIcBZVYMSyQXrghoCNwVOcZwzD7klWbcOwury277oDzut5vpxn2eW/Rf2nApOitmdzlzYTVhjnULt82O/Dci1fW8sdMj7XM4pFFiLAEP6yA5BsjWp94ffT+ClRCcGXO1ydojuEaog0hZK4lmZfzX0qB9r/YJo+oZiQPt5YOBmPRUJ76aro98lD21fzjl+LUpBpE5BiqjsSo4Z83wb4YH8wL9X2ah7YfgJoRGoRcGZSIaTqKHO4lPPX6RaY3qNL3HeOibNMwAixfrtU82LsQcAlSWOJXfvUDcKlhJzZ/kyOofnjIuNhiDRnFGZBxtJmSTCtfO06teCHGaWWRpj1tim4Ua5IXPPsoebJrc/NQGNheIZIr6iYLeXIJFSJZhO+UOdO+V7XOjHoEAyMy/1sAYRySPDFw3s/1UjbNup9TeL4oaayR64BbEws9opquVSETpmX/OEpWvysYatsPjNLC2jaPXw/UGvO+hwUYynsw+JnZMr4FmQqPXyMVTy3GANqtCCoG1J1MG7ZyT1aEjyBN8qSFZIAl9NViy6JTTMeauKrKWuFGaCKvPMMzXqkc+4SkLrlJm3QL0QTU481eyYOjPxg0nnIv8ey3H547BpVz4VEfi+GHjLFIvnJSRRzizWYzbHaKKriWDFNxuMsrn+EUTkO1/Y0CwPBQPqy7CNglvTgj9qm+JGN/88NUQ2Wuv4hvWMouBT3XwizrXVA6ubuQ/pLxM5RNc4RagGNjDeRvLTPJHGA073f9o2foXZDLmO1Wl2+QM2hbReSuM9VribGHhblHcKVhLLQL4t06N5LQAaa3xiXAwZJnQEKp0ggVMgNXlFw2III5Dc3pEC8Vghowp1Gde9QxIDjk5e87NkYhmaUW/HKSXxNLrICgikHajcljzXmEnqffIUnOd/VSGJ4t485w9q7s4MDpo8TxozdVHw/l/A20+7Gl3l2BYxX32y13k+eqnVWykt/zxUJ9A/8mxGGHZZHHCwJFqpCKBrQtR+yi85ozmb3r6/41I96kznUqsqLtzoakGxBaNehXCONNoB/A+bjwjYWE4BaS5IPYqwUMsWBz3CeS7Hw0f0OoEZ16cdXdzEhG2M03ba32qmq27Xil3snZvjGen42FJ2ASCDqK/2asBXedKmESSYQ3Fa4kiY/HUChQ+52A9NgCPuOCcu4GWLWTuQzwFoYt7GChOa8SG478Ex1aAqux6P2ZtxQOC0mtv9eXkATNprt4nlBX39eUbJydlYU2GG3CZ+umT5/DrIPiFBAxMKMrBeU4Wo90/isCM2XPfZH/Hi8Gbc1oHAkqU6km6rH7N19x5qtp/y19qGZLF/Q9dg/PkDvz2BWfCq13jjjNXgPpmupTPV72CIsEW7PtKr0XoCLTQaMueoe/yUO69xquQwQnC8viULdwUxJTqU2HZ0JkN0jm1ByOzubK8y5NQucoLheiNCNmIS+O6N172aPO71xj6tfECx3FWDYcCXhtzBQbygs7oy+IT7wtOStMDjDitFRPR7lirTuLa3IHeFLkAYmVS3cc+St7EhO/3k8qHyuUQwfg7pieFT07KfdDDfAUIDEhp9zQouJnkUXnkS+5OOCE3u9DnQWn/i7x3umTt9b8bbuNkh+82E0ZhzqQW3RtAAQhzNsSotHjZWYNKBH4N7/ULy6sD01UxXFwxSeSqBoP+ePHcnhMBTWJHXY5dA/qEywG/4FQfhVcyxdhGrQxrnUViPN7LJmSzSHrA06u7bVsAF7QkzaMARioASviE5pDnNNq6JDY4vCBA5g8znPSTvwsslZjmoHBRhYHsHg6uWMag9NpLgD0BQNKwYZb9n8wTbhfVDL1/hI5/xU+L5DAybJS2tjg0ywjXwsYvFAx7FP03ZBzM1uEH5f0VmJaqFoU8udKVbeZs8GL3qajm7Yz8sOXWkettbSEBcVAa1RYu6viKAJ6On49YZStIR2Qz2zuPQEkbZYWJjJNgJiovYSYHoaJOLQtiqJBPGrj048I1jz/Fo9XELoydmYC6PD9GNWf6GVnKBjgtoDKosutQVp5ADKyJjNSszvJQkmipClwOofGhc+AHPlDiPBDQgjdg/awISh0xlJpQbwMbs5gpbF9RkALCMXobUKbfqUPR8U6El+6RyqVcH80tiJyaDQpk9iwuNuVMnlyTlrAHJZQEvzjJ/k97KiZOcn0EC+93hZAzWqhbVJszFNGdEytlXrW+HRe9TGDHph1xmeketV4VsdGabO/U7TH1UsJMfs3CMMshrqesvq5KxbdBy4MTAZE7vS2uuxc9omqQjQMlJES00Q2rwzFaVpuHyuuseIZViTRPFEEOD71aiekJA3koU9WFoO7qutDF8+Uv5fM5STlJQW+ErfSrXsuOB8XdhK9k/PGSyb23A2Zt/L5TGeVkiiNr4EoTwn+PT+aHK83h8CKBWMv9Ov/UMpKJMsWSobzDjn/VuqijEp9iymHEHEKGIBwhXyhqpA2j9rJ+enqZ35IFkz0xEVGM5WGe8Ag8xFsG0Z7e3uPUmOx1mluG7z1weCXp0QxWAq5Fq/acIfLqYKIEXsaEMTfaiw05mg/3wf9Xp/+OU1qJ2GBjySzM0E45LlX94bWOHNJ0m0egoSP6Glr42Nbhh3F+ZxW6pBqc4Qqju1PMf2efLas1ZCAZt6tDIuzLOoOumaDElbgW7FXHTHXZ6Tqt6uL5nhdhw/N98wUUY32RxShCgjJDu5bVX5eAoYst0sJUFcOXw0bLZy6r5L4V5XvI/FDWcw3jMDAvIc+GzsTpMpLQggcIAQTouUIZ/yQd4me3+eHC8qyEQIFYGim0xxYtBdCfDZu/YS79DOpB3WzTmUWuz3PirsE7gAdXdd5uRX3R9gLpsK1YQd+r3dlJj/f60iUVbYc7pUfpDn8cfbDxiAX3F5+EB7m+CljPfFK3tVWQ9lARX3uWM7ZTBks6lA2sqNLby5uk31u9c+dvDptPO6zidXNnVaZh9mlHViGYbdyUJTfjp5NLanqOjL/woAB2FcvZzwn0PHor5vhLXoRVi5m6ilpIGx67OnZP9ZytAUukQVoU8n80ItohykvrlZuwV7das+otZDWyEjqOK/sEGi0KoIejoL+86snkGzHSrNYBYMy8Q4EBFRiqPV/ZMkokbIgDIuazBtuZRESU27n1IbZOlZgFsBn0zcGeFQkD/dCGFUKSMtiRCXJXiM9zawkc72wcYUkVeYJWv09WqRTs4JeeQZ1V4TXD8/GvQwB+9O9YQ/cE0AfC4WS6pamzOJOBZkXNSp4z3npsjUnbB7VmwH5vYtiU+8X5wKbhxmHu2xyMW4G+3aWH9tI5GUG6Wg+i0cXGyNLHyVahJrxa8IikCwi+yDY+Y9qwcE7SWvodPv71f8Nec0QTtnlpOlPkxlo8tCLTf8K4jLccJ2VLqY3oNRt2sFHHUOfldxDr/Wdk+MIgz1krf3GPbMJkV1FZzQLXYRhPNrf0ZuCvvjYfWuHHiXKRIBb7D03Kf47v9GA1Oouek8R29g+EnFCTMlXw3aZCO/pET9v2nhqXJtC9iNLBPlpYZgxhwYWAXfKayi38dWa8Fsh/+i+QrJF3PwsXydUTBT7Nsv2dXLs6g1xg0y2SBfeQJhixFr3A/eptFj7gLjTpZfuPJ4hPsd0nTU8RcpeuQT/BOtctpY5NhwmcOnyjVEBHcBUr2JOOrYAxdXZ3J5ow1qfYHNqjxF+5mDvy0iYQDcQC2DhCdu+WjyIKeTns1zJV70R/YRwkqzvg/eikaQsTNs5QWDyKJdJqll6XcixYg2ILLaZwhsYjomyQBP+vWA1e/WE8k4mZg66tyl9zUmasx46ErgHK2H94PPhLcevo1PjiMIPPSZbT74PW1PuNEEsSMBpxImzfk6zpbAxiY1g4ilQfmYe0Ej7QE8Aah4nRXIllKft317DGlTncXcmOI+Bb/sTfRswo+HcniKDai8hHDXy7w7cK2RPpV8huY0Dkja3tXlUJkoSpSq504E5wXU7Gd2uPM0GHMwYBrsw8iE6H+vXOkkoZ+Zki0BSI5rL71nEh7cGVhmZV9CB8AFAzMtxVL2O8qJa5S6sX6CUk1v5TuTpL8DwDlY9d1MzY3mvjxRE2dsQRC2AjhMvDOr8e5nKfOXsYeUOedKRQCXmJEOX+LoJv7ljmfWHJO7wdplptl8NIW4UAEcOhStG5qgXifHMi5KUiGwJ7YeuqcOspeB4q5h2O8nRAmuE9diW74O3ZEnK6IPbMz3GpZkxDG98t+VhSaYH7t1+v9t+wp91SG3tkHPIe2S7Q4Cgv0CMTqdcCvxIDTGNni3trAoROCb3+Wd8mFjT8aW9/dkMqERyJwRJV1xLjMZ8m7o+ON7c12nQgbJd53jL+YqwkkczJeCko772XiwcNLU/SXuS2UJwr3FU76Q06vfGBMcjlS1vRprOJihXU0qe0WHYXymU7UW0TYRIsxLCfSLakBCYbLYg2We2jGIhyd8raofAvQ78/US7YP5ISGvbKl2erYJxoaJSqboUyroXQR5uwPHHYT/1/hyNavcj5GucH2tWqWpQ5FlyXreUYfgnHaqN6K1RLhbrRWg73LqDpwFFfwi5V7GUMCzt9HINx0jWYiNbve6pq89Kx1OH2wgnXgPADUp7QDsA/nuU6ukVmdyZ3pTzSxd2FWau5c1QsSCEX8LxBQnML0gwwt3jm3JVY8MMjgLsygDr/+JNnVp3+LyYbTQqNBunXW+K65kg39CM55r8LZdD1vwl/MLg0Yd3kZuDfu8K9PKHQbuQqe4K6377qvwHAWKJdCfBcvzon0Zk13SJKMFDq3ECblaGr1ho5ocCPRpSAwIZznoI+DtMAbf9M5TPeoLEMMhl9DuGvvUUHvDzPkGz2xrDC1U3k0M+Q5LsWh5uHX4lRrHjB0moA+FAXlr8TecM5M7MEVemSkao0f5czNTFeFU+uAHLQHrb5+ECij86EU0ZSNYiGKEodDmuMLvyCykoSOpORYCu++29kBShwWDKYR4j5z37wLIijZ19O5KAqfIXig1g/+jD8rGMIbma3m0PlS27B3U+gDHzevqxpjCjlj9SXM72E6WZKcsFlrnNya/jort6CmnLYty6WJy8d40ZNDeOalBxy/bjOHt5QwOg8oZLzMvU6iufvalbDchOS65q28AzNsMIQS//82MsZqLbWwXo8DXITzc3Sm6F+53VTSzQH5wJxWJMcH5XlG7Ly55q3IRwYp3BiSKfyPVzIzsDz9EXKXKJJTTPlLTz/a3Q+Ez5eVB2vH6t//iXMuLK+3b5v20pS8Qons63Jx2TaKlDyoGBd+LkkPmWZdNGx2KwruzXwFIGWUKJ0qjNCJAG/pRyRgOzDvZcNpoERCZpuZtN9lLbqMt4z9Y4owAM2q6xpEgpQ2/NKD5f1O8F5PhHDr52ELFL6e9XLKNbhoz7Y3Tz0MTleWT/DdzLfmo/YvI1VABRQXXSXtBCh+F9aehJdickJMFLCjIBfKLbdVRXa8hH5EW+Pz3jh4ztoK9j7YyERHg0XoCJ3i5Y31MxC2vin6l60lEGgUMzv5GS+uL+mWAph/23z4oj2S4pd2XJ1GkJHPpdqHiigYk0oTMsfwudKhyLozoSqx8ADYSJZtd89mluARDcZOIkgFMOf5YojdPTC2iF4cJoB7YLIK38swSGp667nnPYLezSCYh6iIVEPJS4YGS+fWHfQ8V2bQump0ZYuHkOm/xA6vMKxuWObMPV9c5E47iMQyiNfSeIOTfgt0vwRwushm/GIWdRQDvFK5HF/YYIlMj14Qq5Q4j6l/4UDktWq0rwBHXzCT3uQpp340tJjA4xFXJjzS98dd/3JecP86kTvYgWX24CC5soYODsA98mt51ppl2SWqzZD6sEyWnkiZacHZHeieiHRB9S5S61Q/XfUr1oq9Ya0bg/ClwEfNmaj7dMeuzzqCv1wD0OQtg6RrX7EoNKMSAfooZqW+VRf7JKU+yp1foNZ+zno9LP+FvJEFPzSe4j4vGGsga94bVbIx4Dc+R7TEXNqnpGStZ5LeXMOt0vNnNQ90dNU/WqgWB5CuXvR77drzAqYopGh+BwJQSTN82mi1neOmmQJlEYs41JFkQ09zW9FwYarZTTSpUNLeVCgKA8fy7vuB1hfAX6AbqKRry9OZ3y7obEqWSsi69h+sZIChPcbSRoH0gnm/7cvSSOhX6BjlRTs1D9SElj7i4Irzg3Pd4XvkhxQMg9Hs/b9FnU4IbhxsKRItPCMwAuxk5XlHsK2z+XoLJqw0+ufqhwmk4ravLi9a5o8G0xgSMNz6Pyeq4kskJe+OVRLIKHZaG/kmGg2161cUUy6nlCU2vTYn4aFvETIBtfO1BdYubXUKUrwA2/rAdxkizLuBjoeA9zKhdc5vhSWIcBK1S8c1ptwQsySSQuXz0Ipp+mXbZX2eakhhbefkT9iKw2sHlrWwzTTKdkg6RYZIBUfYV3GpClDcqvFFOHu4uKE4AybmWdueX/tCA0esULb5lCDNDQ5w7ypebG1PTv+8eCU6xj3Uo6nKuYh/Fuk6blkLhw9iAZrD3CG4gq4b7RV7yN/1j7WZY/HKwBBqnGzN34SpRvsDp1UQI7ifuGTc2zhvdmFBcx0/11nNskoC9b+4qYfku3tBxRc/wIjwd6y7b1pzvC5yjSAbA7iYAlb5fNjJZbvQl4N95G1ZvUL06KiGN/UBzo1+dHDRtyoG7EI6K8jVp08wF3JnCb8ng3iHAgrjS3JcoJCxRDG4IoC5elN7qP/UUteKJECr8dMmXoJIFTIqtvdyO1RZMNHX+UAJd2lKOrb7COappPOeGEvmu/zUoQNfg8M9bRx4ZHN7hEdqNMLD4SlOlqD3kW+G6tb3fXvzJrYZX6v8/gaGKYqoF4czb+MLi9cdkJKCyUtg06oR/ajTV0ZO04iXNJ2tlTPaA9uxhrgpY/t+SR6cdFSJQ4RbgQ7LWQLaNJsjLRe+QQv7pelho7JfpW3GtMm5rEmSdevPOzzIHo4QmEYSq+7K9b2DmuEAatb/SvA8ArG4sB/FA1AnRqFNSP3kukBGjk9Hv3NR1km15PQvqoHiAzNoZNEFvqziEMNaN4qllZL+HHUyXE+C3bhNu+PnmB4fX/bk4pHjuHelyfuFI64aTMHq0aDFwHBCGVpI/F+sgY8RQutGK3No0CunEowrNa3gQCXqrSPlgQLY6HpbyzYHz4H6cdEk2ZDaX6lQCGh8qGtdhjJvwcREsdBSFohY45HvlRvDLDFLI0OzeAMUIRBt6c26Bw275BKjUsY//a2o4MaABfofGdMKRyGZ3CbgcS1HrF6bsEGAixgKBokUhmEGEaaqGHkS7wvNptSfPRB6TmbOG6Qc7Cwtxqx5On7U0y5ZDngME0fd5hr8Yk7cepjeV1+m7bDGpypmdVpaBFMVtj9vb7r0N0zDN9AOhY89dEyY/zLxWqB7kWYLCt8xF8Bx/THPh0mvxevgnECCUozmv+ge5Oid6g3zA1TnOWqYFsZF9PztEhQ6zPkF6ummkinTq3MVk38OfP1N7GFIHkIABs0zlKVwpEo9gjfbgimumck/Wta5HxLJNSTvnZk8Hb8aFeN9nkQOCnOhJTjXV/sZlt5E80UCK+aYeBMOL/rqXOeS53D2hieat8Ax76s7hRaC2LtJEXHWcfAy3GBsFToHKfoH7euhmxPZFXjMPRfjlDx7F6a8Bvm9KN6XRywe7RRtf2C8nzj3uUMRDZIwW26/E5em4FO5r6Nsi7JHXYrKRDGQuA+hEdzncgsibMrw1icFScL8agtnVigSmcKBj6W8fu0KSLN6lPS4yTviCO9t7yQHK/lrDsPPWXkdJofsy2fnqgoEnhlrGDmK4iMyofAUNzF7+qnAnuUaRic8hq4lwlYGHn5RsaSn0w23fP5ALowsbzNsXS1eN9R4RYIDU3cJy6MbGa9U88hcgIYM5ro5Jem2WCOKuJfAjxDeM47ZNzjzK+EWwVm2b/qnKpfCqvRYl1pVUScPIffzY9zeieQZfqUgGvGL92I1ZDXksFdfGSSWlrdLSBogP8HF+27ixAqd76jVYaILihyMKhtUYV9sdVDmgKg7Lryc6te+xQSe8oi14givdbZBctmjbZIjJQWwV4I+akRxyx+uPupLyvTwcP+fLWlFAZ4HB34WPRPwkcgSsVi93+0IRHiEcaNa8z6zzE2NvGwVgzb1QDmb0Js3/phMz61/0o6w9wCtEUfJIdBsoyMH8N71D8laIWS+ELoK7hWIcD+VXbKTjH9m5KV6T3AfGNzBcoMfAbjCDDQ54HQwdsq1r7hv1XSUz6jqgSHfAbhgYirzpmOqFVO7MHEbFTnjhxNlYn1PWrql8REQxasEWynhKfqUegWfoMSaSIgveD4ng6/QXbY+2rObD2U8Bxtn9kH+G91AZVAtevSwVdA3hJeuJRv2yhym67lDm4EJx0CQETJbL7ydEgGhDOYz9O3cSiPDWBD6rO0U3gtwOkDrEOpZkrnJ/WB/vBwrvRHRBLyFebVC7677BxFc2/rNlI+FT/CN3BAaxS8IWbGjR/tD16JZjauqR3J/yimWc8ROPTEoVBhefrCtAN1jGEw+jE1S7W7eqkeykMw11wLR3G014keCUbIU32gmLHmaownx+h3i32NBaOxmrUMZFjZsNuZ5+LygfzEN7RH8MW+itKgSEChGeSV5wLD+gBLEBLA8B/xKuDyZp6IC3hKZUnpRQha8JfDl7v8YpysTBj6dEjM4EygiKm/EKstVCxclYNfloBET8x3MfETCyBebdeimTmR0GwokKLoPlWi9xRMX+XNwzahLKevQ7nlQfr3e9WpOlU7N2MrhQOeMkYH5AG8u/PFKuarFVwU/oBxCQxCLqrmKV1eCxegDgocQ3TwpqI1MQ9Jl0w6b4ttmeOyqmQQxsjMS1R68WOlFgTWi3H8T6RxyxG9+Yo3Sg9VGW82Q6kt2wxTZkfdED1M3PjWIiWdAW0JDSne0iqet4byYA0pvbf61Z6EAh+AFe5t7YIrCPnfzV+XB8xHyKHpRyJ51eeBiL/Ywep4jhKA5vmH6hgzsGr5EMpyxCVvSgGxd8UN9LKdx3HiU0/PPz9IK+hR0qZbLfA7cFLhhAwX2aqE32JsV+X12SR9DxwEvadkhwih43Fi+Ge+pl/4OkHOW6X6o0kllumIBHZsNG/YA2kqHrD1X86hEYVdFh0yglZaRzO5sCbBwcWcxcpZO/UsYJx51WWDym74oVJLNZPj/PPllA5LxQpLWgBOY+7bbbjSEVtEeFLCGkTNw5xqKKQwDlplT2u/NpVS13RYOjhK8DRy0KxasRjNjZalKg83aK10+7JJ8q8aKP4FBrHaXWusVCUeVSEdrOnhq66IVJqOCMJ0EipblueqmKfG2NAnZI+vAqXKWFDparEnPjs6AV3kYrODP/pO5O2j/w8Uvj9dCMmitJe9/KMx0+Wkp5V+3alOTJ6nFji7m9EWxpvAcP2i6zQFQ4DRlo7bWGCHywu1dYEvZQ03d6aa1mndzFxiMEY7igjfsva/moUqF364np2ArWQl8Mpywk016FFd+T1Uv7818ibd7lkwRX6DcKN/YMuWZZyjM8go6dftLMLNcLCFes6P6y7QerUG/1xUeYQPWgCGRXsoDPZxgUOYjLHk8kqCWj34YcpRnNbS06vgRKzBEg72wOOqzh0k8Kn6EPCX3Lz+BuhScQh+AiJRL1EXzw8sGDdBDlLCOBbSi10bjuYaHGVon7oOdjODkz+DvBwF3HWUOA19nN2TVFFEkh3Xve2B6OgVH0KzpRMeWRl9EAE8RxC5ixzz71ETPzIZf80Nm7PvVtSux7RiSEjWIxwGA9TSnIQZ98YsdLzKLCwvTEWqA7jwshFW9iqGKzFARfQ11/+mjkLA9WlvDvuCif8gzXyOTgEom+K5gj+/hc6ChdQtjZ7fu6ih6JwB+9hPMxMXc6swagziqqMEksUl1fwtwhMib0TZUeTTsB9841aiAglVySnp8H8TfmTCPmaNYJFOj4cO5nzs+KV3OAv1zHFVXH6rJFFY4s3VxmDn1bDxIysVGjvn+usprzcRS1QzEzqYfOQ9NYsdnYLWXQvlGs2J0K8n4mzOhr0MQW1muuusOPn6xBE+uE5BbFk40mEwlJ9XsCcTiNLRQ+D1+7dJy/6Zs0l1szDUOIMk7ti4FQ7H+sD5liUWf8titz70dbUcq1hv3JpS65fFXX2QZ2C6GSnFq9ENZ41z+TOFw5JlHFJOGtMh8ZQHYrhnPF15/MtsnkFLvIwvrmANAWLv+rc4wIlbO4Wr4e/k5Gj3F/rNrf8UpNsV3i+GwE69Vd8CTjveYnM1xcGeNOuqliRwgOjznodhIqtToAiSwJK7qre4IFK6KGFNr6gcEYBo0mqv10qn4TAe9eGswEld3lA21OQnLF7yeC5WkcW1ssLTIggfH/3y8ayOi41fwqIAz5FluNpexUi3kBMVRI/uRyfwGqK7e3ihplacK0xbWj90N/Y1qUfWOPU0hQMmZ0wHuodifgpMcHcD672jtvNdrhvMZyqmgdv47Qv/1JDP1Ke1ALMBWVsJPt1VYvDiYlgyMBEr75M7GN8H6Cq+DjzF68JHge0CUby57frO+0Vl4W/XT79yqJWrbtWyx+bCMZyF3zBswcOQnBqN/YBmReGArk8dc5bKZfY8GWVWik15EOwEyWt/9O5kHvHv1uENDe38GQUINHLvD58ShfGaNl84ePP+Ejgd7POpqIkIeYTrjQdUshdyurXjTrd3pQXkUlsxNdlVodbKPAyXTxPepITxZ9g9ZO4Qpx4C/F+JKYfUeL2ZwE0MMGAZBM5IwXuEYJS3BCtWKFwW/Y8DP5ZIVO01zs2tufKBtN84ysHJpu7mq6yzB33hQ9c/PUeDAK7sYZGNnge3mIEeVPXsyteVG/31OBCIIdMPyvXLmKtjTJkQlASYOgsqIZB230suEXSbo/EA9/dcODGOimzAiO2I2qb6PgNwRKRIxB9oyEqOQ+228+H21lIo6K0HwdsWhD5BnJSN/1ioxZ3o/tRyycRJ5v93Epr+sf9KcXhRxe22mMr1GZHhU0P5nmjj2X3n6+65AGHTQlqjamYkNoIq3CvOa0Q=
`pragma protect end_data_block
`pragma protect digest_block
452a7579bac7c43a25d4cfa5ad9fa7bc839bca756dd1b30d68d90e0f61b773ad
`pragma protect end_digest_block
`pragma protect end_protected
