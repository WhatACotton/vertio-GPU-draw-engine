`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
dpaOUsKHtb+80bVYi3ON+kdblw+W7z54/FvWoCYGcG6b0rZ6Dbg06d2nbrnn/H+WYlwRiuXAcHOZ779iyTJ9n39YRvHGRx25jGUOHeItW2wZS6RfSQFGEsCedO+8oGdoBLDBGn/GwP9T+qkADJDYOZHNOJ0oTI95TLv2d+MeFVHBfJ+Hwzm5KKhPU3wETKD/FRWs/Y08Y+K2xQ+VNi7s74ONrSsjr6YgSj7FpL8quAO1RrPLC6ZACOR754caFKaAgl0z0pxM1fjEjnhDQsDCyXV9PWkcTk6k8cIc2YCF4rAdvO4vK43LBH82jNBMTNUt3qIWk1edKxz2vOppVEOV9IyPCoGYFLwQQ3Gu1TSGmX4Mh+BwrtunZ/UdybMCCtdBY9tI9kJBrj7HGE0a7pJeUTP9+T1khNP45vhr36HvwbmBI1p6bqcfdfBdutoCVkr7ZP3BDqMDIswOOjHvOYF+Kfeev6D5MJtQEg3zdPYWjUsN6jTw9SW8rMpkdqGSg93xAH8O5jTdRXtXH11ZO48GziGJvJeI5Kso2eZ5n3PJS6ffWPDuJHx0YMr7lsFymkwDodi/3sAtYKSXXM1pagX+wjiBfiRggyNn7BypRnYMiUoHsj6BylvuKsifw8lpbpFGkSP+TDZJPgBw8f/FpclL0aXqWbt2HxAbq2ot1V9rfAp51pppQaauUJOMli6ixTKqIz5Gcv+NNE8xRDqcDEPt/4Ao1e2V62NHPz3ut2L50HadEL1+LEzr6OINydY9pnZtMXiyzks90zBepw7yqQLGCQlfswIgJUIxXTeOeoL34BhEw+oKJdPE2MKm4a5Y+JT7iru4+pU2FVRqIglvtwk263qDNi2+LXaeSQMeT9OY3yCkaP/2fYOrSAg8Y9+ML8JNgE7PB3R2kLFtgxJAIHXZm14ihx3DUWgWl2E/CF5++LELmCwrkX2XuNI7N5vVYVjkTEczO7xp7qjcY6AwoQgIVtgIG+cEZYDYKXbd4HvuwqPm14KO5EjQgnKHLZkFHuU4plJuhtT6CDRBcgG0o8yAGOCY6gMkmwOfoWagXzfSv2GEuFuW6gfN2zhidlpXmQ2cwWsocEuG7lnWYXUrNtE2GywKcIF4YKWJ/qVkG8JWFhSnfJl8HFU7AcxEiSFBO2jWeVXqumflewGVoQ/nfJR6fiSeLuMYDxC3yOe0jnDWD/1nrtn86fjuu8ie+AHNtdQMLZh11sQf1KdGj4nVg9/ptT5B4TSlV58hN8ZlJ4l0Kx3Ku3krp2q733ufS9UGwEtaqbp1YjN3Tv2bNlYrqERZ7qL35inpZjBVLlXwcunv/AKmK2IHJT4GroHAjFzVci79X32l/4byExUbXmtdr73vK9acGieLd2X6zr7xTpeqJ7AhTxi/8mWYWFXJiKtlMV8gy9xN4A3zhmOGrLbAn477fjJa4do3ZEcynLIniKjKH8YF76uzSmVYmz3EOqJKV+orwSiXvKQ6k0GmTVYK+HN2JJb/0ryzac9ebS2I0rgjyzpyHZBg1PHEz0WrCv7yE61sQwVbVc0hzso87vnTwrBws+Or3mDpDIqWnizev2pkuZm+sW3vAeeGtx+jANuau5v1/U0zkNzZYNNIhQMa8OP8eCfO+3/nJhGqVjMQ+QjtA5w02ep2pA6UbcXv4KgCKhC0HoizZqwV0++osV8KXWi/CGbzInwetk3e1qjPbQljfihcBVv/Q9VF9yM0c/bnUchA0XEqb6YENKxuIcnMAcFbrWXorlgB1P9oJ7YWyBa6VAgGIA9LU2uAnnUOh8c3AsppBWAxgD38hLIoO6JTCQOgEr0/Gv+py7kgeFPN63L9Xt9BoJoBr9bc7mBy6FWb//iKW3THYOLyqFe4AhRdVZbf14E4MdBJs1TN4qjrHs1fkSlkEVxHRmi8+nlsl8oPUpGYtDpelXufQ7R8MMaNnpz/VRKVPL80Q0KukjkMhzgBPULqIlpBIrpgSATWTLEzqsmk2tdCw+YfG4N2hZ5bEGPZCHkmehgFpySFxOaR3w1XHsTsSO9+s971sHHRKaDGlWjt/Z3N8MF5ASw90UbCQQZjO1IR4dF6qKIFNofDc1gDoYpR+UBQkbjsGusTAA+dY1o87XxFLhROOv7I1pvDjCw4mXlyq0CL/FG+hIBnTehBGW26LCgNMcc/BB+tcZ6dqZGf0LX4A5X6+lJx+BXu4x4lDnMjhD7fJBnmgK9ObzkwsFFe3KGXtOcIzyyckbEmMgR3cl0wLAVbp6obTegICpR6Fjs9+M1b+GCeNNcorz1nBHTmaLo4+fZWYb3qkkU8lsdze70xqqxdDv5bQNBEwd9Mw3h1RmFBjxpKFR1wRlLT0aFD1MSue1lnWSSTIQ9OOA1D0VTQc51JMuXx7NTeurDHmCF3jdV+RoLdR0ubOcvQVElTE9Q6FJngoYYdy2zF9Sk/puLK4SKaW1kJMGjHHC7QbZxdbmchocgwTqvi85NXWp82UruYgrnQOjLsdz/F2P6BHQOUGKw10SSt55GPHiOh6TPoCb/vay/a932CmTqw8PWZ2JPSed+Oy6SkFU/DRBW9ijLfvOG9cBF6RNY7DHkHcG6rFh+cKD52GW+TIOPmzPM0KJwwAXsVutWpvQhRTItYOFaASM5zQbbYVxx7rGYsJSCdrNP2cZ3e2fBU/MbHJd1VYugrNVfSGYKHdVupYJOVAvF0cx0iPScDL1Sd7JSe0/uUNpDtsUjw8IMYUpchYW1ACyAISowO0xHUfiU0RhGPq1V/7OYwsEHSSoXob31bAYC1RlwfdaPpr30a4oPzkQDDqqL3Mlzl1Q5vyTPoWu1bHmele2+yuqomkY3HPWjl6QSCZF8Z+FsqmeFXqaXsmpNqJtrOfSZ8KQCNAJrgiAoN9Wi8mxUp/uEGlB45K7s3bvkVQNn3gGhflMk4ReXEoNosHM8q0ImCbW6svxIrRlzGBxzfdjVtwT0Uf1/BT1n0p9w7ObpR5Pav+OafcUE7XqTNlDSB9Gzgl9DvdIKbVHbr8BsgINngMrHHkC6o4OfYSZO9vrT/UcQmwm0xDbzynQqqJjJtuBz+6e31qznBkJsaNgkqJ3t/sYT0AA6hd/eXyfuP/zx4A6LNGbsHk0s+lAwKBoqM3evZIqhSkE/LFaRXzg576IFpOGuObs0/nj2ES5n2L5zw3D2NjvEQaST1VzmveqTJixzunZPorsA8KdgcoCXs5N3KndtrrFp0q2SITm363rIlbZbCVTg5gFvYlzkjD2BYpY9CynXQAr7v51CQlIrLKdM/Tilq9pie2p/PyXWcEpehM4gQGedRJpyp1xRvQlH1nMIefniEM27IVjySsBCHUgbncpVTygCMGmTozo8v3BlMNIlJX05XWbzurGYtVFxUCyHmV+/blSpfXDk+bfhiTgfIvjlQyE5dUW8i61iUPCBz4fTOdx/zIOYWm/ya9roRJ7Mo/rGia8sQ4/xE3A/ovrwpuvGNBG4IJA2idMtEhqnvyIwxMXlXKvSbxW84z2MNst+WBQUEgvP4+3mJxx+FZDmPjWA85kpZIO4p24BDV+zmeei4g+so9c+h1M1H7evdVX9mCq5DCRbSMQLHAtp0JVwqg/vISEE2VEfTc2ILdSpmgP2u3RWdfl6NyAnr7ksmpYub0NR4xadwv93NKA2i1HoVO0b9i19R2zZeuLm7fFlLOONnMcGOgLwWRpsjgALQRqjzU52t/0ePoz1r1JyylahbjeyjC6Fj308e08TgtSVyyHhAlAn4/vCTORuAmeM3on42jYGH5w4IVtMZIjGzHKPg4Rvbcvs9E5BPxktYe222uhFZlnLYNXxekZ+f2wr2jAZpYHhCbWWGdmowVpbZFoXJWRAn6aYKailkzHXyh4PXyjTT8p2Gzh0ll4IwzymhPXBVK0hFcD8HpLx9l78zWUp7dSNraovreS8ZySeR2oBhMY7o989YV7cYJe+ydf3rqj9FlEXjixdxpxnhGUmkVZ4IH27EUyrQzMxf9wPWmdiNS4P9/BtwPsSTMA8C1Hfk7K0gHu92H34f+gqNV/gLx7W/m702xK1yvc/cWeG5x9XvmVmzUxojOO7fEho6a2HkXhHS1Mop3uujbdetdqj6UasPTzjen6yVfEU1a/66WXUYDxQxUGRaZmCqQZxczQajertXjiDAyTygMTpt6eDIO9Qyde42k7IrHm32BgmoYVMMSgSRGh5sCRePh2YgxlwNpQVJqkWzN1yWpW0NC6K8CG5wVlcvE3Mro/JVvAGKBzTwe+dzJQl7vDAL1xEf/aqFnqDyDz27u6uUtK8x1ZbIZZJPE2X9DZLnEf7BkfSCXqg4R7hzF7VuDx+YFjI//4+JnqrPw95KNMS5UcoIjXanuZZFuHgK+dO1kFwT96iwXhatttWECIRChVhFIxQznnRn3duXYh2DAMcILISaGAKNo97Jdn1kaVw7eInVy+b8vWK3e1tVofizOBSHzuymkyXY44NrhI95o+TpTWWrS62yqiDznI+bmlzL9eaMm0R6K4fw7KrF6W7kQvbXgyh+LGD82QCqKhJs/A0iu2W8CrY02p36INiYJ0LYDy5Vds3rvULQ8wq0bAGUC5NUl/7jSLHg0EWrKxbleqeis0G7C9hEy2qi5pkV/ZfQefN5YnILoqkfIWknE4msiU4qc9ieMQMoEmGhRBtI/Nc2W6tMLom2Fors4tbyEbuZ90URnPxfOHY2UK0P8ogrxmEJtHs2Gom1sl1LYHxPphQ7QzOIkciFwlYliqY/nPo5VRvL8Z3ako8ZmnPaIsembGvuh+hlxvgpCPkZxNis8+ADscHpi/PBcyaE8V60DYL3WE5woWjKCJytwh41Kn5xb5zQ5ZeUmv8LDdMkd+xXXhNCHrq/UecPlrJnpSce39IgyzPkEfy1fgrpDZ2rwvEdijnBQ4+doDhc92sovfRwft7J7tYIjnbEozI8Jm/udzMJRNaHLxGaDQ5l4S+kssOOszDHejfgUpHnJWQ0XnmaxRF49y1DqgG6RSDISyvMyVr/RLmvYEspVHO/Q0eflZdKGs+TNcAZNZ1QsCZa1JfNBlOLU1e/Cp9M5MuHylAhE9HUMp/yugKOHSh8nAHSFNdi03ADqXgrqb7SnzsejpZio86LL+0qXRRZ8ZWKWV2qe7x3ul4T5MiiHUdu/ku6YiwgaWx3OqWc6FQSNmzyvPgbyFUdXfsIoGx/U5HXjpbHr0+C9kJN8QPPh1rKkuea96ZYK5ozXLu+C60RqXyo/h5XQ6OC+hQ/RJPBVH0dJzHQiS+Eg9OrRlJpq7kP2SRLdQd4Josv9KXjBNhYr6fvUHFVd8i8IaSh0RNkrORECmRJJ8kgCKZ9sIJF1WrBfURn/G/qs+uwS+JZmFbFT66R2ROA2kVG7C9BuGvAEkWD6ciPsYLdg3EmqulpvNCMgyZr7zSCRR9jK8QOwvR10ILVMovd8UCJtIldEEcAKNuyjPYEWQrAWadOXn0D6hGoNE1fQKQZF4B/rnleY+P3XsY6NHM0iiCPMnZ+UTpkux8CXoIF5ZSxUHCPV4rKiJAtMRhreztRD/vsgO0hLHe1+no9FgQODoVUfbBzRpgn0jqGDx1N46GL3+zis9OiwBWGrfVlIkza4WNNBF9dwiGGXIUFDRHBpWV0ya0879OgKHFd4ubFRV9lWrrKBmy8gsAZQEw3VemD30TboN83MxqpumzvE5QqJJfHattsmuMazrirIHo5Q2ZNMWQOYa6lA2ui1ldgZHmfLm7FaM4hm84h9xdY5FgJ5PCGy+yDnhNxAFc1kPb+02FHWcdD60mtW+B6q6kXCVjcyz0nLQaLEXE4IrOjMeJIypGa6yEAgiCl1DeplNG8fXMNrUMEd0nv6yuk42Za4kD7tItAgDB71Gzawb2FJ8Z0NIvdvSkTLPKOx0dFrJvmriZxf+PrcxVjwVlPTL9nsfd4iDKUAVYrlWzMLiyu8Xd93FppuIeBpfUBj9O5y7TE7f7Wys9aMDNENAC6cGfV9yph4HLGLAk4peZC2kuJdbJMgA1cpONyc+sKJTS3C1D/p4ZIDWnoiXYOJK2ui6n1V+dv5vKGt3aVORZ9bvWrmjEoEisUEaYNha9Ifv1MQdBRt9LF8J4RWknE3W9+eJjV93P/SH3WNpJJR9/OtXUMaPNXIqGnn2fXpLjtX/PUZepOZ4xWvGpyx7Vy3T1yqcGsvgNS8PwSuEHeOpwa5tILMcqKltI/nHtfwGmHRwZWNLoRBscRCDbzIEGAmvGKF6IRYSmlysCdInZik2C5qqZicrkygduxPPyNUB2EyjNAklB4iWDLJy3X9UXgJMiPOXR1VWHLFIk7YGTmhNtZC4AZ3Ls+8TllWknRFSoXmzmMZ86cgIh3f2WzuBfeOSyXbi10pSxu18wjf7nNWdn9Rq9+u62UFSwmnUgDF3KNjg4NvN/zHfwx3LlRv61OgI5edN1APifJHBkqj7yq9FrNdlpSgHu4e+DoV95ymuBa30A6gxheQ6pGyeubjUfy6pkeOCUWkpB9IIyZ/On+CoCLAnAuI71m+i7MW3k0Y9e6+HhhEFnrJvdanPAkm8lA1nwOHTn4BhhIxbvto8Ccm3ggoUNIft5mgiuPbkffdkyWX4YzmMjH1lDT6+/szXXMKt83eisqD8DYD/UI3De8XpaRoCVqqA0CB+0CGOdP520n2IhdZqFcgD+mnVWQNoPINzpk1HMJImjT1/3Oj3deBpJEpldz0U7TzjOO+JGdh00bXPonoqTArEmxDrTz2NkghCtiMoXB2/lq/Gs1fbLFf4nymP49TrMmLHdM68l7sc7+4T9G6/ej9WzUmZ4yHoZMcrbxOhJx3couh8CO1oFWAFK2o1lrcQMdllwZY601+rc/1vZHhps0Y7Jkm4qayLpB2CI4lu2glNmFIv38QbT59ArzqcJd2l/mOorQHMydryMmLGm4AeDNJ1vA458zIuk6KMTNDZCV1zaP03+9v1re2QO+AqTy+9OGGW/mGeM2oFX+z/lI/Ga1BjNG7WlSgVSgvgRnbv/lp3k0Wll1HEJSIYvcShSSejqqG7zuH1W1xfxao1vFziLCCkymY20ve3wNulcSiWktG3GjHdQNvRCDixC42tmb+aKYDH3eH1KEMetUYEjNd2hbpeMGxcC4hf+Mp6aE4boS+f7v+K2PHHaIIKDPhIx2FJiu9WvGxy3w3Z7m248LquArBhpLcrgqYRFGpb4ke2PIbMCOnzlLdEbVTqyasrfShrbbSrUuSdcomHEvGPeDMtdngiyY++gQXENtXiqM+5oyHvsq2blGZ3C9K8I+EH1XMmD4o87y3+Vj9hv+t3eVuIFBbSGFBWeznr464JaQ0ZjHjKCCke5/rG7Z02ZJ6q8sxW8+6CEx0St3bG3wk+Lc1SQPshgX4FHKJYsJ8+RfAAs0mWEg1ah6yfqlB/BekwcBfz+3RpbdtMD1sVuDzGtUzDvEzlzFpWGdOZRTzuUc5IU+9ePXVl5gD4TLErf4eC0tS+L5ZD0MATgBEBmEVo/RT9usUaqH/hlzHR9ZBP76BuFsB5ArBIWmP/xVgsJ+v1KCyUAS62ByUyLSSi4faDK7eJ945Y0gu2v6zLkORMjn2xU82R9doeeVALNE41Kod1KxJ7ls4LCGQ9c6vPiLxlNcjHJMChS892DEQX1JqbWRZm6xT0RZhssdm+CYdwUPDMpA0FFG3MQ/lvT/gKkrP3MU6FuKwBdV6DOr3IUt0jstchjAxyfShz9iJ0eeHrLcDskO/1srweKmul7tLdTyf0CaaKtUDITabQJ3TByph+BfVBnhiM1Qc1MYxJd3xv0A2MHx8BzGjPKmagHN3jHzwPpRxIpFbYrPFHW6iAlhfyb2w8+JJmmHDSKUCIWRMfBIHLgP3U+SbGOO5DjohS5kvaW4+qqcHIwXpWQ5UakQzRJZBvrK/6/lRgU7W/eEkLKdVIRwvQtyq+jUFUa9W/jra7ws8yw+Yb9rIswNqa/14KXgtUJGeCM/leydS/cVX27kBQpoVN+vO6yNIF4kkYhvI3wJQ9S85sr36QmdAy1NyL/pi6Sd0q10ipr1yXg0Er4jRc1dvFuaiwKdZpgw8PScLdYP0AVv23Go9gDsK0DRojoAeuOWQHmxH6SMoweJLniEMfa/PRXIodkh8P6oIxUL+eHhSH1w1iNhrgmkQKJQomeFvM6FIcvBo+N532ODl0Jb5x1D3yQw0iwASxJKewFFSE2cdxJzqfuXjLS+NrrM0pacg8cD3fonFgSpzu6VEy1RKkBbTlX69S1rNn0LTEWf9bmSwyMVnq0R69XG9e42hEtkF4UcOBS1v561wnXEx/aPjWa6FPugCScifN5+Yqsz41wd1w4KNk5OdZ/+VzhS9vBrKwqUkQwDY03sKuRxdKNuSpRPtcIwQUW/6RN96x8FTJ7RlZuvkpyMN001G1VmKoM0Qft571S3k2zvB3vVU16tZYJcgIXNDmN5hW+tScm996rf/KCgp9/jSh6JouFXE8wODM9GVrtMyf5MU/duMmW+DpziN8DjAJT5bw1v7r+LWPwH/UVLe0XUVGTPHimTYZSHFYbzDt/LSNYKWz0BNi9hAC40KpSJM83NquPaAepoXfgXTqQUlopE9tUK2ZVj7PpvbNxtcDNcczOdzITdSwLKcrUuIjreSmrMFgVrWmrj8oton8TVYlbvyK48ViS2D3VK/+GmzbhlDxgEPjkYKHRdzckSjJbxv+qkeUhTd0zmAb5yx4zY3YZa0ZRF/X6yIHqno9mq6JJM3sSbqP0PBXrH5yx5O+Uo1yK9U2V/KTjl2DEpG1bB487rwqIm52fqpQEixvbzDzuYXeptdadpThrhWKjUnSkfpMXW/vplzZUHgeAzfUCoM3PDLqc2ijO6jIMUAkveVrDCFlcL9l3iasDpNndgiXWBvW3u1i9ZFuSR7b0iPlqdDDqgIzIDh3P/z/3NKne1XfxSVZhOTctce3AF+8LXHoaPtJlMsRMH/9z9IuukAmHPTBoTevoiBfuQMRMb25i7PoWiV9l9A+lzikvig+ZFUiYK8MKfzvO89s5hU4M+KL+MqGuwCUi2iLegrhETzb4QaAeIw2iQRRxABtAK40Fl8f9c/mlOxy3VYTHEGsjKjinlUg1IS6EB0B0eEW0PEiloeK/TeNy23nTgx7fEA5yPTPhVm/uDRWrVIfhTSXF1OkrnLYP723PSzILY32vHm7ioYpyAf2So6jhtrM3Rlba+NvfxoaFGwGf2w4QNvjeUtyCq/hPTQSX1sD7aom6TCJBEAJb5IdOHnEPQ2V1q+pS3mHiuV3YOvyiP/gNXGdCo0E94FAdJ6YMYa1Z85eLuDvvriE5IVrw1pJL0+UOakiyzooZKGDA80FfPzfApqy3LnzC//Qv1WltHMxOAi4caxLI59BMjZC+fY87T9sVUjVxTQLpRFN87jLgZHCekKOcRJoVVjUBrwnb6auF6AnRvwApwBC/2QLDGqizzDq92nZ380FN6hR+wp6yKvFFRXlOtrkxnNRcYfwOm5FIdKF5x/volKVm9goMhRADS1/t79KdP0et6o4UMfoVhyaLgvF1u8nq2kBJT06wuYZWsU85BGArWxZfSzl4KA9WNAMi7oqPMfwK5MXJx/Xzud+XfnpoI5yDOMn8h2l73CDfWnuzc2hpzvwv0PQZXMB+u+5sQNOZ0yqP+GiziXRj99FfXy5dT9T/g1sio2uHhgzoLusA/SkviYQi3bjIgm9fXybSp2xTN0RkcWZNpj/Tvt44V58lOvhs0M7Nn06ZNo+D7N5giwunXCd3eNpO1Yx0T6S9s6RzX3eqDZIq9wsgAkW3i/SUioBTL/YKr8DpBUN3x5ar1WCtd4W60Z1sXOzJcBn5brebtKy8IQmXqHJvVk4RJvcRWcsleK3Whs2py56zFm/U7R+BggbaGQkOMbc0YrwGQk5upEL61uL5Rw5xCy51mKvaSlxfWU0mj1RPQe5R38eOovi1P9rvp7t+IFhlBVJZBoI62zz7futcH3crtLtevu4HSmQ8jWdljSF4hJjuT5NPjUvdjUfLhSV6wHENnXFuduOnJ6/Ue7mM0lMRganyZQ0thIz8H2oHfBtO6dbyqaKW3gE4vNZnbOnY0gakbhb6ypuMAKbN9wA+B8U2NdbLuj5ZNxJc9ARYVolIfD0dntuNIIFJNgD0xD5Eu8mffIcRV/TtXsFrKVn0XXwguDg+zg4LH3J30Fftp06SteT2rZLFBZsjcDHjgCB/MvLw7a4yBw8A+F1QcacTjtoyFhA2VhK2TNZMXLfiCFazmn8U6A5yUC7+B0F+EbJwmUqPBn7SRL20NEmvoSiJdxLGAnx+gXax83bj/PYpopa3U6wDAT5F2tvsJk4Vu5RCkquJ/xCyF6+P1ZbMJYaXTjBWh2ufcsKR3V4y5j8i6ZQHf+b/2Csh0HFy6+d5vOrmunuRQJPK4OiBcs0ixVyTOxmBe5E1O4PHoemp57o/Ctvri2ZVSqpAZEOrKZl6g7VkLgWJqsvfXFx97SQnUm6JS8UfxOj5Pw7IEjv/NUq1p1yZPsf+IO21/YhVmLveHkPGgpIGU+yWKhsc3yIT/wIfUTbsmTulB2ihARX6LlGmbsK72buMUudIdHEbpVWb+0If68NT/K/67eYQhoY3G6eTkP1O06QkBSJlyYc/wiwjNlSXf23c/5ADixq5t+7C05do157z4CBWR/u/Sc32ctcKoi3cCZQ8Dlgy0VKM8+nN+FtBq9mO0ZczCm4Eed/JEDVt5gjlIJMHvIgiQLu8yKdc4lUXZT+BgVD7pBB2aPTN2BrvNN0oUeoddv4WsdMIJ4Xb6NlTJj/W6RoQ1CEh91wg/bgLRxLaoQIsoU7lINb0QZGRMhebBI4v4lelefjqbCWvoVGnrK5vYe7APT+pZesRbuPNhdhUvkTkgOOYxmMzPUqYKd9gcmZtFLE2fFuZw8yNzUoouXabFfkBSBDrvpXeq4Kbn+qtANUPWHee5pcKWewSxJ/C/GrNGny8Y/3m6YxDlv/ycmbaCkDeAiJXlOltm8VWfDSjX/LKATm97zIk3ha68pMl7Gfk84xdyn2xJT8wJHxLngOPi7rIbL0jS0Z8jqnmtb5mBco1Xb5R9g079THNsLomDiIv21KrnW0IWAcvY2j71kTsiuvlMYd/+23WAzsizQyUeju7GpEjeTXPSZeMGcGIQuYrlC+O1lKI8gkdrWpjcVlpgGGPdRvGEVX++ec9PLVJk0dfAtCfl3GHNAEUsLbGBvfFMGb1k6r7iE3bVMa100DJED/cr5rT6sYGQUc6iYaV8P2NBTOe8wdX7udvccmBQux6KaDmTh1qxQ/SjqVcLOQcYS6ILm6F+tvIA+pdByXKEdllzsak105BooqaS2mMhWyp/LqJC44RMEEkf35vM+Iyciwi9hKRR/bigK5qW/FNznjAvvCWjeQmnya7XfUvGjS1tCJEKCtRmZCIWgrdMVih+7eLdCFli8U3p5r2BOuN2VxjPqrY39EN0lErzL4RFwCTBCWFeVPT1msF7lZUJ2YzG7rXF0VhEUSG3glGhsRfmBwJeGL9YTCwXIHvgI+Ol7VeYCUdL8Rxx4jTTyZEh1q0RATk3gY9yDWfFna8L7+YJAyvUB/saKqStMn3YvOapekgdej7/QwCsOgO2hUC6kBMaf2NbizWeeGLyTFZ3l4kvitv2yGNmNYgs+15nVMzLxyy0wM7mXmVKK5BXqwhd8nAyAqRzVoVR3lofp9NKbX5yGBqk5MLkzp70SUTGlQARZc0/+60Xvud3+jcsqMaVoTJEUuQEBs5nlmFxgquZ0Ci8Du/ixTHJNQ/rY2My+pxdssuvUiJ0uKfOhRYK2gQ=
`pragma protect end_data_block
`pragma protect digest_block
e7cce9f62ae4328047f78c9d6bd0941c765987ad57810f7495353a559180e650
`pragma protect end_digest_block
`pragma protect end_protected
