`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
BHZbvg3f0IyDTgkyWiau0pGOvZV+w9z5qt9Eat2om2p1eGNZNaHecKqZVUFV8GBhWH8KEm6LBNuAUwlK5mmWFi5Tj6JWjt7l+2ZeSCqshy1BsWygrcKoMT1AfyRSign8YklpPknwyiAA5g94Va5WDtAWIME/0tXADDi9osFDVMPTpKtBZS7lI0erS/NbbK9QliXGAlapNwZZlmcqNX/kvXjq1qcBK+GmvNUOuEVbixJG+sOx0NIE4ebbGHKHx6OFOO9glmcxrZI5dyPwM3ConjvWp0B0pVLYTssuiknYQ7d9gsXCpTFZrg5OOOJNGVaW5fW/95W9wHipwpvS6/tJH1izcbrpmy3f+WNXbf2+mSe9QTwBizV3w9ZeI7uDcKu7rVMLwF38mAbAfakIc8FF5mOx7s9LVJ5zaDzrQc8SJpnUmyF6Ty3USqDv876RCK2IfktGous5r5CmaJaJBlmfY5YyXyUn7E7jeW0aoubfxssN0884WZ+MGUnsnqJr/0ZTz/BdUOCatCj6b9MjzfHu4HDqje7ExXFx3TX+Ej78DTrsBng4o8qz+x8OF6Eg/2WL0wyxq2w0vv89vd4gWLYs1myesbbKsIOwM8+kXHCspEJyEW+2URTluqE+7S0K8VO8Csihoi0VS/8f/9ZlgkdOOaLGCZzDrOjvfR786n1Jk9dbYZ9T8MS3ndqe54CrNEov5PajL5cALBG8AMxzuozhBX7oWzBvHxpiTP+h9fdn0rxOezXezN/meeo70IaZOuvAOkgJbZvzuZORAWpOsLP6Gc/fsK/eE1cA1ZRwiWbltpqueqY0O72MIdk74pfgPXNt1fn6tbX5H6WDu2rmpt4JiTZNIUyhLBP3+ftxYB51VsTq6WuVVuTjH8MhrumujB8CpXbw/Z/KUa5Mci5v8dGU27j22LAn9kMilNj+zZ94jy4RZU88o0pEpvRQq9vG7QUjyQ72EazcTyMWfW7Q1NHqeg4gRRkP7UPLfpjjQ0fp8nRXf1JZhp50BrUJfjcX8lYXgPmU4KPzBwjblKtDx3uuXdx1hSMXtbYzbwRGF7IbpIxjVkYoR7NqaEh2IaE2LPGvsy9i4NAAyhcgj1whkVJWPseprHhsvHi9nhXAJproBHTO5L5Oo2v0sj4ApnJlXeMxKPsJQUbKx6I6nsktgy4RrQGkxuMsT9kUIOTeygSCgczc3BKlFIbUaEf8VMHsEJ9uwGYQrHr8vlCj2szaWhhxTtHHYzi0NyCDRZHs5ZJR+XLd+LZ9q1CAmJpSqBDfggVk/Ho07ajvat7HFEHiLIfMujvWKbgTlmAspDaJrl6qtZy+uvggIO80iq0LCVTn4C0NcuggOY0WCF+kkp2EwsueQmEqZzGd7+ABqKsxCp7FKvCWDlOba4ue7EpxgkMzJ0qQRYEmp1Z+IK7rsrFfZpRjIgqr5hOz8wuMtluItA8w40UfltLwsYP5gB8ziS2LhTWxupj39IWfBycnAgthlujjTIprQDuYx+iJSyaL2357vHO+NxWoXlsIVAuG7pynfUOgNVyxLGEutBWums7499rPr1uxsBS02+UEZ4IrmwU3FS/NnTO6+4zWsNuCHDFG+qOjdlKo2wddYecTqlwSTIEABJrChByENuar+0FaGO+y1a933dWy3BvBhrihKHvxzrtKr0O2B/cG7qjqRUgBgTJsrSeNSWc217j+rah5I2d4ANru9Fu3cCDLH8Twqe1BpeZiWY2NxdclFg9floMqngvwDbUgOEb+BIXtd+p2BxqK2Tf9QIY6KOxnUO/dgvQ3WDiELONj4SsiA/ruTLajtSJSexXUXmJT81qvlSGccWkGzFT+gbsfL/ba/GoG+lRWhL9Mg37SAMdyiojHLONJMgagUJJFaeq6+aNi96XGFFA09GS4Le6GiavZVguYzxwpAytrBxnWlMc4RCmO24FEWBmNkl4B6RKinQ+jOquzks97xQGwxQtOYu+KeCCMfGClq/mK6sYq8cOGaDumri4sap+Wh8QbZux2rqQJsqvSlHkoT+Bj9Oc7gXFEB1XpCS4aFjj+w4+ZArUhzCdjlmvi3gmo5iDG5B6ILC14Tc8yl7QO96CsvRVgNixQCstGfLqupzNxhkM16UfWaipRWbXL+abJvlfUH9lNtxbLKQLRZviTiWSrTlsaOhQ+e19aiVAO/toEw1NKqsetkCVmwSscnX9jNUBjjFHn9AKqXrlFhmCRj/2NqVFZtFsOX9F+l7VhP5VcXPShrwpRUbCxHHuuC8NdMzxHYHPatZyDYQaMHF0CcHQctuo2rm9g2OhgRwy7q2vAk2vhIH1oPiKDz28FpBcqj1UxuSG8YulfkUfFrpFQYfYbfA2E2rlZ59Aa+E+E6+BqtyACL4gvDD5PXvgOPHa+y9vpRwKbKpfKQ0IGRsQ3C8gjTI+9IwSYI6pMUe7paHXcGBW3DTOE6v8Kl6ty12V25K16cNVlaLB7H6rGKR0goeATmJc0NecYiuiw3Ju1An3THiCh5pvFwfDl4+v3qUpI92fXcekcX3pG4MPrnnhtOBgRQo8jWp0K5/jvYEtlQJW9v82h4v5rZvBeHlRr4fPTGsZdo6EU1BZgFY7aoL1Ngdtaf2vHut6aam7rfjyVtd9KXVFTDUGApz5ZZVUPlAcR51YEztpASnnDQQqiFovQQ9izU+gorFMVuVB0v/Um1oFce5c5Z6q97wg61XmE4fWIYerMnvLPSr23OdZ3objov65TaarHOpzJZ6uPvLaMSSosufNnRsXni/MAxfiUf17EVzx4Vyy3WroUHGFwgeaQHG8pL5tV1/BKvm1bcFEsaxg3BdDhMbd7KmTXZN7KIboWKV5OuzPbMjMNrIIgIC00PSSY82y8ZVg7YxrLFuB99/8fj9PA9SQlFu6X+lJ2zUEcucCz3hdZ1cbjenmUqXGAjQzslHvm4zpatG+um2YzIjUlfdRx+4sMsOdfdmsMvupyk08g//FqxmOcl6dtVoXRj3keyoHJ84dp3zIwGk29Ep+yRMx0LocwQbSqdvPvVW9Qq1OVFHiTHN063ibIGfF+yd1UfIGoSyie5Tn6giHjKC/8LKdehrA/tN5O4c4U3aKys1bLG0Wo0BJp/Q3mi1nhkwx8gacWh+M5HsplTRHPYu87cquvYT6i5SUqWiX9AhA7AQ4hxtHJG1LpEY/RDnjSpa3ncceMY9ygzqt/sywlyd5QtOKM5KYUQj1h2lqlGJO3zy6XtDFxfB8jbz4FkQb6rmkP9wQieHhuwC+XHyDEi4daR/x061CWWuzII3hSPvgVw6Dltv+qI6v0wjTbYQ5FuzZFe+IyRLlNV1opXWofWYfpBTkLJFF/mqnlNs/ls6c8qfBg9Y2Lum5zI0u38K9XQhBWP1VfKVx3v+vSchTTEZ2lQX36FEexTTzvCizAkr9MeVhDACuwYxkJy8vk0PMYpRucfzNO6z3iwLnMYc1eNv2lbEQAbu6/pFB8eRJIUnnCt9zDf0o07I4dwPloURILNRc0OQdI8sRoPOMe5erUZCpjuqKrsNKFlg+3h4ZMa7zrS9YyHF46NQHrlBKsfPGDh8/tUhfZ7sXjkrKRq3XtyQBCbriDjaWiWiQZcBJITmJL1EM7tJ+I+NjCX4Rkvtd5rnPfBDvueWPzcjWsmgsQcWvrxM21qnlCOC5DrfFYbmybVdjxwQwD+5ZQBYd9JYoi6GOBFBeAUNx4kyR5P1k258ZUnMj3M50hhCHrh/kweapbU16wX65kk4J5Wt7PsJT4OX3MbVhs3WwXqFrGWY/ubzKLsbJumsn9pxa+X8LtWLx3Hm6Kaa6gDuUwgY70Ypf4Su1ZVz6h0SjNCz99xZGJIvphuo45eAYy1TA6TZwZVBGqPtTIREPPrGgCl7ARE2TpCKNRqfC65I3X7dRuVeudfqpjLjDJ21/z9Db3T6+jBBLtLQwTn5ArY/CDlvMqsKaiU9nZEncNiLd6iQOXTCiu5zKDxACMWr5GOFTKnDF9eonA0q6r0zUPet+EeLGjH1KZnm7NLUIT/OFtJq9B/VwtzZ0XCDXVeyarMEWnzXdPHBekcI//UZOSF20LfexrFeCuEhx5ABQT8EmKA4wa5ZCdsBYuKpC8X3FyPH1sajqEIUsRE7e2tn/L0cDXnfRzuaWRarz9useSQl0e/4Kx1CbTkHH4qsKWmKjLl5Fi5eILGIziMfsLmgM9ZI8g5TzV2Xp/kJH8KLD9a1dLEpavmdokFtznI2aC+3uk/Wj3ndlmCKBwF3DnVKAujpFgKtUvI0yHAWCXWtacSBXEmnoTucgukdCtvFxiotWJ9ZujHW8sLxMrxTuvvhfaB8Cv9n7JjT6lMSIidevEMo55B16XNhW9BITLqCdSAYOgdflyFYVkiwnHU51sFRo6oVD4RT6t/9lsZqLNQ7+/8fl7gcAeR+R9Xv4gHavG1Jjkz1BiPubPcrf33TVFOBmNe9kgQXcsjhL+GbblplFnJ0/5OmsV+/0osmoko9fGNLHeUbZ5HU7fxQibu/UUZx8ZxuRr6+jyN3mE0m617+H73mVtn2bCdYJI1qMbyfGKLIMs/Nusk+rYk1QILqhjthFpRjcCNpipIFW0/1r7QfiiTVLzn751Rdmbwmkzm1+GmzPFaeAGsLhIA6InKWvv9P2jBS4s6d77u9TIhT6YNCFiwHH8cQZyqBvzLeGcQnQhCFHnVTt9meHFbyl0cK6sABzwWFizlG84VZCLxT2xH2Dn3pHw9kTdyaId3IPRcxyihZuOD5tjLzyZtbXtBJMsTOl1ELO4q0KMh7BlNMNdD3NnOJt2vJ+gE69y3oLuHFTNTM/2mDop4ivwvvaLwo6jUstN7DG2OhAzVu7950ddYVoo4zGt+llRFlUWojj45srK4CHbFsfXN3/+GTtdOGbtKIkZAnfRdjSbSuU+uLo0EgMgt33Sli4YvbcUKmQCvufNt1n36cHECDBIczcwwir+O+C6GydY+gzwcyEgMWSxydLhSvVpNpO0ouS496YRCo25/8bRYEUXXcVAOVj8ugyjf7wcXceXBInmn5oLL/1WgtnSUxU6Z5vb97qT6VmTKb1KKx/DNtoCfALlBXqe9ZLzxIiUkRkAKVNLHVWMyuO96ZgNMiMkwzEyXkxGznVRqmhD4Rvz5BYfTvsKJONZQzvrTR44FiEYdY23mfLsNR21nNEEwq8eDTehzFue2C0JNGpKyf/g1tLzVF1MSRdoZaLhsrI2aNUxHBMm8rCJ3PM0QNc8DoD/C/+PpY3HnKnS5qAkB+0ikV9+9j4Eg8/ch/nB8w2o9dj4v0HJ+D7tBS9F77Lo66PK94agEXVOKNmV0cPWZAiq+t/+uiz5uP7HGyyqBBv2SGw/t7MT/YG+6iNcpZ8FJkw/bTR4fCyV37TQ7i3sU+9Z+fHXYtkajL2SZY5wwLc+AXmVLV0RYxlobGSUEPz7TC6Fp3XLyZ5JLWYpatE7dvPZR6gn0ObjpClfvry0zMO7JEK/73kwCZUFwQ99NtjYBw5VgV3WkpHb8DoMhoPcyRbG2TWriTeImqQX6yBv++4EeYWDZwVKG0cS+OicJ+fsUrdU4pO4NkSENGui6blEYWcb3CpdjbNNtrQDoP6wrgOW91VGGkgG+zugMxuNa9JMaPnxv+KipQJnlqRnL00qC2DLyzkw2forR+D9P+NRKbsfRi6lpfkN8CyXRWyenHhcAvtVUP4mj9Wy46gmDGSGVGU5RqcOq70lDe8T7ijXezCbHyuRZI/oLAvbr6tUnAdlAIGVJ+esOO7ZrzLEW7PW/USmNsywOhG/Q6W2COs7s6ZME033md7eLwFuqHjX7c432uHcZG9TvecRHCltPvGvRnyVl9NWGkg+aiGI8Jxm7K8KkY5TdN8snu0WTxgSD17j9JPSQT5xd1lTU6PznJ5pd5YPTsHCequZGyLWLjO4PwMa1/+HcpSQdFwRL2x7i2U/62h6AZva7nLIoQCaCRzz5koQb7OkI1rkstLkStUkFl0etOLgQqTwvG/MGsvEle7LSGKNDxvyLO9dBaf4tbtWXSGWJYrBWjzT4YHg/g86+ZC8wya0tP5AL1WwujFfaVxn6nHluNfMtns1TXIYzf6Xx7bqlvhJZKgK9nMftBajU+KXmYkfTsB3Np+40yHGsZt7wJKM2KV6IWdAtcW5ORHc/PtSz8s4OKBkXBDBax2DS2vJNL5bP5eVexSjbqi90fdXERHQO8y3DEavpgCE1zPg7a1YXYZjSLV2LnSgbuVGktNWPNMn1BPZRrvymG7Ovbcp01DigHAdlroaADpq15XSbdj/suAQnWWhedGpD0yWDhj0W3BXZLyqiv8xYr/xvmb8dODemapMdV6HnbR9TnImlWOYtjYIVPQOogix22F//RMVaL29lh+7ulGvQyTIkPWVJDaIlrWTmLHY+zUMvkoCq/X5GYMRzh/SFYkYglJiXeoTeq+5SB+1NqY0/kL6dIXyZx9eixa2GU4XwLssDETO1l43yYFgeS++IV45+pV4y79GFcutvOfNF2hsDqbWCI/V/2MEqnlaesM28BKFOnphxMMwvSZ2ksGCV7g7a99Zu87u/ocpI49jj1f1n/a6jSbWM2nx8EW27SbNumucv9dSk31mHmyXKIwkLpBqVH6Q7OEWm3TOTWIO/1tObbRHRoxbYjfGEwxDolC5hMPiPvcIlIP7RXoOw6IooPAPPAoS+MWOtR6653oq6tHh9uTiOjnBdJDvy5qC70tXpi98QgLJ7tR2mpa4ObObmh5f5w==
`pragma protect end_data_block
`pragma protect digest_block
8dce60b4727fec099017349396123c312bc90d6fd246e9b357996c05cab814f5
`pragma protect end_digest_block
`pragma protect end_protected
