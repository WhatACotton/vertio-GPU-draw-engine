`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
DHj5iN1Cnc0eJ7G0hEUlT18Dja3hDFxlPqyZBngoy1a95a0NBl7paf4JG/PkiICI+R1Hp+7KUCWrRBniwlu8EG01DA73mHIdXzR8/2xPUMIqbjjkmQPY2revXHOq3KiiLx1STOPQNNmUrj/svyxVMPjxicysPUxCiZnall/mewECan5wMTMWEXOIWXGQ7M5nQe3JCzX1YhQTNtA/uQJV9LKftwzdiGe+mL3JbbrHkqug1IrG4mcmECTE6rEB/Kh8t6KDmUaktJ8E/1zIVGvpYm1c/2616JtDOYXpTDseSqo3ZmOo4g7rU4cZ/6DplE0A9zuOWlaUl88i6GHzZPcJxtOjb/AnQtwsYLPjcROJLzgnmfz89Yzl3Jyp+JkYgp7hGZr58tEYFJNZsF0nTYSm2UTDz2uA2i67ggRsOj42RWpm4uSAqRUNsRfbpiOyUfx/1BMJ7dd5kkS2nQQb8tGpnX828PM4ylVyWAgnAP/mzt7FRp2NGilQq5BEh01fDWlTxJtIsWXlwkLNMaBcPZhUjxRYpDCl23drtnk+CJLdLc9I9CcI+u+kFpxtw6/1eXwrCMRg9JfKq2sNLswfklcF1A8BXH118aX4E+cNCy9/V+7x4gUNhCE4wgMfH51V4McxjymmWtkt3IPVEtNX3oLJROLKmIlauxdfvnChpI+KD1RRjzinWq1IudqV+Ex+FF3lOIwpJpzz3Stycu6bcDZGVnWqBGVy0LjQblyi5iwAQ54QfXOOPABu/uyma2MQH4HlMskrl54xHKle6rQ1rHkd4UEP7lpmIoZBWRVfMHTKXPStG9c1s0+MG48cz09WitaROk4+bSvKJvA6cKm3edfBoS5u+UMk/cPQDFkz2IywkaJWum/ausWnCbfnzkQ1q6bEaNT52srEvuGwzxa9ph1rmi+sR7hZtZPs76Gya1DGnERTToXZzH4Ei3IUjqQs33iwLjiQ5H4p/t91To8dNXPjnsjIoYxm5gGJmmvudJMIeCew8vHu4K+yl4UUVCLK7P19t66e9PaGzo8qCAZl+OXjI9gth5apPHVcz8pirmMVwwb4/Ywv5s8aB2hpyyMdJAZHraYkO/XciLJwwFKxi+/EYRSPEBqDj/pOsmeFSPdG/Uqt5u0h5w7P2T/tTrcBheM/xGgDwqpYG4YB9n+gTjTKqnmQN476OuTFEPaMdUN7phgwlvDzELsBjII6gHtXMEtIwLsMSvJxk4GVi63MqC62zeeDl5ALDCLWv5y0yjUQ+kRrXJRzKBzdLU3Dx9uhN5RaR4L4+b36hB95/GpC+gJ530eQoK4byaBJ5vkCaBp3Lbr+4538AtESEWVGp5eqG0bkBd41z62poF+nkVmHRCWNf1ZmWJAkGoL5k+vSh1J7ClM3Q6nQ1Hjx7FobfHTR0t4+riZVecn5JigTmQibox4k/IzXSOp2hJ0CsFAIyKE9uw6ATQYaRd4xiudl50yUxud47tHpijsradtpGJ9FRDSdENu0MObSzJp5dyON7jluAy10xxX7JW7ik3/UD/wYzrsKay76IVhXCbL9VheX5QLzutEUvQCCA0mWUWVxlDRj1nhxUgPof1xpEJcP0pn60ooZQGIdRddwEhM0id8Ra+MRaerke7p7yCLyONULaXq5EUS/m2Aw4qhPBRkJcW3GL15uxC8f8WHojE1dKNIsCv9d6dFOW5M/O3BL0T/gKJjNCzB5Ho8mAV0tg+KvNOaXOLTRt6A61zvFUe/fjg2xgpK8CO3m0mXW1kHsfghWpTLn0ovu9ayykgNWVnth2vMpv2SbBE37FqvryVf4r843cKB5yZzgF7E5+dHTs7a5H2tPNNI2kxjEQh0hSlax6DU/JmrNr8NtafJHMvMhzwUhXSBamUGgbiW6HgkuH646t5xZnCdLtNl0HEa+5BHRGWzbNEXsHR6y0RqeoxniGFGs3M9FAu8OuQlyvEfvrcbi7gzVUS8CGuCbIyQ2wu4yQeR7nxYsokTblqpDU+S0VmB+EGF8X6UvAH4DDn35KpHBDKencW/pjCPu1py0QPM1V1BhwoyOfft1fZMWBJbsQGGp7HS8Hl/2hVn8xj5BOaHqVF373gp0xf1I/I+AWi84UHRcFlXzsVmc6DoXO/Qse+tzWXcoTjS4WR1updSthq4oW9CR/L2gHWitRKtfDnc7bM/TcGo/5SC5jfOrvxBdmSsJFTRF3ju5qClo9VODEWzR2mmMQ+Hqe+F3YVRaJ2zNB2rF9qobaNASBM9e1esR0KQ8ddevol1lr4+WZOtsiBV0ca0KRgeaVskoPOpJ6oklJzIeEaKL6lW39h6iZ364WJ3IcHKDAxSQt04VznudqX4ol7w5Oag1ZiJQgifbS5O2fbQrCA9NhgBnMM/seS77kbInFxJBHVM1IRerOf8+tEBR09oa9AqBzUVx/Va3yuK9sfekGAm6sX4wfH3VCBBYODvVX/QCPxDaukIGp+v8H/m1NUyTzgDosL36AapLfK+BbLUZFKM4/tl7Fn3Ch3FBUbzKct+oUqA9a6K6Jo/49b/HllUzqjb2lluErby3ttClloB+jrtlu6rixr9oWOXp5gMAOQ55T5YxNGuqTyFXVvixCWGVRtbegagZYV+CfrC30OqjPj2FbBzDmJyb2+tluSoFR6MHnxXZsQF1v+XgAP1lSQIKsyaCXGjXjM2GV/hCNZJGRF3X7u8P80R7a9fEaszsDCQ+mkClQ64DeYAOAPDfTj+A+4BRj4gvasIR8xpJyEoQ1vZ4bLf8V/oLifPnEJfsZZfW7fYieFNHNNXSTWOmaMBxYe7RktK3WvlQ3DI369t2UgrLAsRXFWxuIKKWaMXl+OrzOYAAOSjGl3nOhjCVQxuCvWdx6GVmJzwOUnNpJxpeOFE7xWpYN+uC/z7JISDbzyapvx5tuWoXf1ixYECLzm2tfif+0SwJtQrskwjrFLDCtamTy+XOqzYqUigqwgLJTxippop93VxhGe8ovPNB+fV+fxvMKKbzIWOVFC2c/qBKdiTMNn8xu/1s/YbLk/jt9VAIGLnUwlCb7AYq45FZ1AuO/rTfONjzfhIBrOaG0sSY2JC+AIAGZ1ZD65HoUpTdyp2ZhQJ1vePoGI0+ZFWpIxfz2I9qFk0TcP0lpkVMEDUuITQGhtEzS+bt/zMndwHuWz8HTQO8sI6w04ywE0iJtosVjInqAP61YWScVqd7cG/PGd2mbyWa39z2/Uojhgb01x0sjX3T29M6oQqqxqXZqKz/+9BVpBC6J/wtdeSkQHi/UWWJWoOscBwIiFbVb+O+93ygL8CWRgu1aVQvrbS6fWIDbjo8TIA0rniF4/+wWSC14+v/nTg31zha1t70PeLqoFSITttd9ukXVIW/tsv8flzUjXTBw0p1l16sARe0oZP12hzdpj6jOnlhUj0ZdNUWeZz1os3OwHQv3hkIl5gR1+5yu/KjJWlJekvDSqX2F3Uhvsqa5lKzQBkq0fQ39Lw126znG6JqU0Z+eO0ITPlu4xdW9Kc3wm2mVP1EHPanutdDFt4bISGih2lyucLbM5iJTKBHGvs/rb+X1pE79MHUNWFEjSP7zD3nhxvisbB2B+IzdMgL5Q2FZKd82c+hX1nsFUIp68IjfTi/jyItGcbatab4ZRQa1gUIW4ogWk/2wCLUf0pYeFBYv6/g1bwPcvfMP3UPdqWGs5q8r3j0n14ohQyc46ku5YU/zJCjFGBjB1iwd9lqr4eTLQ3gx1MGCwZU7hGoil+4ToOdyXEO26/GcVPqtp8TepgJH8z50wAfO16PPI03vyZIfdQtL72Kuod+3/iX17SSg2n4D1WRb3K+ez2HQKafnQZ4k0IUo3MksmvO2XYbsjTCM0oL52D7eU85NCWvniK4zpKz5z0uS1F66EHPciiG8V4QCuQa5gjviJmrA7o5w2a7+y2ldwr+eDE+0FFFyAUVP/bCuBtCehW/M7kX/7GfpujGEdQrZC7W9auKAV8R99lMIWSd9jy3cyVvkgktf0o/RdBHlIFDaJBrWDkT3O2g7nOtCLrZ4vTANNXHPE0nX6UgMIOloJDv33zBGKaBCPBvojbSU0hC0rQe/wr8LyQ9V75tvibWdvE9VxqQEqxUvFvuyvpsSf1IEMjE32HONYdtJhIrw7ufefZtfm1TQ7jc+EGEJDfP0SyAUpGmIPQ6l1SNEOqo/J7/sDWBO1f2qGgEoVrsILBedyCdihrTYI6n9KKDn0Wt5wyoCEPIbblhD6Be7+/HFZ9YXHL4rQVufOdpwO9wtcvpVo/YVfX3PCevyV+080Vwbz04PsHqEbQ6zv1IRPboOhOv2ECr/N2hkR72Yp1M/MuXKC3NOCCJyZQmlGV1BwM2mj30ON+fHtMQ6n+zpUH0xLYSRYzaP5AyqWvYA4qX/IECiLbZP5QuqPcaWtguG+Hzqf095QeshFhrEtyuUYLjRT1xFHweM9YUM9GiELIew1W5TQAZXmgEmbpiW2cE2ocZ6wVc0TrBLRkCtPA+yh3pP5mxWNju8tj5Egc63i+V3MS6ysr2Wdyeizk3hBXMwrabQgMhNGE8+I+0ZisM+FAQlYTjuYpqHkKVvRfLypxu2yZ85JgltJ2IBqbMWHdWebKbh5WyG1A7AmNJCdpQbCtrWptQ54PsoizF0SQm/NwFQzy186skRBEe6qLHiyoXke99ZAGotrWFhnlmRuhOiqkFOB+dt8iAz6ROPtbGWj8YUNKqfx9tD9OXOGLRQmPsdNQaScywQcWckCMQjKApI1RKIsfFj8Z2ViSZ3nY0zNbUgA9blCMpFw0EsijMh+iDqNQ0tKY50Eggmmzr1ovF54WhP3as6AlLsk+rQoQcfZaW6L7Vq+eND7q+b8KFr4m7WARzd+zAmIFLSB9MZfz2vZ4iF4osckaaFplIiYEc2CMpKdGVIERrJEQulARicn18phcWeYSIqFQ99Z5S6xPNkVwsjCXGeA97E0ijKg9XjbMxG2kqMfwf0XoiOO/lnI6FCeKaULwThbOCgXoKYS7AgFSeO8VcFs2wwTOw5RqUjB960/CoPueX3Jaql5qUNm0zOH+HE8ylBFRqSCvb8NIpBGUdfwqaRJVA/MlbKlwzTvqxc1Kf0IWLA3tJBquCBZCG7DDwtRXxg9PlxAPH0XKFaifFf7pnIER1SyPL9+Wp0ljd+lYj9L/PPADy0KzLyXORZK/lNOOZ3QBk6V3yKbLoNC38ZR9HmKvIRmIOQRuVOOo3FQcEavMHXDPw4arcPRFarWzFAAXisbQW+RJHMpJ1rihUZx6cEVZQ7A0YCxMLgPCCYO5KHe62dVO4JVApZ18hZtp75w4+3kROrFLIztBVK/SIiq4mGU7B9LdR9t65wUaoU3+lerA/ulce7+vXV7y19RWtmvxo3iEZLxGg8UYZBxEhFQd0ET4JxqFsHAn8qzfZZ1u9nb/7jJh7sPpLgWNi8h+Esk22FadTt9M1r24y15l/pv6gcRKTDQTkPGRZEv69IogkA/lK6PnMOLXuJRljNhMUR6kAVmZZf2mEe+P9wkfx2qErUhny36K0uAzuAdl2sHDjz1sQQcgrVbpv6ekAO4RdA1qMJ2aWHIRu2umEOKQbJVx0Eh989G0qIWGiaosblN2Z/DW2wvCviPwMBwOVOCKhYiNneArXRKdQMUb6op8q6yBk56PNpzT4ZFNTJ3RthCJ2UZvayWadxapYc0e3offC4ghH+Lbd3tsCgQDD0EPBIOkYKmz6zvvSwx3142mvHRueX3KV5iV/OvLZ31mqfb6q0yl1As4yLhOjEoZ4OelKZVFGhvw4mjO4Iwe+gyAcLbke0ktRKgy5KzOpmP/W3lPp9F/ASZH7+Ev82EbJ73zYnANpzUw1ErI2AFZJp2PVL7Eowu2RAqXFzWzUuUjDWmcLwl36aWF76WGw+gNMoch4XfCdzM75A+4SOl+6c6TTF4/9eW2RQQ2b3qym3aF62Im6hyNZN2bW6dJA1qjsW3qAHb0/rqwQZ9iKiQZWElczeTsw6raMhIzh0Zz1RN12p6rMzkReLWS+4FTEYCtIEk8s4VKhYoG4Ls74qZLaN9ykzsTeFPoswlYPsyjQF/lYtnxtvIO0O7BlMs55SC17i9oOKi9AvS+hZFG48o5ROFcFBB7cWPGNiNSc7tpil7A8N/3IT6e84rFo/79OkbFfc4HQOTYpPHhNcuK8xlgjoE/NBxDXYhhHOfHtXHx/eiqxkNwufddMlSAlmC6ADbCA0Qu4bsipMppaEaBs5AQJs++wIiqvj55DoSo6FfTP3CPEEp35JrD9XZWw0W58eMQ8DRqeueoidVq4HH02SSneyIlgGHuGpZ1JwDnijTJVCdXxnS7J8erw+HQg5JdoS0vXRY34frWb6Vdf8Fqm8GHh6OmonvgvotysFNNp4JbZScmol+QWYtxwZ6G4DQWTCUpDm/Bg8P6MkH39pl4nktdh3BKivgefX8cEwozXKmDJic0O5YopH6KzID3we31oGXU2Xwud0bhfWu6dsbIqYNThUPEADprgb4+SOL521fNY9mU+cFIKi2XxqGfN9wQk05t3iDRzjrG1QrtONnew8W01wh/rDSIrBpPm5jqTvulg7BVXntKggUVW9le3np/3iNUieMuopbGDaQn8c64l89/Dti4f4F3LnplQeJfUYc4AIfSnkFI77tW13Yr//SSy5W9f+kbBn6Zuxr92K4Dqyvvqolwtx1L2fkQGYbXYCaGmJIi+AirDOF4T+DGOX7JhdD0Anfi1mX16JzEy1qTLXodeFesQClWOIkhS6CnqnKp9z4DUCf2CwJ+sjSVtgavT5nM2krdIFcqomqkX+Fl2lFs3GJIxRoaWvqUsMJHxteVav0rNyQ7hwaIxgaEboVTdGcKlQEyus+IdhVGBAzgUrDJ8HEm/+BAZJlbWsPxF3Y+jOX3I4yvkQfSkNkQGGxJ/mwalMbePdnt6D+L8hw3IxoZLXjsLVfyvMSEfP04sge6tAIaRGe9RbZ25WpzOiLGGKhyWSDJgTUBbP+92TvdQixH0cFLddgDSqEe3qaVDeu/cAD/ZDJQv+zynCXGombwpLBmQPFYRRIHlokiXOLtOD3tbuRLbHM+g3fyGrr572/QH3yguVPmfM4Pz25+NDMIDCgXf42BV2NSRCJQRtrUyCWcj6HAD2dog+CtgiG6zOn3jobWzdFLQC4Fdb3PZptyAdbkiuerMQMas0iHVmfehTmS4qEE3riV+1XfcQ3E5iYAG+5iROT8XHjjQ50JxlYlsNAC4nnKbc7+rxP3CJ2G+rYQYY9TjeUV/SrzG7l++HvcstgF0emn/bQZWKksn8wdKrixGEUTD23+oT6QFL4R0q0Ng2lougYgoDtJrYCpH2LgpYkaQbs8F4IaPFvTbyOirDmAlND/pwHY2KtDRblCXASGpHCxQdblx0qQJqqm6/L2LCKtQ2o6MSRGeMwKVDPhBgAoK5+Zl2pyJRU+WDiNN2bp36FUCSWD+gIHZUcH2uRNrA0j8KcBZT/R32tyiDdf4Li8D0+Uz/evfaAPUdudTfUDmxgZQmW8kHbb1sIxvyEF7tH4C/hJ5JHQfKrtNv6PYaCZM5w4z73NL8kRhNaYxnAu4UyxjkegBYKeYMTlDkG1znFaOZc0Yr2gv6UFXDDCqZuKDFIYCavBykWiBhfworoEI3xxKiXT11245i81DAlUSWspO5eN3RTAEthSanb3N46CLYSKuCXs3x4jos3BPR9c6K7h5oNKJ2KtIbwA5pGOIOE7l8n4SMvD4REumVLhEbgvl029GSlOdZ0ayLJxCxBl7jZuuFHi2AoxA4+CmmMRIPqpCQ9KNU6wj/V28OyQTGEW3RcJjGXZyo7XaZ0apj8PEej6PYY5wYf81GUEvCZDRIynC7GVmsWRH6w4ALQ6VoJ5aGqgLwvKIPf0jAa/Quq7VPoA4fJ7FmNXc0XnYxKj2oLErVv4pidzZky7Ai9RNyq+LcAScEX7iiiAxkHHBGZQagsiA2fzbwTn+mUV3EVkDAzMl/m4vpf/+sGZ9sEClreBXnJJk4xSVDjUm2CHF87Zz/TXoCoflyFMSDvNlQpBsNc6k0XuB7fE9iHf9pI15Ehajtvp3Nf2esZBVDub+gDhP5zjzal9N4+viI6wIhc8JPfD2eR+ZwsFIxpW/bz/2XpZtsAcH4RNLPQJ1L6C3U+CBCqqxex+8bft++jhSQ+8JNyS9pOPwug84GMPMNp+OCryUrkT4R1jfpjNxKolDGGlWER7kPMt1zbEs4Ubrg0G+bt7YX7WIUY+gZ0NpNykz7i+X9CBZipH+bqtQ/BfEb0OI0pxS1pifxoTZzrst9yFyP0Uz06hMwVrPa+agc/co7DkzMSD7cIVAlCUL5QTqOepm7weddiCN4rxdyKU3NV9ysBfATQkdkDOxn/l8CgKcVn60lESwYITqid8NtWIUIUub+sBzAHQ72Co/4phfLqXFgW5R+8r/Y94G/3AabRppSrMoiw+Mk0f/4KFcot5B1QITjenKTSGOmoArvveEkvu4OC7ECQoRenKBEXvEDjtd80wWPnvBsMze1xZOglpwswucEuijRpKGG/ugmhZ4d+YMXKYQ1b76cx/i6dlAlxtxPxM9YA5JE/RBA4BxtsqDsIhBmSodBqsc/H2+jL5FgkQipVyMDqzpn81RO1PQMCjnNfDJ0Vf+LA0zrUqBqGI7uKdafDA4tRKcPkoW6zSlRCxJ+D+FwqaWGxVLf8MRx40jC62cYOtuSZT1VOXaUfe3pvybatcAzjvGAP0XDOBtgUmrVg8VaWapTN7/mQO5uBia5eF1lmP2goyumXF00lluT1rxDy/wgcqU5phwIQqwYMhk5lHBKkfg0oZLVdPOuRwAdbdAEJMaoarWXQQxf+u9WROyxLu5oBbOod7Cj+88SOVUdZ+vMxqIupyNflkWgGgQbtcmhiDS4ZAYeWJh8isGtzlnaqzLpqTtQnt8CNnfV/PkwLGnDY0Vv4/vzNV8hQpKgvF7d6IrCMbLhmFZ2u1FQA16Wtn3sGX7mZ7UuG3zooZsfiUnpJZh0xjUJFnPEyZ9n1Wig1XBLQumY4ybNoYIDHnAWEstkqS1tmVEgtSZRYL0FY5DAuRQzlOhBrGa4qmXsHQdbWChxdHppESeJ73NIZ0cdaHkOdtaK+P8tXgf+Q1WXrCeUeNV966PvxG7nSgTBrYZ5kiLaNtkoKNJ7tfktQu6uueaJDR64iIIypGTDynCNhZS4SRCJNh5nmdOrd0sjGZ1om9ch5FanICDEiiyis4+KI03/jbCPifvGtT6pWo0qcy+bHdfpWhBeLxGBg1mSG56I6Rj7FigjzU4NgAmYMIPnX7XXu93Ro8I/jJOFqqijv5XAgEbnddx072azUt0/+LJ7jY5GZUMP9e09Nn/OyJLBCswhqujA0k4Ex5FTzFTApXhwdi2IIF3f+WIo2aO5qbFxXT1pZXw+V+9anAZnaAAG8oJ8bp5aLLqHCnmzyqRpYEXYIp3wFvSxUWPxCy/x+oBt+gcweO7kySjKWyU5iPWhi03YxHBRgxx2K2L694qG/cNyuok5tfG2XDl2JGrDnVuvMTjmkqFOeSoymxRtguCOFC9XSmXjlK2+B6GFrsazjZBOYis3gSQZfYkLW4lRnNYuXfzAsLPwfQdnWGUGtQ+1sxjk+CA5AI3yHFwFRIj8NkzhBB9nF2YT46saLvftAenBh+0u7nJHvGLuMKqocfXxtF/ALrLUpqHIFYmEVxDIUIJzcgodha5RgngVv91nYHTkxW3ykpzsYIhCTMXOrIiShibY0neHX8c8yXUj37PPuh2TjQAZRYAqm0WiwNh7IKVZGBLhpwvyd9Aezen7CT3AqI0kMVcLq9UjzTH40lZTj8k8uPzIpWXHqx6Qpqg8Gj1qLKMX1h8LMkw84JNmjVKExnxJNmDaP7/13/mHqAyTu1TDJJBldAAyijAQzrkUS33bzObfksiE16rOms5rWtoLYWG4mtNtxXpZFDVv13NsGJ/hjlXOoI0yNZE4HO1LwgU7iPkDTYagY/JCje2lsGdGtGeupzH3i2l8VVSE+O9cd2CYfHJ4ZwRlBEv0EPpcY3lvh6OGbQJXuY3pWlbWqTgsyhe8MuiW8vCGcdHklIpOqNU9Q+UnLdzbzqLBbaDptHY3TlbloSyq6Lq3cg70oqYaKYlc73jJohNs0qDbD5e7Zj1O08oyJnT+QbKKjfvQ8mBDnLCm0Mnf+Ep80Majspl3XGjL9+B3N2Phpno5GcqOtpeIgnvwojkEXm26N+jkIaJi67MWUZTAQ6/l4AgA3W0F5KgSIkzt+wq4XPwY7gSDPYQSeCa9BZ/X7qGLwNo3nQavkZ9uo3Jwn+/zf6rZxLIK3mtgWMH1C+hh7MdhGPQCzsL76ROjdxeXw1kMoBXSGQGNq0mOm4N591WFUv3a8koupmLSF3qOIzg8Nk3RZ6+ZZzMz7xGtD0iECSVxkb3G/nhvtwoDoGC4v3Y4jwJtpmdb0V+l9MLZD5C3DziTWlK0yQh24Ve59y5Q85AmRHAhG7HwG0tTqn46bjHYnaC4/7XlzRT3qU+WWi+xEtaURp+qY9QcRpsYgDWobHkHDtxk6pgep6k+jZj39UHOri/szSQVraTEvFKE2tvSjQWzCw3BpTj1Vm5HOX5PHAvSqbKs2u+CLooND2zNlag4AOODDS/SmMxQsVrS8xrYGH/NVD8soIt8IoOoyGZTF+S65mWFhTo9PVrTiuB/M8b98bRO5CBKDJsZKXMo0oWzDHkmvNa2ZJ95zQVxoMFTWfnjpbAW3I0hzmjWm3cnKU8Xa4XLGw9uJkoSbfLrj7DjmzJHLscH7cp2lpv7XgrAbK3IDQxprwfWL/+NxgdBkdL5G6NQyrxGZpo76Vxm4gputApXHYi604MrjhwKxxZlie3rKGQuKpIOWWVGbXsJyPJzguBZ4NbxdlskAm7V1HZijo6pG/dm5FDfEKTvuWyOmhOF/OL3LYIABpnc+DAkt+YuY36OOAQtJpJqZJORkt4P8JTFTEzdJ2rW4uE4vVa6YbIvQvVhDXCer2YayYKc+kVQIrH4uFpCvQ67A2TwTtov21NVOUGj4XAVSSQb/RdkLskmVI0dd3PP36rswnF0YXLreTu+vKNcXPQ3oYhuqFDWFuS94GiVY9HeQIwaJGZFAeCC+3Y0RkcZXjwQO9HRjksF5vF1Fa8BF6/Vh+929roXv9nyPk1F8ZW2fTK7gTHz1w/FuUBiAdsuB5fczJoSLPzElzpF1CIuv4AKwf9axadrApfAuygiMxHTQVVWEQjTuhb82wzuba3+kHQsmCw+qsajPOgeFp0zzoOQMsi8OpanJ2AOtPM9Rt0sKd57uTrLiottph5/nwQAZiwDm11NpdVTUD9E4DEpAbaTv1kdM8p6U3F7IxYvd75BLs4Pew97UqMOks3TqaHaqFI6G9BtX5qpBK90SyqcVcaelHJcjYjSzlh/Cx73IsBLMCIF6/NY7I5x2B1TTe6olZEsIJa6ZIhkuUtZ6LPDJ4VBHlaSfMMdpG3f2ylz7ZbgSe/o9IWP/KzD9D+a9fTl0AGEgfrvzZP3ZAmFzQiqfmkAfDJSkC/YYnmaFdyW9NfoBtN5PzaeRRhjbUf/SH/z+Fc2j1l1IJeD9jikFNfHPgeY43I1+liHDO7bIGth99fhuKtVX5seOPaSMvZbYF6aK6gaHxDOk6Y+2JQ6AyHc77CpnKzMUj9eWU64POMqa6NY2KTtSlZyaW9qcH7tRd86cGC4HJqRWIs2Gzo58TIalv1k90/E9InvYKqX5MiFPUQ5cKv+qToczwUgcCsaaBL0XpYcRrm6HSGi7EYhQ5OdoZDJSBg+xRZYX4ysVpBz9AtVarzGGSkDL9LV2YxP+mT5Xqcf1slz0fIHj3bvbpwHRQwoc8fIFGT4+2ZSj0r323pvw3K7Z0ci7fdr+vO4M/ISqPZhNQR4SYuTMiDxruR0ODpOOqiHopcMa4wiZA08XuSEkRcQlF49O0JgYFlX6HlE46+AIHi6Mt+vIsxBB7HIcBWVgOj9yxTRe3D3QBBv2RF/bDeoHgQv0kke+IUyEPu/WvOwoGXMZU+9QXXZ9MtOkUL9JSM16GSCQz5HLEu+f5/g6HpMg19/Nk1CCgTuWHU7CNLnYwi74PHLsyX2U7nedyfSOuvefoxFYtHgWmKMVkEyZCYY8NVincU0V5IsEafswBdNsnM8qKZa4ZuHfslouRGpsaOL33t/cCR+ai1biTbf2l7lHOjtiNnvUBLiRPYy/9sVDZ3ITdQO7qTtFGrzMyQlnpzCTQihvNV3S7xlQXdWZQF5lc/IDOU6SXBJjnNK+v6STLy7jqWxSNpvLRcxKRgCmSe4/Jvs752CSAYljPFm3zIOr/KyFT4IvIZ06JoqIzfgA4hj9MpbYdQB/CgrA880WEEHLfmHrek5SZJZxuRTf5Yy/A0x9xkoCYMgInFJGjkWfrvSFf+vhm2HcxHcNXlmKRZUCZCk9GPAaJup8ESi1+dr/gMINd+FQKHF1U7G49fIH15K0Vc1yzXgGiVYrhhVQG0uoViuzYKp5eANJZ6YmwvooXrbDpSTmUU8+coeZu6HOq547vL8zx59/yucweF7YgU2prRy0mKitKeQZ9QJUKl1admwUa3tJlO/W2q8xlk2nj2I3HWQuZk6EC5hPtIq4IXzsP7kMQfPV75v1Eiz6sixr5SGOASrUbGCml6ZKE4Eg6jzO+4RtjrDl99Pqb5DEejf5ZWEDgojX5nb43lOVKLWSC/ZWIIrVBHYw1Z3ddATMPNee4AxY3B/9iCwIjUJzB8bxi+fbWTr2Qtqr+5H4OI9RLhy1AVvhQI5ERcse5eaSoOauDJcZgy1ATldTA7UXRt1KzTCW+xgg4=
`pragma protect end_data_block
`pragma protect digest_block
95f99eb51770d93a1acfa5f6d6a19d52c5c42a594a23fd4743c8214a78fc6c55
`pragma protect end_digest_block
`pragma protect end_protected
