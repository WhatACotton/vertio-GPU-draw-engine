`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
Hbzn3QnWJvWJxJzYxnehXgCkhBgW+4CWYyGk3OtC0JZanE2JtAkiqmW8jH4FroCa6CBV/D07xLov7/H6EYKKVh0HLK3IodqBuveEZbw1/bYfqO5JU/HoA9bRvKxVtPToMrT8uCgmTP76Q/J2Qy2RZlN0PUQcYDYidxgySTPGWeMoXv6oeOenv7ke27I9Ld1EqAlaBT4Zbq5HU99jVBryd3G4tJAUFzElVVYOTpL3ifQBgb3+1Umun8ppmKK3ShS3kWsIMPlpXKcGqY4GmWHc1RAXwe7ctdAAQw1m75GwSiW89gKA1+vF2MdCAtcJX6OBs2I3dI1H2C+gXAZBrptIe3DCYaUnR4wy29rvvM7p9jt0DRJdP869qmA+YsivgQjCzOjafbt0sG2tesSCdCd6ORK+XS5cu2ro0AapGB2W6rJMww5NHIbZxGpEKP41t274v54kYaPJm3Vx5cbrRg4WOnpmCx4HozcAoC9MmVHvq+4WsdcCGMYQ0ntbq1EMKMRNHacxQ9l+pasxhsM/NbHo9u412TV+7ofDCFjWXhmTOeSR2ftzpxvWfspJI6vowgqqBF+uXUta+oySoyo34hJZur8Vl+er8qawvmEdpxe+H8g0dVlbjFe7n3g3s6gu8r/qkT0L/6E3wyqb1HkoHHSRDS5x23X+yNWmKSnUGTGb7iwXsAercrBJjGM8IZQh6rwo+/qiclpVSw3n6N2tLb8GvVrRtRAsQX5cHXXcEY0x6M1COHaOcA7c/6XNawR+nu9UGasctPJfywjnXOK6ABYBJ1qObKdkwsUWIRBLBYKQ0fcVWCJfD4Grc7wFBrSizmTpROCb0umW3BD61hrzWfT5Y64fZuHBhSDS3dfJCe0gpvCn585PouRl8+aX5/dw8A1WaGegjgLM9LIgzqWHUo6swGMcKjqS7/hWZTYRjRBpfTAKhzcrvZZ99DDzoyIpE8rDNSmHmEkv9Kf3/U/jY2Knovp1MHyXxsrD7FHaVLdoMMBwSpyqehDC+njOoe4+5gqR1OCbC0kv79DQli0E7ZhnE1ScGJXpvfAM0GH50UpeoTA5U8LIe2wj2uZIu2cW5g1bQb9XXrCco63PC5TrIcCmyBiFqAH/xhqEQZv8vfTE76i4Nms6XJkCOlpdBHtbyl2iIBOmzqtA1swG/Tak0IkGGJUORIfUAGCp06tuDAMK3VhxWJE++atd7jWSv1fOkvO+ZiBlBeqiZ65cdEdgZVGx33DdyvN7ZjZ1SNHqVtXhO84O4hpEd34hdjiOHvPMajNHexck2LWEWy7nTxxnsu15RFd1VXX3OFwJ8cvt16QlQhoZo/TVNYN8VOlR2JJNe4bXg3jNjbpEuDFEtTp8Te10eQ5kGdNCYyrp35BooPpMQB+z4DDGG6qORL/zt6mGAH7ZG5jEZQ+jgfR2nGR6hCP8N/zcFc/mA/8FS+4SWG1WlfVuIekrBCyIaWsLXYWxV0j9X3ShcZ0Aht4fA8I7wFUyNS4nOxGheZJW8gkZnuyy0JDbtcxPkWCtm09XTc0KKWVJNIKuYWQZsZUCB90OqW/mYoyONSgc+Q6ZGdgXeh+DtEuZvk7inu0l6cE1ZSBtnsnwIe6es/itMA+pjbGxBHk4oCqNvp75qugpLay9DM57ew+D0SF676sSnyQ6C5TDPyyMdGwobIJnON3UkfRnW4mLzEzEe7qPp6FBAzEASE0/4E0tXds6hFhtuV343EQV7goEJVBuUwuw7ElUGohLpKu7w6E+H638lZH8fbx81o6lw+KoGH1882DewSRSy1viLvZiK0/qnGq0oFQUH508tJRIloQo6rJva2u/EOp37fZv23t1pKNN9UywgblKNTEbFN3bID5tEEDbD42WTwsD19cQo7hTEIG4llmHqQzFB1K/vqd+Vvj304Rbh9qSzVqE8rh6CnL01EOQyj6kif2rP825vgdab7xw9b6wDNlCVaPmxRk6sxc0Otz10wXzrg5SxFpTeJhT0Vl/QYZdTBoWbfIaBG2G5fBaaWlNfuuy1mRrEC+UiZ7AUWt5hC4PHKXJZxgsy3gxY7RCsv0M2BE/YYb7pSnt+E1gwQQYxHX2YqUMLDAo35kn3t7SnQ34HzvHR1Ib3VtUtphuD6Fq4r8p3uO+SV7TcshFGbZ8JK/04jZd+OUO8OTe8fa7I9vAvBfVlxoUkFvGJU/g/iElPRU6vv6+bC6kdiTHSJ0ZaLVNFyrhonspsYm2YP0eOuOh1mKPntnHxQ1RUYb93mkVBwObvQIHBTgmNLZCbppjitnxR26BPLq/60UsN8m27Jf7HUZ8p88OIyWbGyS2+ewj8WctswCAC3JMx0kD+TQfUIp2lRcoDSUEhIvPxtcaeB83x4W/uBEK8RYORIQG0V4IP+Kj1yvK7qaoxXRuPXukGC33jPpWCVwgavLyG0eEmH13/7JuxOnY+XJqiUWe7/VMrnPA+kYHMy9WZC5NXeFrKLOSvgfPIo3ZnVREZJGaWm3FFokQINa5iNGllzy39la+ljV/+7UIXPv9JEE5gtpzP9Wm+mfy+BeQsq1zsSZ72ipk7B3z2Mw8l5K7t9MNL0ik0iP6G/1gOaKUC3FhI4MkvoTY+bGYzhiuwbs8nV9JeF0mRzcNpMF1fFsHqPqFws3HQF5RGawcDqxTGzgsNcoeJlVaWwgEapKQ2mogQuBaGKa/tVHfZre//FDYOD2kZQph2PVHvwZN0VIIiemHUNarB3rcc167nTnGQU919PzgI35YBfqVQTiSc/iFElJGluSJxfUFqDlU2OMul/2zoAZ49shYIh8giwGZy6kv+jngvwRBBujxkzx0+IU5eVrczoMSI32CsOj2fFiA9FgYoMPiZ5YBLb3U9QvvJXGBeMizF7fUwNTlkYrF3NREeN0oz92AHj+Ach5U4ve8W6PgR3OTltPhObby1sZ1rpkixBZeqzV9mPbdM3p/HdkcEG5SCShKBLQQM/LzXefwk27CIjSgrrlyRTTcDOeWyv5yREXHWJaak6XKazscE8DRfcM6qGF9rrIwlNJXYMdJxhGSOyh4W//vScyCf7Q/2ayfQI3i4wkeoRx2sYhQeWID9q5S1AvRn8YbY+7FnkOj7UKvhF5b5HOc424ju6fXNB4t4YfCjafQVK5gH2E8hQp+eICerB+3hKhEjuZKEvR12pLwFnpGHd97Tqr7lHzxht4YUEt/L72ZpvuAf+RZ0BlYjJ8DDpyeKwwOKGXQ9PebQ/NcMzj1U9YU5GyZBpYILEyU4M67ughhxwzsvumDUnfDNu6oo07gBa5ezaxQgqocIbriGoQuVQsd4hEPeYc5qgxSEzfoZYm6gUjeSRtBTCOD1OLfZUeSMHNwRkm8J5YZhB6V9F5Bv+3UdFVOzGDQ5fhKSNvKl4YWW12S3VUGGPj8nCXHET/PuMbX8dVw4G9u1UIkDv7rkJYpkjjkavLfmam8KPQCsqd1m3oVK1p1qx77vI3nXUebhQ5EE6U5L6FUUlIsZjOS+3em2y8tiNripdW84RSw9GizNKBr7JKBhMAyS9+pPo3hLPy+l6OBD5pOjjEw99aQpIf1emnADDr1r1RZ8XwmL9d7cu5MKDB0SknQfjkyQMJbXWl4ejaD6RmtWd7bx2uBrkE9sGzMqk4ZB4m7w75iqbAiQqh2Vm5d/E/DT9TDsYuk0z56/9cQy1G8/EhlBOfwAWhoRoXEIiaH+se+EwrswUsASt2oryj1JojkPkBNmkqvaxqDXCccS/pbZmU8kc51OR080An5ceTifE4zKi5jf6uZow4boJ9FrPGyU9aUJ2vhd5psETIdInMz6RWauRP+EcNA8MCGRl0mI4ANY8uknwPRbmwOatEFDo3++yLivpWAe7AfHddAhPrl/dqPRXMyN58mh+7GPXix7DoBPHndRxQfYZ9NdfAi+xtQLJgC9kv5stutJuVqRusY9eG4Bddc32PtkVD2Y7wRhZWhrQPQQEG5jJjQ1fCURA+xm0qJJFSf9nb0Jc1VrNhGLHGm0KXHXghRE/WQB6WSiSod3igGvODAVWIIT0DWuDhn4feLWsgRWfsSq8wsBQhJhjeWNEnXEUAyMC0Np/jUoyv3u4YzrZ0bu7Vymu/yYTsApj2MhuS3nlJrQyY8uBzia3j0yQs4JkJniRs5aAEd6gTVBFnRqtHQwDSP5BVhN0cciJmw6pUkZeRL9VLPyNU6c6VtXNCF8r07oVdlhVplufCidMzp6Sv1aeHuVLQ530KPne/nE20JmIT/1glHzpz7IGTs3EvYTFNSpK0ow+X1G1yOufzQgmQ2j6N9Ktw2e6lJBnLaHyKO3HR/y2K18A0DWhEmfLURrrjla9nxV6z9/FqEoIKuLLOss3e4fHpYuqbKLmawSsULnaGIlSEzTuQJhaFXYVHnVJy6xLsIfGXnt5/LLYWiM9vJqKiodlMOyfHngeOFio/aKZhUfQS6c3LfVXb6s9DI+Lx64Qbiit+yA79kGaaWIXOIB/nLsgjUc55xQ+vJwwgS3kZY2xYvx1pYamy7DfuoCOW3FwhZXLKuXZG/ba0yeEJMbzGmw5GRbcz3g6H4/dXG2YHLHf4Z7vyd3j7F+GMOm9v3FNk6hM02w/Cuya1Izg7H12+mHsmfY2kj9DeQtADZUPW2eoHYHIefYIJ8tnaFnJ3YmlKseHRZ/4dLJeN2s1ttIy2HgnHUCFERVt3XhIZGvGpTk7eHpQAZNdNyJ29xS74XfhJgab0sMwavZmkKAQwVUOYhktfGbZHW3KEf7j6X8ito5ce4U4dOrYZCTWvvu7tBGgKa42VMBvXmnLL0r0nlpCCr+Mt/OjLxd3es9Xq+olx41cPhNkdS84U76rrruszdktGgX2fisQlt8anGUf/+AR96b/0OuuV4oVJf/0n/F6E4jxHr9MCsmoamRXtoJfR07cscyD4s8VcGzhS8Pr/l/SJWBPh+So+2OaflbnyDUhVNwg9ejZ1OLKKFaBB1Qx5pUPRxdKiAaXwn1uXKSSSaQnAm9K+tCVHmGOgbs4m+qy1I0i5zVwigV3DZGNRzOsJSFptViAQv6toTJJ3zPUU853v1wXeIeHggADxZ4EAUQNhD6YjzGFh1wIrcWUGmRYyXSnoDpx8tBReMSOn2+O4d0B3P1u38d4apM48LYcN7eveIjdIV4DPnpRO5HXE8uW77mPSsGB1zyFUPoD6Y9kcO96rrGDpzQOgldh9QPSlSgA7n8zIgy6tlX6CmPp+bINXjpaApYxvjtj2U4fD0ZVy0Wb8Ec145kgCS70TRhuxjmItGrX5yA7qNPvHJWWon8fSzJ8YjT2BoLLLfZB4ALaSxOX7j7wuIZ+D0dVCZKel0ZpXGc7oNZkYttkQDuq6OUVDuKB/gQLEpLWKihI1yiJKC5htBQoGtPw9q9kbPDIfXkBodvKiyohUakXrT/smSm2fB6c15PvKqSuC8lH+Iy+44wNRl2MelpbF2m8GoIMAM+eUQvvZA8RmKItxFk3+0PisksfZDpXQiodUTlnvt8uN0cvx9wYGNRm+9ILRPX9EYarAWrszG3CDiOxeuxday96bJipm8yTC9IOgyoi6Xg3KJ++AmKddof0IVPTBhve8kuqRXIM1hKxvn8Xds3CgVzwdaaUAXAIRJE86Qphk7Z/8VD8If/VSxByW245B8wIeDq7aonfpGdQm6hwMJ+SPmior9jnfwmYHuNlLlI9DvXLGF+YTv6SL2TkMfLrHadbYM1feErKBLisUMJWujepiwuyN51g5tpT40lhhBJFy7ehPwc5O0CfELE3OwGP2WWdS5Zyi2Yc/WXWJDW017YpbWFw0GlchAuxUTOXAOTPn8L00cfY83f73BZ8WVcHxqdO+LHf9qycWQ7BoqgTAWHroGj5UHmrMbN2SQAiMdnkK0YMhyKXcBa3oCVugo8+QekDJ0pAtRlZFGkQUaqir3yO9//+8apwnwvotQs6IoArFYKD5wv+jwV9cX0JyB+SnKHqKopc6ulnmWA//CNUtDw/f75pA1effdG/eA6GKVA0xvNUoSsT4J3WYfQQfETfX1Yyq2eKBnpnBdP9a3dWt7x8CypLq4FhtVGTowtqg8oxlBaLpx0dBnXWky163yLv2N1lb9lAlFb+zHEmnPjTjSay05/QBRkStuBggdc3eDpNeUv2LDegV1lZJDRPSfAeDGhwTGKqLrYVJ4zVuvOkuSrvB8Aks66M/zm7HDchm09aMox/G8+IXGthCosqdkhYZsfMErYyl0QVWGyuh0XkcQOjydZwVPpL1TshXHtndo4zI4+bDtDYcX04pwKymh6w+LSoraZpdE+qmvR2FgEwdCUY5df/G1Fb6CDvOB8BcWb5BIIsEyJHnvi09QgJmgMPnqdkK26oWrMYY/u+25+xHV2qr3jenF9qWCCJl/06AxepwiPEw408DOvqbi9goitbPMWRuRXST9V6T/fuJ4aJ0Cm9YCqglbywIrKcZer8WA58MFTLUXKb6kUcYK54cPsWBfAGdruQUavmfBz6gvJIKp6EDbgBhisCIuGelhuh1G2hGBY2Tfz41jUeXwl1kF7kA435h2KCf3qtZeumPX7Et9nyCW1Zrka7re9knWLTS/oL9yBG0M64+S3EjMYX6iJ609qLgr87fzV6V8zUMUf3wBNa+B9SqEwQcmi+Vp/LjT91kCHLRBJTrQZnuvRWW31LmWAkA+OvMWpxIJzM/qZy1gcexjEeSuSUHblikTg8QnW2szA0Yam0tfycFqjas9z52zrBh3OzlAm5I6vg==
`pragma protect end_data_block
`pragma protect digest_block
d7d79d963a8bfddefe8b984247a16ee00d9b116f70b5686499f22efda490941d
`pragma protect end_digest_block
`pragma protect end_protected
