`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
AI4VwXHg71M/l1ulOIlL9+DOurnY60h+Yg1XLkK8J4OZ8uqlG3q6H99QNSkwpRXDUPuVomQ7i8r/yUMoISC9HnuNBYN3MwsW+bq08DN9mQyPHcDdTSQ/eFbL/4X0DUflbg56C9rK0tRgoFeN12W18pG+VJl03xqfIhF3XYx9QQKWsh5b3gc7NIQD3iCGFUngLYlmPXyAOmrfQdbxiefW8oZ7IdNvwhHZdNPuwrLaSRODIp0hTDWAfA1FshEkUTakCI24EIn2Tr2TJ2b0Ys6BxWd6dY8cVUD+CKTT9cBjAScWRBYhbMqmVoVbWESF8TLzuu0fEKhSI9nkSCI0tES9ILHXEuaIMdUey4WgRcrZ62uWy2QFOB4XkhWKhKY7l5RqyRTZA9yBRbIo7VFsiArEBatbqgW2EVaeKC0aLjk0KT6lT0uRLrCXQ75dL0UBvIDEFnVrupuXBrgK5MLkLBOyGSp+SXw3z2U0d2Ui4uMzdRIhCDTzQbxO6tWFdBAeSo4byY4U5Vk5bK1vKDR6oSsOtIDspxxFbuNahuebA+yN33hMiDxSYV74Fzi7rvZFAl8ZAjjizeawRGmNaBnmW3G5kwr92cYEFSb38H2jnJkpNgb37vfMz8XpyyuY2qRucbpoQ2mToY2GBTjPVYiWPjJzrPiUeWyKjYiXfPhjPRHILggFeOCnW8FHbJbnfuoP+CMH0zkKh7KdmiSRCtwylM3tHsplKCK68JRDQO/KMURGuUQCucG3uBtxI1hSL0ezGfcHyox31RTtvBTyoCR7wzq99TaoT2jhzjFJ6Lv7BRCCZPcr9XRFhOs1VppKlu6TpInCt/WIqtvcyKuNxqiidfPSfQ3IaLd5yKwt1vqD3odPhDKHxz1vTJOitWjUcwwR8GaWdX21Lpjl0CC7Ue9kp2NHTBn0zD226IG76RhlW9jJifWuqjcitJTTYrrbTnC3GH5gMLJGr73RWyp6FqIIHC0myFYaOTDzO93OpCoqLJ4qiR/7uua0A1kUnu0sxRAu8hl2B6qDd7NDxhpmNsKni6fPN3yLGXF4xGuxdf4Ede3zB0iBsW1bijSf2Vg0MCTmG+dJ3wt/hgbDmc+WC3FKjfk1t8LyKydlV5HSIxLOMPuUlpM0PWT2rU6hIjGh0v4+9WDv1dsXZyWPm4FWVbyZlSdje+Uu9/87Eorl3tTo58te+5z6FxUcxBH+Eh3igpiorndw1BWNYguNnFXPLALceMRT4eW29vNkMpoSNF7K9grTDZyAOlS0edl/MZNvo+2ihTRfE+Pd0LG+wy0g8f1HKV8A9as1vVv4HxtTuVNqyaTJPoKRaRR0RsNzn5OMh4ArYr2RM0xtQKz8XE5GhhHaT5curoAslILdt88t/nIUI5ljc528l0QMU4vLTSSqDXmxpdBxTew27rZGAGBxFBAoKizOEkzWPCNKYXD6xh2fl7TCMxqAoPofl3AU++bRLoEKM0oA5D4eFGMwc61DPmq58SVjMQbrVpteabj7y8/pZbf6yX4jSTXaad+PCoNnXhZuO4aCh5iUs/UnHHtUvT6KqNHQCvsELZ8RVN2sLoLZIzEvd7JibAz5CeqssxA/NxY9UOQuRLPLLUQQyE6iXICDUpdNBjx9uStQH/fsWVIvyDSyTpJ7x1gdanOUPOCqvcF33v5HvBu1/JCasWrvw/ZKDQjvq6DVo8DcmD5XS32ArnO9fcesUe9UKd6SZ19yQC3jRlqeCfntEYGi+M/JNN1YAh6VuznYXdSHwyoRhSHFAi3CXrxyfzpLqO+FMMseH60AV9P9hgsPAhtcM9b44OboerVUBg==
`pragma protect end_data_block
`pragma protect digest_block
ff4835d2e200e2ad131a29e3e9e3edf0e731c263b735164babcb64ded6535905
`pragma protect end_digest_block
`pragma protect end_protected
