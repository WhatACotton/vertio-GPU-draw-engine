`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
uMDqU7kZGOK+0LjG5DpPSaGylaESJ5rSmeoQuqde0cEYEUsfqBbDxZ+uszyD5frab3TKXMzerVPpwkeJJUzSQw75+ZxfakpJEdoS5DTWGDqcBy+woTLYT4QoVhGt9PZlRVo+pSOs5/3LNe5xTfb+MpXhPVUFvlYa9G33qg1QL5XZDsZBeYF7Fn0K+5f3+fKCokF33qI4Pc3JzW/y5HplzuyWrBiAzquj8BLJZ17xC/T2gZ6Irrpp3f+dq0AIcaoB23FHizRCw/wqyC7hMBhTSjHuAAPgNePb1k8PJ8w/uS/HgxAzvPZSbAaJsrKZBUk4YYKtCCn3xtxCAho2j9YWbdYZAjDzW/75LEJP3r0qzOAEKEEtScTRZj3hMRFy9bF/cjEg5W9MdnMCaqjdzlr9hHpaZKpBF2rQNuLztcHH3LmU9S7xXakTXKDtint8JUKyg+GhzfLroE4Yfe6kDrI8CGj2OZEm7I9qqmbURuVVToLRYrT4bnNgBQsJQUfqwjX/Rq+nI39zk9atheoe+Cpsn7UrMISxUuCUxj8dJHY/7FXrBpXSQVMWP+B78GiY6gSg/+SHVbooPeg5RH9UlU2Ql7rz+e+ZdN2Ch41orTUAKi32IjyuIVruy6xQbXNhnlmWJFE0+DglqwcmfrLAsc+hBAvAFeyG6Q8RdOxoKGAJYXRufguArvwjnekTnHm+05Vbm7hpxj0FH4xJmtapm2pMQ/szv/+vXYEbzlBi8eXv4NHktX3oi8t1AENQgl4KGV1lxPHfmoLeSkMcD4j5Jg0zsBtMNBHVigjNthOlXm6yRVV79Pbk06eOtyhACyZ4JBWRgXCV5nATYhnzAWZ8tUebetdJYzZpRflRd38WauXxDEZg9NC+5RW83FNl0QNl1mETcsOXrkVftxZkEaUnJ9PqnLRvKlCi7ay+49i8f1AO/m05OtYn2RCL14ywxGwJ+dsSQmBn8pTopt9n1jSBMaoLj31/1tMCOlhiYwWtMpV/uWtXIn5jQf/b0NlP25oJDar7mqDYftAhNUdEWPrlGR/y2avMwxm+g3wErnBW02bz18CudMfZwFU/0/UNNHBi006qxNO/b7NnxNIuRQQtel9VKxs8mnRr0JlDdSdQiwOq1flgfKSGl+BuJlYcxpO6dwodcbShtdphVLfafNqVmpDIWBp0m5tTr3SUDbTZV4L5iE93PMb6sMTl1zHgNYH4z49cvP/Ncaf/OPAwjhoSNhc71Yc8oJ2NwNJEe02XrrnJ6P47RHODWsIoz2n6SfJbOervOuk3+5Qg23hw+LNzZNxVVtIvTLJYgvflHNxSUMDChYQMraYPUoEFtnUjXOuroOSN1KLVLYVmj2EO4+LofMiw7igDiW5HJqlIpmRWdS2evWsSC+QdTSwBIeLrDYXJwuNmpFPuu4z+QZTomtneDxzZmXKi5qike79InNqJQ4nEszz3pKvs7Hu5LwNHqIqCu5GOLaB5iwOU6xuYP3262MSndNtFodhZxYQcVNNMqmFO3fWWagtMNj4vCkvjtNbuWvYOCGWiGCYQXMXFmF20iSoeAuV91UOkdJqRWTeHmFQeVI+IlepW78USlb7OK614DX7e+EVbHzIekhgUWxZFG6zgogdOBKTSTBQF2UEDS0Dp/gkACf2wEJ7leTBF9qh7uSn3GdRSKZSSWJrkDrCkpQJhEgj9fV1QqvlgbRGcxvP1laXX+CiwxnPeDPEgt52cz3fc3mA2VqXWRdEDKfLe71JXQIXob84oJiWiIluAc5IT/rOd9FXsGjYmZxVEqfGJhdRfbiI6qJZLET0eF4ZU5zA2dssBOELOAj5VkvmdJxANEkaEr/ztnCLDFMvgB+SyhoyuOCchWsdKD4XyqOMu89PL208CNSPGDpP3Oi4G8hb18fa5hryB5ZJrlHvNZio05YrirAjmu2a24xdF/76dWPRbcnwYs+n74xUwJq59l9NOayLNUYge05aiVUOuOb0YFaZZL79jEetIIX4rPbYP/Dw6W8Mh+spaupe+35Ik7OsxDySQVSDCK/Xk3n/OcKNBFETvquQ6bMluEnHSz18U7vFJqMSkTZ6Ke70fMySZ0GE2B6sWv+Q9PP09CXa15fpscQuWmDv6aTdWe5uXnPzpGcNF/GJpFBhUIMQq8pEqTuTrl0QOAOxj3C8ScZcPxNPShnvj7SITM1NhqFGuODiNwUkF+OpLDGQKenbm4Vkq58vJk0u/AEcORruIfKNPsfvPuLhMdTE/rVQuWJqmZgWZk+T+cxcNZKnw+f+RFvcURuk18gQU4aJesQNfqUpm/4xsrDl3rDUZKl9g7yFqUDKtW8rdR38zoJLvA2/e7TGeKIhPs/pT+yX1KXa5x3AzwagJKQrWj3qdTCkCDfQzMNh4QY3SNyI08/gx+1nlRPYUlWcRibfoQR35ecljA6JdQ4q7f9R9E10SnHSmrKpfPy/FPYHAvLy7rkWrYWlrr4f5G6SgpLXKfT6NoD/NYrkFTTCJmchi6VNmJUwAuQWMSwqzoti7KJ5lND5O65ZswswSIA8K9ajV3LZsyqhnWbEvxyfijr+k7EFI6Ki5FZo71eLaehuIMWkIcZkkkGYV4UH+eo8Jr9S4oO9AJej/CozeycZoB5baBXaI3Lg2mqorf07k0e21TIbcUlTbreRRA0NWIFXhM92T7zI0WLj0wzVcBCaCDyxWNUxVe/4lB2euKny3x+MLoS1fHhcHthTlYH4IRJ0ub6xXUQq4YJ2b6gcqR4F8v8MvwehqUkwBd0hQwkWGFJamWhE7zm/eqFE+IveWoo1bNNhgBFiaCNRykExnaZqYZ9LRsUAF3ABR1xdrt7PGxzMTMtzbSWx4IMruHB4sOL7R4CcCx/k+9FMLC1Dgrd1mzhtDhSg8FIloD+9vYQ1p9cjYUJvqqE7CW4obKhvbhI4gJRhhCg+hihUwYjnVxK73I6qXDIfVpkAc144iI2alP6oL7Br90gDQ9RuwvCqhdKdi8Wd7Zee1jk8RW97d+bzlpFasZGm2Y4scqIIFCCKNLVDvRGeoadbV3dAZiQPUnZYbCiUP4m68ft66sWJS5G+Be7OlhQno1Mnx6XPsN6i64g4vQyvItEsaTJjiVABA1IW1JgzqVAWa1qbd6+oqC62O2ARmcLAFyLviFuKoJaYczVAVhNLcJir3b/9q3tbJUX9izZ9vqAUCJ+0/UTwFtAlJU6BRzm8oHgpc1daAp91MDZnec4LDte8Et1134iv+y5A3jVKslnQyVSAD0U55TYdf8XGiUN+Ftv+0YkDdZ78tbmtRN86Vus4wlNfCZ/VFexAvSclATC09KnoLIcT7ZbPxvUmMuxeGqa5JWkzmhl6srzaUbIvCIHt8z7oScCq5Y7voP/OfZG+cjGnRDx1ywXWV1xAKiMXU7H5hwBQteKVvQjUC8i7fK6kQegN8h0PmQj6xvRiatV3hck0PXwKIoCKqjUr7r0P+eGjfjgQpP2VMxGlPa6Rl9TXSiykR134vZDZu5w26zIinQ2MPy6HS+2g9edkkSx2KCunA7v3Pg2Z5M81puXrqxcAQh0h7V2r5/aZf1h5wlcyZ5dzbimLL+bqIJ7Bqf+h1lFYiVewmfRS0lFkXR4X4PdHl0mHJLD35IHKXfCPXYk+H2/YVrJP83E4wW4EdikcIiF+ETdesURAI+1symkkDFV0/1Yevz1lgGyJ7OwBv4v94HJyFPxNoKPr+hTVSx9hwdXo8pAGXSY4I4Mn4yf7Pw85dLD3ghCd+BIct2Zrd69kC5tTjPUki7ep7Od/HUEoR5/BEyUK8D74IgPia9MZXUFrBxl7vBYhPas8SaTKw5s7sEvVGMq0dmv6Js+evSRXCxtkpyYBoc5hNiIXsPaRJeYHQ0Un57Tt/VMLDpKhPASy+bQgm4o4BnR3WiZY5JUHtZ+wDIy8R7cFjEfotiyPo/iinjwaNOpuYhgUpSq3cUlJkOgLLG1HgmDlg3klydq+liKoObxRRtWfqGdLVwe/Ppo9eG0wB5wkZI1j+CcAGufPfbBnx4YxFsUX68VGcsb8Vf/Zl93WsDL6NljKUmS7MDqmegdrx8t0FQCmSd2X4+Pnx215YhVs71sxj6m/LTC5lbGPurYSl2P5ar0oxThJ21e/exvORyHuPFynEWWEBVmOX+Oe9rdruaYNoPC4teJJ7obqf3vQyZcNPXZlZJ0xCtGmm/7QnxfHKeKidKl6yLmhWMYZk0I184jP1vMzD/rf/30O+ApM8GejEJSfFhuFDuR93xKp9lO/r6X+NJKIh2/uvw6atJ/b+5V+/Maz/gOdRy3kDsOn8mdjFYV1efXGLk2G7gBrJZ89QZi9z/xovyKkfwzAeSaaCCyYh8/Ox82sCDUoUEYQN3HQiRgsyIQLudVbcF+KGtBE08Lxp9IfGSACAndLwDSlkMY3Rf2P2b2Q2au4uZTaVkC7f5parSCMBAsroS+bnnX/FPWX7zjUZf6PYkn9+OA20WfACTQOX3spCmig+yzxG6QJMfVZrI+CkC06t474nk3ejp9M3nFUD6rvBpLfkfQZo2RC4HOYIX5l0hDOMHklqIt9qbUGkFOa1fla+TLT9n6OMIjTYrphHms5SucJkD/IbVgV4ckAzaUoFCIi73vP9Ie2gH3GdbqYQjdL2yClJOof/JdZzey644BNnXaRRdjI0C7wBO+QCLiCU4LnaFJ8rqFSsI6urFpzY1TIwScCID21UR6j4U4XsJnBXU8SSkqOPsQDK16FzHiolVmyL+3jcmFM1E6EmNFoYo5eZ9NdUyCiO0ZWv021ruQ1rIDLwPHQY0V67r+bhjxniTXgkVW3542u8rUAhqn1CQOIDbblLv0OiRSmAzlAQg9HSNaeRs7OJFEAksjLXOWjGekj+raIq4HhQTm8eRG4W18cmg/GJ4x5RUFeAg0voXzEGpPjVyVcbuyiHXpBr6nK4CnP5H7ZJNiBmvAizFMIm9vtMOBoqhtJf8EI4SclrAxMi8yHuFmIs8Wd1KW4bHIeVl+lX+9nI3eZYTjLvY3hNR2OfAzHmLy146q5AReFgi0IMMAH1z54/xzOcQGGM28O3EpnmPNUEU2ikIYewA56PzYzDMR17NhmRDIKn4q4NfBrnxf9yGsMOwzdviuDa8YfIMw9cdHABs8z7GooCxYNuVs+Ql5dVWeCx6TKU2Smn+XV/d/z10kmvXx9EZ3SmpbbHRvUkldEVLkNyHexSKhLxF3t4DYDyd/AhULKG08vFl5Uc3PW765omAKVQDF8rj0GZNzhRa9fr7pj0/uTj2g+p52kGNJrvy03rEIw0kOs9wFjgGc3Bgh3QbkbkdWv/Bk6TyMHPR+/PttXx8UBu+MRuOYVHR4BSpH6ZmCDtIp9tOJRoVGznvaFcL/x2SnUYre6duJLi/Uh4qANE3/+KXIWL0O36UGTvCENYQjBLJ0FgnpyD88qkDfL+RAUMXS8aHrJI9M8aNP98nbyc+CSoW8W1x6QgGsEidyPzFx9ACkoZshjW9qNyO/nVOkcOyrXawVUJ9ISWYhCJeRlnZBGYC/eZGNV1W4YxUd26bn8BJof8M9/5YzGZ5p+BRFI7v+CDg4nOj7Qjq5i8/SR5vIgV9QTnbP+rWc3WFHTEVPW/CNCXuA1UuEwQPaJNd9VaeiurZF3bHGYUEk7VRcWAOSRvirM1I3skM2GhxOSeF79BeEGYRrrFwvchbUcfxvI3pzyYiVlRp/jCews5ig1iLqV+Uh0XyXaZbnZ0yZb401+Tlr8XiyqNNinNKngejqq5IqQdIhcFU9QQEWeim76QmTocw0v6Rxy//D65q7jmOS4q2C79sIm95MSie/eG6oae5aDl5/0GzyAUOkw79uoZMBfZl8dZu37kPNr6sVJVIPxRP9LIMWo6baz6/7bLaFkLDHqspWHGXRmtPpsvgjwGw76Ip8fyn3AA6JrHR/atWsOHY+VVxtfJDYh6Vok9ApxXvQdN6v05DgRDrsBIDzwLtn/IbAjkLLSBKAkrjHX3V23+0g03bT8aGXiICIZMqnPE1NdNXSLAL7Qey/j1Ck5ZDcQjh18Z8X6KJb4mJI/KYW2oam0VR7jpwtzpzn4Vs/QLy1Dv+2jYAByEWpiXvyyuXLyzo+LhMEwgF0DDYlMYa1Uw3/sreL+bfJ192N1UcIH5wcANL1x8FYPtHL9t8sr6lVWnts2FmeJrXpyNu3noSPzDfiO2SUgAVbTjW9skIZKn/58Olprl+yBWw+PqCODLEo15jLIQBfrgKrCthvLOl5iB3zyvkBYg6/IVbB3vM7wVcrJtP8JgnDMBZawnp3V/HPEhQSuchPv/Zk0420gaHfme96cVlNSYu+LKGBi8VGTWm8m0meH+03kkA3jFXDFVVvi+2FmNzVUM7PImxkSqjP5iR4C579pi+6nPCHCG94amzOml3NWUO6aRc4k57ho2e2juWmVJSrOU7yfThOOewT2UAG2Ee9WmhFzcJWGiUagX3ZbofOC0m+WYziAoms1AQ6O8+O0lhsu021rbvuaHmFRGaOg7pkAmoFtMLbcVI0cZ7YEsXYH2WuunL/CQKmyTkhbxRufNMu3pFLXsRYaf75kW8CI5Lc/V+kRnLJReP69UmbGjQghaWIe1R0YXF/NWQCKc5VBO6KKWJm6cOHa9zMqbvy4xgScLw7ff4e8ek56fG/kfEsXBuNdjTQz7zhQ/uG3k0UVh6VGkqyj8NkyvRrd/BEFsbyHyICNFoKg5GxM3iBf4Io8Q668QnXeMAiB/AUMWYgcmo2w/F/aZsJ+LjLi00+76gqrTwjK+i3E6SbeK8GtilVRsOxwL3zvWGpLdkXaOQLvxQJABAvZnqSofyjezGnOBOdZYLINAjfbPIpdF8Q7XhsmiCcC5KWf7zY5nBHOss+HvJfLnZKL1yGC9VmFc5mPrYL/xdnSk6Zx+vvXHlbDzfXJcO0cAUsBU4pINOoWsWpaEbDL+0sytCNRWCKKDbu2+EgZIh6ZgSN3pOTBSiNi4/SRQLVNf0MCSMqlArnvYz+NKgOI24XOqjMTYF2xj6D9jmlVawf8R7RkuhqXIckveA1EjlVZufq8pVYn00LG+zM/ZVdoCWv9wzHwYgbOdY9t4BO3WYoLbolbc2yp/gjEgcHPpJnlxfZ9vN7V93O6EprasKLCIpcNZJQZxD64jlKjc1WmjzzsA/TNSwaMuxLz+hCKcvJpbaXwL2/sHf6AvpYgNPsdrXit4dgT8Cvlu/wb6aSbgqv3cxkfxY4oxj6EFb1ebsdog9A7ptQxEP3x5Zp8xTm4d9yMG0E/K8tW9mu2PsNSOTMidy4yFLGyP4xRouC0PMjaCwkkl/tSBAEnaZgUCVUJDd6er3ZMFbAjVAbaAeCTlM+H+Y0fG+4uSB+vstE7N7mcs6FxX7lsuTD1NtdHS+/sZBk40yQ8VS5hnYu83bclmfkZ8zVBnz4MoSNlRYjLzZBTBBjMVYNHlmUutPbwSb0cjl0ElQzINczoFMZi+1oqH8/5IGp61qn78i7IxMT24SbZHlJ0cWdXUdxm7poAN3lsD/9TZFJvu+t4ZqmaJoczdI4fPy92vrwTCkplrxeE09ZElAC2SL9UuXsppOe+JcJrvpMO9DvVIkncqH4hZj+gCh5cwtu0aPG13kH592cZgkbl7EK8fjxSbQGxkTyaqP6zYZ+87uDgaijvpm3UNrqRhp8Of1d1O+3L21eLkdc/D1XQGPlkWPH7mGo+pw4E4cRNlrjGM2o5iFVM/XQoqin/UulmCt3YvCPQZa7HeFlmV7q3JdqR/6/kXWsNImthkZWoAKM7nX/BrGm51HPQX9rsQevyPS8COW6K3jzyCD9OPQ3gLbj4E5EISxjUAuIvYW0CXGK5Wcr39gBaLQhm1eqaB+eAtMG/K+M8bBFo/RpIItZe+qA43gYX6lFgyEykPdfdDVNDLt5E7EU9R4SxSvtFBNUqGHsDIh15mMC/sBm/qlQinLHoqnJQnuXUkGW98Qjq9UT3FS/xx/FaVIL15Z1ZpkkgrLADyPYXmvHQRKwKzDVLOrkx1QLousvALRGZMuvzpEMos/vJSB3MgmF6AO+prqAi5gJEIDlscnVkRbqoZQhD64nWHyLVyde5w/TFAMWeTNOsRkaXVurocPgsSahQUGUF/kZKbsaUOMHrFIPylDZcVGpv1niP0rPPQt2sdj9PHy9DmraAxrbOnZyXqUCYWUc8Bm0Ot1zGRhh6yXWOaKJp6I2TM1I90sEiw/5OFVoB+lw1KFFlOm54tKBTJIIAV5SFgkjbwn61zudU6VhI73NZex9NQpVz1omZfP5X5RcSHLGqV19cElHiKLjzIlK7bZwGsgWG0fIUCZsGwutApVi9foco7KNR4VAgHZZnL9f7L8sXyEgd0/qGZOJQ2vOddXlvkWHmdRmy4+Lfo56IaN3TNJHpvjp9Bc3f2pYBbfeoO4dw99zexHvpzHwFaVm2w2xUMEohY+x/8XliodIFlp7vfrxIVuwtl8mtHSEmvklH56XjjlP2UDh5rBd9+i4jiknKB7Hn30GP7kGVm6TKFS7FyQSBFAy9vfEd6jAMgb8RvAwWU2f8FaAXvVJ7ngmGTXtGon2baydzPrV6ZT/bBCzMIFXt0gk7LWvBRg2D5frEGzyKYE7kkS/40lLEzn6ZoU3E7HSs3h5z3lm3EghbR9VhFBmS0vEd8mGiCkKVXRlbAKY/HLZpg4N36NDGSWcv5dI+v6+JzXFm6W57CTUwQAeL0WydScsJdAM5jqwv6Jw7FqMQwYMrtyyTluMQUhMiW7oxjHHzPLypDR0O2y28qfamE9gFRYtPB1pACcC/SCG20rNhY1wjmS5WpYpzD9Zb6g+lnUT6NvyLJVFp7x6FKaU62lGWt5OsrNUp30iZq1Z3FMKEHmIffzYnAB8ngBjNF85XcwS+vj0+zNQ4ug8D1bafQNhgIxBhdkKN7kiRNRpR/vOPtHqZVmTXN3V0fj3WhsdtnMCVDACSeFI69AfXYbKJA+izCIF/ISirePe5IxPbFOJwpDpXwbf6LFww2BUKEnCzc9tybpsCJ73I/TpQl1RSrKzVjhcgo7TywSbDiO2rTAzJgUM63slwvMTKLFJKhEOw5ZfmngwyF47tTYUs77GvAK+M/9oH1Y3aog6KxR75aLvu5Otyz2UWUGlQjgGGbcThm22QnZqd0Az/+3Yjjj1gcF/5IoajXa7/O24BU9xlL4yqZi/IiDqbO8iMnxxMV96EOrvgZbX5p4dOWibUY1AvB7bwOqKcz7i4b86e6EnBTYOtFzlm9G1aSl93f/hfTtRTEL50zu4QfYv+b/+TNy9EpQeYHX3hLLjcmFjXZX3OudLemaSGRyCIBcRzRXv3P/ZPqQV0tYpYrWwyojjsQMo1Px9MHf2L5FXVQcUGIW5eHQVxkvi4GBu0/X0UkEs4WwdE97E7zes2r9wh9F4w1S9Z+T9VAPcyCV2bQit0QeNkVgWHIu+TeUvGk3vBuYDt5Znz+JbpjwiM7210A0eX6h/hDZcWojxkHy7KFuU9mpD+yZhv7zx1IaIyVyw4ZmH5cdhTog9MNw1AqS1rL20DjXyxt/7m972lJzPRb22pyVoiX8RWsCFyL4kJIb8femRlCzJOKhagwapHciXq6S6Ib72QKwARgguGz3qZRPZE8Nw2GlfV6LW0yVm6u7UQ/rhEbR+1/i6zzqwW11sFLRJT7MyxibmQ5kb4e5solCXAGeKpQMEqpVQjJRu+lvlSj/o6wJxknIltHwZO/GBaT6v38g16lxJJa5kVhPhDV/PURj57BSf6YUCfev9bY/S+L5hbOmi0+P0wPNR9dgLtFFaoui0g/Xtd32ikENd5F5VQnKXuSO/7JfMunkMT9/649VYuIqH7ik3FspTeD1M6zbLSI1Jdq/fwT6AfFRaDL9aIm4VlNpNDKOEDJlrhbwk0CgQ7hv8z1xktGZ9FcLuOqMspwnGVu9oRGCYmWvaAvD8in737vwrVYspx3R8icvml9L12oFsCpFuRYCs24qih2ekXCANDMMzrMW1SDb/6tNxgU78IE/oZc8yrKizeYo0rRjGeK+D1sOJ6vUK4k5JCT0XiN8+CtGlR4ssxOahTWUTZeJlAincdcmeyfUX4hHsRtfxwoS36Yxyqgo/vcseRXNxS9RYuy7XDJsJpOiaZZv62liZrzGFWE1+41w5jk/lpeYfO5T5grxIFIDbHPhxvCZxLzjcSTU19ILMkUXtx3k9HTd+LHYlhPAz46Bsj4+EDIP2L7ET0mgB9i6L74SGvQshtPZqgeaX5QpuLemx6+Uwy5HO0ewwM5NQYqqjhARr9bebfn7GwYyokerwYVw5zNeiIW0FaugKRCt4d0g96mdrTUPPWxXr5T1y1/sh1iecK1onO14CQhmwVXNMu+C+ftEdglusUcQojAZZvP2y5V/sQdie0KtrPreKeo1RCGSLBtEasmvKzuHv0ceb++SN6DdLRsFlBtJQasdx5KlgwX4YAdIAIMKwpLCoxeGGsfjwGsNqEcopNLa+jB1QV8sY0jcTn8ZaMOLhbsB5e4AnyJmbUYY9eEVkZ5nEJKAn0o1vEVazU4HMh6Fulxp0iEjZlHMQGpAyGZi7Qrxxvg9qYLGdHougvp0y/tdNIGzibXgp+Nuymf7zdoDBLazJFNerSDV40GNS2TcxFNsHAibqMmYUmVmN4jMeeW3V+bwTa3CJ6ZCGGH0SgpVxwqhligZim2phoqzC8aFqzpxezCkNzwSUheqFmm/UoEosUVm10F19uwXDd+nHtEbALuqZLwcvdWUm0alC6RH5raSg8lZs7YvAGAJNvt7jKUVQxzvHTUaCJqPmROWX/3YLAu16MzujHoA8qbcAaBXP/NEGRsfZx9bqenSVLbMmuFMX1fi+cXMPpBivzqggKjnXFabUvA8vcSnHAp/nKqn+vTKVcqPm1u9V7g7j3RKnCz/JUsE9h9ofrCj+0v9xMfPgY46gyRQNT1bPwxN8n5Vh9TDuv192jyHU8YocYqRXUfJ94n1LCWdEdgLnpW4npt9/uahvXPSSTvopD46n0wgkvdOL33KzVF6HwhZkucTv0Dl3xT7YcHhaj4Yrh/yj2SIXO6qxY3BHOwVfb6dz7NNApJYYHLx5agK1wj6IEIZtdXYCAyl0WlcAPshrGBwtu2bBBA2AZUTHpS0MY5wiFrqAmkdjAw+lr0RXa7kISCaBPoTTPYO77ktM/0e12waR4Vgl4vpaqdZ7xGWJsNjLtkIqm5R2acXNUEbvP+wkIcuCYEfIPxCSbxAmZ04rfc5d1tNabusFxX5TYprmypvvqYrilz+1cYmqyBF2jet1i9XirD4IwscVNo+2/wmkK+SeB/4MEhUDP+6pnXWHqPbOAyLEm4MdrZW6Ke2Xu8n/uW5rLZcvLWFcQbWmr+4bbZQcYShC/d8en1OZF910bg+osrR0h5N4KeXBrK6Mm9fHUlLl4qdPI5h2WU9yO2YvYDPblZxpVvHaRaLyS7otgnnTv97fHwBjN9eV6YG+BK3/mrEMIBA+bJ483v9975K3xrLJg6jSMxW+R2P0DiVd9JOol4O24aaLi4DVpfrTpH19CEQkJYHV7UdPiBeQ5eYMjoA4aJyLSJ0AFIatG2T4zIdMG68MlKE9ys0l9MLlY4ReMS93ThVPVspJMONrkFh1I02hEdeZlcx+dTaJLX3vT7e8xzQCjsyUnyNMy7M7gDYjN54piM2ylpXaIlZfc4hshRa5Bf9umtdyAWdMSI6cNaX5u4/zHuhzl9u5sFka38ajNv1v/oFhN4Lfh8n3U8miHbP3V/4sIdK3su2eBTSXO+j9oX1wpOP2mrH4i/EnThKKhTYBYuxNeaJNJ3O2ox2E5mx1RjuXkQxuY5W9srawOq7fktJ0qsK0SyNYOT5wF5VCwkPvpHwtwxwRVcV3hq6wxN8la6B0siMRhorjfawIUxw3+POI3wBHD9NzqZPm8wAeZbrlwquWPvMrnhl/WZenvYVOho/jxBjnzfRuJfK+OE/+c/M8wpgjff+ANlzOtk4De9b5NC8kx7bak9zqvdNGWvikOY8LAEDKIUiFTO053axdYTZT79i7/zOB6i9dqptu7mOT6VQXMtZcy+64U7eTATeyxtmQnsGkIpOGIpBWe1jmjEkOGwZo/uhnNlSOCcZaNk8DPqU7MTbnokU4xM+FNrKcQm/LAuXxgOFYVIg2nEiJsRu0l+0aiNZ59oBTrioG0dk320PqSXjUiVCbKA/+V4sC30Yz1mdHo7lXbM91XRdqgKRRAiZfIXbl7k+P37bgUa9ZHiRMR6JXNseE9yoKIUlMbAuO7B9EGqcYu1Z2FECNFo2QIdsaBHhMkhBUHzStNSHVz+dR0UmmnnMd5JO/BEekqe9/5zsfufdTolFgcA2Y21q8E7K65d1hQfbl1O13rg3Usj2sD9eb8s2Dbk0VLJjGnEcttJljPKVMfMhUSKH0UEUSoSPxVTrITdT7UmeY31n9/Qk2PasW2uh7x/dSez8DUVxbK2tpCKH+PLX4yahArKCEWjgALiEcyPotRhuIGMItROti3svB67jHSnDFOo6G16MazdFw7NFViH+pden/0PBX+wJo12VucKqJsdW+bSDa3JQPtM4jsc+W+kbMQaZEpQmHSGgRrVIsXe+6p/9wBEqAdq/nCCzSocH54oh/rIzN+wk6VOLBzi8pppWvaVeGSJJIcqRFksHZZfo+F1vd3Ax1VhcDC8FQjr3Ktri6mf+v2+0DCeeTasLsVChin7vD9ZWUJTcPpWCD8atfiAdqjWAiGZ2hXJtRFgSjOyZnS6vZieVjnwb/7PApBpUNq7syKzmKOha/C92iMc659C7gxLO2OEl8MVai50qPWegV4LRk7Jtr0GNPf0YAU6ouhGVrIwedp7BpyXsxLNeInX+EfxFWnug8XJBRi7Mik0iDIRkhu7Yos75JIql8J0z1+8wCCZx4iFS67fxUoyXaKcQ97xF+dnJhjvK16OuWpHczvSOGYEzcdQ51CE+VpoLHg+CWGXck4PqTFIH9YmC81fvBcdk+O92OI85XQN0Ey2lIOXwsSI7tqE+18D0z2Rm1/6lHjvkp7KTAZe0t4dHdYVflifsrK96TrXqAsMaWrhVrjBTIlvqEd7UFSvybJnl0X5kcajTc1kcd+6SZU4bc6KRPnwIdCSt+hDCiRSstDYO6UbyKvpWxay43A7Vgk0LHPkfsNs4fZHbEaizBtpSav4ZgdJfQ+oysMedypraGFokOjaJlTpoffmnPkRL1jJv6UNLYwog+ptNEaEz4CwyEnB2k93vkmAXnVtSjHakb4HeI7NKw7hyuED70iINiP5y5a+CkF9O11+J9EsFyjV3flRvzTiMQ8q+d6Yg5RgGRrzIx6c6p3XW8nOBalmQBsPfCY0S+ZXShobeR4f5q2nTmvARIWxDZHTmxuZiDrROnEybqFbqvDmjicoNge4DbEA+H0uY1d+CkBLRoKQXjkp1sImB81WWXNTgtT0JSIJX3ByKoxeB0N/9XqcbBE6UiXGHOlac8mGQL+wrt5kiM0ZLQY4reJ4EPFmcaA169yF8ah5S/6iAdr7Yf19jFQL3fhT4+Wyeg9zoa8Yw+4j/Eku/IaqIC1+/irsIxBdiUDrRt0A4YyOk7ubCR6P7VhbmsglF43lagVjHg2dcI2CdTgoG1m6PEfKwQXnmY1k77xALEv2waWRJ6mgPt0LqkqgXXyBc6j4a+R+xKuID/SBBPyUHww7+MNZb8c5tb7DXNnlT1R37PfIIWZzO3NUPkXBcW8dzYmbuN3d2rWnUtBaz7dzVsIf8lyUxEmHm8/ohphLM6JdW9vZTWPnjs4qaKwjPXW0AEsccX8K70iZbrz47QY+JsPIo3ABp315Ya2poeiS2OraURA7tHoEIvrUyjEFDHtwLu4fQDjmPqD4uKf+1PGWGP1Iz6e3DMMSl1tLSsbs6JogmAFDqb+SH2w4ycxTOI0saMKewt2H9Ph/96XeamfzHH0crntxEKjs4rfZSI9gzCFkmKgTSwIqVSNoYFA2tM82hVcektBUKLDkjKSdWfi4mlWdcHpyqGDVG6cR+aLwhDT40zmnYjiDLiFEc/ilRlqkqhF74DufxhNhHf4Td97eHzmM4FZ9T+jS4TDazDQXQ6YPhYoLFpcfZ5I5MASyBa4F0EjjXYdMK+gsbewnUAQSMeGLVw8gZnMuPKCXzeA7BlimzsxXdSTxWxkKx5jhHkAWZDwhWXQv/HizescyJLKzxRSwN2i82Qb75bWlFwpU5CljzIZMZcpGFXYUdU8yTp2kSfem1E9qkCdF5w2ULMjmKjjYTGkPYBu5uQfE5/qx/Vx7KcgNVHFFYZHk57Ou7qnt8SPzIsLi4hUrBdORzmU1T9lvW8cmtH15eug1UV61qKFWuA+k9qnhEb94KxcCi0IflNeuGezvxZvDtwshijOGSf5KGrSmadaMIgspvwTt1ZIJrd1iGJADMxrHbXNaP6WKdsAlZChLIUB/W4Z+T/aRnrVRYI+yASf3O1TKXCCfVWmveMvfddvlY7dz1EsweuvmM1O874NjBDFm21zQXlCvQrVtXLCl76RNTWjjx8HEI1Znq6CxCKFqdksVqX2YIB9wKqAqwgZg6fo2eeFO8oKlgKXI8wZt1m60aXINkNhEFDX04JUbDQuK0JvR8UUWxa4C4MKqT6Fwq1Duzu1nvpApw3UqFQu5B5Zw6p2qGXgo7V+IpWLMVjLuKYzlJvZiWi+GPhNia0FoqIF39aEeHSG50TySHP4yzG7vP5aibEHBhZhL5jbXe6TCDhXyS1XeyVQprp2Tel7kmh1gqgwRgU+vFYL0tOJIgXLBV1UMJ3BtFCYOR+bANkQ3BGzH/0+bSt7PLHq6Ya3SFQcX+P6bVY2LqNh95fFhgwqNjw+8EqFGdn5Zoqt3JLTTKJoNkPdKx+V0io+Zyf+zsKu3bptUB74v3R1JU13YcHmunoY5dqmpuL69EkNFDiVpyE48rUyBTCC0DNhHUQaYFR+ed9j9lOK4MiVti4BLhEnkreqotPCFDWsTKCnJ6dCM/G4jb9s0yjL7h2GCQZcHPlwYrEeQRYjF3kqA6oq/PJeyn3t8gaJxZSYNJjyScDGPiAT3zSrmMQiaymH9EII0CCjJGZXo0fIm8IODZ4mqhQEXkAUwnEkRGpZ2roLOSMp4In+r1tk6/RoMnYGbX18ILN122sZHviXvUCTqZIKIRz95wt+yYbrXtXMOWfOhgZu/O67YcHAa2MU8ddgeh9mXMHhVWSsbRJ2NoDlt/7Vs43r30EbyAwd2KtBmtb5YHIXh3bpH8mc7oesvBkpIi/eWtSDWJ3dNVqtmaU0hxnYURj5E1hMproBdhjZX3+7pU7Okw7ZdURFv5nY4xqqco8jO9aHwTfvexso/OupxbqALp+Bbo1p6SJlWDdm91rZu9T0ZqIC1tFPynWo4xzvzCzrdIygJflWf98yX/RXpGmFW8JkP5KHa9oo0IzTb7Ei56QnZYoAlvtJuX/rDVHKICGzaTY23rmfx8HUtthCy/YNYgetshL9lVIYpEDSnQQiDBYeKuvpf4Q0UX3Wce3CQ0eIRwKg9pOv/2ewQKd4G2y7cvV7NRRfMEMD8HbzRxc9v411yFzKmxNAqrDg0hFZwDoACZh/wJ9P41PLrZq13WQlp2YA7sRtmEyA0UjEm0/Vee5bkBpBhhEcKo+HvmrSJsn0UHExKLGQGhpFuEUAKgF4AH0UAMgkvZz7+s+KYIrJP85wxVGGdIgyN1a0=
`pragma protect end_data_block
`pragma protect digest_block
d798c6b9d72293cf07ed64ec612a42701b9561d87a1dbd0f6360f2a5c839c50e
`pragma protect end_digest_block
`pragma protect end_protected
