`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
xpTHjsRsvgLKxARpDQYxL6vkzf0r4xn5NIwntizWSRABPdV4QBf3iTCuWeNtn6k52t/k/UGt8K1USaFVv1lN6g3pjUG7+sh92NIN5NIaV8jVH06swz2xcl1dJGGa1Ks6/vzowINkLFWNrvkK9XAAbi4rrNLh1yb0SqTLazj5HqB1ik2fwYJCHXdPdSs1DutG9/4GJfBcM/3DVz4sNWenyGb1EJNw8nmkF4DaPmODVVypiE4ggi+5Dvg+/wtyldoNVI8dS3d3HIVVm/0U0zRmo3cVqvwYk/GhEZQv4PG4vcZCA7N1d+L/52h3OZyx5qdCLsAnxPVMH1RN+5Kdv453aTqoAJTj8syoCBHmecd/iuikBi7q6KjxDWsQSBZN3PNTtDYbiHv6jgWrTD7ipqfql1+i7roEY5o462BUGAtiiFfwAQXqkQ+olSr0dhQ3nyucIFVKSggSiWR5fDdt/GY7wpYBGKrEq/KHhZTkQBvefANEz+6ArItxW3wjx3hPeHc6HYhxDG7aRQa/tcDLjZ/ZPs0KV0OkcHhaTTOF0c40JTeXbdsB+hmhUlFpiz58NhkNVlnQ11fcfitjKjsPQrMYFmyzoC4OK1fV0LeV4sUL5Jqm6PwqppVg5dFNOi27G3MDpv7hkJNYo6k9WGqG38/yTzRnrNYxZvTeCNEiEilKGzmR8FCZ2dfgMTO4Ma/UuaklfDovV6yY2LLuqFpx6xwEeZKDKosSmobvtnDQNjFu/mdA8hUCERnmNR//IoNBc9vSuZfcfs3XorKWWCM0toHMEnJdIrSp+hAa5MQTGePEmp5LZYxlLicixYM1YJxJTzQfKUWUq4xAUICmZiWZkt0YUsFn8vH3g6S55G7IgbuH3VDeQsXLIl3Kwh66zMM6T5SChl4H4nAUxotdHceZL8ABOJmNuQjCTwtm2MBcNHa25Dml6lQ09H4LB+N240BpwYlGLbJSqBOqbe8wHDvZqRyf6gE0e7Xzf/iLbBItkjednu80ct9CV7ATkeVhGqUZ1gZGmkx00Zd7aobIpD4vC+JrwSbfrzFULcx5ukr/m35L3hxElUXq10bN36IgbUgosjLS9g/oUEwx5TZxEZNRzrhV2MqqMuJDPYP+lXulA7PuVHtcNV7OYYxxgqsji98FVSb78eDUGdJoJ2EhMuXgLPzw4JzuKH8MFOfNfAhQUeMlCFdypm85K/0UfxnFWbQPWBLXrQYF2mRj0cS9LVvjmTeWO6WWOTdl34FTuFANzmgRQnhiNlEWWjWfvun84gg8ZQAWulOyBl7kVtTQPY8d10o8bnRHcHqFfghxW/J7pYSSIqdrnFOeYhZhiR3Uq9h3iEafNtIEgQVrm0NHRIuNIAOGjxBm5SwwHsp+HVDf85lQ9yMRC6nt8DltmU0Cwn0XQdY0rCS15RlquOcnKJpJNtrcsFYB4ewXOWDjeIxSLM4eRVPQ9+P3JUyDUzj9akcZiqWMU1d0rqN6abHCjg9HSpaTx6WXZHl/5IK1WUbauuG1h0G69qX0Q0EXFrT+ur/2kRwx2UXjCPNkAr4K3imf9a9+1+iS9wa0KjKDxNzngxpqDP1avFaoDq0LQew9tebnusYJ5iG+X15/0sd0MKeBfeHi1mUSCWPVOu9tMVfT0U0o9s+mk+TO3HpfpVhR2VhumXtAyc7aj5CPOdzL17MRrw3jnil/8N21ioGSuvtZyHLSWrnS4qkZ1socdalEJShgNAPqiqrccEnjDwKG358+lgYKk2Kas/UWfyLE2zhLepHzaOyOy/hkDei7tEz1pCwdCP8R37I47o+Zv3EctchYtxHvuEGNY/kNc16HJzoHfbpKig7YMz7VaVnw5dpu0SdDKRXL5aSnLgroIaFasTfavQcMr1vI/jmyHn+vzcxLvGmI//ua0xP6LBsNEmsF21h2lZsg9/9UNxowCvB/C6rI5RSBXM2XLJ0ZqJGBoqsvtFpZfgpgSnQDvdtqRe8ksNmacr3bslZI2uLlTT2T1t09teIGosF5E36t4OZoSo2DjIRmKRCyuXCv3NNTGq8SmVxY+RL2ZJkQ1+J0DkymoQURAbqhlITFUv+0zHWCRVgT9TpmemR6LQFMf/IsJ0y1Gs554a26Sn54fqkL4Ej/D9IV3lxMt7W/Co2jct1zRAxd/BuxIOZti8XnPIrImMHpGWn6PfIwkm8dbdr4xJCAdZoKDxR3BlHZ0Uwh+D/f4mm614vu8N9GIERNAX5gWojEw26q32Yh0IyD/J0ov06+9D4Be/majhz1jB6rigaXjWf4y4YyrsAzRCnFxrkER+Q94Mu0dhbrwOfzKeb5xMsMV3z9U5PzQh2RPLHT3HK6+nGj6pYyIInLf5eVY7h65d75bZJ5vR9Jjdl3ckz0bpSvs9O78GKN7CChcDAa/TBhe0ZqWbRhbypoEo9y6q1vRj+AeDGzOHtwW2ArtS6jBL5jRo5pxiIIzGQeT4Mfnr/7SBQaVIH2nDJb5Vj8WrPdsST5VBdK6uifI97UhFe+2GTTqXe8+LicUWN3hF4nPwvOyU9NPopNd+Yq3i5U2n5WzyAY7VnbmK2IOEs6GXTcCBGIDv4NyKVqicKfqbQoMza3a0G8Q5ZciiUyUt8tkyGa/KSay1IoAid+D3rQBLTbVQWCE4K5dLgZproEniNcQZbhMWoLo17+wYy2wHxS8Yba6TcwzgUg5YxXHHdTOOQulS6VAVeQupUxId3SDKJpE+GBDI0D/isnvqHR/rWzIkyJNp7Qyhun+oKiaZIOItWntO4eHcdIEkhxKql3KvJh6DhiFWTb8+bbPV3s9OBfX21Rr5JxXdHXAOYkqt9+KPexIIK+BapiMkTtKsBBq3cc4uOyD8IXzUyupanLBzKOqm87l06Y2ff8jFao38lYDYnRhfbDyPGMFn6Nfbb1n874qXwVQr/BgSwV3UuiJ0j7ayQbmd4ceUxAtdLwgT4OHUYRBYjzCzlXhwjxXpFCRm5kmJ/o730lLp94uZiQWhOK/45FcuxUPbVWx/ciym4L4O6+9ksDKJBgCRwe7Tx/c1RYK/I+HL9bd7QhJ53nBJ3sdR9whPawhQqHhgAii+wvvW9sa+iF+EyARf5WzSKFUCyah0sB+OxDD9XfdxrM1uJ0EVRlbr7gy2dN5Ow1tDIdnHVeDorx+yJ4NYgIZ896pdWXI1KcszpHTN4mP51hbIkusiGGQYxeUXXLfEGuMMc6sx/xu4VC2d91KF16NtNxox8d6UOGNfpUGiV2pRc1gTSWhQntkNrQUee5uCkUS8ERu1ld04UbmC0Lwi/Xk64MtEtPskZ+8nGZtxGjaGCmdq1h2Osf9KyzPIwHHknahidRB3atDJWwJ8nSCljrXzN/TuRfDPdcT9dwlLIGQQkxHsnqxa6mROxfJmrNkqA+Ds6tWdBABQ1voNMpy3wf7mnYyCrefkYufkPY4XaITg2Zuiq2pTMo/xWyQs8OQSUERMFSIkfiXf4fsnyMzyWtIYtT7SAiZt6PIUcdJZITxQoV1cayEgYfKB942RA80SREiSnrv8YwJJIx0e6HyridcNTvnZ6SKUjWZPPwvrZdUT7e030u1HtX1N5DTalRVKzrqpXKx8aptpQNXaOryDumjstDtcu4PSPPaRZ0hPmnn0fT9Tvpopw4VqajqerNeA+NYFqvdZ/LuQwY7j6gXtTEQwcSjO4zKE2O9zMJEIV4rtULm1GSfULzZVn4vS8lySjOQHWUh/DUHNFYcEvoZJ3ayNX6NKuBMyheMavqKK9KA7SM5Ab6Gkrd09y2nvo6Gk7465BOaLC93pfloHsb/jkJdbmtS5w9MQNkYSoI0CNVsru9Z+BsGSYNpnVtyZqOh2p/s+VG1peadcWuB+xl2KDnHTAn+x7Urg2S1A2/YZRcNQ49LWIpX5xPbYpCrta8ZO384vE1tqVoAlItQY1YLq0j7bKlo/4TpqR9NGB6BK1iVyxC4fQfIJ3MSlXkLLX1EZUZBIr9dZoOjykbQ7+1LJXsZ+wNq+iV/gBiN+M0bFS0Fbab1KZpYw6Rw9mymD2CyEQnYhJQPX5Hgs1orVhU+QXzhTQzzsn77Ro/YR1FzRZsTaFWGydzR6qY25fkBOW/HcACChz7EqIkUR07/fpFYHfC5jn6on7O7noXSqT3HVdixYIOVQUYZhw83/tG9KfNv8z8+htSmN/aadvPxUuwK7KBzgmZvypi8XKClErf6KBl+fEh4zc9DbXGHKYEWFwmc+fBNkT9te7UIbMXuzp0aH32uypgUT87U1WPHsj6lPwmd9QnbN1Xscysd6Vg8vXyxYcOZohqUFf1b1UcLzWB4jbBdzs9hFCdDmwGg4OoclrIcT6HV6MmSwNe2VqguwxyW71v/2id89ipEHTNIpAXXXMnyPGtUpYLuSVD9ShsvA8GxAVSXskM7AJ7jNXPQxmIccA56f/fr2vD9NpicGH4YfbBTt8xz/0En6VdRRyxUs+gjw/P3kWXf/jjLrdf6C0sK308kHDbUHRZ2NXY6h8eVFJUadR++cwovfEqWmd61Q11xcttWNktLbxBCa21STkCsPpk4V7yj/9X8P3mE/cVkgqQECR1AJc8gr9Db1ConMVcBvC6sOJ8Ykp0RxWzViP3jNnQyS11SEZ+ryk7LUB3yRSh0s5erXJm7ymlqEEHrxbFZgdz3klIP0kRxr28I1FtqhUHPzYIwut5YLu9FI0xW0jqgRSBOcADhb6AQKppGIQd2mutkmX46IluDfvegiDyEmUdds1QRSSHVdmX7UxWu5zYuW+n8yX35+8z8jdkpVaAxTxzQEW+0UgwImoL4KgRfS70SKaDEFSkZok32YwZL32GXBkdgI+x8tiL/m6tpd+TfpDd6dVCgvSwfYMfiwDHYhU5Fd8JbLMci1jEAeEdhmuuh4qs9FX6LbdErRIDv86pg1ly+exxh7uxVlnwmokDfSIQm9D88iSWSPLbAtv0yz/WjkEk0GvtMfICL9xS74G+KGu8BU2xPel5ufwrVQulkhXXxUKh+ixT0Pvroj88+raj52pqoZlESKLFDIkDo2k+WCd7vHmdluVcKOHIHPAEwwBxvkuHI/KRvDqPWQkfR/64CtBwXnyqYGtSZcFyPzl8ametww0jBK4S8/7GOftn6pYAQRtFN+z4MXpOn0cmxyoORDUCGXga03LJoxtodj9TmCEBza9awwaMi7s1b+r8W+eRpdgjwtWT7uC2hFElDiYl82d3sFV2teohnJaDnn4uJF6U7IfBGNV73SXAjoqkNoPhHz6Ywz2O/FPK5DVRaQVae9BsEtwhO+2oht6sMr0tsUjmTazpwCbXI59zbK0hJWD6q6gjkRMec8SwUGn1igb7f1nsgi5hE/PCI6+vMw9TDlDilsRwvph0V+ba3mD51Jldep8mWBzG+C0azOUJi4QSSy2YBBdTlRWQFGvD/ayLiLbxHrGhqGHMew5nhEusXrWn4rVribbfSKYEEa/e1yHsjApWvfup5QU5n3hZZWNlh7HAV9w1SgNWH58jtRBX5suTnRPDMKa/XSoJFEHMC+pD3uma2Jatd6LvEQpo6nhua7eL1YDM3RBo8gJbZeiHOjUATIKiE+lypYvYlrqORL7PU4KQeqgkx0l2Uwnu3x6UYj3+quN1LSBCsKVdVmwSguZgPiijiT2tokdUISU+yBprOZ0hylvEDi3TEAnjxnSSe8fFM42l5klC4SIC0IaraSbIczYKBCfQz8jov6OclnZ8O8I4NCtG7ZurU9nsr1x2NGIu3lfNvmpoBOC+QF6M/6vtQFI5cnwiJc/7zbxVT4yyqmw3chj01D+/jlJe+V387DVzwsOwC6PsLASfHTjjYSGxUsTUp4GzzflGmYp+xCzlaoKIkmJNZmdNlm4WUOw7L3PG79mipbX3bqWE2ZFlnQVGarA4BnMBlSF53YHdSHEwcvBQ31kS4Gh2iwAmOJ32iPGlToDf5W9Bz9ufcQ1yrai4zqPOxz1dT3ZJVizq3Rh6UIPo5QiCySz1qDdXh9z59B+/HHdUKv35Xi8xnRoSQV1suSo3owF61xzLzzruk8cDdGSMCNWfFwokd4TLjhNb/yyh2j1+zy8eWjQwPVANUtlVXPTYP8G1vZM3zZ6/kuN1q1aWRyWE5sjRXZ/V6czVO/feiPwlyy+ePyHpZ1GREuFafmpdqEysJ61zL7dATkwH7FTNqsf7QqN0v9H5fa8Cbsh5Odj42M9GzzFgskujYw017WH4U3Npm2IOGz37Tme0TsMo+YeGqpJa3DE+zSM/H4TKlpKwZaIs9QtO3fZ+8MmMwH1MaSR+rpfdxv8/TJki5Y+GHCQQK4foTdpSKPOhv52VrF0y0LQZvZNd+GtIj2ke7N/X05iZrcwdRnCkik0vD1El+OZ/9xGPIAx/koYrDsaSMLIfVqL2wKWHIHf3btzvMhHPp3ulNNf+oae5lSiNYePdpv5jKjqxeXZ35cNL8pl2FMCLEA+MVQrBFIUe+8JjbMR2rDU/cvUkkJjXSMpn3nVIgRQWeADARUlmEennMzrqjwQO9DTEfYiQEktv5I8xal07vM1sVTvz3DgV4a3xvN4RaZig9aHlmYot+5+QIUL7MTV6DDU23UdkpPI8GVC4gJeAjPFlNGXvJzMDFea73KjiK8Vx3K8fRDggUAPOeRdWdLF5uP/zf5mtQc92Jd+iVWBJ6IewemafQcoASr+Mfa4Q77RVZgFQwwHLw2IRSiZujfYl650PCx0h/At7gFQCSSCrSVxit19chnOWoDfNjrwlXF2X0ihWE3DDR0emPbNo9O7V8juRPY4EwWv+1HupwLdKnyCSQD180tCj+FK3WlDQ/wTP6s0Rx0oIZ+b8mV3hNVXfj6wm16+pM6sQLKQguPGdrclOjTcUFyzpyrsTLB9/oo/6j6R//5mTzQphcV/+fbleBsErBCTVE6uLX0dkkd6Ph5VXA+ZCQ54/ZVpQ7tZT3ysxO2ljHo2iLoa8OgBjSpaL3X6ZtLpbIHMB/16Sl8FUC7BKIVF71JgGzVRLioALuOcoDu7p12qa38m+BiF5cUuJBK489lAK8sB8j04LO758cXUX83PdlqcLsIBppeVA1f0uG53N1C4BATssafKjbM8YhIzcGhhQvGGS8DxZYEZjbwJu7ZH3fIQsNX/H9UfOvt0nhghg+2t8pZgvnLLpz0rM49xXqcaJWP/B1U6lPmvdyAJnpwDjPl+fPdfXI+BC9/531YJG0Xp/ioGf3xHLVTBlrMvcz8aYX3YxbYTepGX74eI24sMLMxxbIzDWooNsE/3k9YVpJKR4Tpm9t/hXavBHACsmpeFRvlYHADvAxdCy4nRp7tEFdaaqVVof58vOwqeEGUqjY8EqxQ+W6nA2IDgvKX4dISU9mORaRSCidgRZaK4lJEZw/yD7pCz9yIMJ8d5a/uZ1bz/OoF5L3HGYOMEpIW/EmIr3Joo0gcAbt2RmfZvwCYf3KB8oC3KDayT7HU9paMk6ZnaA5+hSwBpC9kxOZQV2yL+LXzL4HHwjYcGniyvrFEg04a41XUVWcomyKn4ulMVqyMUIQEnsNzknfw2z/QPpY0cTVf2sKAKWhDqkTtscQwLw7TTgv7PT8R+y1YobpfqHLmHbEhY1L4KHPCeD5gz1lkpR0w0PRDvo5tfy0oO6LHQnea5XN7Vmg6ew25U83ic5hyrWQq7xqYv8mRzncSmbo374MDZ4fSN+y6BxN3s4Omyg1p4vpLSL3YgINEnEMedZ+IVeWmJeDnlGMTqwZdpFPPbKVdsogPhlR/jwplUO1F9to/8h/Is5gqrQI351oQEY94CuWQzKe1HyKaLWPFtmFFgjdLy2f+KpO1Puzb6nyxBOwG4IbFvQnkQmQEc4/+EvuyPmCzL2s6t32BJ2YxWRpFGjfn85LXOqSciRKIUzZ0leV2HHrU3Z5+S4bjEz2tdX0wpBIElXkdjIPHQPSHOE0WUJh9or/hZyS3q/ES4vx9ckT5kJ1MAZC/Qce0IXGO+NbjgaI3dKEec9xOVrbz2flJQsYvklhByuvvoB0SpemgYNF8F5oGvY9BryAYUmBxxhfGpzxze1dsLsYF5ZuMy6gpUCpa/bnpL8NwxvgTM3lMHt9fVi4uPiDB1IbNGVCamgU0fCU/TrgDMGkLnrTD940IyDc5KsZ6cubxLs2EY3uW18Tq3sTR9l4q/AqwA/my5GO1wMUK4+2esyR2FpXLhZxDJg1vXVFcwHOTBLsRhjxaLI3KyWQBrJ3gt4KpDtuVFmFW6xUVQ2PMVYqyiVjNNSXQBLCabj3mblfWxHxrNxSP8I5sZCFZc0S6zLHCujTuRSnV93dkp2agfOsE+qZZiShQCSi4ctY1w4Yw3mJPajcY+7PmFZTZN+L0RhK76ShXDBfCHiJfpdofGSZ0M/smWShPh9FThcLwbvXUXDkhTRbEpFKa39uAFmGo0Em/O6igzLqGPz+BiriIy552z+3ZPKsDJk6PHeJ/046m6c1an7p0VQYWU9jyQwYhlSnnxV3VB6R6wpayND3+oCfWqN1RUAa+WDtZ6bH3+y0Io/ig2S1TUnTINTGA6Ni49JC4ue+iR5k0jiPuS0OmlrP4h/9129Rm0umXL+wc0sgb32S2FifP1KLbVO6S7jodatjEs8cALJpmzzm4cdBjAO9Jt2HHR0knnAapBibh6hdAfptVA3erhR174vWSISBxhlFT4kghHEcrsd6Olzxi4/ODjaaDzKeFmztL+3rSS22FGc6ZJUedlfV4t+us18fj4oyk9fYcsMMcqc3susd5fSV4pECwx/FxRvZVWfZSgPqAXVID1Et2YkBtDNsFKXeCYpFfSFIGmw4Wfskgp33EqI0D9ZOW9s3LOTC7JIu1V0thV89oWJXAWs4VwIbsbeLshB0j/TlVJ6R7qyl/EiRhK9QAJthvQf+9DjEc34WNf43fQQJB/klKhQRojnXONRB6oLxiqD7Lzh5v+dH0q9whHvzfV+bQwI0bDw96y8+OwZF86gPlzav9U/z3RCY2vnMMSx9uRqkohp2h6QH+E1CGYEMrGEH7AsbaN17PHDI3UnG5B18E3mz3wIuX4MI/E5kV8YWld14HMekFu6t/JRJlaJo6wnvcJ4/+MuoeHySKum/w+lq0w3wz/ySRHBlurpwYyeBVtREaWnwGzyR/MULIzwWbaeGLcj3dJugsWU5PJcv7MgT2U2i9OFYdFEMeMmKVZaXC88eKQm+Y28eA0h6d3broBip2JBQTeTv8JwacLlFwuqZbvZg5JoJcwwz7JdvNL91TUn5PsMTR/ctatIb77y7bv9XY2rDfcd5vqqlXEEPQg/FE0XxmbBQOaVyOkzdDETr01E+EI68mp5N7R85GX/nL1ws6h8mZ7EmamqdS4zdTkPlKhoD0oq/zXHoEtWcpJt8OIMUpbXSdlrWi4pyacH7kGEYU+461NcBMO0t1hVl36UOJnDvh0p2QyumgwHbvwSHZ/C123TLodAdBGH0oFlPWI8H0BvcWrzYITHWUjoSybJKG2zjBu5MFRFUYZLJv3lYANBwbQvbzwOJT7pvfHwnkfopOodPgSfjP5ST3E3AyNiajoS911tbtWOtYBmT3fQxnxTXeUZjQDfQJCpXSbhdTmDmEIiH9O7uYHM5vhB1Lfw34rt9H3ymfjs4Mg/YJWALT/0aG1AqAF++GVRiRCHYLA6lD59kuwgjIPLXWD4ij6jr/gqo/esUTqMY6Vier/S415LA/9ZWl1yD6PFN/VTXkS24PsEpie6T45Spwy0/zlEgLM3j/5gfq4oZaYKeRoJbPOInnJCTbt1Ivp4TTZGc3JpyNJn7DIvdjjKLHE9lN1KWrUgcbykGKop2FsHiF74P8HDnkbVEbrwIOFrs1Do97w1uQL6wotMKq42pdIB2/7ZW6L6uWOmqR+Gn91R5nP7SpymTNXHvECPdxUm9mHQoGNL57w0sJuWLy3lui1fOjQIbffyM7OX2je0CtcLqisCrLVc9o3MvCxkmo4A6WFkQ/oqeYUraEjhce3wNoz4kLlHwTsjeXeYJVsHs/xiSSMhxl6RYg8GF5VPWRa4PIPgnVQ6U2X8p7cPV2HS3jxFIuZDW5Pf5g+rUc0H+vo8RHE6nHj/ZcXHZaHgvWdvAKmCPSVNBzV/0SvJX+FAb6H6xtGxHFolRhJ3buL2nusDr9zmJXJbTgO6PbLL7sLW9qwfOL5Pj7MrtPayZuIh0b1rPuYb3tBYwFC7jZystvGax4cJzFOLxKjdP2nqeRw+Yt2MSF0t4OSKi+CexlpbJn3Gs9kdU/CczSWZMSxFxrGnfNjvdpU0kumCGIwK0vJZIsPuHcy9yd7uAbTiT9YyXHmZ6zh0xs/zKYEf6FJDAF1T8GrU/ABvokp2JB1xeOKtIkC5cO34C40MksCMBqWQGNwNOX2hifiuu39xBOrD43xBsz4hFoeofqBl3J8gj4u/r3khbZIREoLZr6m24KBj1QrCj+6rscDLkAeCwFbzTMPvHNc4q40lUAKSpNttUlgg5Eyx9EuPRKdyAiDUO9YcDkEP5osBPqU2up59GtqO1lTT3RymOsz41s4DEdiZ83tx1kjRy9sLBH1YSMzs5L9Ku5OMuZhueRUoZXMkAdeTDBTL33bwP1zomoO4j1vbHLBbX8kbtGQPpMMXSIblf8cA2nVDZsDyvDHAHto95u2MhMHoxu4T8DizUOcAeIQ2T6Elf1vCgGfh2y4I+OdW43qv0xbS8vJKPpn83YaeK6GF2WoaQo6ktTHjS55lZ4YGKAscqOPKae2jaDbUGeFT3QIBrXZQScI0su8A08PJIHv4Y7xTEGVWAwiNYCxujP3pDz+Qy0BPjE08nQAhf61wR53/fvCoCFJpW1JUnv7iCUv7EAc9z2jpYfzJuvS9IC445F2PM2o378nn1e8jY9Eqwb9lBzzvgGm7Ig9xMDNSKQW/O/kZwbLo/nY2TYUxM8cd9SclCCavFq8hzVj+JoFPiOkh+pJ9G9q10Ce4/QQDjT5770c/JdZU8RDVopi0ZBTcemS22tWEW79by7oq+fkRN5YdaaH3uiyv7wNVza28s03UDXHwMK6vsIBhkHqan9/Pank1BzLRJ6lTT1rozv4Yo581w/c7XHU3ECNt8YC1Cqdlqz14bW6ngRXvKx95lUmfib1qJiUPR3byi9vWd6eleojntOj9Y/aDV0YSC4SWOAwDXzbEttaZ+B1uE8piujblVr7ARxCD4pl76SXQD5BXHXq51uHMAeWIwTAYSKQbLdERLjjf8+3wd8ipFQ0QQs5/WokVBWuapi95Yhc6nTUJHFmpV2Ubo2GJmks0yuLSevgNeKMx+XxBiMZWD7Ra59pqxtroWltUrnogDI9SB9FxQoRwSfAccnTcgICl6QywWijOeb64qyBgNdbRao+6lW4G58PxvWuwsagLijN4tt+WoiYGvkL4CS5wrMa1eaXCq4BnDfTcboRoAhRyt7PzSp4GvV6YkHsrSsiZmMuEbQwQNyHW3opIA6ngAmNUP82FIy3V+qQh2thlroPuk3Lr1BFKOcbS+GskbP2ttuC5NcBXie6SEi/0Aztvt62jugDsp3IHqycsTZDw5KifNU9j7pTqAp0ZwKcqGfevLzX12vmKtPRNw9xtZLZMSDKdUDgUojxLkaHmATIdXwIJHLOBL47qLAT3h01SoTukT2a5UMlTrBEQFGN9sjdYljLwlXOelzC0TY6LWs3K0uYD3tk4ArkfMmPDKgmQ9y+Z0HkR4dMdX9tauf0Z9/2wj15hMnKXp7Bt7+jyWbdamCzUPetTdM6uHU63l938q7l7SFxlF+dic+7VBZR65BeOaefBuoLOx4pTUwiJFSfVgfyFvHeWsEg8LgGuSNGuefjT5iZD6SZYevY0wtxSjyVfxMkL4udqOOtTp1pvxXp5mK5uVq4P+rEXUTCUeHQaZ4vV12gjN8BiCVWnY978WS+YnULH1WwIHjL4IqrSSGkGO2GlJqWCZUkw0vKzaIyL23ricHQ1itxRb18l619vg3rFPvWm3x6KaePBWW8NP1MXgqN/UMLZBftSDpPt2UTS0jIdeiw/4JbL0Ha43rA8IcHdKKS4hyQOQxgk2zLKrDZBDAUeBeL2tg5e0EB4a6WHwQES7QDdonfaP3OuT/TV5BWWzCgoGBpjeP//PrJ5/dEJ4TnNAMs6lJgBzEtwZeVJ+/MAzmDQ75r3H+1XwjRID4+DQmIcxwK8UYD2pinbbPKTPhJiclLIf0GfYnMzm1SaoUd4jmamD3UFSQ74IEdJ6LqwpR4SUQsekcqnljcZhFqGTTujNW8lOLd9ZFJPs7ySU/8fDW0AvQgxSexJVp3ZzQCRoqZ6yceLeakoERFT8nQ+SiJHNqJZw7TIMIIWkykGb3SnfQ0ExoMv/D4pa2gecHkV97QVPCTGfRRO1UmDXirKCqe0zEDFPVTHe22ux1aMM558jfs6h7KCam3R9ueGCYu0irTbwG83M5mrcuD0TlPtWEuF91sgMC0ybmpeKtqUMJjQtZIOoM4kztdK4dRMxQjr+6zltM9+NqwJK5tCzlHgHaK52hWfYoSqkSBjU3V2ZFx1KnXfoNywKqs+etViCnMb/+WoKAiaeQd4wFAaPxKnMZMOfiRCE3NmWkeXxOVQGRZXI+zcwCj+BZGMDHv2bzyL5oZGYbK8bkuaVuvrHX883+wuoub1k9VnB0nymFvWQHdTmlyqaaEG0NxSDDiFv+skUJdTrY9y9wPFMz8nHpWIWFFHZu7NEEE2eZeaBpoDmGFRd0hjAVjvANtnsBZyQIcoXGzUUCqz3uyBEgb+0rSvj8O+xqUFARTSBxXhGnax3R/TwrgI2vDgHS9xHNTaHdu50IbSMNBLYxTGMhDUxUvIehTZhvPHAgAms5i/fHn+l0+Qfj3hCSyfxg2sOw3ANErtPh060NjYgfqMhOymLh4jj1jM2i1UGuCI5CUI8kv6NYm8zhLJFRfk+IAP3M2Btuz+FwfsRAPF2EtfnE/Hm9cW308pHXag8F7n5u5idAmWU8l5q+1ojOyqJqFOSvAQYPCE7BCjLWEm5Fkkr3djNRWxrL8J0JnABmJIfS0pRr4Bpt2Bjv/szAhNm6DEB1mcH0S9qz/LfgPwy73dQYQgobG+KK69XJPchIvgozvSboDEquluTJ3eo2D1+Pl1yUP/yk5Pmd/IK8LGDeJX+IqSA7or42hm9+i5gYTufBnfA16UZrsU03niqpiOZYr79OVhK8bWTtCKBRo1jjAhvWJUWDi36Wmjz71PdcPYLgFAMDs6fcusea+ekCGPhfceX/FgS03W1x18mc0onY7tnMlRleEJerD3x37Fg7mc9i8A1IwzP4e2x2C0olRFKj+sSPa7Bivw40rgeSlyqwu2cbj0j07sdNigpal3xmdakN7+6mezLPtWNvtCZ+Aingf5BTIlr5zx3hZNerIiPX7tsL3dcCf67xrMyK/0oPio0XPjR76AMOpxq4GaRwwW84PBSi+nNJ4MiOnfe9HaDspTlyqjE9wE5feKvi1B9wKvA2XXUslw6zbJGLie7s4TsIJlr1im23A+yLZnS5UFg07r/fzPhV2W/1ay6of9bhSw6OTGniA2eUWBS4Ryd9KUSSo4vBtVlpbwFf4yVrD3NhIQ0+xYs1qWg8gmdHE82iVUQW3h/2zKYSdFLdhI8qDGqSzzForK5+nHPwXWeh0SzK40gS3eIlQgNYU7EGniW9uN72Z3jebwxs7J55RrHBymr8fnHSlKmk76+S/eydGAnDNYkNE7PexfYCjKbQin4ZjOKrXJH3mJpFWo8ULgwWYXtMUAsKDxr3FPjZdGJtqEM4s6EaEFhLs+6D4+3DFgrSV7or1cm1P362t2i//O2oz4ZVFmEX3r/RoEPiX3FrQAL0vbCcw4EZYFJpXweyad/yCsHZI8Mob2Ip5pA0ZKo/THfDBZ2oc7IBOzkQL6C9PilNckHvXwRSLNvnuje0iaEdntfBeS1d7/CJGBY+DkABdTP9uDbJ0iFz0ysC9YWo4VFmHXRI3iCQjs3O/DID71Mk1fyt/v5WhAAJDLDw9COqVIzPmo4fxyAQOReB2g1qdD6ALfwkyZhxA54rNCcRxwSKjOvNEXD3U9qv7+Js0od0+KQl96dBjVjDl97ClTD5s2aHqO7hV1tujLF73XRX9Gj4UXLmTg16iktxwnd1VV93M3LjGqxi5RcLGAn0eRe8Z3OGoJb2sX78LVQjPO07mCxpd0cYE5rZGpEbfJ4VVQTTNt1/PogkK1Tef6ff/GP+ks9G/GE+etHBqiKcjbw+H72Lxu4FtIPWK7duJW994ZjK5cbHlx42nAqOhiK4cZ96M45gjXeZnTiZUV0I6l2VLlXUxw5nKsQIFydLFefMGcikhPCfiiZoMJSVjRWPKm4Mdu6HVigjrdj0Mpw4pQVUA9sQUt+2w8ITFDOOeqfCvQiUgNgRdzbm4hj89R92A3kwUjx+rRWSFGlwjyMTzDBOcR67lI0L+e0v2nbbeOeiAU6At1XMbv/2GAMmCH3qOCvSF7VMVzVVadhDhaWlM2DeC+OI7/JSB3oKZ8gJEwl94JBnxIG34F5cBJTIWoU2ALxKRj+UV9MQZT0EwhqfyLMQfFgrmRKfDThUTXUO5LPEvTf72qDlN7twPgyb/fYP4kF0/rF9b91TluXEoNXrg52XWtd0z+IrIh6+nSJj3E6zCPRKZJJ6pmmNpamfTY1ziFroNXKRe/fLiOrHQtKhVPTFggvNI98N/we/cEOM27PUGQN90ySDAcrQzv6DTEoUN+ZIObAuiTaGXg9imtXLoHqfMwmud+FG4LiJRuTwoEvtO0LeIJ/mwwIB+6kun3wIsgnKxGbp+Oa+LlW3H6qajYkipDjGEvNXFMF5WyV31Rh4knaq1nwznU9qr5pcO/NQv/HJOz4EifTPxKvQgb8dvTRAoReUGQL40i5ZuCt4IBqG3VuFTYpObbo2jPJZXdy66wi5WlS0orA6m7BfQLJ3x0Oy+g7iHpU5Vl2ILxUy+c1Ya/AYEssNHn5d/01ljGjbovCvEaP303724Ek2d7Yey4zdDsSX2lJswBF/IMzB5OfIFZSAaziXHhYEzhmwIH7R5Ouh9rd+9qVf8sOjlAn86S0/vnCrhX/TbH7aGNr4vnu4svxn5fJunJEpOsdykDjVR7ELvD7tSn50qo1A==
`pragma protect end_data_block
`pragma protect digest_block
f060403a571a337bd344919e0876e79b5544859929a87c0b0e4f43cf387b58b9
`pragma protect end_digest_block
`pragma protect end_protected
