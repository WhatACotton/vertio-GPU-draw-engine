`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
bKNJs2gRVvye8Q+cWgcEjFPf9FsnMITDrsYK1Hvc04eWbMcr9at5FyoVrWjW5IFzv/OtIPQak47+kQlqVezFbsB28za0iuAr8MCDxjUEbnxgYlQ/j1OApPuKbNG7b8YfCU8TeFZzVD2ufvTBQWFEqP+aLLU+k1nBtLtXobZzb6mGZeGSynh1zOPJ60cTxo5twAxKRziGRrJ4fPV5VDA1u+3eolFZBnRRMJnrS7Vc4C2YDFXy3DOz+b4cmsgTcLx1zY7wy/KQuEc2aVznG0exOu8OGrp0hkw7H4jdwgb0eVllGm1OViWha+WzvSxOo6H/Gyw4xh2VO0ymC1P1k3JWP6kSr9/oJGdMfO9BHqu0om6JJ9r8jK9YzPUtWLXmVHeHATCF1u8DWV6oSDw5KozJyqsVxUk4HVgJu80k+kr4jfQtcBIuY6W0cyiFyQnng9s2WDQe1sRCFFkFGrMfAXLhqTTAh9SFp/2AHyH8yVVYsl0kptMDrm8mk42lrRiN3YTsi2VNqftpzQIsAJ4ZE772WOYA9/Okab3s0kz50qyBNa1lzYKmh72UMAppsVfIlK4aVP/tbDbHpXGuO4RFjsgXJ/GJ7VvNV/AIiNTkROdMOcJOKHL/NTIwfUoKjyTOZaqQk/SKBndb1YC/7HVcgSO/QaIbYL13YBb8nepB/HGMjSCp7+FMy0WifVBIEoZgZzv3JHmTPDY3Mo06z+wREsJBc27R8meHgt7b8Hp6PeKmqN8MLUnsTnix78RaFeSUP8G8zrar66PkAOCFnTHNUI+UYBa3pzKVttJyE7Ch3VCcge8pwnWKXYNzkrBU615gokmDx5uQr75D6dJKGRrt9K+sX8COM6kgOn9Jya+yGjr7wWxZalnNR2jpRZlYedDGFJRY60n5/WOxd/uRsE3OlElMrzMGoA6YESbf6NV1qdMMjxEYs3pOuPhTFtowztt11TqAjcO+9+9tgAKLULIJ6/8jL/B/MYztu30OSz6x1rKE8e9E07hnJOnLi5iZd1qnkwrq4QEdhi6mogu93VxGnl/O18MlhixJl+ebcTbrkxF6JDXU2IvfcN/q8+WqoPuPycQfh6Efy8XVCRC70v1e//l61H/PsIWBWMXCZV21IfM8QfQDtRktDSul4PrcSz6LKnj8fpe4BVZDLMZMUwK5mAKs6HFip7mjhbTZzyMA+Z9JpA/YM4xHxcKRvtAYRbArgaiXjhEST01gAJGI/rpWWokcr5Glh3+ErfY+kaF+HSlh7AUx3QmgaFKyDnilLIKWKhHccxuW0FiQjHK1vRMB5k3GGEzuELTVu4KCPx7K9QPWbV0usARlKNDAcLgtDr3KKaij97FNJLWwZPkllsmtrOYd4gCzqRaWC5syDoojkKzcKNn3Dae2D/bRBvOUFxhgJwc7la96sZuWRF3A9/kRGDczO6rllwvPmUEA+3VF13xvqRxTWp4hnbRigwKu2eZzBH73yvGo7aTp5GmYz0OBX/P+TyB0oi3+tKow02S03GkZFU86j982r64nV22a54aQ7vv9urNXUAZ8onhAx4e4/n1KMgo6DklufKmBIljEmyN31P1u8/LHK7qnFOW3LFGJ7i1dytik88YyIUIbkzB4gke3Od5W2lnyD67KzTmKm4bgweULrCZToMvyTk+26h4puwXQSIEweegna3379liHNYA9n5dTYnzjH8TKidgXcSCEvv+2gCwKF4+2UuO9IZxCoxnK/6KRco43tWWGNxW4nqFmEpyPcpsz6iYbZr1QRIcLjSi6LhVVLWG6U63GiTSSXji1joH1qE1UzV72GXI/rNwgBnNCownl5uy3JEsMAKg+De8DdGa34HrW+vxBSnqPoYUZZ6jOksGWSVVtNi7aZi+8EJVzmhRp89H+0sK1ajRiw4kejHjkrleJbtw11lqMGdV71gr1Oa0uA2312AMwYDvzxwLaTyib0QXl5o7ngXnSBmhAdA9gS7r5iHKxFGtsdQn3A5FRVSyYbxyVz5lEWhPmxW/sl93ImuIqfUuMLgxFMUHNR+xyoDAN7i5A+79w1pVdO1iDhUg/7AuyODMcy37dVZJP4YeNTskAuvU/WBYWsdQevm9smPpDyFFVUs5Mb/3dcEsUP6Ey6lNbNA7QIW/MO6YgAl+iJdt7is4507VkOl0FymmBfa0TLNfUHyBADEK88C23ifPcwKarYtqTMTwOCtIyOZOLsOYVTDz/JW6sHb/4sq+/wYHCluAosO4u4ilgZq3YSqDUuxo33QGZbYqapcVZg89Y2WjY/hZoMP4yUVUr7KkTJAwU7xVZ7Hv+Hi8Mi++nLLp4qOi724qM4x569QIoqr700yXuWOtBHLLuOAtPCDXOvcyuAElshSVWENVj6+83xjF5Yn6+uuZJ1j9hE5CtXJBQjWFuDsmE9mJnuGgKUwcq7ihpydVfUr6QVpkl2OTaGJO4ppr+beO3/RmWxBPxi0rLHN3R36G7sqiAfGJVqt6f/ejbqhPsZLMhPcw2whc65ECa+lV5zsSAD11zwhnFzsI/5b77zobUAIs85ZNOzFvY/Jgnuu54x7CHiq5zhJeu2+7SRFdOfTK4goNMf1X6estqD2awJYthcRRW8wlGnuarpw6hEVv7m605jLHFu+Zey/jEy8O4lW32OEV30AC/DU7iWiRiv7YF4YIWFiMW9HdsxxexXnz0lRxgR574M2ckxe5h+BLMRiANeh8C7OEfTzBGqUBD/Vkjh9lm7siUHaVxC155xX9Fp/+vzK0+zqOsx/MONhzq4xW+UuzalA8cBQtRfVnUnVRLVCDQ5LeYI9GkSreis+zTbZ4OJ9NnYOsRyU/UCUw+7riDj0fPIUVuM/YmG3zk1qf4U8MvZv7i8baV9nMkPsxlHiYx7g3VJAr7NqSWRBKfG5ddGbtHUy9asy49qRPQSmuecut/HTUpwM5lkGJzHL4GVnJnoaFRDM6Kh5MP0o2dcrTqQP38Y1be/oLqA9bRXFE9Ga2J2nHbHydbi2to+wl6e3liuUsoUnSpKZ+9chcNXrLXJrAloO3N0mwf4p3x/R6+xChbznSqMchJij4uj1YlFmLV9GIjx3Ou5ckr7jRm43bTbOUNnr0I88j3z9DaCh/7vgXZsrPekqrMk+UYBByYR8wqbS6IHimxcvdjinEU1Y58uVi10pgJjWAlJzhbviKogeQfloe464WkiUsvKp7xGsRwEPjUqsm5oUFZeQkBn38FU2PM5YzZLsuRvG69QwTLZWE67R645Eky4/6LhcVyXfY67WVRiqbnzV+rfIhWurL8zPqRk1pOo0ustdpn3z9RXGSX1Xb6kg72Jz5N/0DTrOsQFoSTTjBGoQtn/Gu1s4SLL8aBFO/3qwUGBlChOWH3BpE4JNbiGRwOkH/L1B6pjNqXMebdmxLWvH9x2Kc/W68bU5sTvQEbDl+Gu3RgN1PqIgMvcBKypM3Q2M0O3oR0ISzBBgSRFT/okMtNftnHjfzv6LLkJZsZZTDUzBs+QPLSB0rhM0ddaFdEPwY7udzEBHf0SdzWj7AfpvbNnwti17ot6/usTL0As/bfY8b3i1x/23sDzBric+3lb2DK83mysdvjvYGwmbcuraBtwCrPDE01XJ4q6AM0ftIbBtIWMXKtsljERL3oFQ5R3k+Wtpjd9kY5P29jYIGEZcrmIb79alIHnw6He389ocujw3pUEMyW9zAbvoMFdMHj/JXVX7pU8MaDnl4TTz95KIcKHTljWhAxJ9bJ8mwsMbM6ag0x5BSm/q2WNpkezNjsN18REjFxu+JXdKMxYHOrWlLqt527uj8BUxK1WRVByck+7h/PzZlKQJ/39jTEZdOlKrrxTcCp/I5Gt7GYO5qU73LoP8g0e/EgNdp449QELx7nzs312Cl8W9kWJ3OTPryDN62zdrGD3LKW4ka3AfMKKtBi1UybqUoQMEXwJyoMq02iyE3sxZFJ0Q0XAMF/fr3opZAAQliGFCEOTJl2q1AfjlBepFJbpSBK8nyuD9GpAS4lK73l0E13BbS9xJTznR+DYT5arqeQkmIF98FIjVzAFO2Q8APoP/mcf0zEiql3vj7pNh6j33cxYRCKyk3pZG/FvcfhbO6qyW4pGfri7JrYPTyNJ93r9TQ5oGIOVGc72nJA45aS+qS81RcMNKljYKeW+ATdF9oZVqNMIDXfX3HeCatBOV3bdnV/ioukq3OJqbarX4ldqciiUx8Rnzs49L8PhSBjfN3++V8LZ14w5k54TaXelAFIEUUwXkPMYspP1Qa2+wpzx2Lap9ceSOaGcbftG3kHPMNJC2GoUVwgkPBA/V8kduJYxbyxtI/nQUPCYSIR2QO0GUlzhTxQRY3Wb72RnoUR7M+Y4w4ZnRm2ufYP9CdECxwqjN4xQ2J4KSxSVvg8B4nNjlHJJV7WAinf+MoM1roYZk2O/kl8rHyY8dOIgVl5vekHlWVaBKUDoMqz40xtRoOVaF4HQofIIqZwjefWVlyzgc/aA2SVf/YU/oK7DNEpVCqIgdhoidVmW81yTlsSZgFtdFwF3U6eLTI20dNfTbvv+jDdbBGyXZdvWigNpdDpzuWKvBXtZr4pkh1KIl0QiQ0z5EKh6AFCe4eMpgpX2fCl5rjnvf5WBp0LOZB49FWc+9UbQDFFlhrTA+BYfLQa1N+X1TeoDHq9NCptcRayax9E3wpNXyUSnoROhycpWZkNMnSaJxhJ4XZfpu08V55pxx78lOsdSX0CWNRI66ZLxc7zWZ8WSB8xLlah+oZhoFAixbraJjjU/IqPZaJS9k0hIKVZxt4oZ6DP1xBb9uZGbmb9fUjidmzh/lRQBoWfmRzpG6IyzbxFioDz1z2S0WIY48tRiSjzHejoQjT+jLiz02KoHp9waGA7K0Er9EqknGZrsxP5ULJNEfNmtvjJYJPJhFGhFcBhn/2IA7GO068vdpbEfSrAUQhN+R9YVQsDUHLzxuSVL3ZP466kxDsypktwyp7kFW14KTGCGxzGaUhGrpPEqMKCKmCFZqM6cR3n5NF1khSnkTgatLiUEZBCZbztvkq6tPaNOlq7STnAfpP5nv9ppvZdoKsvBOlt8omfUNr5OTE0VRcibez/7FQZ9gXWjy4sjf5FByq4GHHN74Ke8lH2J8f36KbaM23p+xvGjTpUFV8FeIlJP1kpO7tiwgQaTh9i8G2XlEtTwuNtuIN39IWsJaIYZcSOq+35Jfa71LygKYHfzx4OFfajhXyu0ZZ/o6ZOH5vtuxLPQvnlCKBNAGzO9LRsSV+wU0j7cxphTSEV+s3Aevc62KP27TlnFZBoxqj6S8I4R1QQy9CUZVIV8AsVFwqWXTsuXnn+kSjyhD1zw68dRT6qLD+V3YOqy9nYnczNXHBnb6PRlg6O5NKWKUvQIwJ1vAvMvljahgweQhUfJhZYZzhCZnDJQx12U4kZXQaRbT1zsN0wIWIj/1S0Kw26kXMeojVlFSml7mmFrBrxjjiGn+DvxXttF3ipRSyirxOPKU50+65lz1hnE72nPcfPINbXTPnfM1dyeyozFE6gbItGUEybjD3MOkkfOXapbyt2ePhX+RIc10bSsy9ZjjBmboO0tnvdvd3G8hff0LysY+A6n1wMDvF2XR26ayR7Q9LIz3vl8Yw0TlNb5aBkldW0QJxc0dJWgKFFp60OfeU6ZczqU5/Exc1iyD91pLCzyw7EN2NpEsXjmePoYfXGB4AJhjLjwZuk83L4mjBnrLTVJco5ESxpVLH1N/b60+sgToBp4SkjmEGXTBNJ5o+FuriQioqZJYN+ejH4bhVJUPWaid/UucNsHa0PDWEU7PbkKwbdoWmHF9RLX99SJP4hdK9K6NmYVsRHbjIPE8uus+sLwjtcEVnPeOS0oHTdceaKdoeo3ke53rr/sC2HZS2BHAwRO3M5OKjXb5RjZ0IqCinvctan6bI7HRL4Og1wdhJzSu4p6mCVuOMWNRiTiKBYbp/dDURVdxpIzOghc4wvMbJVz/ivbuCO2qjcCDllx4PVwlDHaVOhl+kORgMCSPPuoAZenX7Seno/9pMxpcZg3A+Kb9cm4FR2U9hH6SyEPoA+qIC7v6WzrDYz0DwrcDvaBs3r+AhDCyz9Wy+l03M7vI2sGLw4FvRs7PR1gsR0Jp8EamXXcuqD08Lq5xOGS5CsTPGxft+GhbuXYv9EW7YF/ZtdKxRspWCgnDJhLG1P4QpIC01pe65ypUeqhXnbo9kdXCpJcrXEdupaPYS5QOuNbajnbn6MZ5fqNQHCb1h4lDIaXfrZbN4X8p6FUtudpToneqEH7TkUoRjvFRl4XPUTOYVFtvpsO2vIXxOqhvaQmAFkZGDRiEgmILWAVTX3KJ5BhT6n2uaHz2bo3BGEOhN98OO8yaD8jwadnNOagdG8B1vfcN7wcSQlUr2ayMA2fVWwzQOaliEqBJbIrlao8YypaJSCq7/Qm5LP3TMiP/igd2uAZID+3N/OAfGSPteICs1KEZ4Fv9V+RzTshxdYMxLMSrTQViMjgJNfYC+1UAnX6gwXJg3U5/M0zs5uoXqc81nxJlCID8G+4mOG+g3YtQac8vs7Dxp8QDqQhbxlvHbCZMi0yd+69wOiK4OtRj3wDb+L0Wt84TqzzoPSWRztL1MgRfBZPWZ6cF0WakWUp+crS1TT3IJ4nNL1KrsYAWLKir6NsImo4cx7DfwZa4sjFw3LuQ1iC3d9WwF6t2Z0PoizZnxfM0oA5zidB157z8xXCmULBdpUoLWl/O/5KrZZExbNx1+N9y2bdOJQl+1djj5sK2VeAHYfEiljiyMM4covdwCPTETFtfLcqqHFqU3ZkWd+w7TdrP0t43rvHr01q1oPaUrqnewR0CvGvdJy69RFBYifi4UJJLDqWZCaXtGpifRj1e27i5+IxyJnqT+wWGYyRqRZ0C8cfpEsEpe5MY1/wSg9/HTrkE5f9RdBJLktch57g/EPwOkhXddjh7Bg3Xjwm/LQUr6ENEG/N2KXP1gUHLOYG2tFGf5VNPH8EeXce++y6DYsbGFkBw+QexwJw+MtTEiLGEAo62AjGwMVUGgqLOQoXmydtiCBqsXbP6vumhguj+2T1i+jBjo8iH0WWCYWC9HiwjFU3TDH7fO2LhOhX5c08G2HnxYbIu7knnuOEShsCPD/fRIiLiXe7WKX3yrBrfimDsXjP6EYyf4YQ9SROFqiQiWS8A8F22toFbGLX6cXejOJ74MFeeK3gvkBNMsCy42LDMVWCw84JlUZjOt/xbanJ/oh8IQICKpnGGxcU8uXFO84lvBjQJt3NWUHn1YCgW0F+MsB6670cMLqPEFcRuE6ZoA4FTG58EIx225L4OQ9N6Q4a9eehyiUecoZZFJVdcOa5qtn2PjOmukZA2Ka7TyfrZYe6j4ndOVsTjNCkbCBRFcBXbiaHlRURkVZXE0rvEBSL5caDIv18sqSNzHF2qoGNbqANkmaQakSH/aHtX+81chNZG0KQQriDAl5EWHurTUHx5zJlw0RcemYZrtSaeHedWhIVAhQxc2650fZ9gYPZH7htcWfPN5X79nrNN7LPf3pdoj/zN6h+EDQSemv1KAEE8ykIWVay4GWc2g2d7M6nTgmoVaFb518AkIp0hOJqVssvXfPWQh/qHac9PKttNG58otkHPhWpM0KjvcpTF+h+KhiM76Xct19tRteE43CUaeQ3pAmqtX79/kqveukDKkLBugMZVU5aPsLoXTv3+lOijLXM5Jwt34jMUBD6oS2oRip14iW77f1gXGgFvAhRT2Bw+eavBryhw9ySwEIRoeU3cpfEjdFj3ElyxU20YvbHY6cfrrPsciLiiXTsQY9Dm1JofbkR5FGe5xYK5wd7E00q86d5nhZEoyVMNfzHXofQ4ZO3oLtU0m2dCtFNnLqWPToRgWptBtW1S7TjKieTw2JgNtZPwxT1q9Cf87KBPrRaPrVeTK8GB6yZ5Z4K9lslHTijsK2pmc99R66o+k0AU2AU1Nootbt87qsb68h2l3tg8uPd9V1waKEUnLCw1+AiL2PnlQ9fottiArF2ojLHyD1vM4tH0OCgla1BbUc0Rp75VOeZzFH3RQ8qoermozcX3YROwh5eelBDi+UZlr7Znjjl5Hh07WrlpYDmWNUh/jbha/Gn4yl5r6NEH7JejJDXZ1zAVr51ByfNxQwQ7hEY+QXivVOLSSK/m0GOdXgLrWjJcsZzv4DLh7qLuHLntOyHYeqLBJFNYHz+HuzWQxgrqkvB0c0sWzbM/DzVEm8JPFCalnO+P9oSWQF9A0khT3GC76IB6cCeQIZYvuCADIJT7WUqiEPkoZ69DeW83Fp6IkoMOdyQ0HkYucK3WlE1ni/3+FotuREHniieWbP/251MO5poCpWTSGokSFoPPVZmTiUfR+QWM03n/vfLHehilOXHvCx3ESsQmNEwc4SuxPrskuANtSs/LbmzdYUKUIOc+gZzbb4Gz+G/8CBXaDKTGxFTdX7+trrbxvHJjF3NHO/vjovNaZ6FW3yeq+ywjWYvDfVWiFtI0X1fCW5qYo3ojKd6ChgkZ2Fbj+3g8ro0D16SBsZ2CfyfuSEa3ia2CbqZVmEIFZFmPlIGchuhlOOQYy9PAaZCfADm5wq+p8Tdo5jkFQYL8GkGwwl4NH0+DXZLWnxLxNIJ30X5sqByM8boMeSBVY2WgYYUsyzSu2jGTisMFscSZQjGMKqIMniW1cmiYTHY93BqzKuo22kZ52q41nfiuEYJ6lMUEErHqrSHpP/7wO9ICa3pA7WmkIzPEskF7uMIok1Yon5pskmJJTl9lwRXteqB4lu3N8kIqmfzedq0++hXvzHABBtzJzMhY/cY08gGIyOg5qGDCEU7iaGeebjxlOhiC/a10ka2C9P36/ojJHRD3tl4xid2mDUBRLAMYxHVSt/s9p4NRaTLk+kiK7TVvSberFaP5yF6U2vf0Fv0D9io8dAHYJ0zjnD9JhGGN+UFntulhZo4WUnIbCOhB+pYuKQr3Kzn7a4P4U1sd4mZEiQXaKoRnWcKUu7Z5ymADH7oLJrqdn+fXPykFZXs9UgbZHG+NPv0qMVSiwI6QNcJVfnsWfDBt8pKr4UXmW6XrPQD0SJuVGCAGVCwp1fDKU67HDXfqINm/IuqaduYb0h4d7GyXhmycLT2ogJlJYMEIkyA7iUNoFvOTmwtSEpx51atGeRJ2ct7UDNGnnwkEu1IzWyEYaAPpDjIUcJrBRdGeXDvtkmzpka9qj/xLte9kDNfNU/hZhMuB3xucPPqPxdz0nTSpglngKvdA+am2fRH39OpKIt2o5xua6xBlEloDzkrzCd1wGrtkexuko5Ny05YO2Hlk42X9gtGFIR/qPO6Iq9IUMBSD+5FqMFcedZjXooHxcl5J8ap5yqyVUFOWxN2NZAQnupYG0cRUR5BQd/oZF5IZs0oYstnvnODCUnzaUATWeDBP92CriWgasRJElwnAs7LT3gBnynfAnCvg439CiEBx3D33FepgudJhG1tWFeTpzi/uIYyrkDRN3r26frf+67ZavBIeHYfmPtf+A7KIIKuJ2qqHaAceqT9qR6NVmtHWucGP9/7YVlyX2Wl1qO/YhHM/E7R+dVLoSEojOtypNiiyKLfYeijt/GjFL88Wv1QAb/HS4ekpOTI/vMsgQ40TB2POGYOewnv4i7qJaxYEzk+y98eg1Nj64v2FyfXI5gWNDJ1mqG57yLBQ+6nyYlD26qv4b5bHxbeehYc1pIk8VvjvIr2Co0685/DIygFcuGdPCEbnd2slmkJUS6ZveR6tWmYZCtSFdTCCAcplaDa4OuWLKVdNA3UEuN1rLp/+9kl2Y4drnFRno1StljhRbjK08Di1s/vNOV6Ld1MLWkZ+uV3dHEnja6hfI9vOwuGI4P3Iz9W8VZmkmPVUMHEuOjUCZ68IhFmIk05pW3AKGERMHXPfeRw/kO3JAaxb7vJhkC+7P/DlVEnDTzv/KCsEPyeQKMpm0Rv0VzePJ9jLPe65vZTYrvy0vdRjH20CMVTyCZKzyLOye7qvuGy3Z/GrQu1RStXOf8YyK9qCSQ0csIHD6jPCivQDW5t8AG2D03Tlv5852pHnUSwgrj4/Kz4DWCQEZ+isn8Di3Wb3E02mvyrpKkZMttd3xYiSgkP7xHjRMR1LOgU93Ii86FQnhxEvK6gPJjgK33zJgXsagpmLTnnsA4ArVgtUIkqScpjN12qq/07p2LSBt0T9yYqbMDfbRLrmznjkmlS8UFUNTxneC8OPERfBdTxQaLl/AlKXNBJ0sz6sK9pNFm216XekNfoRTSFGV+rnjCv9kaupKoyrU9VnKARBLujSdp1e4ONgbOlartNIq+MpGKf2DhYkxPVIdfDtsn+FrPRQ1R1gYaEPjSCVKsBCrQ5OjCnUSMywSS8hysdQOVlv/MTVrYcl/lQ1kd7N/R0SGv1zRl2/7tfgKHL3U3QhlrpvNaVmexOves+XXWpMCQLhYyyFNztGxE4Mi9H39h3kGpZXaTXxZGP/JjEH7bzvZWp/x8JI2yaNuEe0YZAsmfjSCb5ok2o/F+wRZkj7l7Pf7XdGGsWa5n86vaXjjYRVCaX0OXlm8RsTmYTKtw2GXESBse7FyAUYcV/548rKE299NbAMOrvcjJL/Exn04feZO91gxF5IZ3A6hhUQi3Jv8dQLKkdJj+F9OYg5q4RHYzcclQgk8e60jUq01UtA8Mt+E6G/GAs4nCPaxAu23RDGV7tYWNz0QvI1YP2xbnb2Migi17AMwP7OUTJu2GmGX0qmxMaV/zCO/FFWvmtgDD4lio2/Gxwg8pl2ej2yozM2ALEFJijzIGdFrACTDjPAmBAVbLi3OsoQWy0JbpdJa3f6k16Pi8bC68T74tCJ5Waq55EfHQwWY0qcFVrM24Rq7Oq9ygW31W5oeyzopqbsJ4WQDxuCXPU0s2gTSQuQMEKsHA5bnXhcfN/oJtbfGTofeZHhJbu6tSfFyg8rpn/4SgC4X7DbzHs2+Q3MUJwoSxWdcCN3+w13TFbuZRqRC6WCPbYe5aCtyBYlxBToEF9vswXiQ2aJyJbwWRkOmNWFhDrXTQFREb7UInXaLo8osvF+hfQvy6GqUJHYuK83UG1oRiAZkWyX/x7r8gfkSb46G3KwCdvYs1nj/v4Qvfgyx1EVRYziBmhc7VmP+0Y+4JYFw8So5mqOM3zhnc/n+A9gGyICcYdEJl6lRyt4rAEEwIXRfWWRtNMREeMZwUlx2m+KXL8eRkfglB7aY26WoaVQ0PCJR/yHD+M5s0bvgcuy1TwIdomw2F42+ghNhAzm0MgzPwO5n9etnMkA6/WP8CfKcWbO6vAkrsLCBDMnHPNklN8uZh4Ok4pdWBhnHrweaSDBF2qRVNi7xP+iQ6ioO2JxXruZ+zqfUxdcomlzTM5N2jKYdsEswnUjDhFtiluAnB7+TwoVlJlXbAISXcyw9ZZ3X5GA4FSAIT4D+5Wu/1w9cD/21asUmxIFtCanJqCYz2uSRLDR1zTppEKlaXX713vWZVPSR/63KhYkGU1TeBoBkE2TexPAbmi4sab9ouPDulqLoOekcl1HOgzmDvdG7E/uuemTiHMuxKCXZT1PoYyU+oQv05wbhOkrihii53D/y0wZwQmAejbk3kWZ6vGmO4tpmIYhmuIiendwGKMYKtkUiNes47Dtn0zPzlxiiLtK2JTbHsJ7XpKJ37VUaGyR4d3RkIdOEnaTKQxjRhwulNpIT8VDMecEzIAb8GtxgxQTMh0nSwrBAFSxcvNIIeRAQUZkhbdkQr+CXXwoOlSaYbQ7nsqXKX5G6hy95F00ROlOhd0bhgXmHK0zCT53X1/KhWUEf8+q7mRDqebkJaR0HK7/gdcOWeWFMLn1ukolRpRzwG1dGPQCRdbN1T54BZpg1VmxWYFpideE8c/DQWQBW/ql6VYEBa6cJ57laYydblMJxaS4RoipnQxzUsiW21upBXVZv+t1RJbwIOACjfR77HHiDouFa/q5OuIseSv5BbpYW2ZRkX+QUE7tQYT7c1ipkBdjn9d6nwmtMnSx8RBMyqy/KfLGN5lxkBpnMb97H1izykylOKLiN8WXkGYsZ+h7OvdXNV5aIV9lX0WsPiq/8xBu2PTpq/cRnXUc3IDyPziKfLAoZJh9tTNxTTSpUA8DTt0n5WlJMFfFld/nkOX+fmYrnhxOu9n0+oGJhIfpmErs5nl44+oo3AQiL5kWh9TQdUOfnHv5PEJkq6PgJ7bwlzWbsNZl0SXjeb0Q9KdHl+2siVMTUR2dAzfXfCbmqwePmshEgKhyFvo//pEm9sOvIoL2huOnKkcZDLtk0BhIGqBron9JzpDPKtMx+mTnqWqOjoANhoRUEhr5vREXvoExcYcdZMEegI8f86iwGpNorgZTQx1e6fHYrGq5A044eUjHxzyfP/Tqbn1dbe7666MT+HiEmDDN9qqvncPtE8BTxMQ9Nb+A1pBMGXnTqpI0NJ6hs/KyE5jaMhifL4dyUHZ3+c0MZtf+BpekDNyFhbQ7HVQ3WXyFXQ8gwiiE+rQAhHlMH5TNo/hi/zgsW7Wir1G/CuuJ4oJfM9w6WU4GbDODeDDrc0XrpPiS0OlvbNwW8mQo11ixX+96MrZkRhLgczmepZsci24Y+dxsdv3CjTs/gqCmFEW8T/8FC9sdtzxmNUblXfVhH3LrVLFo3jNlJeVlEd60JjB9bmmsT/Y8a8BIwvM6jrpAJR1jSZWkubviAZ8684q+WoHpIgbayy3/zDBSxvNPdSFXStVlI6rZQ2WGl0Nk4wV48LPDzfnZNROkJsItu8W4n2W3eK98TFBr4FyWj/pGvZ9aFdvmcWgz0FOl7DpPGzUiGoRkmOJ/Ow6fi3miAFWIiEV48E56EI+bXKzKJIOXozYxV3rDa2532dLIpfNSQ+m3d0VrKTjwvTDcRXrhwHYR0flP/yWd7furiABWHXT8J905gTL2j9R9Yw+lcLocEHQDaEDG1TsNEBcJNve6Q9TlinkJZ4hOe87nLkVrZn5hwz1yP8qU/8xi7bguF59OTmoh84g5siUd306/ib5G1AKMHaSnC2jtw+p6nYDoRYCtTbXcz+ZbPUoKbTT/+jhwwLlaol5pJPyvH6hqc7V8K0u0c770SncZHERpkPuKzEBeSCW8lhZtzbCFcc40oM67u1HUHK9w5I7a13h9rozAimIV8rBzIGgrrpYTGW5Urlh8WQnVfqYcj24xMDQ+R2ZcB+tDH9qiNSdVP1l1/4pA1qF75nfztCS936999wld23IUo0TSAq2tfjlL8Rz38wW6GjxjNWvxxjRYz7FuRUz6Ra1V7uaeieqYVZVirqaDKdPpkkDMt0zBXeIPWKKl5dS4Tl/muVY2hjkiO78gWgkV8kBLXFc2Rb3oMDZn2LD/jV7OhA5hByTpbvtr+gz1e0LhADzWlk1W8oqLytRFCq6V5jsDgnN3f/jz2a/0BPNLYHzoqLNrrIQijQer0nZf4PHiymNJf3qPcwj1JwJmWMBARnU0vCURnUSz9rVZZfUgOJe6leUzrcs45VPBHMCgY1HXTh4nBZ1RNmQI9tLq7oZWT/rvKDIeD9Fn25GA7mcAFijRASAj6XruGg5/LtzO0UcgTNjOO7mSGP9/vMe6g5X8bEbXGft3uklYXacgv6HE8tsGRYJNyy+dpIOYgmR3HIB14J7elxIZbTtMivkQ9Bi/vHXkZdzfshHCHR5C5PAqE0jtQ0t7ErsQQ9bOxCsq31cbTbw/oaA0V/ykqMPrBYB7UJFdFt0uMXA9IrY9zPZ/MDpjaSOVAEZtMekC9cH4EneyKCmUaKC+34h2/pxb2eOHWqQ9kJ5X5ESKn5c2biL0CN0x8yKzFDpTGiCan1sUi5l5dNpkvTPCR/UIMqK/YEydXg2cMcEYBU0gYpaU4NIap78XhbZvTp4GA5iSljcmr5XCJAbOqTdeDVasno+OmXzWPsQDLH1ca8h29Y3Wm1v1uDXwIY3zYoogmX2a6KVipaNR0Pb/uxeVV0akL22GM2k91GCWr6RZx/ra1s5GWu3cZKkXdGUbXXlmAk7iOhri0FNzBUD6jUqJvyYTH7kNjoOtEmAF/YWH8ToyyGcs6+VndZSEbI9QhXlbxMfi6J+nVUUpKvOWIatcxoqfIaHBaE+kSmIT7FYStjgysysj1D7RYdzuWOLr1MTfzBFLG5sDAIv/nV3cuLM70nSEjS6P6XRFbVSrD3hs00HmoMwX53r+jJX2TH0sGW0XEuINHDxpl/IVKAarnlkAWMZp6hA+AJvKa8HNlCadMeylVj8cxJvbbxXWVu6eteOlBW+OC/YMxPfZ2MjfvuT3pH6AqN0fHHEuzTitRYmiJV62w6XGC5Wr4KrY1dfAijTiKufJYMY7zmPzk9nkd1BVTt/csteEjFsVjZ5GBOVQGdQPOO5JWHrJ205y+PMrjr17sV+8weTr3OB2jLIi3QTbn2ip5FasVJkrasFq+/NHwiLSVy+TuNnGvcBa09+Njlm048cd3bmGMmo/igFSE2L+uOdzNbbuik1OA2ZtHLjjCG6fYn9HW3uAXD5DDGihZD3H6ysEhaOlw6vcp+shXbBwIgL7+Jj7Nh8C6d24UmB0XZVH6HYcnqJWlkCnDsKBTnU40eRL29UeHJVxXzN3sL7+xrC47Xi6FT1CefS53G6vT0G6MkSpgCzLTUm0EuNaAFwwL0niyJW0rTPhX3K/weIdl8zMuC+1e8Sfxlit4XDDUC2xq+KEdGaxE99qPIe5xA4uwJuoyoLeEv1EMGWQ0mQjJ3OWITGBheuNPEbTG7d8Z7mT4ZGnBceYe4BJQIurValLaNbIzEq4ISlBnwZUXDmYP/jYaZSSUV94ti5xg/gJkBWakvj1XfdyTzkhZXjzu2fPDB6WpBvJ5gnji1Nf8+dRx1T36Zznda7Ie0mV7Xz8iMW/YCULastTboNdTE37lnk+XrtihhGfijcga9I0T780w2bR6k2LHYoKHLFhH1zajkx1sWD+yB4luTzqmfQUFaqycYy4vLYFJqvlFsmsP71S6aRFhVUn2TSTiWQhcfdoZIFeW9A2f8eaaGSjvxtPwmI1Y7xWg2LNMliTl3vtw5PRQrlQ6zM6Uyi7hAvEP1VPSju8z0kqOHoxwz6HtFJTT0RxzYiRg0wS4J5BMuSpj08CYnBYR1xRBdEeiRSNbhqI7n+E86l7w5LdZc1hcxSdC+zpANaNJEcETI161hGjC0hmIg8R1e5G1WLbdDFCrjWnVRlDcMZjlsIs1Xh9PIxuDiytQfCATsKQb22adCszJWZWjnTnD1Rhe/LWlvsjiRHbsu3lc4sIfVW4flYY0AHMa5HzBJ6qISqdAYbDiI2FN9S+n/Df3o4tN/bGCHC+cVSNFfUhpmFeE4lMul0zerUxAQGeKOoPRuJKQKkvn5JPMdPinqRDgTkJZ8MoeX0ixLvMIPEWKDjpem+MAgEqYA3Ojn31vt8PzeMQj9RJWrsYPCirnEt5YHIMr9WCaolLaz0h9uDgcXAmVfPOu+4Oydh7Ya52fILaalW094VEea+sLYEn1xNGXt1PNvv0q7cBi3LdwgRhvrT+/wGgr6Q08kawxbuohUR9Td3hFsHkzoYE+uhX3vECJM6wwmel7YzyMcBUc1jZPaVWE7+/s8Z6vBcNP6ZCMqHSmcZ7owlGJMGpw0zvgVwTILaFFmarLuWc//AlaWwv9GaCXgO5sYzUIUcNZCR7WbdMAJWe1zAH26UTD0WyjsPcV+F6sdCnD6VRRir1RpmqnXaGNjnO3pWPBXyAnNQUF1XCvV7gk5bJ3byHDEr/staNIG//FIMeSu2mfR0ZNN+gW0X/qb22xkvE09JxypWrIVwfGo5HRFIwUAciaMK03wgodlKFhxdxR5UAx2eJyWiFJcJ6vkU70SSIjD64Npjjb8h6n9jiHAyXKKAVQ7Y7NAlWJnjb2xJbDI/eLJ1JcGGEWqWKWYkMSrWe/A3AJeJE4jFcxqh8qMOh/iSdN6MIA45N+IHMoZOvporLeqVAWrRssJmib/bOYGh/l/EfzyYHLfKKSyuPidu1utBskoYZkHv4W3K150Cm/JD2HXbDhNcQUrS272N91TP+iyEQkYyHpf+9BnEsvow+dsmHK9+VABTetHrNUp4qF+VN45vcTAqpNI+Nw5IQq5pBYOCqiQGKNv29xo0tZhdLXuZ6XAj633ir5k5hrj+umG92MDYo4yKJgHnZrBMNby0Crzwf9t3m98zsV+NhUl0U1kJrWGEK60M2Dq1GGDpoF5lIQIvCzmXUqvlbwdVFfD+iJs69QZmf0I/hChokqZUV4VYuKW775Nhg+x6rJlk1RMlQ4p55QLF+LexLBtaUHu8T/7C5fCh5y94iVpgehhlBBWHUsl+3z2fga+b/wRI7rsDJPdwdbzSZJFdQ+SzDgCM2n6fuHOxl88ONSXAT70kb/NkdEZzFkYGMoVNxwUlKVXXZdld6fSYN3MLnhkCs2vcArkPvUZOe9foblUTvRm0ZlJJXPwAKrKPn8mYjxLMZ0ggDRV/xpvFG1WZx9o4SSyI9SWEfcxJu32/CdP7wJ3FahEm4B6DO/v/bofTOnKYqVQGEgjsOv77Nx39MP5iGOhuFILvyZABHp9ZkAU7AI3i9BQWE9ZvTY01vuYXGKjfxc2+w/IXnG0WeSA1QsItH07PNSsTQNeKODhjTu1VTIdmyppGUa8h3cdTci1lIT8RCUWqs64gAYWY2dmApz7ppTWc44rEn9LQYVfJj0XMvN009a6ccF//Ci3dG9O35KvHvFOX60f5TO7OeTQ2yAu+xebzPpf2usbFU/RUSkveirSfsUlY7j6H324iqchFEK0eGnGN4CyOTwBMhxsA/WfsP2gPgh/ZMN+PLNwMSMq4944q47CMxeUZktGHnxrp6UtVNNvnz2pZqWSNmU/QjcGXP17V+mp07o2gMyi8MoYS7i3v3dWZZT9vEtwtJxTtM/1kyXwkvp4cWnpkAyeRuU/BP29xCFhz3WMdQGInnq9K8QndnoNVBsAX/PPGAmOcFNQtJblYH1NdxB5aY1RK0AJNaY//luqlqC4nUVaNGumhH7AhS4M4G9BIy/nn9daXWoFDxWOHIXwkGqO8g6D58LSQj56KwvF6dDbus2BmdCjkDdiJjzRED1RSUZSjv1uYjUr05qFUrbHNwXzkVyiJ3wD7hDoq/T5z5Aklxk6l7hmJMChB5iXYZ15eQBSQZ8B+ynndOT719gSFtP9cqwDk2Mxj8sZHrMpMkOm9dpKQecG9lzXw7iIZYL5u+C22gnKi5tRbwnbYGF62HjjNnM4HVct5cGFqD3pQaaDsoz7T5mt+rggBbygWO2POrur5r8Xiuc11nzdTbt3l+0iMmApCB5xWYae/i1g7DhsLZYUo7pqm2g3XTKhtlUqzTNawAHH3542EE0Bhfkxb7SPGfjs8eHH6bylrtqD3QotvgPxyBPqNlDmikni8A4mD2hUROuQ5yfTygmBVBymjSU+qc5iotxcH2+3Wiq0/1gdXRil+SoG52czvbAYOgcKTPhBCmCi2eEpLdLgrq66pALAmPsMTkM5BdAhtbnsp/9x4qznr5+9LcWDjdCJzZSZ9ZiLdPuFCjEvenfPs2ANZ4kbzXATzKyxYn6GEFspKFv/Ry36yh9VLBPV2MFvNaGSeoMvqvOuSi/Gw2H4AoX8mHUannv6IuRgv6V/DXdGR8ojGZU4psED9QwUhhjZsoz1CFABwDy+8cElsBZCJBc48LtLpYvVg/qq1PiqUfKuk8yAf1jL/im84NnGmTR3jhI0slaA3Ch+JWj9IzAe0e4fX5+n8grENNbcMtvvszccvi/HDAmsL7uJ/on94L/q2dUKJYgSk5n3UX9syGUZsMkZN+iT/r4PgJz35spd+ZYnY1tb1wubm00Hiu62BSaTavkaA0yboJXwB4P3+qQmIXP7iOdYgjFGZz933cbuh+0bPgQWGylVZL+vInWmVxIl1g7E6IVWe1LLhrmVaCBwPiPI5sQt0tPtZqAp1aYUh2fVwuZQhaiybGcBSmpsOgtcd4TIpnsakZ6AkjTSyfAHCfIe0DL1aOfrl0ymHgDcvAlEQXYe5P5RqHXKNbsuQIx7dFCC0UJ1zX2iTJb6thuBaR297yhnO6mCB5lQpDlgU7HxdRNoWsq4MEQCzFSbjwwooAkkCaSJInn0e95zCoGPYhMoRKh5dpu/eRtpEC8CUUJu1GxjYYRHIYv9FKl3Q5IYPLIJuwUjNuDkZqraK3cLOM/X9RfwxDHxvFVXkhXuae7r/gvSPQf3h4PgOdbpPW3rKaEoc/srgWEd2EiacUaqALDdrWj/Ku0YNk9AMwcLB/zOGL1zvER+lCnt3cchuBJa1UhEaULgCwSZGtf7y4TbERel3riBEaa/l+zI8k9XqxGfS/W+eUi32TvPQt25cc7TNFB/j1a503s6Nk5VLQdd6C7LPi3fLhwNYn+t+Ndk2GejO7SAbZKqTMe962g9DtAuNlRtELr8ecV0TnM3NG0VMfgO+zzNg5LhfctDUXc5XxT5jEApvFBFpTUnh61hf6lCm73Fh1joO60cXr3ybrt21UAVJOyzrZGpA1hz58svpGvyt1rNCE/7zpXiVT9JSRb3k3tzWpjbyA6mQismlM1BaV3HLWPudWETWx6EqFYGlhRyqhidEKUnIJw1YjN5BKXAb90+V16gDHul70GELifyght1CCT02s887dlqY4O/CKkXsQEyzusHtdF4CFJdbmrTijoOxSiwP2sG6IbCFNE9qi+L21SQC66AkCh8AUMPwZufCxMxR6cxONDwXcbCrEXP2Ko4m04PDKWQ9lrsxU63yk4P3dVHYWCcg3tkc1fYn3tWxHRfAMGlpzaVupIU4LbZcndcqKQ7E4tgIQEWAYPrlPzqkQMa3BEsP4ukG49i05siWcFbPhYmXEbpTfhpgc2sKu1NEwG2V1d5oEPjtnfoGq2oXDWY7cEfeTepl6LkOyZyDbEVM5n/t7aXKFAfuNNcSaYmJZxMMZ3qgwBlW1pxs/2Svr9wkkNdBWfH2c4ZkVoAHxEml8N6NNUdJ02tKPyM1deInVnu8J0Q5sfFG6UF9aUd9FFp65HyU0c2DBkW/dau8Ll3cvblKz7E1ODr9dBXA8CQdnf8qWwZSJC4GqkeaQSMErOPgJr95Lyf1XK6c3hTLgjKwPNAHF5dtDsKvFXEMZPwaJas5itytJXZR5CklgAAwvZhSJiLon1qtxrAqbwINuak8av4k3f/AmDTiqe3IexdYDlGPx4q6rlaytAEoOB2c4Bue6NPIfVSdmlSB+d2xsA8PyEQmSf4LhT0+Wy50QDC67+5MDRJEM91E8dLIb7hB15iXd4hQFzvBVje03ahcFlxVqPYTwRQGf2p+NBVzgbzjjmPIOdUeoqmJvfq1tle0SU2qpdF3zuv8EIBzjeipm3ApjDXoNlxLFiBm7lCG51TtSDQHg2YHNoLiVN8VGPs+NJrWOkNpE6yxcOSeC7SbqHQd38rzblDFtG+BTqr011y5ynxEJmPLwivwkO9RCT1ReUYMx3EOun2dGlwxdjGOTmfC6M75qJ9W0isVWkI43bCO20eTvsTpPlZ650WgP+v2s8va33ZC+Sli8Ba4VM994EYDBVcdpxBxPCqDch9F9eJD70W15eVhu3eixw4WF7gRCc1tHEm6foIcs/6STXOq/Kgsx+/NGx8E8gjp9UN6Wc7m0q/c9Kw4QKzPTYctM0BRn7pfxGshrpMu9t5rkYEWfoHLyTTnLrXRixig4Ia0yQFrMUvfI9Y6/wUInb/RON47xJtKeW1QY3imWipIIOlqoauJeg0V3dGoV5Jn0gGT0t1Ys6/90VvofCzNjVFddT9HsbOJChtu4mS2qZofdKJI3qZKsapP17lds2izw4DkojQMkVqlxwrge0YTW+wWTUP5QClu99ts1T4cHL7iyMfaa0elCHCD7RuORatoK93zY5Dso6ugG0+IlCYIj8Esrur0WbZ59saYISLWhGvb38VUgTeTJl7EwzhEOxwivozwGcO9hL0iGhUe+RTVDt80I3RmwE5gI/1HRXnuesHYZ2SwydMjEkJp/AyDqduhjTMlxRe7mo7bQR1q7Gbf/6NboWwXwcA+XyCiuBMWHuBlR11vLI3febcWZnMJpbHDQ1+nK3ToywzvoaUY+kS358BzZFGrgzIMeg5mv3FEF/dBeRU7TBK2XlhxO8ISa6bC8ZJigSYPc8UDzrZAbaq6NARLHgIlA0++ERufv5cvTrGlRCyKRDShh3FUzc/uUAxQZB7VkV2coJ+rSJKg2L/vTVmQOdbdjkaN4fHcVIfhOBdF9A1pQ5vAPK2CD2xPmIE50d+gOecpkVT8IBWZb2XV/57BGHWauX6Me+hLBp+sCtGiG4g0oHzYsuvXQbLdaEKA47jFa8Zuwkm7KZZPh0bg5jFMJrdhp3HJF+IF7subxUC4qxk3VmtX2FnATYDlDsu54U+4tc9w/azUBC5xfU4oFhfIW8a04sODFJiCqGHEjNdXnFnnXy2s+XJNIDtfQ1NuD8IAJFvhkRzOWsYptTmLGCUwIHotecw3KbaI+JeK5+SH/N5qkotsFcV61jmt/xtZpE+Dklzd9ZfnT+G/pG2dvHk6eFQGDepEJ3D4HrqeTtCdei7IUc0I0vH7LR/ME+n0S9Ydu4MC9BSxB/IKqIiB0dcLojzKmwhoIGm1i0c+Fb3yG/YD8cBzCwt+dvPDoARPZEW75raTUgNv9zdCITbcDu4SjobQOtgZIVL30QdJ7w0igDHfQFkrMOjoD/zgRejP2DrPm+AqpVgZPV1jHJtywfv9nmU5QTGX5GdohWMZJZpA/s666Co9Mlpuu65BaJxfDFT89+Ojq4bRtp5es0Qdjr67FyH/+BwVXf4HFDWmtg4Kd9LxL69Lkgl1Ul+KIJez3JjRpkcSMv8FRhHSRtO/D4Gv1xJQ2x0I7P5f0LeTdtd5dXW2ujIih0x0y761ayNQguykwA2fZN0uP2c9bOc2KFN0anuar5Ls+YE1QTexHfRLqmDQPLYc80/0SSom1aBpx60b04ObgApwsVpYGfQZ40U9pEpjLkHxRT02TyB/+oC6B1sw2IkUDnfMQY/Y0GUT2iEa+oiIdWvCGGG5KGf0L2UXrcChpU8F70RZEgGU/32lfh25h+1tyDfJSwKiEyW3hn9KKmBu+tEijVNOzU4xodxdJ+FbGIfWCqfVXmh/2tBxc991qfdvn1QySGfmv36Wd+1GYJkVm9j8OsaqtHM+wUYbE9oQPsqHvx0s0mqViuW04R57guWI9ThMk1SqjCEpOcLVZqBU4bffo4+gvHUxB7FHvytxcixoVMA4IoLQID1G3AXiLIOXCCFpASCU0QiZ4quSGzVJDIyJUn9x7fl7NAJd4fBYEL/13k+EToqB/Qgzim4V0VCASqunI9E1sJMkiGh8pNvD7GkrMMDW1K43vKAh+FE4Wmj4Gjl2IEwwACUr+HGpCv2tB/PKASEzLGNJikqkc8xosRpO5b8nJZlR2nwoKuudhDhej6a6CDxXC+DKOCVVoL38lf3Iyaf+FgkgE8vVYrHJzQxR/QMOd4stxE0xxEiRbtS49rZ/mVqj/zI22hn9GkgUIfvjsRJ0+1abWBE4DitNKWXEkwhBMWDqDWk7UrHcl4p48Bqao3QD0N7GxfpQsBUk+QWHy3IECsH53JgJBzfsv+MIXrv7qsTgIL5kUpy2YXaonmi9eP3FvhKc1XdJVD6ABRqqy2BgCcwHplY2HhyilGYiS9cMSC5zeKHJ/v/IbFNXp+6k97gyURk/6PnE49BlQ+LpEJdEgK39sTAfkj3/WGiHhpcOCtV18TiZUd5WfL5ZMMt9S4tbJol/PO9RZSUlzIHW7nDnqtK4RRd4t4Ab+nLsrm/0Eo7MqcYxPRVPMNfYJpFalipLrz69IsGo+dM5M9YJVT1w8omE4GEE4LWpymaAxLoZah+Fjn4gN1r7APNnwKmdTyzmXF8gIt+yfy7U8QuKCJPKkOqsBQr7y5yBQKITohU/UuSmXOvMjswtWh6Tr4klviAOpR2A6HPcLzlnhHagvN2mN2gsmdJqxuBCucTF7e+i5e5zvjB05+lvpa6wLJ+CKhf1rQA/QVxY8YAkJfHJERLym0/Sd7Y6lcgCpGhtxI8bmAkX+ddrL8idrm4z6dVHTsQ0F+IAN72MFS2BAecWz25f5TogBYQZCORR/wKOcd9IKDKAlC5n/8w5uEGZ7hjga7vEJJooBts11y6v3wON+OHIEzBIRwnw7dfhL3pKwyHB6lFomDZN9T7ejNZ5NvofrmKk/NpWdQtNU2X/gJVbH3drO3c+EtVmIRDthnzdm/51bC5lR7r2b7h7yIMuzO3yOVLHiYAQ+s4Elov6lMrVP/Hc85aHFS1MqBKvqrqCPfKuufMVqV7PDieKXEjfeNZVty25xS8ztwFBzoBsxQkVTCe8Q6aNOUIaTv4/Vrp9bwpfhd2M72b5oAFi8d5XQAJak3xb4hFHKCQpXK0rQApIzMkMMdzui/j6aHbCwiagRD9tVonOGH8VxobjC5nU1HFY81+LiVL6SBu6uP4Hubbe8mbfll7ilfw5NpMAe6k307/k998rsNcGI2Gmkw0Q54jp/jriCoFZGEWKZY6+Yo+A/aYutiL1Vt0O/6RkQhmzV0mIlT5GY0oOopufLvyPwCwgCslvb4XRUzRxFswTIXca6MxSUUE9fvgNfzhVYZZ7z7oELUKnByvkjWxxgJmY+SrC9X3qDVsphsh/39lOSHq2u9SY4nzaymGTWV3+KjbfnfafGXdtt5tTMfBfDsYvxtcoHalKvVql4tb6raoBp+TwNwPWhKOESc66M/N0PMulPfw+nXqJML/uWytUUGLshWLFN0RmAVwN1D23Lx/uf58Pk+kUb3kJNJBWJpCRwQyc6s4d13xMZhXtJr6bJgotc6rK6MbVnxNjMJALHH+CpUi/ld2OuwRcnIbphYdEWphAqJfhxMoRywouftCnV/NSBeR5/wAY+JosGIuRtt7Nh/lW3saIt2yF503p67m6uqOC8ygSRfW8lCKfAWXkuAE/t0vcJLHjdBlc4uW7Ie7GrQCkXEuE77O/mCffd8+hUJFNaHPkLy9xj6fCbs2YTYrx5nUaEn/Ru8c4oIyG2VUKHysUQDio+fzLA0ATTxyubQShQJ25j9XzL7+cW1qC8yz1+i32BkohGayFnHYKezfKjF4mCzR4cEKijWZuQU4HhkCAtnduFMHC0CbXFLQOQY6Np3itwt2px7GaiKvW/YZxKymuwQGC5uZlhz0QWKGVd8xB3nujiwuhKnOMxKRz3ItalJTeLZqVrLgVtZ5hqh1sXSVpXZHMaLoh3sx+pd+U1BEHWQPjH9n58s/HyPfmM7i87/r8388NVLH/OaG4MnemObbbeIJzwxMgcvs61wpLxCNjwyaCTaiMOElWvCD9p1uVI6k8QC8HQ1YSKu3ihQ9EdmbkOkQxjsDj1quUgAkrNCLvk/uNI/YQa5e7KXdB3dxiQeRM42OL9X+FMSQIx+rk2b1TY/DiP67Hj18CmgA/bye5qz/+bjog/BJkhTtj/1kPrRekkqnYZ2UzJNTSeydZObGh2U5rpOHaoiJNTe28LDCbUX7TN7etaDYx2TZom6T8EBOF6kz1EvHmihSscCSTbKfUbBd+CqzcXDuEOdh9Rh1T0TjqLLn3R+CJGxB66DYNlYcrLA42Qxz0knWccodPDzEsI/oKF7OqQLWTWlytXCy4Xj7aAEA9bd47VS3WkLu3dp9087CuzzWRrLfELpNOnJdsMym8cgAMar0pogSX80++HMv8YgwNXdtdp6eulZoKR+tZ2MEXTawH4T/eaqO7T2MQzqEPYqrY5/WYJTO1tz8nCu5cjCr1QtD/ma4/F/ZRz/tCagBdI1OlyQxUmDprecJOIcfIC3mltZ02wMNoMDYTAImve8Bqn6M93U5ZOFa08T/CiI2xsKZUGLvcQoiHGR5s01MPXbWWVv3u7zq4Op2yElm74y36CHW6EwvrtDRZ+uBxjbDrD0srqWHioXjbBfrcQEZo8CNvU7AJDx5YAJIcpknnme/744oRBqfz6y6W3bDK0lExMDK03Cuux6kYY3AYGnpBFyeAQCQRZB1oJD/1wYqg43WjNHo3f01r4pXHCW3Q9HxYiKjzOpSrs6jO3OEHmXbZzE4hDAUlyl/8KPjBi6xLbpCk75SmHnCLbHXdTBzb1OFx/IuA/QAqvMDs7Cc27NgB3mjA9/x1NlMMzfLmbtpQSSxjAS8fgl2NbEZt0/t237jJxjfaW2WWJFqd3a7kXjlnjNkGiaXqKi2Qs793EDG5arCzB0K+rATsqpvAPN/PZN+lTZOeFlQG4DCPh8dEVe/NTIWZYLn7nCwpD1luuISb6ss3poBNqrV15QobTR19uieeYd/CFIw/YHZ8rReBh56SwgKJdh/+AbShNM/f5RoRZHmM8MoRg8pCo307Lg00JvXQff58oGchyrAMcwPSxJRTTBGhUq0BUEC9ORUlrY5VQ6rTz8aJZui4dGonFN/Oyr+tJRRs6UHDRAHcSPUNQbpGFC2hTQUsNOssDFfHyO3QQOPzyZhNPTnrw7srFQjzYi0MPPdL5gH/sNK2284NwbB3tC1qFfqNioXYyut+qZICK21iYaXhY1VlIxh7HKqCmJs+7jAcW0xQKLVg7yBzLwl6zLZ4SyR8Byg3IXQZoqWTXZxFtY53hMn3H0EzQ2CZ6yvC9gNdpRMiM5vT36wP0243GW32/0mSekSmPA9l7ZnieRwVEXEzdIsnbwRB7ryQ2r2CkDwEBsYsBJGjA6gvTeBtUc7xNHX0FCSnuJp1anXVXvnsgrqIW1APHTQUjbU3pjVuKB5cbX3Hbj1/tJ1V26H+xtav4eaMKPCgxIN7RjIgdN9ZJZYhYHt15ndpAvi3FNgPSws9s/ZlYbee8K+imYwXHLy1XNUe05c7ymhHH4LmfgwdRc9fyC2NoWqNN8iFWPIRyLYLxo+MAysZvu1gScLyZecyjRROHM7D8LDIvkl8ned/aERYZ+MqnrdosoqTyLnciqqV/EtZyDw3ukbH2IfBre5VwuwsqcwiuGotx7VMI5xY04j5yLhIdWVzFyFt630fo+D7RqPMNeTmZWBZbrgZdAbjfmViFjvx41T4zI7zW7nxpa3i5CpkAIcBDI/GT4V/h8FFwCkOIjnrTnuVfv6YUpKOwYvy5+1FXNdyYqkMYRykcm/wkfdw5IMWheR1895XPbHybk3piyJ/AB1fcZdSCQfVQ87XLqdbvvppJvCWVz2pOourDf+zMpLScjyFf6HsLPBpd0I3DchZTL3FUusIs4i6GKzBfJnv4dKqQTwIi2mQIiJSr6cEsuNE2dVi9f7zdcw2+JXaDKRo1JA3KkqWsEJ07eUmGa/ZpaqA41eVTedSAk3wOr30dSisQoM7MozKpB1B5wwpX/IdSJKcSM3MQ2uHQOWC8vrjBGf5Ey3wnuQeEqaNmH6UfTsy0Jayqsa/JpjhVTFLpl33/OPDIZAJ191AU/LfOIcOg9o7snY4Od4eeRdKyQ6rNipjqR1ZgmqH6hiurOCdakwH5gnUENUHoUVePnKDTufIRq0NCE1Cqaaf6PP2autLvKzqL5byQ9Vftzq8T/jDrQhHf1Xe5+EVK6Q2rrDrbd71B25zV7+WGd/U37huu8qsDXnI+hvp/MTsj3r04mLnwn29j0X53W0sk31IBPq9xZ0cRoAYwa6Dl97RrOj6drfv/yuzRir1NslQpcByokjKvfxMs4f8Yc9pDgOjGEcWApt4brKIX6q9kWlxjCwnVRIoP812JMBhyl8LWPj+fbJWJibP0VqQF+H6TsYqX3vpbUUOnfmbRS2CW4F5p2UWBBj33QELaOnObbK4k5wpwiKtvVwFaRW+Z/6ab+CMCIKlC/j0UFjka6dzhegW4pQEv5FxcxvNUFMv7xHTV9AfXqP9505+pC50HGPixBRBwXpplSTD9Hrg+GZAz0IQWC/85NMNjEKy6euCpEhVO5HvH2ktOgTF0QT4o68aQXTxklXrPDydLCn4zGjwfZUi+t5iSYq6beok87Kaq4OzIs5ucXT0+7AKE7lAtI7Ge6/1avswwuSKTVzCbw2lQ22P63Mm2CBOVLP93ujh6j5JZQY/Wv1njoD7ySKjWKhs5EVXkpDxlaWsUJxnxlGsSuFer+xgQD5a8zRQfoyBfvAwxe4SjEL4Z/To1myPTRbJavsLcF6XDkLlTTN5RieSluuKnYilrvYuKTd55FEqweMCbMg3HIR+Gb+DFvAWJ1LF+5A2dExyx286clBuXNHwn4ydIeezjMX+7DENVkAoeQ8rSYkfmfKuxb1WkgoaMk1ertla+vm+5tMmiB3kAZr/BukUTvMSxLd9+xwKvJKasKuWRvax+4KtZ+W8gUSQ4LoQeMdqi9VstkhNjcbd8Skak5LuAAANaHb3RqAEXepftpR8Lhx+7Vef63fSI+bwPACs7rzWCTY/hPyMQNDqOUNx7yuu4wQs54ss65M+OPRp+kMK05gML6+oId1DiiukejrwLV2jCIM/4ojERrIR5gG+4EHDk4GBJ6bi+kBbzzKsGHUrSaZyo4cP52rliH6yp+/pRo1jeAGplSPgCMayGuWjrslAvvkBXdH2ejgVynL70oIZWnqzwL1uJ2d57JPADqkfbm4sZue7K06evN4cMLdQ8nyr6nboZCmRv1EypVpR/dNvlWfoF9bgkJqpjqu5xwIylj7c+bHeu9+eZ74YufCcNg8S38EkxS3cfeIYgHHpMfYI9Bad7SSxY717tickrqi2bVAIaLfRt+h1nfqU2F0nZWOGJvACutertu96mz1cpUT8axe7mafR9V3kd1RbzHfnLEEMKn54WDbxwGDVUl8whBi+znFDKYTB4bfAzvpxSAVyrmASKPi/295JrU+KDhANTAPGHAA/dbRkfQkyPkZeGZD/cMqoTrihy21iqg48oMMxFn7Zs/uYry8+2p06uNrfk9yJ4xptD5PWxJD9TWqc5bLXcSwJWwvpQMIYTZVzIi16jYsN/UBQ75ayvFTIWhv8Z6WbufXOTU2e6kvzTLbtw6JvKGKTe8vX5Is9EPQ1I3d0YctDKgiDVjNoxHWyGMvZ8PyvG3AHC9ZU+BCzSXDahEx3mxcSXnYlp+UF9pOL7CR8IlsgBK9ZCw92W9g8FYWzwLWCnrwqBZHMDcjP0zBwdBrvmQGxzSLUXjjJ7xqEmXwB2hQnmB7gcDfk3/Gji/JyTXoC/P1rRhuZnatdjDmgSmOf0XwEplTMzyM5iZGmCOub3+DO1awAZXz4UMNuPb7sniLrzXZci012jgRhcLNHxkFjCU60X329QbTIjKw1auaAVYhFYm9xwOcYEpNwSp9dQJDYf3ZI78JE0YaForM2KhDDattDAsjEAB+KbxeZLwOQw6UyhgZ8i53jT7AbcoZAcxfyrioT1ASvwQrsnaUVRknVeBnroq/TGtHdiI9kSgJA5Pv/lykk80DGF9n6qg0ZnE6KyvugbpWaBgq6tTHPzz5+DzXgB/v/8mj1KDuTTjz2I6tH3kWS4CU50mMZ7u33tLHhvoXrNEc1gy7T7aB8pH0gZYnbjCLMHcWkWRJ/wvHgfPy58f/YdhFLI/3isz7DqTsRRV0sAVyH8Es/Qc2bUxaVv5nkKdPDnk/y3+8qdWDKSpNyxoyi5ZC1nkIXVp7CoFcwzvCBDM3/N0W6ynM0p0bUKzGsXJw+Ch4QbASZi1smoxAtB6c4xsaubjKoDBaCGQw9Il6aArLFM/upo3icM26mx8QDvHdViETGB70LaloVQZ9j+DmrQAoBliBIFXzt9LkXMZ0Gdix4l3QYxHJ03iIj+4qECiQ9GYegvNFFe5tX7R9ft0E325SxCds8NeD7WD09K9TV40KU40APCMAGnS0MdQMY7M6uSK1kkngP/kpkBuYmq3cmW1qdjb0sFgDozIib7qalCMngPupRG824MnYOSefOgGYipqt/aHOzkir62BARMvp3KFSREskf/1f2Zg53kWtXSmZRBgqoDKco2slsvVckcUdre8F4BBJ7YaQpQCdbDG9cAfo9+aQQI3kV56Kw4jX/IPiGQAMYKqUB3/M+uUDj5xYa5zB12ITqDqJ6AHGvaKE1cuI2Ab0RCM0NKL50Znd5a04D8srGxBZMggpR8AWdPMO1MroS9l7ETOFKGAB3E1d2Ox6Cih2BpSmfbg8f+XL62lcyJMcs3jAGK7/Py3dw/l251i6cQFBsLg7C2F959acF7NaEUkxHkXQXJqD1+T2R3Md114GNtPPAbblDP2Hizsd0Rpmvnv1jCUQCeja2xGFqVdjWqeIdAawguZvBdr4990719MxTXbcGmw6h0qkB7Hktvu4nQgdjPn87W9VjeflCt0F6wVfDaqFPhtmV5Uge4jebWpYBxRPizQA91H74YUUusUIskeA0ZnP7Y1lWrqPuvg4tTuGvZZMu/OayYH93w9WolFRkdjpo62l2CK3iQgxvWXKgvX8+l79gW+YcJZZDe/uOCRL7pEuB1Y+iZXN2iaT9JgYCNRM87+KRZbLmXpufI1FKZCSxyETdqJkh/HhhHgfU8dMUQkdgVlJfv29Egzjy6rLJ0gZhEg2mJVf8Fz6Brsdj7rYfwYzOu47gEc2sivDTAsy2doV4VSHUo9LHWETN+I4XG6lHyxDVCCbgIjnhsaJqNTsxWC2Syg/cF2Bw0jPkeh2p41S/y5Juk7bZd7tN9qg9xeTuU8SDw6we3+S+4yrwGA2S44jV0PsekfMqRdjtOCbfxshuow7fqEqTIe58heHZOuPkr3vKWHKQ6+qW1cNWRzmxGSQmWkXXe0qOkKbyG+3F011CvUUnc/GZmI/uDpF8oGRnKtJEVav5jnAnG9DBqcve4oskp/G17BhwpFGIrCahYCKNzH2WfrBXY7JixwjQCmMYEzyCVHPU8aPcPCY3fD52CkbO6b9NI95dQRWGm3FEzM9Ek37ClaxImO1R1kH5dpH2ZgJZq7VCU1/1ZVxncm3YoEgboBmSM0CFAfN9gMcEofAoUi+u0c9r4royEw3MUROp4WaVVlQkddrfU2KXwz4wC/09VGPUSM319SSHILWhQSmSif+6Zsp952So02bp+KNvi2QnmmByFnLns5sfjGIOv28TFEP5RLI1pZQgKmPMWWvD0X2T0g3FpPwTHZr5RzP7znjSrtBCIv1SN4XSEmhzA3RXIBl10Y/aQl2DAfKR2LEHVvxIjpLeBMoIcWqTWjJkiBGEPTslh26ENN3NhVwUBhLTtcTWPDrEUM6rh+TXQp2MPrshZH3/qnqcGJccpLTbO32cqEIQfWBNbACpi+i6tpFN9AGRGFcvSydIQc1zJ8Ew1+m8XotSxgB3ALPHBRIUOAWma7y6/0yl/z9PIIjKnnUhO5HNyPJX/TL4G9dWSPRj2Wk2mst/HWcjs/f74qbRQQ2IrNDb8jGz6llS9MrMPIa2RGeZ6N+i6qYEslWRmHGn9lTTwpIZsSR6BIDKTWfjw0GnfQc911qsE76dPYsU/uxhiDP3cEo+2O5C/GmVKRZJQixMYVfRF36Z/DOpfWC3svJc2uNy2d1jT+ezP+4nUpAwEC9OMDUmEsFzh1UoJTxC6Ep/X8GE1fWTdJnBbQLygzc6yO6Zo7IGSnaU5MxHOcT8EyKieX1ddnLBzBs5jLM11t/HD3lmPFglQnC9ELDEoOdxPrXS6QFSG9iYAUNP65FhZDMIjPfDRXsNgILkjrqqud0DNtHSyvS7v3iqDz1hdwGnnaPlssjSpcKkp1dwOVl6vkpLN9VTV38eQL2n+XUEeAQXA7+EVXQTU+wFGR4dYoU90fXU+hk4doxtlS/B3VztHr/UK+EynYvxnI2+vh9iTnbARLNquee5eRosu581VjL2DSyfbHM277EkJweDCxySET/wAzWHcLJhPoeCKrtAJPUYzvuNhjdbY0W0Y5x8dqH5r/ViGmQGS+McDiMPowc++Xto+my4CzAxG7Dnw7/MhV7ZmlIlPPiBEbGmWUkWLMkd19DkvqqidNhxKKS/or4j5Mjn+srAPajBdJa+E+4bpVeB9iJ4c178F71rnx/YEMiOdVp2MEyO9ivA2B5gD9Yy/wcXIlNXQa9Vf/7/YmgY7pE3u95e8pClnzeHMwnTydj1AlpTH/xb+AXCCj7QA+7QnI1iW/GLiJJkCwDsPoNaDlRW3gTLL9eRaSYc5ooTsGYplLx9qJwBHYwFuJvs0b2tujKdKoQJmJuraghgBIN1GzlJiypb8ruK3mXcNBzM8xbYThS3fC0zrhmk3VI0iZgLiidH8A4CfTyPJq8iQMW6czaiNW4KfZpuOJEDuRFYSJbxwF5u46U7f3anRb95SgMxEXfCMoGV3i0ihZSrAO2SwcHnwCtlaurzM4MvoknmeN/9mHJdj8cjAL4V7qDIOXtuUBkNSGYiW3ZPRje23IPp43J9IShM+LEDVbtzlDeiSbSJ3Xk1pfdugTGLXWCFHsy8OLs/QNtshBTTZnr65tyM6EvHOqaxENOYr+GXHuSAGvJ04zI0XZxJv1ec8detUMgCOYOwAUk1aFMho2E5fKYxGAPF0ernyEUKP+TDZMyhegjAAndoKJUwqn25hJ181uNiBOb6xtVd2mr4HHeiKplb2RW+OlG/cVDuCfGa7BcAXqlNSCanAQ2LgBZyqtgwTIa01aWRNabKfenCmOxsCUJ2Jr3+prM8Q7lcWKTeuCcc14AeGugWB003UtD0Yew6lxetLppoVLclV85lfTbG6S+X5athrliQEF69DfOE7O1e1gNDOG44PPtbqCmjs3IbFy15+JYKqCeqxDmGTBxwcq8bqHHjfUD9k4PuNLFONo9hNAKcm0A83Pcg9oZT15GOFuefdXZDmwqxpfwnDsg291AsYI/ecEgZC/tMl2w+nZDHbTGuHUC7ba96F9XqmiGV6eH3poigCqGEAjywYbtzH6m7hKvIa8cZVAoDp2X2sSgWM2I1pbA24p3LyJTLUK+NXRtNL8YLRoA3w3AJfIvBlypYv3IEisqsdJFjile6VnzL9VZxpJGDHHLO+WAwAzv7NvbDI5lIis/6uOhADb9++2jZD6c+Z1UKI0l6utwJFlApV9biICAQykRPqkE7P7ZLF7893fA1OIeOToBisSYmcU0ZN+oEaYCMZNox1DUFgC5kgRToAzz7FLi8i0suu4RyeHyFfPUAeEaHyjKk4efLwQhwIAmx+bbxBAffwUPEbjiR0gaox4FnBZieqdiWfSyRl9BB4rdxmcncxHGUFVVsyLyC1GUQL/8TJg5t73KzQtDihzPozVk+gF1F5dAv/UXoNk4CShxos9oTrpb9jRONlJSVU+k150rVjFtrO8oy2U7NP1J92XSxw6IMHoxh8sTOLpBe5x9MPHp1fMHaJc+vn/qsTWZBV+5EeYpBqB1HOIriSkUoMrQs6tYKYMXrB+pGW3IbTQmL2f+6d+t13ZuRU4RI5pydbWiqWxYEsRhiYgavGW1CMWbAgFZ/AtqyvcZDxZReOC3QnI9YSu22CzbfTMj+MMLtvVgRbxJ/hv+3JzSiwG7X/rjEvWDrT+uN9AIlr84Ycoj33CQSe5CcI5Xt+02c/+syAyN0BLz79GauvEVeyTWzW13RNhJXyBUlp/ccdvI3BZQ8u71lcngAxnlX+KIHkPVqi7YQlvTqI+1UKS9MW+9hEcnjj1J7lWXs05pYiGFwTpsXLvaK1pr5DGP4uJ5gYQj5pRSczAF8OdElXj+Q0Gt7n3BdhIwYcDuTT2Go4t7TZQoFMyXtVLEV6AdA+kzFPNOhZiCBwXbPOmu6rsuJzxRS0swrrRpWm8EDxtBwIrTpQivyty6BTuA4PWXALaxRJEv1YlFmFA4dDwXO3wcFqvSI/ejVH7qMdPH8UlP8NZs7ceXiq88e8ziYSIjs9Ua/dAa4NTefkwaxSEcIPwjmwnT1xsEE4zgfGEvJNz7S9AyURYWHkfVtDJfYWBGQ/NwxqbWYq8VQDGrR71YIJD2FZjSsp/pKQT55XHhqM/j5m7adwcgprQpv/oMOCS23+pkLYBgpF+nOFY1F4Rdl8tSwuFxL3d7vs53tMH8doVUYLe2G25tCua1XV4FqJfoej3inhvQ1jWrhKD9mMpku2CQtlDInlPwlkppRFIiGxXLI4B2MwoxswnrIcAEL5wQPU7E83YXFmddmFD5inXv6jPI1m4eupZ4sI2yaMlk0LtrJm9yVhFe48jarHmHny2cBtYWEkXk/WHYVPtcMJT4QaKTgg1aI2VFgXtfpXDuITYdPcobDCp6tizefQvaOuuVNi4Tnl2VTEgs1deoarrv49BfsLzG4iSv6TN4Y15NsdSS/3AZo2uxhkXyDROaUg6973qSwSHvPjEqD622agaQ5gTTVTTr3xnTtPG7f1WHbGiREPn4AqHyXVBWqRSEY+Mm2OAkU/5bKsnazCCBdaylpyZ78tLlqLkT8nea0DB/WSdljxeQl9l0TRVXzdXAnkDBBtk/HnjLjYBfzjBbxHD6IaIqVCdyujGwuQmzqxlj4f80U5o0QHHnBrlMTEjlODIGeaI5u6VH3RqHA21qywN4IW0x5+KK1joUUMMxhsSwFwXCL5K3xIssc7747kKcwAw9nMccmRAi27M1OQAbmpZEiNVi0Oy0DWra+3LIKqK9DAgUU3UpEQlnY6fCUyxVmFxVQb+9VCC7ldrUlNxkCEHrIYvnipq5zFPIcYm/TeJahbiDiXcjIAXoYFtn61v13lxKtD/R+GQ/5XgflEwflp5sIV9CCxPrwrZgyA4LOQqJW0GOsAoCKkF0M0tAQQltym44PRnS18QLToMzHx8tZerv/Bh0gI48ZXSREQdyFP9EN/j337B4i7x4EHlGxRN90U0kWYZdtB6qAzuSEJoWHW/BVUhfLkIQv4opNGB83EVEIrNsf/MZ0k/CgG2knOs/8sd7SLDX4C6DCGqm1cELXFrwkWCGm8rgmyj8yeirEmcbNBJM8//lsYNlcTkPIDwbNCkrGh/kVC2v6Q8o1EQFqwoLl8w/SIl4RG4U88C+57lKNtm9BCaEFPAD5FrzatyqUyCo8CB9sTZP3mUan5/YdmwVs3mP5b/3bKbcfF0ancUldP8/HR8FYG26PX3md0TIkXJUcak1wbNDWj0vPW8DH8VneegD4kBMcBnF40tfIEddVNcqtPYlKiVKpBq2KhVgu6rStpSnO1hoCV33L/VNdufpKnK/DHKq9IygkYv7XaqQyKRgwOWDJKeAtPeBg0OkbsYc0mu31+9ny2jZW6xoycYMA2/RD1G4PpW6rNRYRkik5ELiV9eCQn0XWuf8FpPIZesYqOOsu3GbcpJEWGpVQLN2FnSgPckeaQ3I0XIBJkqN883jsJV7XIXaomFURUeuCK88G+GGZOERjryro5/nRsFM99BnDOzg0eKI7jfGlaru8XpjAoqp73MIiDtREW0MNsfFpqjO4fZwoQjV/zEZ+/k+X9DO1qe/upnUq0rI6U2HF1FCAMDIVipCHYZH9i9WCkKseZctxjwXMosZRopEek23EktrXFxkMdg4ky62nWiMegKGLVR+wJ9OJTldU8TT7PP/rPaFwDMzwU4zwPsB2ZPkNxqx0WhH6Fk763RhiFRiXITsUzZSTwVwG7INm7mgftjIhs2UvYLA74b8vuuu7imJfk2siFmZFUCmybV2LB8IkoUASz14SBj5JVMmsiEIoNwISlnjWCPOH1u/cRIsIdtykcnJBwHE5gvS0ltTABvIrvZBlAUboyh0ENg9Luuw/iPv2pMkWG3o/9i7rb5PZA+laSWU9XtQfiXQW24k6bVfLM8rWpwjyK6CxdU3J7EkDBej4cKDAubOtBFvZE77ERDhVlDVBQi0qGyCtIVYFHZ9BkWQGXAXT9wU5DezuhVbDkVCEhisedGpKABS4zSDloVsLjK+yEfkKOMIWux7Imn68V/6/h3sSZpobVRsbmPNnfwT2PjBDekcIMTLLpTnrtAapYRdYvwD4/9FSbVQnwmXYr0MTI+B3vns5JpjMcO3ikrlAnxmlNrWEnJUHXs7aQV4frlqAlMYMwzxGpJFOCmEd1StoSbHl+eHOpMBOOWtl6MdUSwQ/4vpQGK/l/TzWo2jE/vN/al9NEKA2rsPLmAPWBWkjeSTvto5BMG2JF9NbLc1mJ+C+7XuZu5JEVeLs2tttZtXRaPAme/5GrT6qLnK1z75hZaurc5kMj9LwFsAMyjtSbMkcOOXtFIhqFp1y8cru1kwtZIxptbbr8wL0tz0Mo11TkzAF/PKkAEaYXcAtUsnjNdKjXrq0gpIizIN5J4y0CedTPORf8ROvdjeuutla/61fq7EJDGThwfF8musuv17PmRDfFjO3D7HSr2jp6egrnQYxQXhTZnDcMSZFxZiYcEUX8nIoFJQpg3BF5n+taALAGDuoktdEuP/C+s2MVg2r0hgwFe4pSoScgJCynCHJw3ulaXfoUkeR0isrJX4BNhgvWD5mx4N9j+gBDgrRjdmWMODOp6suaX9vGiKqIpBNI1Y3krm0B1jbzd9sa0BFtqWLpesBxWIEAanlaPLBX+6dWBm5EyTosAmdJ3lQ9Cz+eGr3zMIKOb3ttD+8PP86YBAwOKOBRMfOrRJJMkCSVD5nvA1k7ZIxkqGRBl3a+oQyOfpKKoNMNznPejAOUX0F6PK+EQCY5AyKLpBVvQ/jbDWArhNDIpt6Gx7zu9x9EVhhiE9evMEsIvJ2nRTN4Q6xtFze47j9czk0BaW4kDbBxpkMaQM9GyM/NORVwygil0nRdjKKn7JrL5+e5qTkGkBRq8Pv0ieOIMGRXwXicIKft2lEIvs1XIX4OjsrlVr1/FeCuD1gzIGLIuf/PDG3mp71HUoAYfsvR5c7jHq3P89l3Kog2Guc2z/lWrz8Tbou3UPpMqXHKss4tR7djCAujyAZWaOWqMUtMe+wI4u5PfIS7aIfV7JFngUNSBeaRDx9Bb32aM+n0QxaYUzCR6PtF3jATC4z+MlGarp2knDRhroj315QMQ7vVUtUrWb6FTzvP6iomoJFC2k9m92N1KFe2VKQyC2ymgQmPmsYlYeiJxmFNWWWHSNAAg8UwpBfDDrTrlXrLRLKQeRM9EmuxL3IOU6eXRLj/kNDSLbbYtlW16WiI70PY8cBEFJbyNYAcuRwiyRD1YvIQtA8hLHKKRXuMfUrO3QB84Bf8R74XY7o3GsZzxYsMV+6lLgnYx116GYyIpY4/5y5SWFkIxqWbxb0aSvvOVzTxbbdrrDV/7ZTHhyZNjyvxOoKsJIUdYYxVU0Tlt7N2p+yj4Xd2o9MmQnP3hmOKHMnXUp/m/dv6Kx6NnguCfj7odmmDcNWBOaEe8yDWjbTHrLkymXxKxI3lqBiyiEKqN5Vi+dWGnpZ0QrxqNI/Ci4ATtMWeXnMv1h8XcMWmdeCeeHZFFg/XkhQb7AE8ssKb+Xpm8o/1og0E2hQ/uzjjoGOBTCjUL67DecVaY1TLVH/MgKFZeQai5kop6j0DG233JdBO1UjP/eWLuOifAW+7vcMhyKghFk9uPeaJxkwEwbv7kCC3/bQOHOMYPkDMCOM2/f1XMlTB8IPJemgol27puS4hysAlUB87wor/FQigx0UWWpknzchvf+D+PblUlosHZsCoI1//KdEyW6zyqEgeXupsmfeDnulUuX8xTEtRnPsd80j1GGucUj3JFXv2iIyCVFIj0MNdZs/kDdxkThZp5NuBT96ORYe1WtcRXb4gAbWiF4LEXjmMDn8S06ikcgjlmcc8XkZoCZfCu3583lulkSWKPIUTF1LDQdVfWJMYwKzQLRLhOw299Y+ZINTq1zIYUwNULJQeFQ63X6WXjYvEPU8nCSqzLfMcM8MNgygpWMX9ICRCKdJrV7RW9pOemkyq8teItK4OF1nYtVZQt6YPvZ4OpJGZ6NSkqVfBm0whUAQEfqjXGUN90akhetcEkmiztFSXxobNv7zpJR0eQmAS/v9gXk/gs+byxQFMZeqKT/LsTNnzc7NP+2fqpksAPiLMOR9lXU6vJfsQbz4vcNtSnlY9UluebuVajibIh2kXZ2ujXnpGtv8bj/3EjZnxI1m0GA7KOc9ExDop8Y+lCH9/3G9Ey/pb/C75I3MDKxPEA0zu71za0HVikQPAYlivpCysbfYiSmukZh73YSELYP/Gewy787UTYCWZStLdcYgyIos5ujNxO3Fj3kpSzw63WtoViiKMIMiwb9JxMxConZWNA800Dh9vi8MOIUOvfMJ4HfH/2aZjsPAxJzlV8Wo29y3d2nKaRxouL+JOCK2Nl+9j1wQnAwyZQRmx4uUGfp7TGy6x+11jKjn8wz1Kah5Zo/cQ83Xo+WsakQ4L2ROVSvgnAPY/Ub9KEBvrKFn1W+xKRwLXjhAWEkKxr46Yow3cFt2e1enwjQ/8UMgflalqmbPmlhRpDwfXpD9dWDQy9gPGCEzto32P/Q5cGiE+1awjycymXTcQR/fHavhH3BNR0v8ajQ386B2jCBadfMqiBRDD8NjoztdsboQ+no/kOAScSpHIMr0TE0LWGz8qdMs3bipEcpR5suzAK7ZEKR/Aizf22juBImXFABYWZ6jZn0KkGwjXJ1XoEDUuKorfguGo2ZiNXOtPQajhBdLtDlUtr97yGMGqcj0U49WAButZVmdjtGGn/+ut1OERkJzCpyEAbWWqSUcf8oXQ514wQGELvY+lU8ElLLeQfYeIg//R57x67jtpw9CnoL+3k0DWywUJaNEO9hEQO7AT9/4QXtVkx+cC7a6Scwa2JTFJPoivvb47BKxcXhvybzof/9UsxgQkIEdPMReENqAM+lB/HIjeJeE7RoqgmEPbn3HTcPIA/rUilsITDlRAD64kfRUcv39PvoyPtItTO31EmqUw6XTn9kxqp1JhegL7nj0GmqXLHtE2H7CZQM0iLVT1NT8kPs1GdqC+J04xWqYs/a8zNndI/+iusMLjPVcQasu8bKs3HMdWJnAApvzsA7b20r7rEYNIJaZRW1WgglNs7+0Opqz3cOYOyAfpiHC617MQ6IkImfycNYR3aKWAJ2/ilZOOgaiRQQuxR2EKYy3ezUqustxr1cMX9IXEJ5kvJn04h5cOE+pdxNWB310stTYPBKzBDq/VG6mWrcFobfnn/tKwxwOLyynFSLRirIikp55D7Ngged2lU+15NzrHMoN8veWFGZyiYF9GShXPEYes0PT4dcij3Dn1POdeWe0PS9ahHVGAKC9NGCRZVE/+1sfuHcN7jY6dAtvilinMu/WYu3mT+B5+A7WYWz0ljmSloiflyKiGnt8XU8eY7jhwhv+qoSYbMf7UxIflNapKj7U5/oOP9Z66A4vxtsSO7uMblbFPOb4rf21OFoxnEMLX15aXFi5DABPkHbILkieGT/nL0THMD8ang7oFdUakrFc9SV+tSGII4YViCkvEgQ8CofckqN7mjah1XEZhk/B57hU+gcxtub+L+3nE5giTBlsrvyOa+e4rXiof7UJhnVO0zL6EnN5wkRZunzC8L3QlI8CsDaoY/eTRlft9ozU2epIedmIBDG3BWRii6xNC4p4AWwB+CBEzNz35eda2Vw3v13+aDqHQtUeZgCDwl61clZx69+UqWmcq33+xuPWWshzUXsDEFNSXZRjC8Ea50dpt6KtPD30w3hbXQ3iVO6ll1WU556wkE574k4rzomQbkMPkA244PWKl9MDChPVaKfL7drWAaEgCOrFFqfFbULZcf+n0Hrk9CajORw1uN0suHdGQubfVCq2rBPYTqQEywVju80SVtrHQgvMwqFnFoRq8HMx9Gj4NYz7QQkUCF75XGcS/+GcS4WAAkZTcxQAxa+hXr3PqEI8bjIWZC+3HwZzbYMr2o2c/KHVmGM2CL5AihMTmwflYUczvaXrddqYZlxCbggH19wEhAnFBIZSq1lz9A7ESu+vuy5utnz9Xr2bzhATbGtIridHPhPzP8UKhe1YLa+AWjoSHOhq+d0fAg0SkFxQLCE9rREwAStjlqnbESIeffbnH81Swrlw2RxUVwPFrfO+xoup+0/1HugHen9d/oCzaeTz9sPhqQOIB9tA8ZKeL6KpuAZWFTSz6AAKAOwBuJs90EVyb8pNRjqJnuItVpgTRXgnHgTCZulU77JO/SDWmphYtse87ATn2wrRiys6z0zAQ66iR9TaSGjvgPJEmAjevfAcR5iuJWgY/2mMXNnCvaMXNTkEzhS47sjO8WKg44NIj5bgh8b7fIdUTerzBOwCwAy+Hg8CEXVPQRs/AJV6J4Bw0qGe4bmKLCNfH8h13ZgjHvmufZ/qJg1yYkAcCOteeTXg1JGqIjuYOQ3xlSeXbQgUlW+0sdGM6WOO+4ARi/lAVFfFeCDp8uB3BUV6Pz/ID/0/rn0UBKXJPIChPmh/Y2Z4SpYBISlWvps2bPTSN/SODn0VPKOjmrFMubFEe4ewcwRvg5hqpSA0gr/di5CHsW4+ZV0IwdL912K/l7d1KZZ4AT5/dstsEEyuZePXZJQ4ftZH0wqsw3JDhbDHkmY97pA2cSdJbuuPvypNGruRJfJwyodmkqZP45YImYhSe5RYn+KpbyRwcqT0U7PUcd1w8Mxso+KoMjQDIIbmuhDfNolx+P6ivO532R2uGBSKniYpLetFUBNcJTCHIrYxS4ET7cxjLVLVyF3IOiPUxQ7uVxM++IUi9DfCvaMW0crsVCSQho9TSv731wuAP9JAipS1zWbYUDwy/w3rMstbuJ45hn8fmIXXgTovAYcy74pswTrGScLNO8BV3dR4VkIZGkmn9Hu9lPcLoDEEAeEPjcGyGHp0F4DqHa69kO0Um2udp5b4BpP99plDpT1r+YmetrxJnvlxG3blvlImD42SU9GG0bX9tGSdI2KdDzc0/gccVhGBMFKYsLJMyaC47reGIKhSMOGWkcrmYaMT5kKo2pns03ZHOATxW0aXjnMvv52wKCW/9zvx9WuPYWMmAOcvmZecIjOZoqcAuiEsOEgBTmatb96AkACW263a4k5j18avMV4FRD1IsD+RkR5Gu+fuv1g50F/sE/SaO/a0PIMfHJEITleR1p6K1jdeyyw/vhaN948tjzTW6JtTTrsGwr2lJjM9+90YDziSN9AI1OPYxG4DXcoypbmoQ5pGeF7Ti02twEndxgr58UMmCp6GklHwqO72TsXHtqH9JFsalxNsk3HyU6Kp7JoMseNB9rkXC8VkNQ3uSJZ62xaONzVLPANNAk6UIkBK0KgksVPLZQdsQjSkR4G41SkCLai8bdR4zCF2/kTEJxC+jNjNDelYKexpp1k7Mv8rUhLoz5aeB149cM8FfiAgyPMcY7i9eIENjYVCTysFVULRgzJhlcTvFLdiudJeaKn374u5myRfplXR3P8Vj2Rs7hMfP/C87D7JFitXo/im6wWCeTiVfgk6pofIqhHrpOYDbrIHGm8dqsu0gMbI2L4ga1S2OfmQTUOeXeqLz2uE4bk8tVUH8x/M6Gm3+urqP99ThOng6THc51KIP6taesLQ4pwjC6wgyl1ZmpfWiFj7u6WV8GCfU+oNRYJfvlGbThaCQRtq5teQvyoSKI6ShB9J/6YNqciPQwMv07AiramHs6uZ+tA3yl5v+eoY1LzULOAOWXQ0ScayrMMCVL1y0whgttW/x+hvSyvnxo/7tVH/PmRGrZUfhylcrjI/zz6H5ecnFkbi9zLwuIBIl6w/z7R+0q4OER8u6PSeiF6Gyuy4rGGbWAayTjOvW9Ea1k1FUCOCihNL3cecHPkTzWipxMZZ0s0lbv9jU9vBD3srzcOkNdZA4rPWSol+llYpu4gYo2ABXI3OKhKcsmyx4u2l5K9oR36qexLc/2dzpVHlZEmb15DGJL93zPjd5NZTdQYN/tgP/leZxun03mYcbhBdTMAImLCywyxWVH65XthWr6j2R+wdVbOcX5Pf8POIHiGZfsvLXwI62ZKqENzyEGpTUTtREpob4SWx1EUD2k3D/w85VuL+W/XrKgBksGSJu4OJBOzDZE5nBI2kt6nP7IuR/AewEqhBFQUTknTfGNvAsdBpN+YBqFM2+mFWUC1+Ffk0tG20EzL8XKAxy4FctDLe6M7BZOSjoCvswEQ0pCaVzWAQrcufUodjwnvX8c/LMUIcqN3VP6k6ltp33lP+RwSGH+g+HHZuL3gaIb+ddtGBjSTYBqUg2GqQYQZrTI7eYDmKRnNxEYJZimAtQE0n0x1UhLy2T07EII2VAVQrd2vAFtWtP+KfiwA0QBDOKE5O5obEHAXLHsN63xQSQHnRJ8mOsFE/WJpiz3+FH3S
`pragma protect end_data_block
`pragma protect digest_block
7fb315fb680fbf39d2011d73d96b48c672cace7f964e597db805d65b23209aa2
`pragma protect end_digest_block
`pragma protect end_protected
