`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
u6Qo1O81yw0UtaQ7kD1dr16rJp0QuCtdMB8QE/g3sOnV+8xf7+/LP+5axFpBWslOi+mE5a3RhYypvw3JcxdenI0WIEKhJUJ4a6mUaPVspXh3BX4e+JmQuWmIsqjc+2PbFd9rBphdtJXeCQUuKLlWyw1Qr3Tz01QRl0nTrS61Ed61VTyGEhfbfGkSPYltwEmRKPcF91gjWbnY4nNZyH5XObjMcLmHywG3XVUsDglHkj3mYjJnYjT4LEkdl8D58w9Y1ZvV55V0nwjTGot3QSEbURHv0b0RVsOCCRQvOuyNSnPZhH5T9hHVuMmjhufk0S4iNkJGjfxLgVz58Zq2osdqfba1HCZ+d1euIe41huUXlNLZAhPJxlP4/rlNSir6Vli7BuCKy+rhT5H0VzhVvfeYrSIqO9iO23C57FB92vLhcWOfZyCeEP7qYJgrj8Y7bz+qPNgCl2Ug031yfP4EwsglnsGNMl3DgyxXgRV9yR7lolAEOMg0ozG9dMYgodEn+CJalt0NaCpBgzMr4C8hWAzl16IhlJnRglermZOIfVrMwddWGH+xGZIjtEgYPoDmBIu0BS+Rm9rUGZ2UCyYKagRyT74Cglh2FwVv+uVVfmoqcGu7J3JSzTdsu7SeMtmKJvD/smIb19EUob5Vx5RTMIQGNlEUVOmqa7UWtfPNBtMqkQFvkQfsK+3nI3NwHcZXcLcFF24/qbLNzAvAVVS8K8IaFa4tT62+7lq19AVBybtDRNntUay/jnoGkMIHzTx9kAkU4PLnIulupBzmqo4kqFu7D23qvCwttzYxN7p+S6d+YR1IanxCkvNIS0CQfBq8ineKFmp1wTn20jdQ/FvauUg8yORvps8kaor0RZ2eqLikFGfOixVlvxg2AHxQ0IAgtBkzXlul03MLhlg4SuCiYMAiNd6bu17L/Vc/WR1CqJMOsnVBvBIsL3MiBzDxeexX3RSJKeE+/EBbE2WC+8RiM/+0vaTnyEU7BT79HMHR3pCrGZipY2Py/Yv9l503fsisNY+Vye0zgqmjb2QxEjtHh6WDfrrbzFiHHhV0IqfV6mz3aE3w1JqRZENCKC2XcpvLdsi6dxc+knDd/nfrL5SPqD2s0FhHWXlzVdIImiAQoloZXYQjqC5xKjkvaVo1yuX2EB7xhdAJBjchi86nGNJmaq29Xx5xeX91r7Gxby/px4B4k+8wTmrZPKx5rxlm5AZW9Qd7jyNI4tF9+3MHlYjHJC+189mcrmuFWrjBf/QMVbEnGNx0kzvfX/psnR15MeSl0D0nrLuy477lpivwjflv1mTH73eLFjYIMBgtHD2p68zAH/PLOrMKFy+vUBp/oWr3546a3A61NRRSGs+So0Tg+A1YZ5FFH4bFvBXXdVjMNuZ5FdXVeXQkfuIwDmEyhu6HXfd/jScAP9fjln9MZCNHrxdbh/TtTqW409GBeGXqcx/7p2DQCNPfCLu2H/PcuSmGiPRg73G/IXkymOjqhi2VuPcvSm8ooXziQR7NNwIyGQjkYxGXSkpTECVJs1VrOWppArztpr8J5iB8j+dDx49A6hfFmBb2tLsV83ViXslJrQ8MOpza6ttwMjfBMWGvD0K6BQ0batSiKjfBESa7GvemKjC72O93o0SmlVEhwCm+poKHBec/Q3LggMNFSgPLFyzKBh6ucbC5zVFkFoCEdaLzkZenvRyrnEvswJO+zXCelMQiqW75NjLk6wM2uVXIie/A6a4LULfQILRNWVtNKgoW6nFsKUlkjkmxPHPF563+W3Ma3fXj51OEMDKHJXXlxjCMdSIYG/noxJ1vJ2HfZszCtPUMiebhFsPnxomv7fQJFljcB5SKJ1s1tszCDdJIIobUwefrigDMOPRH9n915lBET4ialYVDcr8zDtVDjCBgwOqZKCJMdFgB1vy01uixIa/AU6BxkcpFGhrtcmeDxan4KML1NJYQd7BAla9Q2Dag6LCrt8HzAt8IGkG0HAlJzQF7u0BGHo48lIV3HHKiHfkpocx/t5dJUcefNEjTuTLj5l7XF0WqlKC3+Mi/ZxGTLu5jsfx9ozZT5PuOTinyG83a1SdPfu3MQ64Ihnee9qMbMdYw1yU5uVffUA3Vy7hBn8xSDObl2l24bVfcgRr98NHKQs07aMJDrXNij2ByYgo/XYamFzQsCn2v6MG48BJLagdVtCfeNZD7/SPGwJfyxbxwTwF9+43Rtfwz9vWQLXPzGtI67tmM/AbO0oKiQIn4tyIHIFp1dVBcqNZlL8sKDR9FvK+qDgpolgeSWKAxFWopCcxOOyCNI4L2HhfFaoRWjIF/QgiUWyqFvk0FHWlxSRJ0G3Pmu7P5DP2fR67ZNcc+WE/Rjlj+jwgCJc8N64abxFf0swNZUihSDlNr/xInfB8bW767M037zefzNwIvL+12jz576A7DpNGff6lV50Jic4dcaUBQ11kAyiLUpeDaTUb6C5JMffW6wxBx2taGNrjTDl8khrPH0nYyhYdXketNDEhIwteAPIknT166f0jFkMtZ164Kp4IgtT61BHC8xxkSq5T0KRBYbRfPy653Nj/xKoHS5dtVg6tW4HfeyGEdGuZ+sw3PQRzBks0XZDxxo8qbG8rcgTJZv3rVtBV7CDkJw5UyNEyCb8m5rtJtHRPD7RchTJ6NBQ0OBQ7lsEAC4aUi8b8Zuvi3Zj5ZLPA77VgK0sNlqfO6sRfno90wxG6iPblZ8W5KFonPHGWAvfH1zk7dSiJtykmzIncNubKYbSXr4Vw7biazK4z21m/VXhYd6yYKvhNXj6jnUzSmPSurfnQFXnynieyyeTZBQU4qQ6GGiF8SYZ3F0f3n7VJzWm6QR4NFUW9Ne1TF+IAsfKDqUeRVqrVwedZssZ1xNdEPYqMxR8yfYaPMfKZKvO0K5/M8pPcI17rl/gJTh2NnJAea1PY4pPinEqCZRsJuWygn4mLx1kZnnS1xCh+6LyZfAhf5kkPF6TvKObBZKpwBg4RkbBMgoFcEWqiGsAXll9IZJmsr0niCR9wdxmf9+JvDtORYbkLZLr0pXh1IBIYiEaWHoB8MMF1iirt31zdQK9x0G21H4fTm+e88G4IuS+KaHswedznbGvXvNqQFhOY2GsFIX9dy1XaAlHVCoyqmNtJSBjWmjpGzWoNJTJ+iLzsdu0+bEyNp0SyrZYCiNzcLSf6eLTxNB+k8bBA2On79A8ZxhP7yzldZZ+TvQBkj2KXSsLxLLISZ3X3QgDbO/OVitO+wV/fEWGeTa17lh1CU9jqZjH1jwCWllCRexCViiHV2cW8LyRLwUCpzd3EhtiVLr/PhrANttLlNKI8LccWQqt3YBlm4eVxUOm3+uA+zSQpxnbD0d9yuW2jDNNtpXqxJmwbr/rHbt2CMuQlS/isdsaVLAt1WHc6ETVw33ykYvQmFnG+pao7m0QB1wGz/7z0TsCQe/4nFyhJGLY6Yx2XKoP+OwpygufWoyHfr5S0EWB13N0/ux7yH8ROQYblPiJpI5Q2/r1NGNcYya0ix76Q3fmAGAkJVBIHIqSzQc8CfMRg8plZWQQ4Knfne9biPkYtrQQ/m42tC/Vq2woFGGE7d4a6iLLf31HGKwLT56RsHECIdkrp058/PYC1vkCHQbMLzIMHU1oP385od6gyUuF4jrhfFtGab8yGUMViCokTT0mb0HStqF+KSEfM6RRqgNEv0MAbNyWoFUjjQrZvIF/bTVodmeySmcm1BfMcSeM411V5TO2APkki4ezlVDh1oDxaxxxr26Zyt0Gdl7vcbmGKUN8SIdxDPGXIQY9ieNu7gz1bagbHxn9U6+5E5BNkqxJRzqG7ZJ3qx45g+MocMjjRwrB681vcCz5iWTnE+BHOYydWDLIMYI8+OF//FOxzN9wllbyudjHLsCdEaMr4yrR0aDuTjVWLtJjw/t1h/9Gj9PACkeLjbz8HcWQKhXKJZoUzd2SBGgGYj6HNfjJ/siox1k+farfBOwLr4McuY2KSVgFTxxXJdvWVR+u9BGrnfWnzo/lgeXPPuksT8ZQakaa0WXHLzaEVO7lUMrLjNfXzRy4XZ5GY4d6XTLXM+0dvMdtPqC7VWFfMWitV3m2TT1qL8Aam7MXxuqXNdEORAO+buY+Id2duRemlYstDr6nhJ43qZaoFy9aN7lHVgf1wchlY6i/pNztezrdVjYcNeF+HMP0zPxys3nTFFPnEfNQKRZEPhlkNO94PRNRwEJacDO6tGtF7HG5wl1Q+Ic4X2lT67yMwncJ0HJqvRyrz4Z8tORKLq3g0GfMoZjov1Moz0KKce/uBqYawUquD3AUzbt3q7UUxhmZzE7TO3mnqduXda+7YLaZBwrydernRwKM7ylawbIeThBUld+WJBFCC+WmhZpep44CzD7oFm1H35UEwOnm59Ni+fC7wVyK4mRtICDPFLEfUMHr/1JWnKKBqfm7MrSYkQyq1nnJABMz+AXjAwdBLgT+dx6pi8R5E00zqH8RlNhQNOsRR4VJN6mQyyNZsaRLFy03lDiZsrSscSoITReeA/E4sBT+wPmUIs4ehCs2JXLaHCqHcwtuUmDD7a8LXvh2+XwEa/3v2luE98LxDx9gUgAN6tpRgbPpCYIyheIEE10As7GgTBEcYE0juk5+Q063TDC7W/vEa76OVk4JwiJLb6gYE5R/GKZLZEbP1kLgpzSzR50FsyWN0IyD6SDU+u9v132P2BqGipUST4quRGZOxn3JUOZJMrWoBi02nK8FcwJGfwu7hjZM3hRfH3PK9G5qf2Cm6ulnC2AR0/vzhdxTz1CUjhc4ncGjcRCg5MpXExUE1U1jTREV2OktA1/FG1JV99zbjzfFZikJ/vObnZ352qzeRPK8xIPSG+hcDR51Fy5EcuMvdbCFMd+Jwhyxh48994pB6zzMMgYMmg8FbteYWpu24E+njq0Jv0/Oawga8yzSbVlDf5gXfzlbq9+y1mKHLudAP9IyLtcGu2Sj8Lav8zNgeoNkfGcUBm/RYCfhkQWnxTbE/zrnqxTCdnDlnBIjcmqTJNsi+ApQoLm/vUracWNU6wGZrDJa0Nd30dSSxZeVhxyQ4NQHa//Hq0mGXntN5h5hBM1FKroeDVODinerSrTOOx0UdwRFwZbBtqRje/08gcuInVUrnAdmQfW7rllprnaVfZYLkDyYksNJ7UUYrDzCZXyvO5jLAEuYE+XdTwyeaaMHE1eAGYyGfF8dQWL+81z9Yp7VzjRBhkDaPjjTC5TcRgVwqhAY0a9CKXkPG43I9zZT+zz0GJvP+Xyw6xFPY9k/KBJeMdmyrk3AB7qM7ogvn222v3jNIT7Hz0MbSVbc2NbTePyUnRGD1ks3K+95A1pbtDqGp5Plmw27vZLsCKb8Xag/loTD6W/riSCsjU4ekj1FDtPY6PEFMkADw1AuwEigtSvpZdmRog4yXUydJRhbheTi1XxogbnjvspWoHWYKj8z8vXcfrRcGG717CKxyfeIN8Be2StYMPGbTLzhWfwx30EOFJO46hlbcGXVayWZ9XgdAwS/qX4nkU8aZ/oTQOS0P6kQ50HEE6kGdxTL5oxocSVINEglkIuDw+Sfj/WFU0OS84xo6uwrAtAmmIyePCPQq8RGz6UMzOBoXmCfcmIt85EBLAfa1+P7JOiw3df79QxzZtEIEyk44RcjMgBMjBQaNqBwWmb+BWxKd+3X6VN5bAqcCRy/WNp15h6FecsKmmfEb60HKJJS20sB1eACPiYSVL2pRpbmtY7EgJRqc6MEAjnxgBlJmQvQ65cxoTtNuXKO/4EUJp9sQwzN0mnok69nlhG4XNSwk1X8ShSWO3jwtFJr2e4X+tch8/j8McvKY29szVXzuB2AGA8VFGxBpHffaujFepCz+C2h2nBuSBqmjLUSuwZX94YMbMDBlwARiuSguVEuEtRtlV7J+ZaPQ0jxmKB1MIzPNyh8yZPgZXextwvoiyNEwa+Zx0+nM2zBKIMvK+geJDZb4OhoeqRiSIpcLsZ+yL0u6LPwifD7YbYd8cAvnNpH6/Fk87PbjBN8rDgM+VJ9oWbIKWbxJSqKa5wFXA0y/+O/sLOCbyygrwQmGjN0Es7JXeMvD8uwGHxAk8HnTW2W0cmKfY9IACyukGoZFPk/7un9GjtQmOs6TKD/TY7gGqP9NfOzjBF9oypGUdUzLp3J5eXof5ya+VNC/BfvLCRGrQfItuWQpgd577xmt+ps6B58XCEH5nbv6518V5gjdvR0dv904zi1HlBbjN2W0zRKpOtJaoc+A6nT3y0FwIOxhha9nJPu8pl2eP3zdJSZrtTKIxQHIhN6p+Ne+YyRtTW56OPCyWFe4bXfZ0l8DIoQTOKMXPOexbILfl0qYlElaAQTmc8hoq7FhiVnTpeGQovvt5oGihGwtv3S+nPawF0Zz88lQup0WV3+86u/ndpOiMB9/c/oH2ypQ2BPb0qhFoW8jIA8Tko5EJfLX7fDjrQfOYAjAxmAx2NK/v9mxzFzvUkddgD6Gq1Tr52dBMHmPbAqDfZWPXrPD311fjUt7XJ0l1eYsbtEQ/HPXxwgZMOc6gG1GTV5STCd2myqcy+8Sj5HaiTX6+pWhBYLdyvC0Yi5cahzMd/O/ZUWir02YBHA8p7NCv8chZyGFLpOtnv4wFKWsF0+MAvJ7D4I6Qfjg+jcWBacpYYbe7xhwHtoshm6cBbGg6VO6lKjuYKpcqVGbnhGJiAUELZP4dkjBmzszOMhl7PNI7meiycVp6jUd56F5OCl34GTQz0jRmv1O0cRstVJEAye4bQkmXsBS6bH4R39bzFA+CUW8pyDYPX+F7Jfbg9VGOxtdBt1OxnbOOGvQkfVDIgim+S4XOsWcJteodyqN5Ug/yWe0ZxSJVTM+IyuUgoQMUZvnGu/J8az/4Pr8uWQ2OGth0Zv/ljXctCgiPN0Cllm2O1QLCNsckyCGhMp2MZ5UVBoY9ybSpDbThCsClkEFq2KGn6DCDcxJoTQPQRPgTLfMdSmAic1iXjfg3IWoX0/skOY//KhilszUZPGeTPFnvcHIZScW070y1rQial/LCLapgsHlT/l1o3nHzzsVkBXpAoe5ernjUTA5OgBR41iMeVLvXWtrfD9cT2OVTWROVR3DMGXUOHl4hc5UEph1ojZYjY14YMDzkMrQagODYafJ2HlCAeHSnPokv5eb+ySJuu+t+ODbUJCcXm5pYy4b7olm/PUEuN0c0qkVSSccixZBMrF5b3XWwvcfpniZvO4mT7wIsPwauVJB7Ph9WjVRc+JqjJhPLPmccUh79uDkEATsdY/wbmZ1KrN9T+LBY6YoAjn/Zl3OjsVcPFpyTvc6unE6avHRzeXksQaWu9BCAU+ZNaQISOCMW7hPJSn45vIzM4yEhnkzUbqcxk0Smwe9AcGIDqPe6Q6WJqnr0X6Ccv0FCZUugqL+HRaGqZl+VffkR51GJcFnomizdIc2Uz21WCrScxXgZQYUKI0mmV7+Xk/QT2G1i6duXpNa6qmnteW8wgKnE7A58koqlK+w4+wAigaaw0AoDCkCzX9Q+43q0l5K86JQrLCAVe+ibL/kR+NrmWSzWm2z2od4v5Z/cVqLelLZA24tzBIs/7SbGNIEgg3u439CEP6Tfp/YnropsWR1OL5OkHOB/CLb/1T/HszBfg2qsAtsTHNwTj3/zc6J0yEXmNPv37TeMi7qyomjCMukFaiOgJaEIy+wcGk0nQTpIaBi0bLbiV5yeGWlWJnYSBqvFM7sSIA6yCyvy54r8y9xkSdsbXAdIE2x3LCm5tsfFScb2T8mCBg4Zsc2861b4o+B3pvrh+Dz0UMPCLUsI+3EIfSwEsCnaPd88p/v8AkIYhO/Gr2WT3LpFxCIdrtB6NOeTWX7XC6dXDMZz3lF+0OC/2f5N6EMUKgOuS0a7+cpSNGLy7TkTGA/sdvzHQwfatMPsvQQ3L2FSJfwm28T6OY8EWvIG+NLZvyP4XHj/n/MJuaJEe7baPRshTM08SoKGTooLhNmHQ/QV1CofddG+WqPKMVHdCWPLbN3QIiUF6ls77lTQN4NJZRK19NDnzbuzG9H9LCxsAVbLQ7xdV08l6d4ey/6yI2QvpAbncnjzDPoW/O2QF4f35F+JJMonLzmJYvMyBZCXFrEub8Q6tCcfRXzCxxKeEdBijNSdd1+iPn4VXjUJ/dlLFm/y8Xa7BxiD1//w9YIGbMsMcjGK1PC/RUyfkcNsmJuPS5jRRgVNufLwHP7sjSx9pOxjeAS8NQESX0pupK3tem8rgO4XXDkET9xpiOfr2Oyp5emqIrTgXFohuUbV42543DKcmcp95tSDZtvvpK3OrKHmhfatoNkv34ejUMzBMQAKhC+OZgNUy6O5ZmNsyL4XuxLpi+Twb9VGyOd0xknRNWXnICfQv/LmfaWQOrL7Z3/6yMpBFfxWXbe0MO3GycJPEJrDkjvZHKRGF5WV5CO8fZlb05eiArHyf/owpvTJNxeqGQj/9zjsx4W6Jc04AebLsFHEL8y73M2xbkWVc3QKHq4vXY+WueIcwkAR8vaR8qokeNMIM0PvzeiaJu10CXRbXjrbJz7Hw1FUg4PjLNFZCH7yjLok+yh9Ji3aJc7iUIIcrpqocZx4XzIw4Tu8VvQFZOpAEUG/B+hCcyZPTb5YuW1nfoALsS+ljxIx3BvPdsvp9KRaAF0EV5/E+nkJPczNk1XTkG0TDrlPoBkgZAvZGOJuLJXVuogR9noJlvjJMH8h54e80fNnkOgzMYNs7X8UfXc/lI6HygHOESZKQyVxznF1gVUyc4JwHp7WyUn0gs3XQDBj6q/e+sgps8/7obIgb3cc0T9OSOR6zPHhRUzpXdTNC5HOamKh+PXRTdJcxDIn4hUeHoPUJVz+td8AcHZmH/xzxiacqJCyZ02Jdn+6f5iQMWziXWKYl8RtCZpJqDpdqx0ctJrnt8vS6I77HU/6BrMbokJVDxuNSZn348yIeyrAelNjHD1o0pOPATsC6COzkZWiAU2Xhd/mPPQUXvmhYl60DWvzVbgdvL23QPy4RjeAM6QVNoDvrkWmRInXWX+Ewv1L/QWFOfHloNWoVXTpKhAy9ily6fzBTRDpIOThDyN3p0iuHkM0ZRwgcVZwD5j+uiNcDFiPVNNPeLyBCZtjZUX5NI2B6JLzLA8WIUmP3PJ/yscIKmumcNSKnyis7Glt5nVAieCdFfl1sYT0Z3npZfnZPLYunDzhDs8xI1wYE6MqMAbD6zlAH4dFXMnk8GfAKTLIOvUGHIUbInpm/ehkxRy/V0PnqUrxaOmrT7QkM4DJda/zpRT1YJVRKOdFGsgFfa5+rowde+8iNiKeBMXL6t+nMLwAx05oyNwqq5D4Do7vFoYrdbEL7dvYoC9BuqNkZyGPuObqvaWDGK6bIXipp2ZWWIcuOAl1mJocx4mws8G9koIfoYOXaXm0vgmGrzS0t2OI597GcRumPPu4mCFQelMQDj4pkwrpj7vMWPush/jBfOSoe1/GA/yrds4ONF4AScMfZr0TJPw09OAeiVPUfmpyhI74h5ptExNTfxUIQh4hUltROgmLR97w1DrP4gaso/8XLEVgYSLXnN30AMsTIjhQEXX7bScSjcdCrhwJzhtGJiAamb/4Fni+1j+f9ZPoz24vkCF1ItT9ywTNstvjKelExjHMkaRaGqhqa/nLvAvQZnvomXd239XQs+RQTbBJdNgpZc4X2Wqheriq4qYH657f0zpsnWCgMfJOlIX3nRSTpEg0n+NC1e+BBlZX+dZwqVGFhLi1TrGs1oeQg8Dqukjp48jDXk8ydxBvx9tklbpBLUEH8Qx3U585uSRHHjj2HG3Q0tuTEsvmByzAvZddsa87UYa33StScEOoKWqRDLh4eZbIDHcChNv1YeunADEey02VhPzg0XypaEq7GnymYjko5fczQrhylOW8X1kYZFRvA56l/Oj1YHZbEd0y8bIZ5lj0cld8AUqs16Eg282QsKLNE/NGZAaga8LJVDCH4aREUs719e/JjllkkuoH/E/g7zU0QHQ7lAO/5xkns5MA396hHAGxHGgHbe0QVeq8xDl3mTv3SONioIc+kOElYkAsl2EkOhD3EyCuSaTXddJFO5QmH4DYcUW40rQZdS5VdBc130CzjiuwFr3I6ey/AS9zg4NbSvt6uJiLVdSAfCgeiAq72Pwf2ahmimvb43wDE4U1sP7OmcZQH8A1ulvWJdjnnCpUIrv5VCPN2e+QPHJuRnvM0doglKNIkbyOJudiYK34+IgcE/rpxmMDL7KG4O6pBLmZwe0IxYFWVSVpIge7NRnIp1LWHYxD93HyAoMjJnzUqVxG6nsn/cyUmJcqDd1Ls9Gb9Jrw01WcOfmKk5O/Z8ZNzdIXZQRsBO+I3cwFGlkmX92vAKvxzfoBkqDncZ2NnlYNSejhNuAfTB750RASa+TGtuIxFlczzYtxHu6AZ2vWdJVjAhRjet81FHllVIPCO5V4x/H9esDAFdEgFXgd+dciE5JvUkbO+LmiByR2XS43zoa5AUBy+plQXiIl18xJFl1yVhNqerQ1wAzslxlPRsT7NQUzDExvYrk7enRWsQMeGSZVpYlad5YUGCWSzvmc1ENuB6TI//oS5tDKXMlKlXZGdz8PkHqGkpnBL64b2MUj30PwIli2zYrrdrDjajnQZ1bJbASb0KukwAKntQz0DuFTPEbp8i2/ur4RoZNlgYMgqJUwlzZDrMFuTqDg8wbQrJc3+UuGWfkg1z+XtKyLkyO0Dbehv3qxA26jGKdTSZHhMF15XxSBSitKdm7yymU2hqpjMPkuQbu9PRlQtVTh6/bylpMcZNYJn1p8l/eVw+w/1fGCARt/rjJUZnTPeOfIyo4RFUmvVm2qDu+yuZb51/fPzZjyg+QrbwEJvlhctoh9nvC9ohsogLfo3WWeMjJ3o/MObNK9EWe/yiyA+uELYvj2f5ekgi9Qak6xFyafzxd0b/aPkj940SkacrdXewWjgkegJAzw+zgsop14CqmabDqBZdl051UXeiVMRq7MminySakmoX8vxas++yrNdmCpuFNn9id6qpaFRShklk44XkCgYo9E41YsvqKKPKcvkE/X208nFYtMgALwt1/AsEdyr4xCu6bijBtUg6LfwKGPKgw0yxsXCRKTt3xGBEL+f6GLe/14TLF1AAYsMGlykaSLb44zhlcXst3EZerpqaIJjh6ymdBoDThNI1sT36ncE6jLhNkE1/3ZzjDNsbEAQmqLrZ46dBxltpjP7bRmPCpVQAcNkMcw5ZGar+x+CCnsh3yx9pe6pbouxdaFMtFlHW7Qw62lYCnEWhf89PC1ZaGyIKyu3r3pZi+3xYsc008JIClVuJJ4WsgGfMU+uFw/t5M+FthkTYoNsXnykbrBfAwhUFCqSXtXeFs+aFgTmUifVBBy9oO5dfOROwB92pQpTq9JJNGQNg1nQY0ZA8NmMEYbIU3tw+LZfeLpqoR1G2lIUpZ5DIBbMP1M1viXFjWPIgofVZ4q7zAPprz7vxgf/g6LwbnJE8aCQWMVWljrfkCpvsk3NP9FfDNO3P/PqccFdddsNxHIHG2H3wFS3/jMg25HwuUTAw4/e4v7nosz33ySvHVUv6FCEIa11vC3MDd8TcPIxVtSJB8KMdpKtqq2wt/bkz5I911hR1r5G5nWMpCx10FAiu7E5Ek7akq3LycGvQGQOnZTMjpk1JuzzX356nDrUyXRXZeG0Gb8wI0d9QLyhJj5D+u/35lSFEFw61p3NBAPJyZqrErvfoxqegAgmkcbQW9lewetMOmjQY2aGMlUhen0MGcRJ4o/bOitUFv/Irta23QKClvghK2JcqxOv4LkOGkc6E+E7RARAqhwQ0Z5tLI51zX3M9A0Lluw9yFhwSlxFsBzhnxFPbFoKo0eYH4M4WDUv8naSnrBiTWrpiLUKB3iFlkuzUxZS7UIWZnuUuj7KadxeTYLJKzwLjhiYETx8elVHkN2cUhzUwEv12Zzbr6EE5M/46cuHXU+E97vVudwp8oToCGQvmZdVa/5UXBfM9aqXBrm/NSS84gwvMDICtMKmpBa/I8kfrj77vOJZWT/UBzjwqXhfRSZDsnat7gsJKm1HCYCFCYTNbj8GapMPOeFaDGzejbRU5SDGxa6eVvx5nlvRp6xqAmufDhXg97HH6IMG8UYmQoxCl0XsLh1uh654Qh9zA6G9mFBcAzeMnafRkFHh3diK32tqeWG92APNvS7roMEnxSINId7gt0I2iHpRMSg9YAS94R5KhjAtNFBe+jSIm7Mhx0PRq/12IKZjCdfyboClOZS26ZZ77tduQUKeyTSFlMuguX1NDm15ylfZiYqPWiMOiGkgA3NP2cqCIcjAnzMEzsVc5D4T6BHlmO1sA66Zhd5jQdTo9Fz62UXxXHwiK7p2Bc+9siP+2J/iJpPRiA0B+fEO1WKwBQcu07BtvnVl0ePguISIoL2V48WAE0p+ePUT3cO2EkLfDhBs9Oo/sRjjHW8NhwsMtzq4EMe81bKwr29zvpQQr1tf2Zaor64hR2Wy47Zo6A+KI6zjVbNZqHW6khRaNSFBs7nmsLZX6zRdt/cyE1fE2MLKxfe7TRh4RZrEl3fhK4SDvOWi16e374uCDMllH66CjpPD22lQYOuiUbatKQcmg4m67FUtFfeUL22TQNOi6HRZozztS18APZjZgtltPGC26+kYYmVl9VFRnFdSUxDLBngIIy+N6mfw4F7nWEQdusiEkOo2dIlXhXez1svnxCk/SFQL1rZiwugmJpcyaLDSpXFowcUp0yqphX5ly8B88myCj/f5ZjXbXnAvaAOb5SsvrDdVJltK6UoN70gLYHEjmBhWP2k15SmaLHB9Gq0qNun+0DHkj0DHDE4/BZ9vK2Cx+4beXP1P1GMbfyn21u79wUxH1qyci+qSVIpklPNPUaU831NylYmuPvDH5jSGTc/3WohTm8LoSM7rAICeNUXoWTxg55vVkHi8gxFUUU4s9IondQA5OoTdIVs5LfNz81OnztAu1oNVWGWvYwUNl3SUG5v6xAyz4oWn+HpO327YoLdOI1h0IHCjkVfevgmOEVRBKpahfzYUSewT4+kOspF79TjlX2sxC3eRBkvdSOVoX62MXqLyuImxNmR9Ef0M1GTrKn6Tzsz+p25BFlogh1TrIObr5NY1SIKd+Hqv+fwVU0+yUOoBB4HKebQwbY1D8JsaqDMIeIRcat8GytVs+aXgB8D6yI4iLXv6ryKMB3zFQLh2fvsqnRJIuKdUowCEDXCDykTfi5tvLAHPhOhbzq+15mcsAo0IsNAWm1xUnYDNJRAt2bCmY/UACowCkae2zfPz+9gE2qIJuHSzNcDodSixu2QVZBsLH2bIwHWVcEOb/TEcv/ZmUIETnoZwuXhKP9IpOcbEe0BFD4JCjtKd/ICda6a+ymIBey94vxmVnnZJ6Hu30XjhBxcR0mQPdI+nR1Ho9kQsaXBNpUXNl6go5v2PkaQ5XG9p/fBfhf6KylRS82iAis0+8/INnLD/CRTdP8c8LH3WTp2fNG+3+PMWzbzZmPstxzDwQ68ormMYqGd7PNcskfEOAYncRZHkon2KxeLej3dzjPJ/BEw2Z7PNvgRZr+nEA/FWDsREYEmTr6WrseKd5t3ET0ZwsTesJHH/eW1B/ntMFmLC5vl1uzj6wna8AXvOIt8GUkdoHNTUxp6Ah9MvAQYo/ML3+1YoFGUtIO7jBpK6I2h1HdNhsLdb5xMqdFEdoR96ANKm/1+axzURD03gwDxUKx6gU1W+cZHxXdOP9C4AuYCsRRZ6wTw1wZu0JVGQ71D+FUrg3YnCiwVPEonvgqhABV0Su9lGPvH7ixwsvH6PUPd4VplPFb6+Xz5CPAlNDoZ2+yi/qEWxdXxbNxAF+9inhFwdndifWgLzim2FBVJfZ9Ann3mDZGaoyYOTbzmvA/RFGwRDBQKuqTl/Hmom6z58R+WahJZiI9CwBcHCUBDF+8QcodEQ9F2Pq13Vgv15MdRjzRbzHaydgEv6/LU8kRu/atI/sL3YKip3UkRtKcrbqoVzwOrudBCU/dT0AKl6ua4wV3ezG/zoutzfzTMoU5UAQTPgXo8dColVHFpOTLupKPt9B14o+YnxJbERDDowWM6ctmu1kyaJM9dbDgzKv7a7ekt2v7GsCmdbwRi9ayJDuI2piq4xUUuzSZDJdim0ZAdXsB2/cQnRBkXu8479pNw5o8RHWishx6asV6wdc8Vt49M53T5czC/wcFHHi49x6IApiCzAf6Qi+osQBHvcpmtEMG+4X+ftCyENyU1e03wqn9fVBdWYR4iHTK71oytEucKv1phq/9/ZBJH8j/ysLiODJICgBzLeAd5LjFbnsWqjgplvTwUXLQQo0tboRBFcyNbyARrMW/+WPK9VRgHyJaoD2Q5PTAnqDuO6ceBZrc6KBcg9GYKFHPQ5ydt0HxmjY+l2a5wjT1TLSptzw7QrSNHegwgHIIRK3QGuqHwELeQe8EBZ+D/BdaEWPCZes7Ykj2dgghkalQrrcFJub3C6X2joI4lZpwWmgtKrMXM3AWIUsx6bNscf+7xDwUzeOPjrP1hsd0CFviDa9iuJqo4bFydI+MlQRE4dqn/S7sh2VTAbDej5KPErddq+Ujkx0TuXb1NSXiUUYu6cZfyq+k0tSlh0qEY8O+Prlk8VIrd9NNFG8aynIt4p1c/Payf2tWDWOIy/kNFH3uxgDL07eSMfF31w1O+9NZqRCE/ICWlumru7n3He5vBfqyPkDrs4dxVx1Tq3bt39BOWPrUFvhI7f3Acqjlo5vIJNJu/zWoeuEM9cB9nrPGMlNPy38PM0k1Tle5+cPFtMa3hg7d5So583GoArDOKXO+EqvErOHIeAIr5L/C+jzVEY2vKdGK3C/1SMHRNxya3C5movn2jyof/8SJfB+eepINJhOtTcKtbRSSioXZIS0RUkg28GKI2TtJuF0XIhcAgKZEF4mrw+prOXedDYwIRlfIYcj05/Ch0sMxp0SkdcVc5wYHTKSLLpnuYWpo++2nAmGm74KjqNVDHPH3DhPe50oJG8FLlihLuUEAJSQIlN0NR1MXzfW2yod71lgq8T+EtoXDVpLTlIcZIMwbHYlwGYAqlnE7vn0JQyONR1q2tWcIAkKUIFvEWGqQmA9x6SmevgO1v2MEfEJZHD4EG+idQ052FgWPOaUZieFn33o+EUHWiqTqgsbB4SZadBE7Kd+5GSu6T2T4I2TTGxalIpujBbwONZH4dce3ew0rnuCmBd+RSzpEoe+CMQSFreLVkEN+ojSN5iK6HsO+ppoN10lhurhANs8HLl/WvyBU7bmtkWUK7VGMXfPrk2XzN+KA1qNJ+0fPdRhG+2uvqpS5pavhRZrvH4IGAONzJuWa/LbEJPd7As0fGBPxeMqJwdz/6ns3zSGgOoLf9m2YCLKfSPD1XqFH+qL0LisAXq0Mtvfv1KKkGH42bMe2yYT76ht77t1GMzYBfe5jLGLdBDqfRf6+AcL7QkL49veqf4rpsoPTbgSe95x336+8GtK7kSrE95Cxe/B8oVK5iw2cKHzGwNVohz/zIDITt+j8brLFezilPsI/VvQm2U41aQAQPtvgqJwDKTi3a6eF57ws+W3Y1ZkGwxFeZXsaU2UnOhkJLBk2l4pUZmQWWgWbb+R0fqz6jXfWgaHz4yEclnuMkfi9BtjqC0hUyy5pMC8I2ETmrafFlYJYCeatsB+TaIttCvHK63ziWM/cGgv73QtXyeVLzHVOo6m/2VEsQs5DZp2NkQ0RMZjIMNnL+AzL2OUnZOFc=
`pragma protect end_data_block
`pragma protect digest_block
b878545b7cd477b36969513633c655a370b99328b63941d244954e2c84edb96b
`pragma protect end_digest_block
`pragma protect end_protected
