`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
pbvvpuYY8NHd39Iob7gEMbsrUg2o/eFFmRgtjromH3JLPVPr096NzgVgRGzCVMCCmIjrOai69eAYBPTnqPglm5t27b526ukuSBxMJsZw0fGw9M/pVAhHO9AUCf6kRfu7BvQoVKBCeJ6muwjf0bYJprea4WRNZ0QP0fwNj7lMcDLFqlsOXJBxe2M47bFwwWjrUmzm6gK6E+VqHdaYPHPV1oFugI2QoEo9EmdLsOL3UEikIOu6I3IuXoz3NiDYzx0GGSZeQdp9RVbq+fhgKDjQR4lx1YbgNf9lU4zlG0L7Ywl0V5Vv5am5hfBzWgKpDtE6NRZLACMEalsZauqZySFrZvcCR/QUWQsi1vfa9EESUan063r/ibYB4fik7VNBVgvhO1YssNy2EbLZ7IELJS9KrpF/vgbMk2AVrbxnis7CIgWVekKnxm8/vQuOsOhDidfsmBAm/QWXmG9benk+ElFSKnl5CCALJFVt+4L8HfudrWvFWHNom3e+I2KJUlz2ramhT/r79oGADLUQaYLSWfLSyyoJF/84ZGeEL5OI4OMW0N6Id24OZKX4yBJVB2L6g6C4Yv7vXG+siM65agYuwUW7NYYahfP/m6Nl11a347TrjpwW9sR4Jfz662u94noe6wuMxI9XMpX87qENa7Lx8dw6caMumSD8WNTX6ezTej8Ov7CT3jby09AqUtn6m9FTiaza/aMuUyzGH6eYJgfvMDVut6JRhRgE/JNAdz79QhJaCrbx3sOXSsFLhAd2Ixy/DKbJZinVHmwxe2T/QKq3ibyGZVYPTtSeLkJp1gPVPGqkvfaKkm3QtEpZPytV6u8xk+9K8GEbvJYqlbGWpZPsRp8q7BLyDfgQWaBFMRF6FbdeWeJYkUJ9WQvJv+ChGNbTKePpQTOWRJ++PSyAsxUcoMSnNqK1i8Ru9ZiSnWZte6F1JvzIykFKQRVmQJSF2EFPcMVN6O+455aviMhQ2hAgKuLQFD7VVTtyf6aTN3GvkFuvkZbHdPcvD3MoJCgyVNW41V9FOlsRLvDHDIn/W8Fi7NmCjv2owJd81rTZQDaF+AjPCbik3kT+HYS7Y9TFTF8SeZYQdc881Fuv1443pVA1pcHUli0pXDI+WM7+SN3ivbxZn6jek78rTDz8YjwliFAvll4CeXX49tGv3tgx7wvzmm4C4C1BrT8KSgcqkG2CKmGzSUxKnwICbY1pjH2bonGKooGa1e+Zsl2ND+5cMABNugRv8ER/Cibx7/VlZraCIwHpJFQGFn+bCGRkEFdUMgUyR6gMOrBvktCn2JNlvnRnUD2OzG860bQ6iEDBqSfi/duNXrSBUlGdsRQ1vt2AUO++SeVnehdC0pLUHtTkRvDELgYqC4rQLFB61EdeokXFR4SufaRZy7ZCaIaI0og/Z82dWwrmKHo3t34IcTZolDLs0n+2WnjDISiSSbDDnUVsgvORUjQBhNeNphbLlvKfU2XSsiVd9dmgzfZwyckc1161g36fS+zDCV2pRBeSSSiXoXBkOWxANbiPI/rvijCPldoxQSgc+a2TR8LhokA0XDRlL+a3etmKIfUzOPw/j6gVrJwCdZ258iny2mDUf5Hgz42KY3hh24nehklizShlQWtvDNTSEt/BIFz1OBGLgb1yRuPKUfhhDub93rdXQpzRvFUf68tCGWkJG7bBBd+m4+naRoq98PkrPzbyXtiwQ/27EBPoG94MKmLSvSJbwR0Bn9IjfWCzBLuzxH4SAiWIwS8xzjcoqpVVFYM61x46DmQf+vm2L2DKSQLgP0+UVvSK4QJTFCZUKvroWfYlLAZWhLwzZ0MOOxNQvBAFXZvEcp3ri35CTvJs7C/mThn9IF4Q7YnJv9bbDOsnaB5Bk/TFI6j4NZJZvQpIM1ll+0//ZJbaA3Uvv7dVEwCoIHKVpqj1kSAf7MTS57tR2yOYk7hoKoaQT86tLycvoUjkwfoQU1q0x93Vpb21fJ57pz0aAaM0gnCdbNQ8nJpi5ockuqwS633wS49qplXZPU2wPhZHWDhKy5/DUDvV7E+7bMdM2WsCpbijwK0wOWZvC8q15L1eakis4FqRSKj8EFghw47Q30v7ml9BHLF++rhlKo4OgwOyiMJWhtNSv8/C8QoLrLt9PIE7nlBURcmMH7m5LYbDW5WWBJfGG7WT+iLYeP2hbmzEdPfNcbDFkkcai4EhcQr9IhOCfS4pv278p+E8DJ0f8zjzxUN1W8eAObmy1pllTmoT7/TKRC3Q4VKG2+299G8RoLvuqeUXVcNMYM9pvZNrBzZcWVQa+Lvu5W9E+JB8QX9CibWhCzQUl42k7i9SYX52Kl/WU2yTqxoJTAibX1D9wOskTFUQHoc+FdAqI7GNF3jbDDSwbrVTxSHw/LAg0IlhCxwWyqRzeiWrkuMM9BmBAX04Q6BwfzTm+wEkCEQ1zk84RFVMZK540gjCE8zv2kBq7j8iRs6gN1HvPIkg98C/0dQ1RCXFOkjfVYsXNrUedrOT3IAZ2+YmD43jBw52cXg5YdtbSEbd8BLvPXLOfdcn6jd9s0rK4R2zJ9dXNsGTAoXbd0nT0BuBhnHlaoCy0qMepgdPaixGvm+ooEu6YeldNH9AhwtmUm1We+/TQIDLV7L/XOA4lMEivM53PadUL2N5uD8axqBokxqhru7cdVSmOCrYnmnpb7B6Mgv/39U9YLsz0UGiXevx5zJZOCRxHnqMg+KHiT7Bs/lK31WbKQPZSl5AfPdyuuFoA4iZD4BIoIAvo++c64gpUIhUp/xiakIibP+jlsFD6tuf4h6sVu22Yl7ejN0huzevSVxdOcRlEYj4/2JfOUpR2iPJ5a56TJwKptmkODeAQ3sio2LIxQ8wS/klDJ6Lq66tdKnFUtml6ckywkhuhW5bYDnAwDbhbysXy3DvIdKO2SvJXombwZv7DM+b//BP+To8siXKq9T3BOXTT4biyQigoXA/bmKkrx4VUuWFtWYyV7K+XGSIoLMNItGvtBKJUJI4aO+MZQUOWydUBrlIpzuO9YUWhaLUy90uAfibvjZsdOL013y2ZV3xb84jcHj+ArMiDPa1DqZZuTeIynCNAZ/o5ezIsY9DcliX78l4nOZTOTvY3zidOkTAPyd2exzRQRy8Dx6638Iiw/F/zZU9P42Bfpqq5xldXXdJDkeFFHiDXUFOGciriSpXPcrnRWGBbq7B1gPhkcKj7fYhJyqWdLjXbVskOg0drBSqZ83782xC082CMumDCN6AR2HCvS0MsCaGuNPV4uiMw0fhgL8varQkgcr+u8Yh4Grth+Wh47hVqWxklKo2WAag/2FSwWpdeTM1gS9I9MpJF+mhAgNXPPIIlc225HVokxz/MA9SL1L3RZlSUpVTfYSYolklwSVa+8M8uzSl+dca54pPHLOGaxXRrOT/NXf1BNgsaBiFIMsMb57tXX8YWhpMuiYfGL+uHdZqZJU/pwKVwyIn+eZ+zr+mvUeH90he3upepF4bu8jiMNXFBrw7iJLRz8x76WCyIU0vp57BL5lpgE9yuaVsOtN+lkjlAF+mfh7OH3dGq8/6E7rzGa9kx9GfV6UjfY+dFGclFMWvaIRN+qGOmc9u6cMaFZYky5v0KaaTuCJo7iszIyfdl30A2nRonTUTB+qG2fxs+6qgPUFz6jK9v4xsziPoN+5iMiOCstcShEXSxgw6PZXDn2AF8L3Ku8iZYj92AwvBPIbjW/Xr9XiHcYvDS7oLynJaIKnqKJJtIbF/9ttughtyW6MD9YilPBocaRCvhsNTAj3v9d8v2kZX4TL4W/fNKl0FZkFLagN2vZWFyjesSNZi3I3nqc3qwJivHZy50Mb12+Fc48uh09IW/UJPnLSZkDOHanT99LRTt1g/qG/ibUONomW/siCsHXkWYWsV24wb1ZlysCSgX1YFOhxZoWmxmRSHuVs8xMhKVA+GNV2M2aCxKScNp/f+TpR2O9Sqga2o2w4VJUI/QL2NAiH9Z5RNsphKTFA6myy/nr1gTTJmpFZRIIvfZhpTNmnmHa0Sv4qvWK6GJkmrU1mIG46ziBpPhIRqrUwesS7iiUnEuf7Ers3ptjj1CM75mKZspnUC+8AVyMX2Kp30BJrqJExrpOvFcH1trH1eoDsS4xX3ar9A/+Zqu6OW4muHwfyCmzmlbf51x9ihWDgDSuPGYYE+a90hyVjKZ0G+63aknTjJLq5yq4dEkzwInfTvvJrq/32ujNMAbM4zWCjzxoxbEOXWsIE+9XjlhBOTEusU1yjKv5mFC+pT9pxqfLTFViwwuS1mMZ4RoRfGjWJ7o4ATHor2TbMZkiNc7aEvEymbRz+KT0GzYd8WQSTjjSi2mB0YGfQULaZTRfC27+y3q+Nndm7084p7X7e5mrxDSOFrLFO5z/VCytGpJj3VZidI3t3QCconihSBjl2B5MPZG4lyTNV1VLwTgI14hydlHMENhjQk/nkYLvwTUZYyVdYu/zq17so04uBmdTVjfhXAgwr2KL2iuHmvRki9SK9ib1FkoN+1f/M3JH3kA3a5rJ9XVEvNm2K1EY7bn8FEFg49s31D8XZ3pJ2Od0iMtUi5XrepXuNlgb9I97zdKNWvW24c6MT2Q6ltuCKQViigv6dCowHow8M6exGgQpq0udCR+JWsceU89GjqnbzWS7DK1Pp+oggSUp2BN9V8WV2a++W/bIWlh2NAcezFN6TKjXn6Rkay+rKEdlBkWNA8YaGzl4bJKltLoyPCHpZF1v0ZuGnccRfdEEoOdXeJzEQ47fkdd0JBplWgg8vHBdpWL/mfD1FtftVu7j1ZvwdxjnlmAU5FmLnM8KWst94/HvhrIK2HRznBtx1GTzwSWXIkkCAolFzS23j9qnRcG1YPEc6kP7rk/me0MVkUu6OpwEnZJLc9DhaQbDAKM3Gdq71V9PSOcHVhBiA1FO98PMLgfXCr0E88cZxgctIsG95ZSdkqTb0gKKa94dp8yKe8RFAd1FmmqHRReHuNmQpm0TCfryqbXEsND9I/jeUtQF/pKKcVtDj02yqltzi7tiB4pLBvgEwQ+FmBTA+U3I29GmJ1bZV7RIJ5ygVuqQbqKeOa2YaP/eWDtQR8ycLwfSkqzMbr4fEjzvHBZaNtqWTWqzOX3BfHhkjauT9dPKU+LCT8AfT1KHWjJCMTBwvI0Q5bPcl3dfFy0d+WYAGVoTRII2n0pQ2XvNyoipQY1ipPXDzwx8oBEr0ag0LReDBQRjHRnT6SDeVO+sGxFCB9o3/278tNurt0RZGGE1vw7Bi6UOmozEfzzfq0FjJi7DEBTDVr2zESyoRuar2AmMSgIgpqTZ43SOiyCst4MDKRon7uv91ik9QXKHMqhjQpE3nRTbgmE3bqfBJORYCD51zhVgHhdkhaTccgqh1Eh3zX/jrp2EdvDRPbW9Mg+KKpjqYTrSUsYMvp8DOpLlCyNLz2d/iVaedqoehYvfV/hlMGjYi4YhY3GN6o7WQGeE5xykFPHZY1Sg4zQPLB3sV1NDy7d/cYHLr4zAjM/O7e6D2e31KgxHtFXddvv54HWcXF0C9DlhPzi74wZ7ZS9fkgNLgWfbYmuqeyjxi/qW5zirTYyEWQ8x4rhExJzZr1mcydRL2EQJtLbPdyUYY2hkhb8QXRjbzjXe8kEtH+fWEG9wFN4yoaBzvwpeVjShTO91eeiN3e6ugOh0krVZB73Ny0kCh4Kp5YgQWnVk/DdL7fN1QcOhjr9ahpuhGe0jsVCc6UcLNvCGOtXA4EuDzPqF/EhhQpFl+iv99FwfDTbAJdJr61lkaUADhtMSo7RvzO0wlsmRHS1j/hvmQecwJP2m61r7osI9r0F168sbJHxRdb8dBi/36yx0NHd8fOb7gdT56bPwbJuHtPuTkdn9ezLbxoPkpC2gK8L3KK/vMrgcCWqrg2yGQ425BNv+EMaU0QINqqGAWHdwssaxf86A3epHSmLHKizU/r3EIy7jVTUDfrN06BII1T/+ZSCiE94g2XKqqbvMyANT7GOBH/iKqQ9osW4cLPBwpr5NE3qidZDcpRIOqm4YLMGlDGo64j6RDPNz0Hkt+hDRg6u3sW0L/fWZ9UfXUGcmYTiXuHyGgFDn2jwprn/zmaGgplsoB6RgULzVKEcMGcFn0xemC4WVMMdVVPiMeJiq7jlDVIcaSMuXCNIR/mHHg32jltPq11NdmsCUAf8oT+7jXUw33ehMN3OsBHkCU5jPaalsfYXMmYZy9Fo0epMfZYF6Qp8NBktnlcN7Bi/hirqIppzalE4BIXZTFJWy7kmBTQ84bNxZgyGUYrhH+UjVLvYY4tNRotgiZKR0nuNMSHcO7PiKmp9W4A/6iZoYTYnkZIwt183G5e82oDikvKP9IFuTMFAx1Vav95P3BN8JEOrJSOY2eO8EaWVMST6UNPf/MsQS0FuuT0LIJKnounL933CXAV8jXRCT9xqT1qrdnUHbwhb5UinUsMclCpNMocHK8PS21xLNkB4k2kqbrZEvt3tOubzkHB1mP9VpUjZ5qfxmgimCIa7zWJXXyQBnJRg5nTCthK9V/DZENae201yLlQ199sGsQhKy5wWAW7Xy4vdBzRlCbzzc7QRaqf1lB2fiG9KkrpQy4o53ejKtrQuwThfuzA54cd9APSefoZPdTcT0LMCGaQ9ZJRmUjqMTrohIUbEkUbPTE7iVL7ZLTFM9jjhTXRRvkJH8aUV6rtG7VEG/X2y83ewjhDUUD7A0XcBG6813VpJLlPwIBXaKsRhnKSPG5SstcMWgdh9MQCT21NEINl3j1s24wxocQ7f/Q1CITUshex1h3LL0bRJ2KstZjPq3R34B0qAjcL9+aEksrb4Tbl70VkOup1VFy4m24yj3V+rrxGC7oUgLIUFdyIjO+B8fgQTt0lqYFNs3VeZYebQOv4E7OKenjNFKCCcnmquWRCW3S8tLVHrweEjDm1Zmpzy34CxGvjsSisu38IHAk9SbZiPNUeBCQsWdC0SYfe2viKI7BDj8CzdmI+EFnjS7Z2bE7FSWWKW5ePS6O13+PKkzIJn6b/b6SoDIXM/SHvI/xQbH0D5RbVJiPhevkvf81j5Q9LlWD/gvrzcm0NzRHNM6ucM4DNwToBjLO/sYE6y0TlBNAJavsfuOdtI/YrQ/7C/ykYNJUptCEEdYps0pGrwi89X2/iPoF+aFCu5Z9BwMgaOjof/z0C/wuF4+Uy6jhkii3g04PNIxkNT+7DmkF3srW2xsK8o9x7q/gt6nPdYIFzZxC/mwhjtVd8CgV3je/bunb/XbRgAjrqlFtbiTK5mw80qQsTF80hcVUEwH1WEjQQ8bsHY0v4Hn6aVowdhBQ1az7ZCBvjMaGnoy5YdfKTMCA+J2jGlEplEWTLv8eZ72fS+fqlTs2l4UCFTtLr6Qo7qSsdJyREei247P+WFOjfROgcK+avShmAQz7y6sCjBPTrXiBvgQ9pbPOqEKJpwuNmsGl1g4bamlCi3T6q1F3AdA7ljHX5RW+myvxtSAjqhhPInAjcph7cwE4axnwMbtQyjWFcm+N4bqG8mMPLhi8NRTXZ7dzSlllqRO/vHvuHUmfsxvcG9IIDKC8XNGABwErKmrA6g27KJHaYwiwHqEdHm4swuAH9nUuZhv7yy8qG7nrddtgsP23ohURMOHbFza4Aek3/RyLuf81kLJowm+sO3E8T5cLYoF0SfaAf9nygiKjanNqCoW81VBA72tn1zDdn4/oRCtaAP6HNbp2hjQKP78RFHSBqsRVNCuAD113p6O/c14crYfCFhxeIud4yS3LOprbpMCgx8/FkEcHpC8eFjrLkZ48o9DZxcGyWOSkKRnyEokOrGoFHB2FziExMLB4GleonjFM7rUXOLg1SUwasrrWiKXvUjBvj6y+8coD4DjY17oGIORThX+SE5dZGvQXG17wfrvbqtMBQxBq2PjTguwWTs6P3w4R+8LDOR9QAPLXVNMdQ3GpoJkXjOI7sKDGS4LJJzqZq/6PHpC5tUi0MDkxKI2fiZyl4VCZJFH0QHXrWB6lnzxigsAuJ6iA3xWen1VvZqM5RKpXaiYX7WMJHyTRCdPmtAZ8ZiFhB6+7bfBKojyQ35WgE3X56/9druZC8SlRv+ndzrloxm3vRKv0NNYGAoTEvF6KJx9Urw+t+V4L1awmfICIzoVoxia94YA4OrhDpduXp+3Dzh+yrK9R5Ccz4Ip7rZaOiY+pI0Z1+gpGjiHDd8/pDGgOqMu3LyBsMYe4ohEIX5yGuhHWMeS0guIUEGLvvhZk8I1rF4dk9wGvwD3f8aICL/E4dLsNzjWkpFuuqxJmY0fxmr2tXLZgC4si9Mfy2ON/2fFzpjUlN8e6pP+XWn8OGr4Og6jPeGsOzpvJCBK1ZihMEwym3QI5PsRD6BYpo1jkJW/1e4VLw/TJr01NTvrwwfMKme3+mG96BIUYNOm7mqJUNeHHv2PIgpi49SQbCs3UrRLTcs05as2FYgXvmrEu9V6lzSEZYY/lsg4gHxO92+q/pM0QmLOExtsBcCJCrddUU4A3FlZG9FM98a60hW67RzJ5DBFoj04GnWs3riUhEqQt5bMSekAhhXxymGHyB0oWS48UGCE0AQhIEW+e3/8XC/ZOFOr2cOayYiuDiA7fcHWbPEDwlo7iicgEUmWVNPYCjNVqpFOuW0bwWWY9iRnaJRhITjhJgWCEe1FlwPmuZKfsbm8CW8r7GDC6lxZtm24R4oEC31DXiQMK8am+rUFXybxXq9NABLx+F6ATkccd7HoWmVr24ypCdmcWiVwOn7/+9lOg/paMITmS6gRZIK6dyHUUN/HVgO1YZbjVBjftZvElVqE9r+eUrtrAHXwxthw7HytnIbeiEZ4hRZBTv7hEKvyQojfulqO/K7jGgwhj6q1TsEAF9wUyFQIDBlVblmFGa9mpfrP8yDeOzgjutXZ9zfDHbShwcDBCQTcbzyaK2xlLcG7pzLziR+ZAw2h+fZNjGcPZDvY56MVbO7CSgYLom6tlZDMt423jH1DQx0j+i1u9ZDO6VP2pY6UtDOqvqLeFTg2d3hse+F6O5DRBaGqkn2RolF078xZcjQkMAxuehxoJBNRWwR8XdcwNjBpffgmGU1i733HkKlvbZrJ1rcox6luaPqdJ/jGg9tjfCuJ23j/wutnjKO6fO3e4AoXPa2PRvvRHdTzDBDetgrSflhJ4fJyMOgl6NM/mEtzuk8SM4cvswMtF2ucTZmDY0CdMr1gXJWYnJEFFE1bRj9oUUBUrt+5WU4nCOHZ/GezysLPuMMZ8f6ekUg9DvYCq+CRB7iJwLEY5zoLjeJFfKYY4tcrCvk+yqgQ3m6m2VUKP3cWoBofuFVTzB6yd358DRwatM62RNQWF75uFZy47FPkQ5TxkhFz4xVlV8UzVwxM1anAgbMMfTGttbmoHf3Bea+h/Ej5yldxt7opi56V0oKYFwhDeI0DG4c1Th9It134fGnNBN1AoZmgPSsDwdJlUTsBGoZt9EBBAgjhHV528++GGpzbfi1HTRxJY2CuFBV4jO4LjkPGgdYT66CzQC8n9ycbteGOACDtUvxt9sVlMumWEwsPWv/HP/XzIX0ys/EN5BDgZIDXzO/CtaNxV2R37q8+N6iV+/QnhpiFQbTwSSKwtymB7sbs0ZPTVeI5g4ypp7drtThtL9xCsoJ8EunlkGvRaTrFa6pqdudQuVR9LsME3GjTRYwe2H1vnxgKzNbmDb+OdmUSTDjtsI4QMiQrLtzEykkP4BXVJh6A5amhMoG+9GKXyq8awlidi2hbemYsPY3pjkC5HZleBIl8qMD1/HUMICGyT56mrI5aIuWk/TKTjNX5VgHo2KGJc3lB4S2rGJkDaLwNzr8MCAZBegwKn8k/Lkldjtsgb6bgHJqAPNa3z4/XWu08qsXK3ljCsV2VRWxgNjNzTqtO0mFqGCiKIrtX+RFFAGj0k/ODyEayTu+yZ9nv3vzK3iAEHix2NLIHT8CT5JWguYqEw4fpsFIIKJ16XC+T5eoH5+8juaK9fTlFvYPGZzPopx7g2VTAvFnNjAjlq2RlPaxKCdEbsW0pcxf6Es87x48R2g+yX4+Zx61gicV90xb/BUMH1aRpWNbXjR8zv6YO3ZwQZt0YGmkjXoh2P8+3mETbQF/rgn3azkjpgCx9FNR7J9j6mHRnfwEVY1p2sTusUfu+0i3CI5GqV+cPk5ir4M3WSpx+eij3qJcsJ3Ys/xOVfpXHq0JOAu9F1fYlguA+XBlOD1iR3YTNLkVMoBw0k1t9ZVywhc2pGGmvG8Ku11uVIgmxj1kQSy5dthAXy3tpROK7fWubKadq2b87+TCMoEkceRheCkySlGPYCf9SOIl8IyAFDoixTl3J9VwafpRELpRq/XDJQiFRzDzE6teH6LDkz8mLVHRMe08Wknz/3w8Qi3dbGVqtpLpxcOwmZSWQm74V7iDj5n01SZ13fCbZwtR0ZbAZnNXmERoqSG9rpHTHDles3p5mBLBHz5U6kKLdN88m9udRK5bKL13Kxc9E8fZvViFLGxG6TrkZZTHGEoAbO520YgD1hkpAlerPMcQMT0NELa7kccBcsOe8RHn/zodGan0Vy8KH27zNoDkzSLnT6VZdDNFwgnjMT5XezmuD/CmfgNWCh3kfVrjJSSWeJJfmAfUIZZOp0unZDzuswmavGH2hpEhQkU+3W362a5B7dU6kr5KtzzTAFlKgiEUfb2kwrRTgU+v2jId4N0yktVlcWBuoc3u4TQauPK/8vXLsUXm4MRBEmm3E+l401e2MJxtR0XCTk577UETMZKaj/T6P+H10aQ5TfkLUfHqhe3K822XhJAZzJ/2qIU9+SxjeaiVCFExdwO0n5ZQqw6yhVMi7qKnJijfsAGeqMIPmRH8BgRDrsRTpm2Q9UDY16tkPCPfOt6m6KfKOWazfgWM9v742IiJr/ZOGj9Tanw/vkni5pRr1ARkC7YU7XcT+oyMLw84eVb4q+iCkWYxkwb71YBQ0rq9PWpq86UlyLTCJtl9GDHkPxzwOM4HTD9kC+rLLTYBz7csRNirdBgMTX0Aq9zYNsWg2sFMBU8v58GYrMFq3SdMysludGfWkafLz86mzE3rLBo5edONU2SKoYqdFKFZr2L0WWhg2SOqx7GqV1ihzAHBAO+jJfS5JZH3q89aQjSSXRNT6ZMiwUgQ8hETlbjEjwpK8jeXWc/kvo6o2excQBHLLzK2XAX64npYdqnS0yDH0p3frCKNbiPliMu1CRipo3sxsgawzzXXIS9wNTt5ylfLsQQRAVB/OEfGbNkHvd9XTD4rZ+lFfasrAmEOLYKemBmtzqMiNuY/zzvg99aqFBID8QJmiR5sFDIwx4efgDyPY2AVXL/q/3ZKVIFwXwUkp8khqICe3lajHoKV6RVG8jyk2dmOGDWctPql2y8Ulqhb75h70W7tbjneMfGBiP0WIMwJGuyvFL5WoI+Ax9GcMnr9FCdZGqZDWLLgJy47jEs5kFIj2P/OXEmBdRwYePYAVmSNKlxVvx6lcNOORncLHBg5frYEy3eOB1M5iIxYt0NHOFIMFwRwBbgCGW7p3TT42jkgHoDW7mYKdYnP91dGAfJ9Ryuq5uctUhd4d6PfXvXUKIk9vqEkoiAeBL6jXvdBXWF2UPDihdOqDVzNPMckO52pAFxqsXj9CMyfvSaeCRwxNKnhK9P5S1YtyJx3/CXthAXvOjMbmf5szaZjOFZy5qInecOR2hBQfa5nGekmBMCRh5dyuzgtTdaTr7qKi+6xiJOOdwlb9482hd+sGwWWZL76byqcSc8in/kq+igmqvcskmnUfL3n/xnT9Xu6eDteydbrn3jlkgTDFWxpa5vVojmabDzDHKxCqLjIu3ZIDeMDhEaBpn3+H9A/KD1SSHMlh9Yd7+/Js+vgQ8zVap/YamwJVPepmTzzD0Jd+RDUc5fCDmqfHvYseS1gMh+72hBhtTc4LWamabGJ4sVsQNGnacutj/5wrAIo7AblOfYCV6Rjs/p4UWi1Mry8OnXgFA1oBMUcGdQCS7Ax8VMxDE+JBFt+tvNRsyYs5V/I86vUNsDani6XNwlK+7FiUsrFm4TcbZJV8934Y6Zf/kNmgWm93xrTwHSDcRI2M2KOv7h3TUppdKgyzLeBUOu0HW9CH7dt2kuKU5sIQfxDWeSgBNHj9pp07y4HyTAOobyPzY8Sff9FNGmsJGrEsW2tSGOMf3gAldAdUpgfQNf8lwKKrLdw8xG5K062dMMaHZuhcjVb/6s1SqNRhpwT7ih/cMQzEpNgWf3zZcSCBbvpSNY2cBwA1KnEGKwG0FKNeVwR8dSJzkGIfV1CFyy+9dc2OsnO5sgKpxqa0jawsgZ6oGr+fLYEMtCXrP23gvQwGRi0WP2GAmCQHKeiSmE5tWBalHvqHdPQpcoTBvkIwXj8m0RFngJYwow1A0colEVtvIO8d1P/LqXxk2clWe3xgR8W4SNAIaLTGqlzbPJCrxsw66yxbR/1e0Oz6cCG+yevj/U7Fm+QnTaHPSGO+yuM5d+ngz0RzFdthR6uTSmTds1K9U/nw7n9ivPK2pWlP+C2JwHA2CajveuKU/yANcJRdHwx9xt9NnGc0qeDSsKnIVcFQE6IdM6jq8i537/Eq0ta4SIuNKJpNdDj/KGtkyd8D7vAvBVHu4vwUjp9dval5Y1mJk7D0RXFVFWQHLv2O8Zct0phUxWizGEJ5ff4609Vsv4un2mshiMAnGTmqBHzOABvkXT4WpWAsa4k57ETQCvTkGTwbAAnBFp9pDlcgYwvx7uKK7hxOExCezBr1Nqm8VP0eHYK8QMDPwK7NQgwA4964o3WQj8Sxasg+GQBU9aePsG7EYc5Q7qNkACy2id4ick7U7pqzQ1Vu2G1nF4xcHeH48gfSZjvgEu/5XTAaIxpg1DITM6VorspX7kd0R+2HDhkLmmjafpDj3gNTSUViGPEG2gmYbtq0Givt6wL7j6KtgvPfsULum0U9OaNv1Yi+TGVaQEIvSQn/OTbrElTRNW6Mg+hKwti1op3T/Ody2hWzRH/EgcJtTCmd08Fpl2qcfG1bysHbdQFtY1diJrEnqqOkWCC+TnQ/r2i+ASGvoFIBEhlArs85DqAhkFcP0drhfTWvQAzOySdSnmWdY2uisLo2QQu+jyosFXhxK33o1qtlrFu3PMRiaat36ogcW1waFrx3fi/AGbe6p4pK3HggSgtR+jPOTjiaWfwQyBGGuJR6AzqQWnA6I0sw86SveMw3t2v1Qk17xTDBi5+FFXTMmFt1ndfnT+LlZcnF814EndHL4iHMLoXDhrJDCVZOiXX90tc5fnitVSYb1dyORB068TjIt88nVfZ40H1P0sm+OdSPAZzxue4OMP9WcSnI4L3iQYSjgElbbfaSbBa6vgQ+WI471ZNtQP7JQ33IVoKQf4AVJsYoK7IWcghH6/bI25W5TZy0PUHmFoh7qqB4zIwSDTFja+HkLdfNsmlzPrgmT/LLmyX7x0506Wvu5US7dq7/kSyMKe0z32nVlLmcucXfIJrMqdNfElzQpAdQR6baQWq2FmwSlX53XzUSTkvlo5dhSXRGjmxmRz0koKtxNQZHOAOVVKcjTPBB1SVaY2zQ1AEeEXOgKkHcJ6gdNqlfgs6FkOjaqxYwpmMSOt3l0IxgwPTqurp+KsENh24EOw29yfC056+rDZ95p0rMTNxoazm7XuDOCc5q0kjfrhk2d0AllJpr+P7mnvB4sl8Vh7BsO3s0NMrTsOvgdW/YCaNSYgZldFioKj+NCEvlekULp/Zuk6hOOKD31CmRHokjHOHAy4jw5qoHMIt6WqYwYzevWNxdjEgLLXogtU+Pt1yOR2IaqHyF7qsAzTQrB4sb9FFiKdDuarDHKWDaiAEM0OkriTuTtI6uos8Zv+UDmpYQK1zsBehyaThT9UT3VQ/cLnQM06MrWoBTvTQA9PagGqVOOxOUkrJre5lTcQJp3UyWoBp7KpwAaTBRSkrcvazInWcnW+0SuqBXtfC0S3UEdaawGqWDnUhGjvNzHmgHTRfM1iNooVtA4hBPcKgts6SS3kpyBUgkgugIdC+5ioM7PCUjnu9EwOPe2qpcwiu8MIr0mICkithQU4+8dXSpplXvpCnGO79FQcriVf/I3Sw9OO7607dqh7JJrCMNeMK4wLEVkg0Ach9aTziDgh6Q+kii2iXjZsyPp8kpIzDu7CpCbORL9AGL7MoMdpd16wRSG3zs9CTgZTKhSDEHamhV1EmZur6snh2b/XiReaDjMpCmszGDGQR+Ese33811ZSlvUmCZaue6TG6iTBkk3G3CHsQogsxMEEYia/Z5ytj/kCoUNV1XAWrMQB7jVt4TMH+EXHNDFyYV/xDSXnGy+IhhsKsKCBurbxPeG62Wb45SLyNMzWX6cRf2GNw7yWNdnKEBMy/h9eIDpAm04jGqDfazhCf7c3kvJ9rNchB1NXSmeTCUbjo6lN9bTBGiaDg8i1yehTLtd2OvLEOpXv2/BDcgm2o1RMGS+66utiJJYguKLmSVViZ1Wct0QmfNzyYvgiAPtIuB35xM0NbzG33pJ1RW5QSgkFaAlrKXgMLfRFwHdzHTAvudtuC6yp8Tv/Btq0TX76lNjy1yb80O9+bEs7z+cd2v4l57L7yZkh4M1qJWUYvlxz1omzB8IRCm2JQ3TTr8v7uzQqLlx5oLKmuA98KOYFwhSmELmWR8jwNKyIyRhqUK2C98w1UnUf0SA3EnISR0BUdBhJxr71OSATrDxDNyydwPaFOyhCybXwg0jdty+BsK2wpkuYRIA11QUu5eGHwhEp+B/6/j4YtmJSjuGvvgxruN1Lg8lt3i+Qizxe0Y+gHcM2euLsOBQtsw5hXlK2KzMEdcAkQBjqKVaWeCi/9PpVN5FDOtlZisDRuHT86M94pOGQFaCo3xW4fu1ZLqm+feN3SZa6HSz2l4SEFtJEhl0fBt5jil6akfWvZHcOk/rja7EVTO5oLc32x93Kr7cEJ2UPC+A6hZYNfxJ8Xp4Z7V0Hw86H5AoxnWbBtFFVndJ7BnXPBgpCrSUeFuaSWb3xlH6qdkJzERyLHW/bx+yg1llhZTNNmoqz0OVDgaF7ePytrN6wsB4U4bYtKIzfVLYPDxfomMERAjd9qZc8j+JX9oGraNoZ7J1XgALYEhMjugHIFNFt5rrYp2wfToueUzHH+mR4J9NtH45DTXil9ccz7hi/CclIO5cxKzFyPOocDmhCCkXw6DgnlL4FutHoS+niuEsnpdtWXekAiFRN7cEUNFAVX91iCRjZLyQ0tBpIm23PxBggYGGrDAk/2pziri4nMYZSBOhbMyLWB0V7qsHAYtxqjE2EMdUsv3PS/JGHLvIfCSZFYOHF8m9QFhOugGxKV5ZIrlRimorNsOBAheZznf07DzWYxz9e0OVRnmzanZw9VX5v99XPstdiXad35+OdJChmqXwQgXDzNPuyBEZlIj3N1RuKZTibYvcE4gShcrpNa4bgIZhmfKfCULuovzA1A427h5HbTBnXCQzN3Ro5Ym9MOs0szrtqZ2FollSHnGcp7BAVp4vExzzeB+NPXJaQN/30wXtNlmK+SG9LYE+kVszPv6riUBkOis6H6f0MctOq33DZbMK8N13ZK0N/LTLn/xNGTunQbA1T5hCbpFJj0mwVr4whfIh1Xtf/cOCO34T9ajazyD9ZWLXa1rPd2bdpmllC76gRa34+H/HQtAV3RNtEISKQ8TRtXWGh0C5nFoUwEe2Ifze3pkZRaqblXNjqj7+KvbFh0YvnU90v+Ul2wPOy+aeSDUn/++i2NJLgZhPsaPyIAyEzTD88BVX2Uw1yV7X9HIzVQpnxlrozceLyrJq37vt6jWGk2X0w2R33ikngtKA1KihiGGFMcPlc3XzIq388CHrG5x/VgAVryY4ckFXXgNkg3hQlnZfYEE6EPwDPKvrClMsU/vNH3s266pkBSQjNaRl6xSCfgcFfK7r5DDUfsbjWRE9+XVPwo9YvsSresJzIY1DNa0jok/z74JnUq4pb/VDfSVV2FmiIr1HFfq5EdG5zP96f/erbdAMVXaEapOGK5iYZ+fteJ5Begzf8E/6xfJ+7zlWL5ThFlaYjekEoMK8QtUqXvtY7cBqXvo2ENKjlVFwgH7FXCR+agF6b0b284J20ZVQgl9OcMvvvIiIGEZKdbPX1dOlW5pwUotCs1KAfN7CvOXJ1CyD6CIg2bxVIiwu9am8iLP9ms3vdr1v47IpwFZSPc6yMwgozF7TXLa0NriLkRBb2xpyAdzU9YFoNEseqPlTxRaQ2MlTPjasCZtlumwpWjag06XNnw5wjTrgtpXD9+qow6uUE1ie3yrp8rezAoZczbh7jVoSMJE8T4o59iWPmKHix62xRLox03k17MztpS5bg1e1n27NMzkosbEzZI8E2iJnrcMinu7vXWQz23148mx3nv38Z/1MPm91dzeGl5yAjbIDd1NJxUyNQdNMO3RqlVfz8wh5NZL7m0MI8IylHNWsBJCXHjN6d/A1CaQU2FH3R3UoSigCzlLd+femAZqTQGj2J+zFOoxTQGa2bJ0IGNnnneDPCpyyecsQOZXCFXumfjqqGaNnS32/iWm8nYsQgn+sdAUk6G8jQWm6P88zuH9Qyr1dL90k3oPDh/tsgtdT+b4g/jgLncXym1UykkyBvjrBsRMhRAx5dqR1TEcO71Rg/VovlIj5jVZAnCtCuy5l+OAOgvSrtX862H7AQ1Mu9HWvEBDnTnIiAO/OqN1vv72AFHo9O+m8TU3skM0DBJCEbOmCeOjskFepkqAD6FZ3HF96T2maNuzE6Qfx2wBG8pnj//8VTTtawQA2OhtSzZSNWfu0ViqxUSL9F26ITJsXL5ptaJ6SXtBpc9f2CFvQSt4RURCTrYNytgEDKAUJ91MjPj+9w4k3bh2E0NEgQ7Q3nXxWfQJYUwGznJgRLhA2YNSeBHespKAmh+drem3wxGLuViY5AaptpsOxIE7HT4yCc/52ncopllf4b1Q60xfApp6npTRrYELInP4BeesVRniqhMydBSxyVqV1LQb7YWppRMmo3/CgkZIJP9dZnbzXYVKpXTGPN2m4qJPqcG8MpC+D/nMzR9SJqbOIeL4KjVgdI2X2NvwFU8pPd6ywyOjDutiDpkRrgn9wq57Rb6Pf0v2ukjdned5dFw3ehE0B9rh8dDR8sgrzoZ5Ow0dhRVw+nPEz5f1PV3qWpkbNhqhFG3MpQuirzZ3/4++1PzEul45gY5Sh+YOSmew3U4DlmULfkpnU3SWiEkfUeCWSHSoWbr9/VNfeLByP22qoqOOnS+LLnKheufsNOubdXATV19lTP5nVwc1KQrXh5089y/A/b+zAKESyCuI5zeQijzL3NNNlmLcDU4khOi7B+HQhUejzywBLTALpiqprlLfkLhfEwW/686BnytRhMM8g3XgJonbyYgToLAgMn01yLNOYOg9MOKqt7OJDQfxqVv+h/4eZjf8zIjI5vlVlxyNd/Mte+mtzqtId8KBM8yzEfOqLAcqDDAnVEfIEiZuIncWJFLrorEXelmwB/9/qJIjilNVEJ3THTzqFu6WvkLo9d2WGIHFNnsV+A1sLvFBYCKnP/QKfhBImk8Oz34yyuYZirFb8szyAmPezx06lsxsH5472squNbw0UdESNv5JyXFBCv8VxSWrJLGGYoaGWvGziFXXIPGeUAwSuDHc8Z4/7+EqFCRcOZ6pS4xDv8S6l/w96KdovxMhpqr3O9czb/F9ALQ6EQMusjeKR/+q7wvs+MRyMA0BjT2L3MZET/G0UYLtnHbKexjTeGemScb+eMxPajK2J0bGj2rUZIwEXMS9S4G425b1ePtdFbzmzW6F3wcKcLgywmkemZ0TDZg0Nt6/+5pZ2iTWZfvs1Xt9WfAZhRrLfB00brb90iVScVM9o1mzmrO+Bh8jsxaRgO5MXS8ctOL0EUxdN13UdoZP0SL6ZO5njudVYM5E+Dk6eQ+DQr+xhM82Y7ukJYDfknFvImwiiQWjoDA/apMf0gQSgGGRKlU9QpwRsPUzh7HDb2fpgsblUYaiWjIDthPbkpkXqvYeRQrGWqkFSxweeKTW+MSBUUU3JJtBQxa3ggCJGTfOhlrghdoZI6pISSCMjDLlvQlfG82236PRH+dEfz5Jy7etqtU2gtjlKXs70+0xZsyqMO9EWa56vMYnNPO2g+dUleGK8vPgrkIRMyzUr0Ix8l8S/dV5ODyyXf9Vy3MH9XEsrA53SLpXOdZtq0ZPQr+5Q51qNfkwOtXz1SQQpy1cZE4Q25feCSmrS7Ke2F9pMRQf/CIEFl4HbRcOMw/S22jy6b+yXpSt8yjliEIXobxgL7qxXrueol6ezBUD+n2Pwx+lrTRV50V4CoVQkO/0P7kqJF7sgo21LvEvaarCsnL8lsbQwRblzLLz1kpC+2OrfRUZI4tpoxEoAWj0a7P58/JfIb93X4vZ0yzMC46kKCInZQkrWgwsSR8nm782/xbjFhGvDbQ+PeQUOVCgoGvTsoVM7Z5HZlxl3u6s6TdmZRhhEt/whQTR6ieWcWYfxwtWiZ9PgkAzOcn2kCF7/8xtybvwmeFYB9FT7UYR3pPuuer79PJQRkHrmIw1em51bbpOAtb20H8mw2Ez1EWzz3K/rlI+hXdMAiwtWe7Mb56NTNcqSm4Qk7de+sF4o5fz192QKydLV7QIVmZ6UYxEELJ4sVK/3W2HD5Y3aDrBGOUdKYWW7WRe8RO9q+8yzRASNITxlhRxRx0XXHyrID9QBs+GW9swAWpJdJXIMu8YDf9doSwXBMNaezbxG/ZH3TVEwleSO74h/9JHP8OuTt4higsZq1dmUiMb6vf9lApJK7dcTkAefhaX0l7JLmqMM4CQ/gK78HVmevv5onDbMLlhAmF0c3xIQ3dT5JpTj1SQw4WtxP+V4s3cfJX+jR4PBg3Aelzrd1Z+EhjgoRAVnpks5uNxNiYSf9uwJykFcG7QtLKgChC1pQ7SLZ3e69u3CyN2aTgQbwoy8aU01J/ekUMzh+Z4GyciHEUPZdsLav7gW/ybFDMHf73G4QBPtMYFMdTV+3bsowkZrptG1IsaEiDkvj+X5nyA9Mt2BNoW+rPGVzxC4xytP1qS1tXNTOwuqDuXbTgtP9i6TgrSHn5tTqx1Ja2gjVuZGKrRBLMF7vftRTtCFBuS4L5vQXyjpY22+X5ZagjP8E5VnLtOR3cfyX3ISD0pXdWxXdfGCRhvY+SZnokLO7OQ/rWJxN2zdHRHC4r4taXmf7bpFcpV/JBz4lrCBev3SfY1xn4c1BSnXCc4Gi/DWL+q0ofwJW8Utzs7MHUJqddkvyyz0HOOYHqG6qaTB2ha/Wl7Bm+3wAic0przKDqTdVyBAl59FN0PaV8dOKVeDqL3TJj8g2ElXjK0d8xPEFxN+SYoXO3XjhBP0PtJCzT3IUlch8Q46z5r3ND3u1YK7fCYwFQUlCSGNInKhaE8aoiLYHm6hmvo3L/USr2B1lQNKA5jKWBbNVPvUlIOHgOZdwgPjtZMbFJfmfH4CydY5VeEXI5keQv6uZR9uc2trfj+o240LZ9dWlM2c6YMz6FSDWa6KN8Z+C2ISDawZjTQd7qgfbbRQzNoDdlsh7RgbBnhU6hzRt+arGdIiMgHuUn6+fod7+obaS8cyRRs9cUJfIQTtUcN0DtCJZJBRkh4J5Ig4Q7C45BqzpNItIdU2h2/V+LNiIvqYXpz6GX1Atr46wlMtvrERuRtHGUwRXnJAnIsNRvMg/+TNljL7LZJpk5/TRqn8mHZoyMnB2uw+De8X/jpkg2gT4nhQNgOiv1UgzghcOI8uTVIlmJa6dpdtZzZlkbSZcTBVqNRzQZRCu4VrqUXoe5xAfqG8QpM2CFEgtuzA/TdUROsFHTTN9ugDMS6FL1zFpjAIHtSeeu4J1J/HDmiZtWYlwBy2uljhsWSAtIWfSF2emsG2OHpIABW7OIoFn3AxL0X9M/ieua1jhFGodBuQEDaeWf3fTBoocPcA/rxdqnBxvQM1fYZRo7+qB8raNBCjPyH0XL0BMJno499V5yLJFOIvy+Bl1PiHNfli/Pnxt7MAZ3hH7xbKEftCHmBiZVThmqh2Sx6g+/Npp9dSyHUmJFjpuoZwtkBs56iOecJIPkjgMILCvrLY2wOsg6lMrl4uxue6UwjcGZ9+etV4Q8iAXuuqaQy0FVlv/Ylfw7bpOTr6cdOA5wSlR3BLzjYnjVLU8eOib3r2mZX54BiQ/EPA6OHodRI3/XU6+QDc4YOk0MjEGC2FHyDIHt/QVLanI4EzzPfEjvbJ87G4chYeu4VYhWMq2wAnaMHImwM7l4WSkmo5invEHhTxyYy7iQrkQf9GLlR0mm8V1Yv3G4fASCCWnKJwh5dfxzCMTLg5LD7InwRGj1leowlzj27OX7bM7dTEtrdktcNvKxlccndPX0apiZbQYE6wl4Cww0RirZcx0f+MpwMdoXEZgvDtOWheLt5sA709eiSGGhbckOcOXSxfmCMbdHh1FBuGPuAxfNYtIhhorSshPThyf62hgMBI1USg3YolVtygSsif/ctrRDeN1uce5wxvhdcr0QI2O5enHOCF6Jru+hQBZJIeS0y6Lc5f6a9S7KmhlCJJjEh3ckBaN3YSPtgr1B3NSdfs6bOqY8hoQEzVmbJIUbHs5sq1zje0tJGnFR+VykAB68AzRc92LKo7nhR1YgiwyrzZ2c+Zrsgx3mGJ2T0FteaDzNAKEKGyQIuqanykCzyxWJE6/9Dt+BUJfMBwV3w4xRAYg1QmyyAHXO2feAGMypzgsSjQZBcclZyqMXrI/iguI/s5pjNFSam96tj+hMWYjpzO1I0y7EjEA9GqYRy1b7xUJ6X7e3yTQgZq7dVnGCIuVJ2RdKzP1GDvV/v8wLio2/BQl00SLOf4z2XbIflxoLfeJFOMPV7uxPYnrfka44YQ2upnbtyhI/BDnfzARWummpGvqTWGy0TP1gSonOqzA8dh8W1w//PXbLnzeNaxctRcnQMYByIu/dYXsU4+MWYGYVfTzxBRk8UqS/dNhGAt7K6/k54wssaBmStE7FmLC+gEsGsEA8HhZsOqrgRixpj4gep8sVEW7LnwIZLRCzKjW9F7spqltnakW8seJhzh7A72dbNgG3s2gv5Lir/n8OsLOoyxxf1drcyk+GmGC9H0p9OroeIJ/hiNbnTVLIzthzkntKGT8g6NIzSV8baTeQ+iEkfWLdq5SmwfofTkKNCqFIiq7gYlL6Ly3QlpxrdKsRFZNR8Qfc6jaVL9zXPrPEvhGrLGvKTxC9XmP15oTSYku4tolLbu9SAma5njRKfSAQSfGhtFGFftuyCOdqOk+yVHl1uCl+c9VxjfZTSDme2pYdjJ1h9vi9SBhD++y1P6MAEm3JpZjbrDa+scJDfZmIRPgzb2XjT8LIOgaNd6B9r15BW0DxGyfhC79pCWm2HKTxOVLqRJoReTQdIdftIAtMNnyivdrNHx+aaBVUwR0m6AHjwsD9Ca3rp0Gf07HHoXcXCyJbQlRPQ1HZMva/rrYyHg5kVV11hXaeolh4c0NfoIP8INIQZAeYPHHL+fqEXKTkioDFpVfoL9l3KDDGNW7Ayu8HJ3qtN+Ry5Wf1LjYKMrrDH71nkqdKOFrjcjyR1o3+ksHQ5A67Ba2yXvS5UbcQ0z8t3jWTAMFdNzeT9vzFA97BckNubLWSXbAUFvEGppZ743rbj4f0C8mfwHMu8YyTdH2QuscbVADGp7UyTJoWcKsMFGIvreBQoBJzSyIOHyGo2UgUuKCkzUvMG6HHanQinYA3bMeKojnDMvFzqXYWB8OR/eTWDxSm8kDBcx+ll9xhbqiMpTcwuV7B+c2B4F+5fCwIDs9ekd0uRS0K6lW0KKxLZ6+BjgINRTDqmHunh5M2kLPmADzpdjpWbQz+GeAjs4K/UI6QbHYT78X9zPDZnd1AaC/6yaWVb+W498YF+uvOggVChLU9nwNbNf8reOt3o4zb6VID4Jgij0kz0NFk+WsF+JafkXaGvEXAafgcti3oImKIuCOFaPwbTu3gc9uGIDxKSIwIaLnuUcHnDRwV6HKVsVY9mDCkBgaX3v1LtCLRkKL8cds46XIOSrN5Zt8Ee8gNaGMy/75roL6skNuk1TdV6EZmGgPaTCLRwFycmnI1RgI/71v56pWQM4n9oH3dl2IKl2ekGyt0+Vl2X0VAqQJdNgqJvg4a8DQraYqJWaCIvAMpfYeUxCkt7PYqMQAed4UtyMTMw/col/lLFDfiPPCwSv+KQh9G1+4nzvf+x4SDLY63HRz6hPWV5GwtY5ew3iUbKatjGdEtZk9agbtEC0Kca9KT1i4YC6NqWOMVLXNiysySRfJKSHhihyhJ3dWjxC5P43UeaXwlW7DrCRLNfRFhMVJGJaf/ngWn3NUW5D6f9Y3rT7GudEkCXJBVPCzIirSjimuedb3qrbBG3HUIEVTC6JjmtX7ImCs9jTAa49Lijh2jnRmqgXj8PuBRhBnMadZL4MpVg/+KRs7371Y7B71gkP+fLoVyYSmSJaHeCsSCKqcpLEDR6vpnIMsy4cb8dD1TPKxs2JYba/NYMkaxnNPskvScXHTSNxY3jzJDzqFDg5bXnFuCDJ/m4VQg+OziWiF0Qbul6G6gp6bgxz+YtdebYZVdtE+dKO4MNBkQtn+DDmsaYm+ESiKAHeTaDhLPGX7kMeTRtiErVAg4q2WQKQYasMqN/zmyb8S4MOoTCyMvPNkLJZXCu2qYoyaMhulrkX+rTFE5aTASr6yjOyXIKJtGZr8M4B2Q22j/i4DBVwPowS/NFIimuwWL5tlqxGYhP0BBOOWgvlCF/yE8QzmFBiTu0FW+4vN//ztemvtPOElJYxr7Vq8ujOG8VS+d/hgg+0AVauIgZYYiChCuKyFpTQ/rakRc7R/IT6iSRWSmnEXxkWen+BPk3WINIrBhVGcUOXWLw1+eg/dLsHzTqeeGm/eQ79fZMrLDKCkcfGqwdShxuO2Gp5gpCFbnHLv3RWPx/9XwOGl3ijYwNlWZ1fBIl38diBtPLCwBAyfUZ6DGogGJUxLqGUYV0Kf+cgPyRcYx/AhX1b1RxfOmoL+El1kYu8Z48HZjUFrVketC5wzT/xnDTjYmmTOONo1nhCN+oEr1+zg/RFL5Z3kj/BLkjHDK5gYIh3sW1EL1kxOWis8ONVHGjZPr3ilw1JV1lAPxsvSN2Do2bfC4nx0ZpGxrbJyYaTjNqLozdIo4Ugomp0NNcYQNJFhooUPPpr6OVnDPfPS4pSHR5k8xaVVHjtAp5iv4tFzguolwPhwz6o9zh61ul6lBPNukCUAOkJPXCy0RtnZQr79badilHYgB4JFvaDnte4OeRZQeesJepU7JAiT9ZUieT6gRg5VrjOKagHiMTGhFNQ7htDu455aY7IrKlisc9TZlYOz1xNQP+lQzL+kdgQxpAyeIhrnOW4/Jcwxt/8AzfzGWGOeL2pw0yE1ChohzySnHsbBHqfnNVgxBAkKtET/Es0uVrdHoSP+YqhPcCmdeBR1D1z1V7sSxy00FdiOEXWjaVtnV5qIQVIGRkAhYO0GqIfKqTqh889nqIfV0CFQEMklmM9tDaLutUXSx/+x8fki/T+Dm1adyNbgevmt1d6AJhRB25yV7+wg52PJJDVOwH9h+J4CbmjkL3mqDtXRQmsptLrwZl79bpVTxUNNv5K7DIilrVgtQGkF95aNGbfvjKb5RuKJSGTRQONzQ89P8jBqclV6h9XrJ97V5qG8L4OEE6Yy9+GXkb/+xFcSQiL8N5pvGBBpVNvEpQ8WJMxdtT1b1g0PYOKuy6lG/4UhzNSOQaNQdI9G5ViVN4bJpS0xUt9PFXNuRTAGAHIGnpTk8j5V1EowdkTNSJILAs2NHadd/r02y4YLVyZ1WjhQOIYXt58prncougPnqQYexPZhPqtzV+At9QGpPMY7AGjsY0zxlz+tu56/5atRyq2IohBdr+hcRATrM0HgGDNP8cpicM8866BYp+xFwEia5ZaNtxmTQ0wRWnfGCs3Bx4QUd2eozJ+CZfOwnLLVv1x/PH+5CpWWSZ7OLlKoACnpHj4kkKzpNW95VMNfHKxEciBD2yqk6avNdJ4MOVTzGAquJSd3VWLGD4fBisyBAeoZc+hJWFHJcgZsGz01m2gbbIWFcSdTfUMlae8PfLaKcGbNAQ/k7ArupKYldQGmm9p4PKx7F8HVwymfd4mZLHNZUVhU4RT6LYOVSzYKEPIWwIC2AYyrEm24TETrb0lZ0Wz+qlJ2pFxrCxfl5Gyyr0TUjwFsvD/OJbbQtQA3nQkpgeumi/V6CCg9pt7frHMovcHok0cHHwc3rzhacul2yV5x1e4NoIAlOD9hBR2rZvVxnmF4qsh0vmDi1aQamj0b0Tiqe6WHV8YgKAAvX5Kjs7ChWAXb0Ly5wjuDG68zGIEo6PL4fXD5U6G2MTrEzQJ6zTegqUh/c3IC/Q0Zz42/Brlpgi8r7eCO8VHEyOPT4Jiie3LE0AvtzVPgG6hObDh49784JZ+58KnCXWbTfv3sA028ueTCae68KR18iTmfM+jpJUoWHIpLMIyVvkkfP4nfnEBiJ/o0juCOXx1uENHl2vpuUQkfFskXQW9V/Z6IwivH/O4WR+MCS7hzj8NAKfMd0oiifwBRAA+8XVqfbcTj5RoL34EVVmnrPYJqSm38ht4u9vbwMRnfwTkXRoMkGo1Q5vIWKaBsXTwdiIA5+PIwaejnd3HhNPesC3viHSD+pdQRmKTl1n0QIwU+W1Xe+nSHr4awQMt0btJWtzPgPtKYHq4LwVeo2jGIbv9VFEBJiMaJgHMzz1vpWKxzATm3RfXjNdTDodfeVxEwxAvCcvtTuog0WcCajqKM2CBcLNr+wuBhXI+30XeAfr3kk6H2k85m6HN7PD2+grCoPOJyHRdJiezhd4hDl74R3bOcrOvK5YWz0qg0hQpUsLiKYvIaAkeos1G15NUkIIfPYbVIDO53f202Ug2yANQIT+rf6TgiB3rlsFsChPb4w7GGsawbD9g1cI5DFySsxfwWoC2bHjRAe03srhKnrD5lHm8FB4fUYuZwEgaWpAA1Vynl2ht0Z279swRvRt3fLguArG/BYAuL3fTtYQAbFj+g9bRUN3jd/RM7Ydneui8UCH3W6rH2WEAIypCbN7+neOQ9gRZpLHDZW2pM/++Yu6q9GN2CBErib7j+tEF+VeXWR2JE9t47k1aALcX5BlGCIdzLQeDsax/QmxJfIwb1u5KQrJF8e/QyCzLQWSgc7ZUcvZbKzO9Sf88hth5iGRH5Gdtl5tg2+4KUS5HEUidxAz5SpDTiV4LT3dleohtkcGrt0PgSmgi19ZMp2s0/fpVow2oEWKo0rUTmvOC7y5hWE1KJMNS2pSvhO8gZUtGWnBwkGF6wQoAaSIGOoviMQzXF4UWuo1NOSJbHyDqIaWuDqK9cGDJimbvs7XzwHeVNgNFC38FXiec5DBKLPpmwAa/sVq9LgI1FRqctafhCAtCvqF3z0nMn410/muPFxcz5LKCum2cxddXjV+JdhwXOP9f4drZI3PjrUlumWZACHcyyd894waaAl0dsB+tIaElKLIaubnfMzFLdrew9JWUt2Arg6RCGO4GRD97uBEbSl4RGrImUNaxG2AlEqTk32+CNq1VsE0N3oBJ8hfuNfRCYl5yeyEoWnpXYRIGozMKozQEfVeEVe+I0fD1D5QiUaW3W6co0bM3tIzWtHKOc12jGRhdR0ndHEP2mYY3fYui0LwFB7lqak9LBanddLma4ixH6xFuU+rLSZcylo5AERyHgGGvimr2H6udfEi0pSD76PWcUmnDl+AjG1QBHSyP8xX0kW6MfcqyKCPiA99shsrEiAOFKL1k5/3x+2UIjL9atBWQlxWHELAU5N/LjBVudu3TGex2+WMYiJ7GGgNZnHSffglZxsb1avkYXp4qqhccIe3j2Sqg+C0FE7hPO/tpD4BYW9MRjFbSKPAxfhm3Kd9TPGjURmVYNDCx4mSAjvaDWivYERd1QxatvBTTSbzWz3RoPISOigPR1Suqe/IrtShz7hl632xeRb3A7oKFthZH8oX9ocb/u5JKaT5koImbx3rZrFH/z0YAltbi5BsTQa2Eddi7AzYWy5zBRddsSZsOa/Md62mvzl5qOrufifFbqhIKPDYq1oNMiLD6JBOHQqRRcEOvtyZF4AnRpnyzgYgo0YqL82YakPmuvmGa+I4uRj3z4oCBmCFRuU68Ya9cctsV3PSfsJc/lATHIqvk9ViZgLG195HGQx1k1fkFvTnbzxbUnAERX9hNKyMHfUiOLGy5BvjZyLm2o6FWcPgj/hq+dc+6fXik7/xOVWTaNlOXvhoxTHm9oVs1RvYizr4XBJPwdpN/mjDncxMA6nD/JhPCL57KzJoprb+pzTRf3EvpRJaH+kR8bfJ+m11CBtbvpGlrhdqIhz+kGxz+kzEI8FEsV+X4Ng1ug2CSJJglZTr5jAantpqF/7drcirjFUbNOm8oSQK443hEq//+Ve9NG++JEMyxSOdz0aJ1mvJGGqWpLIqQmnDPbI01n605/KCW/Vzv2uA5JNN67BtpjmUeW7gS4q9rzppOr+xoaQGo0QAwCofx3E++88ZTn8QeunjFwaAS4L/2U6230lBBkFaWu6gDBcWw3ivJyxa2ZDjZvAqdQkiiVav0+PnT5EdVNaB9asRLinhfI88UWucd1L3CYepF/NV3GeT99Zg4y9Q2eBU9yDYljl6lUwUCiJkq2fRjy1zQqEvQxE1b9FySboZ5W/J+XfBfrXxVLR6XYMoN7SshAH/F+XfN4N84T+S0x4XtpRJEyiKZ5ewLXWkbxpMfRiZsK/RVb9LHiVHHbPGiQfpWQOhDzIw6jaXn+wDtVzemZg6bTkqdqUXHqSmCAw9IPruShnyFlWiynsYV39OlOoXOlOM4CujZllhc6mEsAu1Fs/nA2M3I2WFyECFyQnAwZsyZZoV/O94S1iIT8pGxv4u2DLkpCyxJ4mIGX5Svx2vaOrc03P4bE48MZghqKlog4+QqhNJto5nYg+DmyZRv0NSrBIgyXFxrdiWr0lDbtjObZbcDSn878D/AXAXjrbFHAkxRRZuX404bM/DUm5uLVhIfokEuykFZ4rH0YfB0LaMVePW8cWdZDTuWabhgb9sMSAThg6FT/Js0qqhtHZvkZqYBswweD+xA5pjZqs41YIkf98swxqgcQxCpBRQZJhGDJJrtZ147c1WQQ2We8dVXsw54pFMe8OQpKVU+uEq6Cyw/2s5DFqIzRVqHELgMrAYsSK2wwsoPn9m8RxA5vfs/RrTsrjWdU5QDrv0KFouWIf/7Xww+xCCzBooX04TKEriL0d9GvNQUxYEKBwY8GmcoY/GHSxciSzDXguSOt9efOcyIgmgcccS8h9xXQhvpAsn+ttWJJlGwah17YmneKMnHDa/1VqCiVgt+zMQMra52+ApvnGLOAGRWoCddHnsNJnzMDfgodL/x3TxzrX+TqsOTve+X+e8Qp2ecbWdY5ozTKQvk3Ov1AIAb9UsTDM/K3Ej1GaOzDeBNLO8i50K5MmZbSPAwjzA3W18Er9bdLPe7M9s+vSQF2lU40WojuXsFuD1ZLat+nJuwZpLA+4uQuTsr6+/jPEmVpkm2ftfN7G5Cy9YhnC+YupTpigDwNZP9n3FkwwGTnvCvVAG4ozA/sWMFle0LUUIrg+GeFHBp+dsAsvFYp0PtF713g1H51e/e3AZK4eBRDqjiFTzUGJHEV5J82pV247pPLogFlbcw/xnER9zyXyxlZjaZL+nDx9X2qsHetxNPo5uXzjXI+Q1GuiN0bIH/HvXpUvuDj7scE7egQKXG1yRs9N8WjfmlpOfZBcKWVF0uAjBdkWeQM7XqAxnPrTJadfFs88tsEGdmemtn0SIhWSKeAP1TosZZJJYlWdKOXfiiObP//eswXXBha30/z5o1LHWf4XFuRMre+/486xrZS2JWvK4PHOFjWw8TPK0rLAzuax3xIBmGQ4U8AEZ7iFKfJKI9yTvDdO4MG14h7ZvezzpxqGLQU6qbqSpuYAzyB7tJR5dgzaP9ayOJU0fWyysIvF50bUCMDicQqmoAE6zU5m4qVGBq5DSnx7qUcmbwgRpbI9/6cQrhih+IzacjLO3nxknKW/StkA7Ia2NZeLOLXoTsE+/zGil4d0Fd0QPF1Kkcs7p1iCG6KNW6yi4SwnxlX6kFPFwytns00x1JvrYJ1hQH1CQnkGxBwD2tKpyJB27+VAsj1XBTQNqqObjDWTcQr3aH7JN8LEI2X8Pk+HK5cjr6Dssd+2dAHT63eQ+QPNzNRfM9Kss7wsWyzOEj8bW55DT850YPSDoWvaYJ87ktcX/kaa//VZFAYW6ZB+oVMYuBfis+VmngOqC3bHXfEBZVC6jMvkBRlBlgGaqvz5pjulj9Nkp7SA+9kLbLHICn1NsWUGQXrJaTIZZSNYCgBK6mj3CqXHcD++OCrDyMtFuW6jPjwezEFIOLJrkWA/IhjfbtTL9x7gPmj1ZB03Bnc3ObY321gLeZorj7OnSSbOCjkTIi5rR+TmK+wY7HbGjR1xZG1U9nS8rWXwcuzvD2NqbKpk5XIiSItfyFmcA+UwixN2nu9PzBEGeBC41W2a399yZ2mDTf2fGp9DaiQfAQ0WW/VMl5CkGDLYAJLhsS5COvGQ9wZEr80N0GF3x4k+6BbD31nCXjol7OtRATgTPMZ8UcTbXKt4q3OpcggK/QJpC5SyW5IgN9k2qmmIEqdapCRg3yr37GUkzjm7oqXXokxUlxFhLktUVuuYqPEtA1ifY+gjXkXwGxG1k/EsWT+OQdoPXNL6tMgzCjqYUmglnHXnRbhGNR0HUttphJTJmMtJriFnLjO7DPbkoqfSxF/cixkNf8EZ1ckrycZJ+hqnvNN+DNl+HYwS02k3RnrUbKyaE0WekDHfB3e8IVMYHrjy8ZlZ7bvmkFmBswbkG2pwQ4j0dHkpBX8H5GAR5JNIpvDba4uSyxh17/PUFMEsx5Xb0/iuEtlytd53brzDCQCu+E97XPok36Lp0OPqF6EQId/e0h1LRHWupUj5bP2Yj1KI9JwKA5SxOQOr5SiSLb2YhAleoH2U3tRlKixcG7Lxbr0bhlbSBhmkHoqrabSm7ek31dbsdGRJ4QDz4ZfQkuXDNXxhn13CEfU85wJNQENbpL4vaxbSuWhqmMbRBJCQweFSrjGKbTQT/WigHXsuKCgs02DB95mHEpDqNsyhgvu0rTnoi+J7kjK0UDPWEPeMhUbur60CjQqDCvjWJmU6mcCFyjVVgPnIAVGxlF7h+9FGw1I9JOtrKyklI0cwW6iQXzW1xGHSg40O1Vh35NTrKc78i03MHr/gRUN7oal7pDviYozL5jf/fgo4zm/2fVtqwzlLozP8mM51g8zbiYzO1V5AP9nUFA8m4sTyoHnC4oOhjb99R3U5jiTnO+7xlqwjK80b5NL8PG+pVb+2BlH1DM+Gn2H2mAqBafO6CzHhxQAYuppcsCE8OrPyfKL5JVBII+PfBwqQgoZ8i+cgJ6BuCvj1CbuKDb0551IJDFsYS0o5s/ATi+8PewwtRQzKk9tltxhwvfpDYGNCADa0HMF3G8RB/RMNM8NMLFLxeHZCCBITDIARPB3bXarT83OYBnkYBJ3XqjdeMACqn85pzivR6Aj26pZYjt8abd474jNEVwJaBg03LBjbQ1uAqilHPDx3FB+pfPF6GrThURYwnfscHgUW6N4yaoONBanSbTiczY+9YTtlPPRpP6l28jzDkhuPOUoWydAFIqm5mZBSS+lljOrGo90SctJt2xXDjRSU9eIJLQT9avm6vFFS784VwyJ8UlfTeN/GkxuGPPFEzM8kv4AqyNDcLCzJrLf4BzHdBdJ1gaSAght+hyOi2obwGslpynxbBTXFuVjB4GLr5uKErf55Ac8CR1sppW8yGGfgmzszdEtvr2J33J5kzL4Ftx+Cq52zXAfiUIUC9LBKZyHRWaPrm8huR+m4vEOoYugvY7mjMV68i/4/+L6tFqxH5kAHIe+zG2b96IG4Vwq9GxXC1gj1TyOJ79mvdCR2VuZGkEwVLh8xzsmT6FEXG3cQmXTVqXeq4t66RYgFoYYLQmE5za+nsX9fqPiUwsTRUNGBy967ApgP2uRGpxZdH0T1OKB+QdcKmJ0KQUw9xwvNSTg/x320F834OVsHCJiEq8/XApbyL3Oaqp/DbuUE3xcC2SXvi3Xgk4ht+dL4CCOK63Iga2Lx2g2oTzvfSqLVMCqUgDkh10fWXycmJAziff0V+uEr/DpF9Mem3ecPhrhpL8sFdX5CE79jqwtJRmjp0kVNAqliLvtFV4/Xh66Aow8uH4zwMMRBv7Vj378ApUgMAiWi/m4sXgBppz6fNK6xYr18bCOCpW6bsFBdECVfxrppOslrbUfvtJIYt7/x9QejnCVzp3JyqEN3LahLlAdJxNMmIAfy+TJ5F7VNkYIUJ9nlYRZlsNNF1AK2winHnsHTsgberPpnaXwaQcs7odUPPRUoqk/Hxku7Md2tWQc1Fd7Xczi7awWRvESQLuqNVymvCpLmSzwU601AT4pPUi8DiisshZybuZrleo8lbC8Q8z0NKG1NcGEeCSBp47fHhsbVtgrMVBLk/eoF/RrGfHv0BmxUF81q/xbbl9ZLxZztK12QOUqePweCAuBNlw02Wm5e52yncDBpxZeWDX1WtyOTnluAoa73DUYSPDynY94ixbVaicR7TcIjnHIDokrKyivednALnrXeCKMhCosD17seTqGVXdZR4pdGkXXKbaAfSmynIPB53Bdv+3bdNFVlzO6KWMG+vKLqxb0g5thJQb5wETdkjFGweioAhtTs1gNTqX4JsJhJQ/jwLDqP8q2VZmrJDunA0YdJa3c+7LBkK2g5vMps09Dr3de0N1asAcvKFA0mCqlw+RHSUo/o5NnccfsTbK/mWfeOzS7Gsmx+RV0+RKJzOISKsIvBS6Nf8gvUKsu2EghNFs8wUNAYRygRYBgyJ81hTMzE7ugznNWnA7ffwhiX5I8m5a/7FUrNlfkW5G+1EO7+2uGx4DNwDMpkyeZ1RjpW9u2TcOZSDh0E/b2/kESc9QCF5spmBjr2Eyw6S0RwWeYep7WKGOSfABMF0jugujQ0C7nfM3zV+3QUocEi5c5Ck44MBFTxMgpJL+anxa1jeI7Kx4rUFSx2VU1J3n1c4z4wNs2FWCgGVb6y7v3xb+lu7w2PG9u+UVAWlaP4OIgGZYDFsRAdikSF6zUj6QZ+qYUMk9ryEMZjNt2iPo5uj2md1oDMJQa0Ds49MolnA9Z6LuZPtZzCMWxd7oj+LW5fJpsK/PiuDURnnNee0BsCjLzYKuJkA7n+/hDMP8Mid1bK9PHhlVl8TJoiVUq0hjVxeRgdaCDDWeXLsv1a3vRyQKuB9t3bI4BefZE8KWFxNkbk++w5P2IXlNmr71w3esxj8WjX2UrpwCLKGoUXTlqCcpTXPLvfu0mbTqDfa8Ddt3KYCbh0yhlsWJR0lOlOdeL6nD+0Fng9GtpVhw+5dbHZaf+1kKKUXjQmRWmvtBCR0us1OQmdwi1nJ52H2ynUs7/oVyqn9MmsNGGrLPbLKYJedGz+O9+8migiVYWaL/ncP8nJy/8WHEmguW1Ae8vZVSWVWFZk/FR5hgEjNWIBb3XTsHsb+7XuE83zl7ctVJlKWwlbS+IzDnIGwzX0ISoT3P07WD+JxNho3YEKLL5NsybbaWUIWhVnbSSVN8/e6Nuu7vOrH8Ap65RhPnHCDCRavn9t1MKe15M7sfQXrqdL0F4fBOc/as4Tvc+mAV9DQWNSwUjJgLJMFSp7UNXaiLuJIrUQVoqCzu2xH9DYlJ+coFvFCkP4DWSHXoWS/VK9cv22Ybfnmmud7/fMjwnTQ2NnZ/d7xu3l/QU+kftVYW5cv/BAfdNmZUB889g+tU3C/kHWr/q7jZwJUarJSB72G9ECABtpB8rN0I/wW8mLrFYzX4BhXBqrd3YunI92jPBg93w9UWHmQErT9wAPPJ07UcNNRuylwPSYZ+cidKn6qNeCNs8thZ+7ukE15daJiHo9Ea4FR/mDYnSZJovRvjr/XyWtbBXqwnvSguopjBI9AAjOf4mC6UesDG05mqW/+eblK6d2h5VxSooeubG/cpVc06lsuM5QQcUz//BgMXxNeDvjirm40DbIrc/uxu9uHsrOgINq5EA2jMljSIyWUAcu3AOi63CFfKz7eASPP1+SO/AU+gO4wuhiuTLBCIa7O8LWuAza9dpKInP+UiqJox8s//Aq6tMCA5fr8fGbeC/bmE2FNbi8aFcRojAY8IsD6P6jzRusz+DeNVbKj1UXkP3IexKXAAdRm2RYiWlCaULNciKCf6yWzakTPIakGlqbv3DHzg9gD7ceXz7uthQ1cxll7N+JySol7NF/jWEoUkp1ud/7qroAE9/DR4K0sZZp4qpJnKgfBnXvABlJxymbKcthJUQ7GXLCxKRkd1gbzngYHsyMolQYUtP8vT7eEKGd3NySp10DZFv00p0G4w3K48vTGsTxZsc4U23I3KoHHRpS9eq4tJjZ2w6+Fsbj7K0v1aJ5Y6fWGTDUm694LLdIhER1Vbg8FmaK5CJud9aptSQ36vS1l+q1pMbBRO7bDlXrb+CJZIuHjz5wUmnvK8nhKFYqLpEk9fxKpGkMSlUpyWIAvS9l52ybCJ0GgD3tmB2wKB0LIgYf4QYLkwok0ZrB6jZkl8C0zzoaDev17cjgVp/1T4rZ+ruiGPPcj6aigEVOLrC99skEBd2SgdaAyZKCx98J4HeMx3kuzoxYpKGOuQWPWBHucbp+Kd1T7AtjzpV/M+gDZrsvqaY0DQt9YLqWLm7jYWwgpyH1M6XmxHTQ3qLz53LrjCx1qdi35YmyhCkjGFhAvJAseejVcsdpcpG6cBSPH8b1VzZC7G/63Q+gx59C36HYTDnc1Q/0qN6UgnYVtVsdG5pDfP9au3qgJfu6Ab2z+PJ40o1Ur4e4bWSF+H0b07wBfjnf06C7ZZvTLEzddkO1hus5d55zVMgMoKM8/E83bafzpjinNR1Q4NSqzlqvycIUSvoBvvsuQ1GknAz0rht6cGV9rHgPoiiYddYNmFxtbROQ0M1BxzwYoLxE6U9w0Wb2RQuvhXlYFZaaEttCpfimSgy6ZPcgOBR5cc1hs3H0kiJGpVrgVYH4Ohdxf2PSMn+EgSCtRq96TGgiYoapaATaXtBmoIxYbyQfDxBK9IIC+740Gi50887HxYMSQmIGIYfydqd1n+b57VBDBalFb2L7IYNUaJ2SFJvquvLoE1SSA0Jv/Ben6p8+CXSXjVdVxh4016Dvo1MJcH5zt0/YJx7gSaY49eP6Cv5rhWzhe6mAiDKHhMGDxw5dvzMK6TrHUvdyQjoBowFfckIcse7TpxetTBUXis2oJW+qzd36MAA9LlEk5qQoJRP82ojE6aohn8wQYrGehe95r3EyQmWZ5VboKryFqG1sx1+edujyBGSraRXUEDde2EZ8FrieKURAgd3E1pKUrCcgIpafNDdIJS3CwMYsO9b+TwE3/Vb63e58qtt9rqvU+HVWa+gQ1GYf0CH4EDp9Zcirv8zDpcrQiD8SuC1qkltcJjrb2NWatO/Cet3Xw0cNF0V98aoW5S9x8t6doqqVdVnvFYAEpUN5jtDuoFvOySIBmvnOYIErQESHJn/p+RpWUd6k3GWcI6m/nWfTG5IeLfCxS1qO/XhXO0Mg1UiNUQRfOx1zm9KEt9c7cv0Qkd2/5ZcjzIqEQA7XBkg2BKPBtHcopQ07ZfHfmFvzh2s1IbbQ59qUbBVtAN+qbMtUYT36G0P6nVHvCjh1clPGLGBJ1bUFZ/3LB5dSjdNEwASmBfHgO/xT0SSRLmUVm6GFB/wNYybczkG4/hgIkAo2VMD3m/2YOIHFwaxL+nTCZ0xLvXJuK/uoTpGcj1utLPenUTiGOKxFGemDVSqV4qrJTFcqBAMtP3xxBCd2VAbJMxqWNj2mVVGmQismOcIOHxOzKK2q/fBcsra0s3Ap59n1urvggsWUjbIOn62O7dm17ARSBwcQe5mZ4rf0P8BhhbwsG7uZ90S+PawMHA1A7WLRT1dyBnFgyySQmASSXV71/5qoarghhUb2yy/JPzAlEjSWRqsRU4a0lRQfYIIKpfHO2VdNRhMQwKfRs7hiL8e9kCRsOFOtLgWcGmjf8hmA46KpoVs/QDG+Ts1OVaPDoJckeNy2Ni/Ljf/ZSNsycBWgmQrcKq1PCI9A5amldX4ULHD4WdAAWdQHlZPKgTlF2YX3ywSDx7fm80lwUH045jcRZxfwpEs1EyfTRuTFlTvshVKrJ0kwJVOmLwyufnpWkfFEWroVazN39Gh5lKRdXkWaVHSnQoaAf3/J58pHXwvNa+B12fJ/XtRNAAB0LuCqFmAF0dlkxY86kt/L6bwr1e+SIJC6fpTHtOoPlnQrWQQRtAqromY9vh1znIbqMfOzm7aJ1ebxJxE+CREHUsR7NqIK3aM1By1fgxTsD/GmhkYB6c4QN2NxfWaK2HrYsKpUrNRbjsnBZwW3UFNPVNH9D9z6qLIerv8EIWv3qI0ruQVaJHf5ucMRz2W/qay2SQtitC+P4RLNhQ1EWAXOxZidGIbm/86sYd4+6NBM3iYHgSpFhhF5amYMkUvGeDA7qk4zu3nRm0SD814fCnF09j6stXXnq5WHhvMY5b2eJjNLx10PUWVVmCqBVtpVPc/0vXvB7aesR+pRG8BRksdjarILAe+lZHa1E+3Y5sOSd08cWbSJzwkq4Up6weKGgmt7S4WJTWn/OtaiYpXJqgVJ0mVRgiUqF4y/OZQNVRd1OW7lsSVEya7K/HmbvzKpnDHivnTGTUmoIwzflTYE3MrjkXHqYNAPFAH31u6EGdIkuC6pYy5i0WQ26FCjpT3ojOfB5xtql7dHyWrg3SdpvLWD/ZXsywuRHuT09RTPxkhyR4dbal7GO6CQxOvu7SxI5/K0iYOJ8sHlRt6i1bZCzgkMgdY3xV/w3qUAqTwpiyny0VOwWxXE7fS/laUa1u/aWJGjYrqdPWShgPwsvxRUBjH2FTumsxlhGmw4JbQBR6ZhvyEECm3nmBHeOby+TdCLr2SF0BLEb0NhUt6T2toqHgtVwDLHugsLWy7Z2uiux2YZSsuerJNdBAXximligFxxQGh09tRYNRajDB2FoJB6BSWz2FWV95FxLZTvGRvUqcdu0CvMekleHjFtrxOOyQlaOXSCT97n+fUDLdFGjDJia9NA+JuWtGGKxRyEwr31Xy/WgXcZYnxgIRxgb8SDADcNjMj+bOtv9st6mqVZn5Gn05dpFjRGFMfJqvF09XSTQdAY6GfztrnwApx/AZVrD1kO5pkHkuvkh1ZaVsge3RKUmpEJkd3nCtJHpCx8YRt28D4Ku3rjZRYHYgb/a1Jz5AUT04I+ZRB2j1hCLx9lf2TSLodqWcBe9njPjYOK/oIE9/nN9/f4+aTMyW+Ggef8DGU+jcwjOCuozeZtPNu24GvrbCwV7PobJsmIDte1bZ1E8eAcsLktao+FGVkm2eJwvQNI9sdNum6zvItPgguc9w7tH0CL+NKRxYhFgjLVWORFCPfXdwgBtFqAxb7NU6Mbt1knBl1ghncxwVP6U4KfeA5ScpK/O11Qf1OSDU+P0LBo6iqRcvXUsTXuvnhtzJo8sus1syNGZ6H+qpi805Q+bcVmj5ZEdbT+EVj9fO4cMlevYtdZsu2AdbTcAQr9HjGp0e/gHMGtd9QtzUVABnQbuiejYFTg/YjnhsPAve/YUGbZOKxvLLOfNuWmukBWgimfXZCjBkUFVQUrEdP3IbLRzt1SsN4HMx+CuYnjRxlHlyxUl5pBGBYii5qCa2IhS5cPMhtlzZdwI7enQLHszdVXfCa0lQ2ioCJmI7QwZ8cv4xR0wEune3DOx7XvHFWS+XSsP0VkSAuUm6GtLab7MYwM2OwxrJr6sLB1gEmFgtpL6iQy2QqJnwKAnOLorNMLl9JgXPIBY/Yz4Zu+wJ7oe7htrUxhjadaLwoHbWPDeeK2FuBInqpoYkKvUqfSCKzROH91UUPQ4R+cCzzhK31hvtIQqP2X1PZGA2+8t/inFdlgW/0XwLClNO1ZZdZ4/88pkjtoursOZ1Wm0ucSuMjHsEWjsMuDUfYr/oYi8NVcdexMHbduuD6HuhP24Jo+n7A76jIOHwdPJsXhalmGoOxDnIe+MjkI9nUm6jqU75UHSe9CsmXoy9pGCcmirBbjndS2LOT5BSHXUL6otB94s1u6qL89wt3asbkXDw/OZXACCe7fdf5l7/wy/Lh6hmrak5ISmBR9gBFrpkaDwFxzcZq1ivhT1TQYqr2vkxkQ6C2QlaKK0iaN9VKLi1A7RyNIFOxWWrDgO22zq4HzXqu0V0lu5SkJ8ndqTgK54b+ufhUKaxBm1v4PTVL/q4FsO7nAMD5ssAnYL1Py69GBqHfyjqrOSqQnvldb9qxihfl3qv3TNXL7R3N72RYVdRd4DO8zAUnHP67uM8fZsrtmMEAJj3igjj8yfH/ynXsMmnTMQ3ufm+lS3XQRjDFR3csGfHizODZ7zRiLYNEIPKbHnMoifZU2UD506STh3iFyjVYF2gFBRNxT0HVcHr8ZBMpIVzpN7FvGpqL8DNagPKbRgULA6GZwGKA7+SNX3pHLPRf0+Yy9wuvkWoUVTWAOgsh5piWh1EsiRBYE/CbFG3Os7cGkaopkj4ojWSZvB6CeSilWgwZXxxYce7mJ9TuTH1bvvHVPGe/2HaHYUSFf2fMGU67vCS9xz84JeNAAsYZTdsVCyFISuT4aP9YVc7KAOQ6b11FAbsbwP9tqjkLXZOBO3aJHRUnIQ9DqzJDLA7+MnXP6cK0OPP6dZpyD/cnGh1XkFykdgb8GwHt/8/NUiSbn/xyspsLC3BeXP1tdmhAsrmD60W7wpzrJejTX0EmC2mUOh1473CE6ev08i8lKiacEnhufjJY0HM+h8JtM+FxCwanmWxUcOxXujoxcheny+VRHC49MaDonadMp84ugN/an9YhhJp9BFAQS0LYwsFQU/TZwEWHRNhyu1Ji0RtJWlNuN+ClZe96mpE0kNnBzAsUzwN1pmTcaLonnk8cDFeOCznEbOUGQZf8F4J78LDmlN6+GUUfAai8EuvUNY/605OjmC6bYUNy/PshPubghdDxrA1ZhZ5Db34lXyI2xG43Vgn3dUBa0x7gXpAvxiz9VpgH5471b+K1wTMZ/bn9q/+pcRMftGej4vjlhGqi3OHiXxl7ZPtv1wYg6BKzbCJtU5vSGhr2pmDOjrhuBqLPv7Iugn5e4kuMRbcowVMbcaGG6Z6tqo4CrfgW7+mjAzct6o2OZm8vwRzX4f4QlHsL+jPMAEGqk9sgu78to6Ad1QVTVRL/3MCYyBGKfzBnFeHqM9xre/zcEx1eV0Aqr8otj7CmTgKRZdqCT2rUGa//X9bArwa5lgKNJmm4GUMUZFNpbHRcWUxwPu1XjXqCcvPvd4XJ+pLxKty1KYv5HX8lyPIGuIfyY0X+Gtp1d+RiSoxVESM1uperkRELk5wkNy2zDAMYlgZroix0ECQmxCxeDcnWqYjwQFGJrjR/rGQmhRtFRDs61ACXYl93wAKj8OLnhitCyAJdK4Sdvx/bzrFRE3AWByeSUQ+DSI9YMJt8L/mJOyamJU86qstiKk69bvF2ucI/7yDRCC0ujGS/cl6RvywIgzCKBsH50xJQI+rvzeR2o9mWpvIrfY83EQKHqKl9nPzAiSWgdbkFA1W9tIPGNesFpoBLLDw4mtTY9YeRMWm3q9A8GcdX1g7vqK2bCX6oSuXBE6Zm8suW1MNNpK5CZprlYcl6gdwsU9jCvVY117topD86SM9OIHTcZhDuxt0LUAEiIT+W+LfFIiTmNXX/8RZXwIlKVSTYA31Ot2Xa48yhyo1/aHT8c/ms4M5K6ekandAB2uWcXvBaMdlvfilXlYnLgw2kHboRv/LdKty3a5g++6udQDwmguC1WQ23C7Or81b2smjCYAmyJkoaLPId0wOsWmCbdYH/2ANDUph4AV42ojCIjyQB4db1gxRPKa95mexR4zZjiowyLQN/YS7wMdkgOhqhu5fPmT4yoaGE2PO996SQ7EqRvoeH27qXbmfhnZESRTzvLtmufV1Cw7UZxaxZIhwfVW/NikyJuu4Wy5SkEOaaOvs10lOGJtchAAyNptN10nXevKdxiM9nB4ZFAHodjhgWq7M0p5dYo1BPeVSWCbtY4DEWv5R2n2DbhAzoz7ytSGbN3m93zPRNJobkqBOJUwDsPaLltbZXGRQojWY35m+YFgdNODgAeV3+jeEMrH9OnvtxGCMTqEyco9rEbhFYQdZZSqv/KDDvMSOR7VBNZo6zlidvODG1jI+1oIfRfFnlzRiqnOCYqptWOySqGWhhCAax+7n088LnTA+JXNwWc4HACWX9pgDECTTL0GZVbTybD/jXIZ6qtw38Q/8rFKkHJ2C8DfUgzjNZ5jcnzH48rw8qaZ3iUQGLet3/3PLive8hgZETbSWvYLydrb5zJN88rMvtOqCM4Elm1FQ4BrECJ6wyqSpvqUyEewUSG7Knr81IU489ZCK8WjLTs81/rs7Kr8jcz3h81GRQr/R0PQn+EV4Pbyl5Hw3dByiVadKI+X6MBwFs8gCRO7If5hsG/Be1/VFRQiw9xY91lIBG3Yg/ssBRsffmjDljDXfDQrpYfaw1YX/mVduUqRqs5JuxEAGwBMA+248WvxxK1QyDrH2chufCmH1f9C7YzRA6YuZzGuPwjFU7mWJ7fKofUhlQl+G1mvCkRIaF+EUJfeiBEjTzsW53tqvbWnlTN2qvX4Bt8up7uhsz55g2fkyrbncaTcpOHIy/uEO/KkeaA6O99X93XgVcJS5qXkyLarx2jTBO6R6GgtaD92znbXFhiMS1jm/7N2ZYdMz75ilGgZjN/GIeg4r902M1HE4LUdfJHWDemmwqTQbmS873TCWkSJk9c9glvTNFSZgDQoziUtW2tO5HS1DBYkNgtu7juACPkV5p+w4GRtwI39ZkhO40l4B9mTAFxmomWoqVFGPHOPZ2UyJnsyo6DFE3ExD8EHaXb3Yqm2DvqYaJv3acY8ko2hgIFqiYIzgVoDYU4C+iJTW/wda4nFvxXuyoTmIuu2BAUzCoBLyo0yzvYvx3xREWRvZPmncYsm4Pfdp/Wf80gS+zOqC4Uw/bGZZQIUyHldSoSz3hScqXs2eGeilTeZLeud77UKL7JeeoxK6hxCfDYoJIhnNSIHkCxPvtKN9dGHOzoZqP183oYrZAyflsg4vGLXxa7J9/GE/NXw/RX55mnngG/WYXSwsy2NJBc4EmazqVCjHibjbYmIbTYHZm9hZZKh6l9abXRPoqkRLlbZy6I3g+mcqSNkQpyYmZGVblr7g1NQ/PhX4W3lU1IfETrG4h58IRu91veXRVPW8q4nnLyXoeUVh4sx4LA3QzOtNxXrX1cly7H2twfuh9dyBaS6hno++tWdEK135/BOkhjhC4h87i8sJj/wc23VXu5Xb84al63ZsQ/05odrloaGH0R/SnVza9t0LDGdSXU5xycIy7HFJb5ww8uRXmbjJKn/hrvuxH9QN8MP/r+4fBdv2W9Vhu8wnsTFqwsmNUOMx864mlr1NP1WkS7y+AgIXpZzipzN5L6ma4w03uKk8unyulD+Khu13PvxjKZOiNujJrvwuB+UM7A8clW4neAr52ZmS0K3cfbGCwsZqvowC2Z6n0SU4SJTBY2qPLtX00rqLeWqGqYl0+naC1KYOJxx40FYMvBjTQ4EPk4cpstlHg60Y5kIvH6/DvxQdfU4Rgr38wintlzKI9ft9W7GDxNqf4UiaJ4Ke8cOSNrt55EFic03+on76IRjQaxtj0G22cxHZ/W9hKAvC+DGbb2trfsjPkxKGInqhe3KtjLq/2p+GKrInO7Jg0UT9eR+0nJgjDBHWaqjljIg29x2AdAEc/o9raehwVTFZ6Mn7/UAnB3ZgVYc2JJoIliQN+w6Yewob+Hy4wkI+joZN4ewTJZlMHNskiDnvqIU6pz4rATabISPjStBuRjuvbbU+U4/rEtbnkywJ5EwZbWOMU/Pls9eMfFWSftCk2umLg8P14yjctu7pP2jvtnmzf8Hocbxy0YW/ugiEfq50YWXIRPXeVhJuz16E61Yss3JREr0+E7sbLBJyrjXzbxVpiPIfMgs4oES7jaMIvpeivsbJY6w/ap2ycwpMZn8jOf7i7My1JwL+fwbS23dGGhC5BR4QUNDhZLmk+wuIWK7A7xbY1IEDcXOqLbggl71GRJFNjhbHDfhlvzKZIrz4PoaZaUKMI/6iW1kPRO6Jz86srTaoJ0Q428AeUljr/XIa96Bw2TmffVU+z5Ht/Bx2LDcKiVQ4gWly7o1sAwLgz1zelM+X1FjAtzVNF/Ah45lc0QfsXHlKrRY7rpbun4ZqSvOhwY33k0V6kl1mVd+f7BrslNsF3zI46nL4ry3edoPr6g9ebFWdp0orEGu9PGew1QBMb0q+uFNp4dSreC2wjVPGq3igmin8Sy7p+B+qzXdGESkM1IxpZAAnmcqWjdunzqw8OUidVu8/0NW/OgfBSdgWrpgHcTy7pQNjNR9ZN7WMOhDIwEvYP+UqEH05830DbfYGEy87Jhgh9QkdpKdG2MURBChFaaQ8CUy1+R51KldcIOKi3YOZsaMoyNypy8N4+cYkHi8IfJ+6hqNTbdMpJ0tpVp+o/JZnBNIKkIMCDLI7Z4aQpExwvyGTkp4VZY1FFqvO733Y8XUTOWzoTFura7v9DrDpqCeZ35F72MsKetVwFjQuk7YLGdCh7k5CnYXzGIGqaR6emswrmF2heOta4gL/F1EjKubejtE8/XeYeCuHKAfuQtgKlXbP2+X09qwIk0aBw2RMw0lIdS+X3+8eEWl5+Dy5tqaVHbGsl05gzw55Ud0SBigJz0oOb/UXZutEO2vu8CNL7dA6GweEqAlhFshw5OWBEZoLby++45sT+5dDFkotc1XEPdSKqPch/H0voNQX8BPJ1IZ4IywNt09E2924Z4NFffs+8J8+hptOu1oq6IiINc5I8+jpTMnCfB/re+nMLEi3MFClDkzQfYXxEBte1YqUMAYW2tTUqjp7yCWocwDgi+ndRorST/Z3+ISZVNzLWD8tHod4k88soW9It/07/nQ+w5uFq8TqZX49pgoPMOATnPnPi37lQ5W9RfIDhNwvFQzh5W2/PGAzxoYkxEayRBsnp/ogqw0RTauqHDEM4aI7QhE4NLtSrHmYiyNf1b7s/H78t9I3xyTYWF+syAlo4ptWq6f1IoNBcslIAaUwjENG/TWGtLcEnOvyGeL6s8PQhYZVGhBuH95etyZZi4o6FcRgoPNbu0CcacWUmVvueZ4qqBPkUUTVPfhCZYlt0Bpychs8JhGdoJmpmVLW2yfpfeJvOspLUhBEqcCFBaM2ws3arisc00G1IEsART7l0nCAqFm5YpdCBRqsOWq4zbuv2gkJCKQfm2z98VMozCQd5P9VP/2T5LO6ooVB+1s1h5DDc4P6WWLMQO/4LLzsa4LeIm5zhj1dJ8Dhfc2uTWUA22ElzTJp4/G8y114VG4TBMPDCnAnOs0pRu6T0yo2MJS5xGDcdJ0qQhYyZakywL3Af4OGlau7j7oRtJd+jvq/x11E4PpvQaadeyH1CkruQP5//epIryZhrFA6O7HjpW0wWhMHXpy7WREgBScr0wAPu1eZIE0CWieecgdgtzfE8P3ZecT3osc2oqMg/iDPLs0Gg1mtIZ0qNU3w8K8jYATK8JFbjVfJU4Q4vpzY5+joyRqgrZaeJXEM2J180Oz+CQMQPjL2tiSDmXTTDGLz4V0L+wO0EE8mGMbLC5i54EfkMql9jcHhQMWf6b1YNG6Ve7/ygWeHqA8WKEuNYGMh0QGwISBWtRBLqsSWabi+UeVyLvcQXD4N5xdlbUq5pS65z6/slrBNxQiYkw5Pk79fe58ODHR3rbLMv1DWVReU0+49TbS+aRP/bWNfoVsIBSfyEeQfZqERa5vHfag6KoqNIC8f/OW/OOAv5k7TX1DmIGwmUXhmGBMZS0j0/JcUhrgTqPB34Qw7UNe5lGK6CFuqH+tAmJiJPeiE5T9WOm70rzTglrjg2B1DLl6p8aqpKYGsi6EFilPdu/LUh0KqAqo79gtleuxizhxXS8DvLa0nGUMYK0cXhM53EHTY9fkGn0wvEVCJM5J9dDM95jDq/p5atZsbzvWpSUOsBus+ttOUvX5i1uSGSCiNtqT9Qux1EdnjhwwzxVMQUJUF8CxLADl9kwdk+UESDhZ+GQvCt2PykEGhONtpfYvVSVG6Owfr72nDvoD4nZ9G8sc1rmTwo9KOPiQiijlTHXLopT+DBZ9p7LPBfhZydnpEhlHNQ5dsDNRgm1IzkDimFZejEzG/sMGrH3BJKLI9B7uHuHmbuNA789XJe6fG+577Q7S9FGx75kt29bM8aRaGUysIQyW7aQMTwrhsyk08EwPdLOCPL08qeMDih4S7trxAYCB2UJim+hsguB+hsseBciVzTN23BBMJR8uMFZes7N/kA6xCIfvm2VJdUARzwRPX6Ulx1vN2NJpI6dvI/W4RttQVOyvBpWappW0NQEG6vTR8qDZyFtg9nEEoJNIvGdQHUcU2nkcHH12UXTtIsnp5qt1X2O4uDGiEqSgGsrK7iXHysD65Ldkqa3QngpmTANLOYfU32woKi89zfDP7i6UjAPl7575FgNWj/+Z+ZGui9u15dJikeZ4465/a+Zs79dGIwDQDRVT5kryRCvYLPbBJ9i7cb6C8JtQa0TBb+uhHFHmkjm+UKe3WXZU9Hz3nil8R3Y5unO9l0RkkP3HdX1yoB7hZLFDPk3s/5B3MwClHr0ZCECaTvsL9nq3qPNKI9Jw4m56RDbxczed/fayui8dUD1DYZ+T31l31rLvigIRtaBRdvjPnsdG93gseVZhRKziSyFT0tsojt8MjeNhF76byBTfsy144Rr4oFs5hco9srUFtlPNC5SvvE3Enw0/wWQI3mXRa58uXqK6VUXMRGYWj5Yr8CPPzFckvtyuTXJpP3/TjpNxWdkjXKBtg6kFXxDjlZ6t2UgnQIara1qHe/UUbcnJUZvR4K8uGFEWfdL03bzKlw2kcyJbb0upxyIInOnHazzNlH6L58s3oj4xISKfxe6M4hBwt3LQE1X9DZ5ZQ57G6QY+3lm0ZIW2nsA8sfNGkMXS7BkEnu4bUW5LdvnMGgdd/7ltBepPPTWzCTka+aMkNz9s6oh+OyF/u4nZiHK6OY6FtNRHwx2v42m3xhNIubz3ba7/YfPkgMloDiDDOvydwaV3zhM7nneW64ILOLQHbEnJ9cVYeGffkIzyp1JfH2LJt9Zg7EoTZd2ekH58OZpvKfdnVWpUgKnSHu+NHRi/qq0KOsr7uJ/jQVaznjNNeTZt+7vNbHndSM8DQMRvIKv2KJqZrd0Nm61g74PxLbEldf0R94pN/LFx18h7GssD167UEt1lm4ixOchxGZlZN49NckG+NVrx8CiXWLAlwAcyGjvaIYxkGiqEZ5E2EtZYCj7QBomRrW5stMXy3k2hVjByQqXtnCNeCYH7oXjm3QkmGYVd8dNOoBAZIQfaxSdtQCUlkW19kuH73VMv1NXKQpdbvf63pcTn0KOV9N9injnzOJcZlMgZ4c3Un9VZ17v+6i4M68rZajEmv4krqIXFv1IX9j+sHGldx0BbOpT7QbnHqfGSvMYXz8wcvAcu1vsHk9Lk5HuZZKTy6i0SDDSyzL7uR7wv0Od+4MbUODOdWdJzcDF45iYRZPrR/w698AA12pI3vYbxBWvgHrVEHYydbE82EpAl2GRSSyaLWxZD6QnoHiSMc353pSijEDNuKrRWJUbhlovkgXRdrEB4RV9hZG7h6sXdXw2zztGbuXahCVh+tgdp4j7gvVNa+fHwbYiDF2T9xgaKNIdi4aO4E2WC1Y10P+pMC9V5Y10UPO7X6r+bSS5sOwy8r5t6wlxQdg+UGN68gq4TDgRLcNYt9mVxG0B2KGuQ8FreIRCONZyL9jUL3PcIZmlS7CMabe1IEXT5qxMMTAYguDoSB6lfoRqDH4nK7f4aFO04PikNRU23oE9Wi8sAEmQxRLTn3IzI95elKGwufZUoQRWuCJHIiQBM6kjD2tqYMSUlnoyCqpwYXRa+rBABCcz3mtVTgw3m2DtEIUU6Vx09r4Nq7RDVQykljNYtb/UkG4+nWZvzFr1b3bvrLXpXWwyG4GApAriapJHeZhuzX09wVDP97+lu4FG9BqMdsKrsv1EwogwjWSrG+6Is7VJkk9WdfRJZH18wmNtBpmt8a0XuGmqRmT8fCQvAupqD3zq5P1m4jOLi08Y0TcI7T/Tj/MQypk+DKH2sWrQUyEssW0AmifM7uANmgIFrizZGNQBUecZi8RB7Lq4TRb0bTARhXDnkDmeQkVNiGhZ5HQwRM+cDKHy6GxE1UTw3h7kYAuiSuz72KifYmFhgMjAVPnbIKGyuCenR0UaSlU3zo8vgTbbUXh1G0YVOH8Ei0yXONirlGKNIMpvRXQvo5s7RkjT/cnz0sW5NbbtuDg5S9h/HKqqLDSBQLwdvGyONSYa6oqjtzqPzFqLoxkYORgyWNKD6jn1O1zitMj02VWQV5cYmCoLUA0ocIYkwBD4W7lkSJqmc81cE/wHwOJy83RmENqos5fco8z1MQRSkqNaHw9gT++yQXXnhpRE6PhCv4HRYLl6G+kHoEyvre2cOwl4PHPDluiaFenuQXX4Y9Z8WjatF1g4TvgLgPQics7wew+ZpUN4ZOsBF0i9Rn41B2DUE9psXb4/0ZRieSSOWnCL7LXcC1zS+elo3u09pDHBA/5ZCsVLm8YkLspmSC3r5EMoOlzTCUk7iglzyj5Q8hKPo4jS6XDOLCuGZVhQwFxFNJXnJcn/SoxTdmAI96RNqofxMzJ4A6Co149bbP8VJkaDYBuCCCxkHn5j4vwaMzu6/dIH2hXMagpt9OhbC+V7FN/V1VJoSJxu3lsYVE6fBSOClOEwZTJkqFyCm62W69yMGcz1CQtT/cNsA2GkA/CH5nO+qUyNG+neMhzNrCW9/mFzpoItz9za3l8VR3LZhxV8VkeABlBXfUCP8XE7VPeN+9hH64PzItDIU4tbXB+bLJfUuh65gr/7BCYJOBdyrDSLMkm2Ld6/iyRMR4gvFX3qT3sK2yBi3hrVEQUsKOwgkhOHqrY+R/NQ0DPCAJa/QVeiydvZ3QFezeDt9RWC6W5bUMRBoWVEs6isykLjHNfe47olBEro1xUsQwklh/AbrzkIbvOTW1OeoU56uzq8goWZpesZS89M9uwWAp0QwIO0O6sYwNcUYTEwUILPgxJYDyzicDZKtmTwGhabzPIFIiTe3uQODejaUhBzVlQGGYv8o4tsim1Ihz6ClZJptdyH1PQsw1CK2vYwBkyqPKkqZL+aqW22VTMVzF2LZfanMCcnezxdYBFZkf/uoKbbancFl6QD/vyJEJTLI5UYQTf41DBC3SeHfD8bChNTyvxZZkdklpbucUTvlkQyPcv3KRHxmVqH8wX8DQ+FVSsr5TJtwtVzbXOcyqpt1XAiwEQfPnzzxyhdqHjpruocV+Wj27Bp5HpRZobcLXUe+3ocM2TsYc63Z/k5XBXV1U2SUPNChxZqdE8tMbzkYra2ZOLHNODw7Xd5tyjA1P1cpgE+rSyfy3VeR8j3jt8XjAUdRdfrLQBDIkgTe1EvV8L0mtvKsqj3hepkp9Yrq+8bnfVZNQWP1a8k9P5hQ/61bVwCgY8WBXZMF/5gfcn1eoxPcAAvmWVvsnSGavyjFrdmx8Dv1SkV0S3rMEAVWgNnADYldNiF3QJNfUwARjX+YJppNSwBnuoCuDtcKzs5a4RoEF0VDVHAZTrFhKDx9tochoIyaXUQIUxi/fScJ+nfqswqtulCZ4PLeqGWFJ9KYJYSlI/O/H2rPBsFzi5E3baMPV99LPLlLDIlc1Puapu8rt3jnW8y8K3lnCBq/MY8ytiE6avNh24lnMfdp9Tz/JdNzSQHL72umGQEdI6X/X1G9ItBYUygaE1fEo9nHl9MC3cr4U9i89FCuHvoVr/0u8/oAaciihXzL15XiAt5mcnvktIAJ2PpEe3pNKdONITSSFyTyktAtQBDLqC/AlHYpeZppFlrNwZ1DhIQc5BgxNZkjEpoN9/qewBW+aIcdht0/V+NTA1gm+lhVXA57ep7UNxno8zbMJ+1VqXEs2suzjRaQHbJVJk6EwPOWv3QpnlKs8iTzHEd7INfxiz6iyLYloPXCYmiORog2Xv1BxaFso8AgWWmY4Hzf/k5bTYUdt+Uxq6TThY4bXlflVqf6ahGNZ4kv6IeXjPWtxybUZt5FS4W7K+iYVQcNkp3qz8jgmHnv6PdOmW6nMA8Ns3rQqXhFC6DcVwGbyS8vYOB/Mhl+Q3jmFTXq7LN13hUE8/mJoDsnTk/Nv2mkZ27aLd0381DAeaiFFzfd8hKQg8zqOWExWBbpddcy1YMgBCiHmX4Z5proczi6Ma+liFHpSBB6pVNnfFzOfNIdL+E+/h6P0Oc2kG02bvH5btoewDRDFQYrwCrdl3deXMOtNopspd9ArD0T2/pH8w+tszV/jbsY+9XYXcEmzkYL1wkkeN8Mnc8djeOHd+Qex1uM2sySJWHAA7s9iUpc2N6zbTZ1I2UMDJcVZfiSBXmlN6Md6ek1ts27bDszHWIUtZ8bz0Br0VE/spH1E2YeOdSz1qiF2pb7H97fWlOwFYspoArouk7FuCWEG6alxBv5laKlbMpSgtjNw9hRM/QtF1h79zAkQaNvM/STyq1HC+WBzAQPJkbEz/qKXkdUsUDb503/smz2VI8w4TGME3A+XuzwMesd5HcIvwuM+L+ozpH3NuwR3s4RQITTBsSsnBCs7hg0iVs5S4Kdd69ONkRiN1zQOADr+3GtSSc2RZdzCrBNPB4mHJWDH3k6pdQaZRLYVAu6UcoopU2HSExXPGVTtakBcG7cBcOkhBnxwwioRPXwXQVsd9pycwi0Yz1tOuRgaxPTv9Qa04m451oJx/M44N2DRfGV1oFEtoX/k7CKPfDslca42fR6JSoJrDlG9+qeHaFFW7wTKVJ/PlMt4LXLwLWQVeAfr6SDYdNsHscL5BlW7MKrE5I/Elm7ElAwLJWpm5sdRkMoC3cYA/mNdxXCfCU/ObicmFUkVRP1e+M+BrNuydQiBvI6ZGRXX/ax5uM50YogETsq7I/vHm4MJSOxxiV2ncDCvyHz70JhX/9D/gMUOfP//qvstAH3Zn1aMw+2z/MPkUdDy9Oi3pNR6KCslP21mccUqjG2o3L0JogXbBMWQsFqWOJS+WpUwA7x7D02vjRHPulqt6ML+tj2gW8/moT59GwKf2Fe3nly4TmZtEgkzEWGcZzD+Rxt202WByPFUtpCc5nEUUuuiStF0GO5afAv0jIexXH0EW5y+Fm9AcFriZ9ff1E0PO9lJdZrwZxJJs27uSZ/69vHTYqRPGqnVTIM8ZLcvcEO73iPZh6EwBAqNS4Y3GfuG7fcVE4UDSH09Syrpa+g8yn6LZoLKZtGkibuqu0vAHGX+Uind9EKPmouYTE+mQ8s1Z5XQiyZWEC4qCKvZNrVLRjyKtmySodFaTpOmP3u3GCcrFwhMrwL2SFytzIpl1OvpdzKec3DneyDu0EBexo+z5UF+86pz0etG8f0VFyNEDMZOhImjGXy2KBkMn/lUwWzwxH5/FBBT9BfAcdC7pOXfn9PhslisIayn/MPkcO1cu4BT2kfK/pJDDZpgJzdOOiAOD+mtkTCh1/BhyzLzqQkNS/MoLqniPo5IChWZBavRYtenWo1/O6MIj5QdCs3qH76fLmDSZ3YBf6Hwh73kxkqZAOnQrj4KLZ/bz3VeCuiWQd72q4bZbc9/kPlXyAfh8wPyeqCm79rRQdgRIPZ1y0eOh+GsVrvyFqAAVV4cSIEfc5dJtchfSOiYNe44CvV0+kMvh7ixSXGHjNi+acUWrBnBzpfeJZYeWtkjFp6JUMheQ2R714oCOrX4+9LEkhANA4y/iLX1wwAPSZjSHKVxIdxYBbWFoG/XzpVJH8sAxhpu//NhqgQzNc8v41gI+GsUcHNSc5bZ4X85uOLzUIIgZsnu3k22TYd42NWmbvu/JGWnzVtkloOhZ1zFEKehL/bwqdjH+WOcvxOMcSzGw9J6jKLpY+a19Wu8WVpl4HQLQDwbRtdqB9T4yUUKfDp78HaNK7t6tf/Vz3ETRezvqPJNKYejEkve6erqBOVtdwwfduy2eWVc7tpflOZ99T7XTlw1blN6vwAU9872HuyiQ9txe5gQ7KZ1eH3aQQKwSGtCoHtGk4xwaSC4vsr5907yoZH2whpOjSdIIRJd7ivfnzcCRzXtDpbRJ+6VR1sExko+vkgNyjDQbnnYw7uLR6m01zgPYwka85Xiia4oQpjWtahfNwxpG90QLWjbq1V6OtN9DEkNSt1JIm2agSbxWbcTimHiMn2b4GX6+uDuYgQxTrBeQGOsdXs2Ta+Kn9jG9BjxH5TtQIiO20cE58SbJUd00IqayHPkxtVYhGf4wPeyMj9pGAG/vb0zm1VWpx1bn2Tz7NcacLsoYxIO1QQQ2ViUGMO3Q4IzuDC4qHoieNZ6l8PHVoTOCMgmDwp2sV404MlmSc2h1LDJv2Gqf+E4L/rgEVS9Jn3960IDZhSXyE85yXlErNywTgKK9agJDXjnzvHKYQj3TAEB739n9fgMeBbyA9L7ejb/K3CY9+KGdExmfYBW9Ec7rtxjh7IHrjYZ9LrQiWqCsGXhK4GVK9nRqr1eJp8uulZ9019LrQGxOtM7tmB8Ih2ObQOrsjaG1cuoEplOU5m6BcLoc9z7+APjThtv4XTlrKQXG7evNhQH+At4kBkCyWcgYTDpkuRjebFrw7eYvz+SUlgvh4QmJZBSN2Poh50E7Ma1KMr4t/Jdswaxd54+vwp7hHLb7Vr/UcTpWh7e0DZ9eSf3fABbwHT/3seyCacTf2IYIsirf2666EZHbHz7Q5PDZaRZA2cFUdFq4WwU2iyfJgNav6eo9xWDLl+tauhDUGdE1zJD4FtyspjcR4eK55PAqI8kfbT/WiqMBKf1/nyJ+2WOWaMuloPFJ8q/iZhHcd9s0Z9pPjbgumB8gEp6amFqfNq3wnoH4IdnSo1QlfdPbCegV66RJLo4bydQSIVAabJAK8ZGP1UNxLRlrM7u1tVL9pLLIS8rZddL4onGfT/txPMJFu1jBCLr0S4C7JRd49bwnUNg5MOdERcDj9zTnAmjnYRjBBQjeznVN9OhLwwt/UsMGPUt1XHVD1VCJLv0SdqkrvwiPEDOe3N2G5AysFbA2rHyjTPvqbXXGCVs6nAtP5lr6GqMCNgnJ+eoMPtjApw37gBme7/1IT/CHoMtKMv6wMtCnZxHfKWsLD+siGwnWUthWZxJPHXq3PU/+n1zpXRAi1zRjyX80s3dTRSJIZsQrVDJxyY13FYUqpyQk6LiyQVlfgkCKbb5GrIIQuE7MQsxR6cfTMx6+qIdzRlRGYPLOmoJDtL3v4GBOBUXGckciMthUe2n9ZItSKtyyJ16hSPlm0hrx/Vcewi0MZWOH5c8iv0gpYzUmzfsZ5Do3Qebdl7JDYYEBal9Shvi/48xfHs08JBYjoz9+sqwAFpS5mhIhN/5lD3tM6qHOG+BaeEJK1206YfeEiVdBsutJ4ROfAHHppahUhROkGZGQRpISBa7TB/NY7aC3t72TtYRvcVMxGFX07lkFVVzlGOeO/FRdS9wBTG4H+4K+LnVQZlJKdWukKITGwfFvfnpnvBpwThK4RxKuxEpCNweID1wKfaQldb8WdwGGnyBQE5F7ybarmjRBlW0dYNla/I6GHmyBYKPffQELm8EcKH4ndfgWQ7MQi2JBB17bDPqyJJXJaYK31Vc/BGQdmGE3N/wgNKnPSVOYKRFfnEdcuK2Ua2PT2HzRPUvm3iVqpbN/m6EQJXhcrQ7ynqY+H6d5B0ff0A4Lf/EP9uMDzMj0oxeJoBAftrCubGH8QwwTZh3ELTsE5x2zVpN2xClPJqvJGK3gfAFcR+7+QpGeq3hoLxkkkqaE0GEeidLARM3pevUUWevvk/x05MDe7//OzfIXioJn5CzKa+v7dFYBTZkRUzQd61gRDl83+cbg0Hyg5KUm6VLowV7kpTme38i4SnMfsJJAcIN4nlyUxUoGvN2xfbQ659JC8IwXNZfEuIWZh5+LFGX48uypHpNS6bmmRY7SFZuFAbDH8nN5XgTGVbuVl5+zh7feKt3KfdPDxEqe6cOHQh2WGkqNgw92tRCCgHdPZDFsWVLhJYibb48vEKnYydX6nJBh2vde84GmjBTisRj4QwGGfuF8bz0cl+ACF76Qb8ibWYt2KpL2LcGQygdRXBnBVUDo7wwgVXQKJb+W1+CC+ljnXHuw2Hc2HF5IMlbsQU/FNDQH5gbNV5Z5o/ZyWcFMVS+sgvmWC6lr7GqgKIlFgI/EL2Cnl0isDFypqeYUfMq1QnKPE1WncjGl5VfC4IVvAnf/05ar8ZofUhTRZxZ/WMQ3lUw6JIpNPLWuIitqLvXi0YOsn3wR6m1Kt2n86o0gkXwFdrfz8Fp4wIgjm+hrzHR3N9VR1PvzB2TJSxoBRlp+T62oBn03nzU8qKb2KJp1c1XRqqkBwPqC1yLzArfrvAvw7IEitB5G6s5b1TYpGgZeJnmRXofyZ0KpXRyNS8l33sFsMTRgV4G0xcexyO3qL0JVPs6K4MlgDh9rBBtKBt0BaYK9uqkymg5mN3EvGUA8G5WjtQSth5Ucl1MFNfn4Tv6Ya5VyObFu6z+aF6b8+ktZ8imQUDWrywUFZ9ZWRw8qcQrXITMcD/GWG4QmOkS7T56D+TlQAhjnJOjexrKiwMa8cTMtuDGK+ArrNXebfqmv9I8lQDC7+rwNOlwHvTBxbgMO4EkHdq3ShX1cAEwc8wUuYWW3sWotJcpeFVbo8xJlRq32m3Irth6ybZSwP0Rcmh0VPUW1O8qTwSDNpAnhJLt7d+EXzJHkODe3ns6yVFDsNiu/3IVhssyzG+JOErzZgFsdBhU+6/ySpClCexlabJaB6eWiU0u5Gl2ZLuJZtjfZO/g2hAXdrCeRAYNQssJ06ltj5VZgB1DHtic+GGt5oke34HMeb+0OaECT+swbY/GfFznmqyiGMeT+Kn5FBZaK6UxKF8fWsETUBT5nHDb8KBY4J2jTd0tzzWNmjdd1Chjau88Z27WNmLrld28hm+i3VdkX6XehzACYGvDb/ykArw4hIbd88PHyTMHgK7fDD/lsO6a32fOz3BPJycavD5TNVpvPL6QWSuMHU10oXXOzjE/kayIaRXR8nLtTbwUU2otejeOH7pb3oKqU0E1NtvYj3SypMJrxqbJRi6q0TTysBBNw2XpuAZF7tUiHIVqnoqRLdP2HFTkU4MbU5rdj+ruMf+5fdz0+2zWkFV+R6GGr0QLXk8FinsKHYW6J6/skV2EuOJ1vsn6x5b76bcpwFFpd2KS2miMFfRRbeL2t8+aWfO+1+PHKW2NgGaDtgX469dbsBh00gc+/6544difKVtqVwV5QydG91/R77m0cVTPONPXCCbNOtB6WorbbDePjcmnzIDl7MPprch8k3e0OhKayhQlRgDk2Xp5/+qXT+IlKPwVzdBGIoBgebRZS+pJnqYxFReApPFYVe7/rUzVUogjlF9IjbNi5hCYQdWzI8hdzZPtcPqW40HjkEpxdBVqnBKaAWcKLGUtZ30lSqKuaQBv6HG5zcooi6zBuy6yyarpLuL7foyRQb9atTsozgPb5l1KSaqGTWsrdKLF+/CNiyQaQ5VxDJClhbqHeQ2YLTStbSNxLFXP4r4D7YuCqtjGy/kE95ZQVNn/k25dMrt/JE2BycPfozYlS1WHRnvu9lqIiTSLrvTmKToO4mQxa5nSJBJwMAydzu4fm52xhYdTIGvM+edXhJGThHN8XmHvdTDE+bdfknk4EDFTGZgYtip5Z8r68m0Z5/Wq5kLAXXNxKOhw4Oe/DXknoGYs6CaFwFGUpinLN9qUxaJTaEvBhRM7XiMAKURIpCIoywUF0GOTTVxAHCcfyGHirZnpp3mqSlbjXGBhwVt7t2h7rjz632yXns2svSOnaDFp0E+mNKqMrx07pGaV2WID7t0phKqy42tU7YQsrL4OnO2OkUSMGpzywN3qwuUNbJyXFMOS2geZBcLQYhGxONr9hNIF11FWBO8ycg5x7wzjxafAEcC7w0FUYpGIHxJfOYk4ytyG+a5L2lex86y8NaPe58SwgPbFDCfo4VLKgELTf70UdYFW29grXmqVG7a59lIKaSKPyl23+ZSEhhrgTC3pbQU5/DG/Hc/ou+LNhZTFshjQ6UexkHux1YPmnT7EkOM0dBTupqinBFvcNeHQH2Z2Xa2t0/M28ghjlfg7CcKt57K/rgK2QpGfLzJhHMojwX/wA4ckiUGskNl2YRsj6sDPjc6asYGF9tV77UUd+8gg80F/EOkpVI/Y/Z/+Bgt6A3F2YYqiKc62UfDDV2BSXdStLbM8Ne7PZ2BLUYdgjhMdu6VD1brw9myOK9K3mUmHZy22GQfM7Ar9RmDsysVkSqO839Ooo1MYz8rs/D0UnEptuq8cjOx1Zig9oigKYV593hDhVHixtVtRs/xm4sXr/FWobkzzOSUdkz/wesDqrCXnnl/MoOvcPCskVbI0T8idkIPyjloDYzE+nr0crsNae1Oyu/kZk08ff2CCL+gKPxtpixnDIslxQxLvW3tMtalnollLzy+iKEn0a3vT9S93ZjyVBGLi1O22+MglJENPUZR2WtjttaaEHZcO9szvRNhMINqWLVXadGLzTWnI2AA9uwx6QG5qBzpKI4oLu48spVdelmVEE+zN+ggm9D66ZHtb5qErsB1gXQK76ZOGxDCZOP5n8J6+zDkgTLHgz1fV8walglw9Oqb3rrNJa5TZUeojOjJAde7QERh2dWZOM+OvKcxEndWHkAx6tUcd6j/EOnCMfyGgCjkWlCG6STTzG2ROCRfh4AIizxiUSgSeR+TCcWwST1DZihvgGxmnCttzftnojL4XxeLzoih4QxTdNlFvMyqJg75FP2sUdl1Gd9yZNNTgAyqP0xwL03bUboQnpE3CfM9lFgv70PBMpZ8V8dVx/wKx801ZKYVY4mnsek7p6UEABoIS05wcW8RDOQSRaJVHaS5pXpLlQ4jgftTafVB5wZE4EBJ1iuwL7CrZwFDPlRy9w5qDHfmNemYCkfopSLEu+w8bANew6WjAsQP+u58ECOLzjDZuZAl1pPzfEyyp9rcX3VHJwMWoSm88MC8py00g5DDId5TVlv1hyEq/8uCjqzCXvSQ9d0+j+JMhCSVYJClx1UUVT8WUleYSpPhg6gZ0ME/pbvvFEXm+kZVVA6jEh2C230mfx0bfQY20Y7kVa+FDBT7WINTi3Vy7hQvZxF8zENJt5ASktNUaJhWPFSBTaeArJMNJa3XU7w687Wuqc99/HigJnC0maKNutzfmCI5MAh4GG0SEikun8JRLdvJd5/wKhDnHCrFWjJXQYDSRuk7g9TPt/x2LakVtmxiAU7S3t/6zHVw1ADo6UiCIhDC5YQ/VtasREblPPXrgMryz4s+UtxqRcD3JgCpeixl5xkalpSe3Gn/hGnXLwOdLhUvVk7+WkRq7YrOWF9uhwj8D7B/55hu3nRpk0l1wdw33heiLs+/i8RzcdGYvP8wkVO8oBQs10Ul+AGR25+8qLwzc2HVotv5LozrNq7vFYiKGIUysnUh5Zlb+lBsjf1BtJAiTA5kiPdTlHEiKRuY764RFm41YRQYx1lRXZbJcJHXzwFyomPpDsfrxNgH0kHpO4Afl4feV05c+Xq8JbaDff92+CNA6ShT6XjBEgHBi3WzMt3UfSELGimavatLHbjz5OtBWLD54QT2J1hJppr8VBQ11D3IkXuWPnwx5cgoImShLUkviyxrj2YV9g8EfoK98Zn4VQsOcEOgeuby7HuYbKYJTCevUDHuaYQPDiU8uQ50fcmP7jj48nq1Lk+h2rGCCDgFRZwIzEyZj2ndQgjAj4sjyMSu2qpxfJRZEh1mLrcEdnMFjNhNyJ4qZPHpQcPZzV/zz6PXhqP8CD6RbnpGUHW+2qW4XZI/YsQk12DbV/FrKW+AOfqOC0nHYwQBgVdY/TiwSt/mA/ODOlN4nocOwLASOaoPOlekwVAsjo8vUOp4bkxotSh27ZYZt8V7S9pzmHwucfS0iJx5LpCd6eb/t1of1RLCv2HMd/0VIVRKp0P+FvlApWNorRA8hp3x1jg7/piXeHsj4gZI1W2K8=
`pragma protect end_data_block
`pragma protect digest_block
7056c7dd956dcc632fce8f9f6fa98329057d7cf435ff1400bb9c5b42c58e1a77
`pragma protect end_digest_block
`pragma protect end_protected
