`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
FO3nDdqByTghGgQPOrWdB4kJsrcf/BJdJDDLuO8v3frKYacXe05c6CSGdS65roqXa4u6Ldyeak2Lti9RhCcM15mJvNn90aUO8faN+QtPIJtlizV7IoHVVGcpzN2ZtBlrzTe9K2jVbSyOklJiSiJPuT7uGQh7XVoXbVA31S5dpOlavUVQQAmhoJB2kZ6dbUMQSNp/5KzYOXsn+39SZJq8rZi11g41mKG7uT5Wg0Q5T/hAYB3IpTgf7CU7pBIEuCOcEnI81dFkONPr2bgadNK3WJJrTSHcdTD9Lq0iwdVRdsoXQYyV03/0hXpHqVNAUtiRMM11jQNb5VLK/dqBRSBhoWPuBN5HVnWc5pq5bO4+Wsk46gvItMjOJSpDAlyv52VFFX87KWGVxVFMfndTWZcgW6O1/OA6gvgp/Mwg4z19alwkRbLWqBoQTT1ylmjDfRDfbhFboNRvUTFOkgoX8zkTv5JSx7TdiUnJWw/T7V+JLFGzmc8QLoVs62OckAx7eQTLu6YYFmCHGxp3aSxlIPk3bS7boiRdwcqZ4RY4CShqHjmoChwZpPnMvqU6E1kDji4IWzgfFmqYb+P/4rat5pcAG2g+p1KRZZ3a8KU16MWvrcCGic40D0yMyMcjAqxgUbcNjrAeQ1gAHQU37hthQMhUdzL0/xca+zUNUUX72li5VCQ9qumyAYxIw3+ZzjdMO9EqnoMcWqiKs6dkTiE77p2PINEl/nYwY78Fy1CBBTp6CHXEC8uwIHahrmaJ4fZbiYECDQos/7Zc6s29K5VCxs1DM8zt2OeksEWz6sBCi2HUX9EF6zAWguvh2sg7P4yxLvO0E14sI5ZkPmfzBsQ7I9tph9bw0nnfT6bxDczWXIjFFjwXGAV+VN2OQJV214hkS66wSzex0WIQPifgWHu4OVmHwVPKqDgpIHCy/3CJ+1qtfTTT3Os/nQRn0tYcSP93QL4wF4xWjJ+DRUe5BYYVBV9X6y6l81BEVLWmJBQQoZLdqCGw7Ewi1eRBbZIGATcGNloUFJknTosxzc7F53cB+9M2LTw6rlIZzuvV+5vgE005BysWQlqlvtA5lgIQfUUlW4nGzJgNOF9GKF/GUO1B2YTtYfLANSFNcjd8eREiVI/Q1tbDI5tNMPsrgzuFg2AHbrBYQIWGEX7QVQik0I+d6Wf8fLpW1wzIMp9M1zr8aQ226KsbcHgpu7t+1JIBruAxw9ZjDMiYMDm9YNy+Wx+yFiMxFJcshI8w4xypQZcF73pSX8xH3ngVhJPdX31MgFkkBwS+dJX/n3wRYKSv6nEN4a75bAWyiS0qsdpg7YBKIs4q76P9ZlsAag2m3m5iPHwU/rhRvrDgqH+Y+gvAC4hqAUzdsi1cNkrydCD44rP4Yn1Qt1JPMqnD/wFxuvnhwYMmmKW9J3TzWEBetyCZgR7Bp4/FLfgIbMWEeZn4wqLwuMOcX7EOIYCgy3XJL9eitse/2b3sp71YONLqXS/QDmzbcu2EjI1sznl4Cvo09Yu3Js8XvPheYBRXdeMUilE8iylU6+m/AtC4zTNiUES3y98c55I/OE/lMqU9bBz/CMY/KF/uBLlche7KTPX+RV6w5cbnBJdtfyHT+LYfa+JY9KiuqFniHcD1O5fwuKTraRb8q47R7r2CdRpJy0dfe8oUXk9skrWyJ6qyWTuo1c/X8YdOy/HDR3wZL8EkbUZXela3PoTifiXDA2T1yqRbfxN0OvWO4znYyOhr1rz90ZRh9Ht6IpabMAgI3ZN7KpoWZKFR42RmuKFi8U1olD+KmrrpX+VUu90XTOZInpUtq5pb9+h3bWfwG9gqAF1qZar7/ASZSIPAtEPklBZpO7YmvLY2VNXy9yRkSwpzvohaI9yVTmr7sQ9rFJR3TDompazkrYT0Zcf/2KDrX3lhSmKhNVVff+SwQLJS8I6C4U2Btmg/0/dscjmtDUF0XgLcUpRYYiQGJ7JZKnsFtnaWByKoAoxzggFOMMkwyIE+maIN8s7Nvl+LcxSFQG0vOgu2+T/Sh0JVCUMRGnF4kKOtMd/rJIUHdmjUlIBenGClGBVolRyFEypuW5c8U8pNiNmDPb/LD2sOI/LWhD64EbQaW6cAfciEHpghTawknoLzF+SLoUqLUnvHe9jrn+PbXGiPVVfFzBC6TX5wPanoLBZDRhOZMBAwgW0tcob89+n98Fz5xC9xU0F8LAvFnbp7AjA7UpDZjbzSsmWdR+1GQ3nJX1I37V0Jtv2xOEioAdBSMQf4d8ie6JSqnuk3lk1J8upFeV46S4wTyePyKurmShfuAH0rCy/XjlWcjYr7EPAXTlp5Yc4F07D4VayyrqNdYgGMf4PCRZgubFVG5O4vC5e55daiaFxQ5WBKPqj9Xi/I+/GUNqXDKYIKcTQzC/XHNSGQkQ/8GHqc0PEePyMFNMp8bwB3x81+kwaO0+b5z561SxbVv5CRCesOqTKlVQAtV9tEWsbnpLB+wXgDpq+VUH5FV2Ss0v6U2QRO1Vtiv4ghG2pxFWILaa3Ldi5PbNwtET22AaIDxgntAC4dRFyawsH+MOY392bu1sye/uy64FyhMe7xS9pk1bxJJAKQeQMeV5+mSZkkKXZSUPiYjLBPZOD+69xjN83Fx9u5z2jc6ghK4OSi7XpDOgCN7mqri8Sk4AEtzT95qVu2MU/fuEzWONqCOV9calS+EgzeCuEGPl7X1vO5neBoHDnpt5It2OhNrvsOYVCypVVCkWx7gy9IqDGIlie45yTKzxgFTS+dPjoi8MbfOrPdJ2sxxWco9IBbtQWtL8qhhXMWL/j+Oto6PU22cZFqRPTVfrI7LberRN4OMr8kyEat80ZED8vUPWrG6A8R2vuWpWwwzCiYptFngl8+KokwBLFwdDcnDo66Hb1a2rdAy22xdyMtKYaY+5b94554d8+vbB6Y3HTpJFXX/wrfjnJeLQjGK5M/9PN2FKXhnFsWccE9KjDDIFQg6xhadtmAiy2M8ujQm4Mq1t/yqkWX9UcfQK5T4OI+qLGipYoMEO7HVN3SbVsRj8Rn0jHxf9IMBoeyQJSmFMKcIUcEn1E+RTeCw3uWeWeBI2ie7ZSImq9vFFgN4kLQrzYjNQbxwyp6qiE8dsmfzCLYdAyj+MQ8D1XhOymimWf5NkFfGM2mKyQPzsxI6ksF0JB9rhZXpOfrUJoFH5Tjc62khZ0ZZXJTJBnG0asml3XUpRUjLeBdJyowvaxoMt+RIaj/P630fjvdoMK5+fDZjGZhPcwVSzHX4/h/ds/OEtPN/GZENOvTV0hutlJHGOt5q+2RekTXlNgQXubQL8ayWc6B5rWUWf46BzO+Q8K2sMv5DtQomW7XrMOO1ESnlIGQRQJY8qq/gRIju4rYAKV/vjk06DPJpFApJBl+0zx2TqdAMlNvwvMEEbKuSj6zcKSOhwt4bOkd1TOFSAUsWuW5tnPrBunP51HnKf3gRYE7fjChEl5W8hFzPP59BsWSASmplJ9QsOIPD0LWZE+V4+gq4ACmbPLA9saXLvz5aeu4kdgOfSlBSnTsnw0akunc8M31qADcitbkgNKZn6b60c3rpr84Ghyho0muyHsdyeKNV8uo/HbgErag5gYnwVFi64ZEumOVJE46s+akYwoNfdRBc4z10+lbDg0HyX4rAyIDfUNN/PYQe+C0zsPH1Jnf5vkoIGHgSCfoXrIHUwYQfrHp3QtSypTqaJjXlYzPIHrDfjiMi/92Yacq2m7BfCVVqyWSqWT1BTNNFjU9VmXYrZY8UQlGEOePvtjgTmPSdNu8DNlmmi7VNL+ANxLi6hHZqJyVyEm0tlgKblEPBlF47Ii43wgVlm4/e4nDKLg9UpePPivpBspZHBKVwcVwSO0JoI81W4ceRW/18iFwDeonuANS8DEdUShNR468ycIAfLHCLFFcMhWWiuKVV3aT5fg3NJcxxVHZiI/6xgCZRM1Xu7BOhsOO7oAtclSf8dSSxy3e7Ok8gkTHEk30VFc2Bb5Yixalca3vxVqd5RiSSBCOMON4rIdXk1KbKeJk749WmDjb6IfCylKoNOcPiLgCcTqQqAEwgrxxo61p32i6OvDyOjMG+sUmtUNXv1/C1LWMdL0SKIVBFlfXGOCr4P3PfC9XmHpWGh1pITOm5VuqxQWV/Ln/krr7NND1JBKYIhkUu26vTqkWBIgAD9itrwm3u4G0SCPqBgmNtjyg4gXadmz+SLsutkobONZm5XMP6IOMfPHQBVvs1073Vr3Zd2HTTxsLdaMfLck3nd+Qwyi5/JH4EQx/2nDX/KhCmJCnZbdXD4jqJDglaAypSv2eL/LezsMmtlyjTNk3hB9rX0hlCxdRifI9OcK1lhglvXVUYdDag4OviDmL+JuWFH4dFkMOr/Rj8Tl5e8C90L/9vcg5t1spVM6U2UbSqKKT77PHvWDjY4tfo+61g5TnKM99pYb5Hn6ISyqrfFLg6CtzQLNwFRbXYRhwWXyvG2I/tdIbIyqWfF0LvpTzkvvq2kHRzYBJYvBdNqLnh/QhUPv9JDXTcOcWyhfJbLGy5UixwYLTqnZl83rNqWZLVtvecvSO543cMchWjAbpxYTSniuPnweE6TxutMU80euaMi7eN6UjMWiXTZk92sSigO6aMqUl4yWJsBrwLokD2SFUoEs+lRy9oDTs2uAk3gmWRb9IxpcZEj5nQJJPARnjIRpnalHicvgNPGqWI3rasDHMxYOyBMq0c7AuhJENIb4DU4xagtnyEp1y7Ekj2wnq/ry4aZOZrvoieRje5ZhSRMdkFNcrd6CaZ/gv7GAHztHlm1ZbyHvXzhhKVgp/KKqzcLUVYOI1dK6yx5BBq/i0rKxsLmUTYXoHNx4eLv416TT/piUP2EShSyhMlEA63smTYvhjXaIg3FsMZAbSam1DkSBpic2a5jHhqm+AVuEmR5XNW/kIWDAKktuIdzBXHKXpYNA912q7BY1ea8aSPPNuoGVMbjMsiWmpaFnJphaDwc2J5s3apQIVIJp7Z+xqrIf4zKFYVgZyYr3PpNwkwE6VY07wrHkRMUT23/KccLwby2zfwsT+llHcRH1gC/IcimdubHfe7CUuBcpT4BgAfmUtYeEu9h7qqbTmjCMiZU3HX40MGRgvIfp3Q2QbfC8Ke2u+ihnaT0yEF7gMxaGHIkKXZR9lLDUkHSeSFAVRQcqhLFhwx4DHB7MNlZVFF/ZY6pjZTSXR6mRUMKxRpHHluiNcn/dY1XKhD1XGvObv79VluFnN29aKtz3wkMvUIpbpFqX5jkArOn70crl6YxSP/LD+sDZTvKMTkXIsWe6brTlZ3E6tYo1Q6ILB3wbtatc0VWB/nVSy9kvYSYsAoZhM614sPc6CdXICC6YUfe/ZBuDmSwJbWu+W/WUw6v5womdOW/nE8fGuK3bq6YERpydgCBu9z9r1zMEf5gcgJ+g1igwRpMBB+XyhmVhWTqzsp2z9/oHaVd6UPe9997syuKQQ2kSadU1HMlpxzvtHAj4wKUpaCqfAMoc9vcpWAU1fSx4FL17GizDJaqi3QLiGS2pdNzgHDrHXZSPEMhYr6EuI8LAr4DDVCZrAKYnu3u9cAgC7txSsmtkOSUyJ5HsS5mHZPehXkQyvyInwg80TjOveUSWN1Z9fk9ew2FxndbfTwtMh23mU7cUhkoWV02oxFe/m3HIqCvVfpjePIeADJZWZE4AaRGf/E9RhoMlzM9YsSz+F4mn7NLzgRDrKNY9fxAPK6f/wi7yTXRCS1IYSZJKSUre+WLKX7RUOwk03N11gsK4RokZzOcTY+e707HMxr9eWxlgTW9krFMonB43GPLQRFLwenePlzunZf8yDB8WB0LJ82xHwXv9bAGtxrZerAVrlaqNGQJc0yOi9C9JmOjV4e3DmC3ZzuKRTAlxTtXXs/FRNiGME2GMUSEEqjeJuIHBQ5k6Lw/W7SNcU9pOQalCf09f6NhXoDU+pFMmc6Fm8u0GhJy2KmkTJf61vap9yT8+aNS5q9tjhXsJCn9GPo9egPYP5nYiJRlhmPkyTq6Eh0Ejw0cWitXO4m3qxEwDSAnRO6Ss9NwPR0/9SpMflN38zsFMUcfy+K3ZjCwV18wwaOiiSsip1KQsLjiIliCL6BCQ47gnfKbE9gsP/0QpvWni32cpeE2e7mSKZgpQCzIBYH+jqawsDkkjH0py+sgqHSzIoBIbt39v4CTJkrdmyK1syUsyitUMNhakiPs3Toial4rKNpvM8z1upRoTzb1xqnodhqhZ3LH/MF+nfGtoSiKwLE5ANoTS4mp+WeyH9RW47VXoBL3msl4TvHTLIKso8sdiuxhf6WtN2D628l5Ip5aXEitxIVJKEazQAXkPFBNVrMSnYrShQd/9NBldWFvnXLKyge8mCqy1acjVdagvgOfZwqUTB3N92iVQyCWM0st0voR57VsAjxaMKTdTttWq9b9Fd0caOlNEKRekbVnIr+ht4NJ4YqJ0U8qk2tiBQuLyVJ1CGn5jHIuOLUsylA783bDTXRhIwMAGRnA1vc7mP0AwXw/hqtp7qRflXZbc9qLEHl/W9gAiePVdD7XfoSQ3HzqfPKRd7YAGQPQR7G+7+upaSuptGH/Z4IO+c2SBPOOIv4WpNfxL93QwsQ0I5jYnQfsEVDyKUJb27P3Ere/xEj0CdF9toahXpldrRjaWbr93OecK72PA4xJXIdE5ExvsiIVq0QsJ0rEDQqz08X8qDUkVKlEB9J/HtNuS/4kKGSaVJuN0dGpStoMOnGRL8L2HU0mbBi3kV8oVxRd9tNk4ZfyuBKcSEHNq2/SZkNB36YXboVznpSiFnGGQ4xps5DXAxFe6ke8C7um0NZRqdelxgyEfHrY6GpMqfImj3ri1UkowyXpxjT0cUL9B4b/9q/dTQmA8WWWqESuUjFkkuidLUfLCm3nwW7QmqpknX7eQ9D4DRgNsU5acWHE/kHATF7vdcL2AmJT8ozul3nm/BCyENKhjED96kRyAY8hczOaLl4K6HhXpjaZTm+I2nHZUL0f//yvbaIPzRuvXkUiBryF4HgpJvVcEsbQQu5CdZ3ADo8cN2QjjySsX80ZmYyvcMtkYL6CTeAZ1oN7yykX5F/XbHoTphjYxdsAFXqv/wpKLZx3dG8zWvFmyp09ekMfFoNIviebxB6fV7e00tENcX1CpPOeqj6fZyiT64luzIWYV6FELa29KPmozqZZJuj2EJR0oeJvgctv8ZGQ2ChmZ2XSLD4aQX8pqu4TbuEkw0bhrfVxzluAURoAydxlet2QFBBpb292y4sUsawk1vzFfI97+s8RGPMB0nL0ApblSIfeFKtIewo9lI9cJhqQ93c1CZtjaKyBYMpmQAWvZkoREt0MhzTGFxKTVTqZCy04XsYdyi10KXa1w2lez+pY4syIA13WU7n5WMqicfKFNtLxYlPPH1FDffkGeurM8juakk+JZ5DPFdA8oiUUXH/q1qrWK+g3WwK5YN2qOLfLoOhv1qO67/hd8DnygqC8eL0UFfbrTwklnSC9zpVi5oNdcU8KKtzpUEnVtMZiy3qFOc9s0MOWMnBbX8yW3eR3FwibdDbvCTu98f1F/4rT+To4iLD6x4ZCx1uFF8bDNMSfvfwyNODb8nPA5R7VXBXnz6YrU2UAn5CodpGDZe7IAiA0Q86lZ89CDx7l0YEwmj5TKxRgzMYk5Pl6wy6MwwEwqpi9rQ6/jmTkg+CllABITiI9lNMutDMjoV0tZpL6HT5IDG4q+Sp6aweb2l3fbfwkM6hUqs/wLSs1GULqnBowtjwSSUoxX5yf5BHKjjMA/mYsF3ZgEhUZ4zUEmUtXrOLFBznmNx/KRFnjMfmbopBNpTuuvIVgQtnav4ln0W7gJjdys4Ow1A7ZUb6DazAFEWdICpKNim4je//4dOMaYA0XnsB38ExKk3DlnYJ8L1Jwk3z7UvGxuQvZ80OOTawkXZFDwxQdd46kwYDkBxGqLzQ9nTkz19Vt3TOahVmEHpQnzUrm9prQFKeqQrcr7y5fM5JNxwj0uM/905oSmEM5wZmnOJAteZui43LDklkY7LF3nn18Z71x2/TOKMHkmnkMQXiwuiOeOSt+MUnXBQWA179Iyj0wAmuBhqAK+1YkOYfrRy26xXqnvSIL0E/pyNvaxfo27LDeZh0cGxqNHaCwHL+1qHa+hiyL2go0HPNgRgOLrHoz6p0aQOW7r3SHjQ+nnWLGNmBQE6AnJEEFiy9RAPOAYTHve/TuOGhk7+PLhr5ur6+v1QUQIQZgSZQOWThn3zcpf3n32rStVIldHYqMslguZP0c60e4oY0oHx+b6JS2bdBqh3FuTgYjQNCydaj/0/5JX0ITcYXMt3xAxDbPO+TkxyZoq9ZvTxun00PjNtCNM1XBsTzQ9Z8jtD46eAlX1udLmwiVoWFvNhAaM9Gn8bhKHpL9NygJBtZ5D5vHoIaeFfXkLmaTAJvQQhm+ObDv+s4Nc6CGWHuDhAJPDBMi/fFvES+4hw8YBLZ3qJdpGVborKbBZu2mN9Lkc5gdi42iFl27dHrl6vJgpYH7/ruDZ6U9IrRlNiqjPvJReSjdTCcIaF4e47SMYfnnMhd6AJd5bTUOJA+l/S8m0k6xmZ3XrwsZAQoQ2VMgUIKcTLOB/29YRvZBOfhf8ZLM2zeDUCPkIOH1eq3/vDg+4txnpr/a7oH/A5xApBbjhXbVoOpx0tshk3taTs3Fe+HPan4/7w2ycbVEVv66Mrd51XBPXH19ACiwGwx82lA2fLUwg7RK2nmrze+hE+1WOTeifrIQeRmfQA2kEuvwj4wFzKys1ZB9XYEfEPKmIo807HeYZG7j3E3leLlF3dOTER6E959z0bd11FqQAJ8kNwF9msZ6CclBcPBMvMTSfB2GQdJ53HQukZX+UkH0iErV4sVpqZKqdXAPnaur7gj52Kjeq0tQScz7rzDS85ZIrnhko8e0ki6cbfEnbmfsfCJni59ed6402qgwUCLoFvrMMfjLe3aJt0DP+TCeSEC8qcsDlfP1hbVqKQ/NXJsgUWsQJ0nv1J0gL47cY30pT4bO1ncqPMu3EFQaPoEIwRHxxMpx1xR0OjE5Gm0EIfQ4mmYFCMBrNMwe2wr82q8MoEJKV3q/CspUYuI2NiZLAjsnpXDMnal2JyokoBKq5Tog6RjyJSM/aEZgM/gUy2f/YSoVmF0Abx2T7iiN6ClPgJRiSlQJ1vvUFQNwBfKzqUOMsJh/Jg0QGnZtirCMICzn1BtP5R0KWaoPzWTWr9BLrUzDbUIsxaY0qceMai1dW+nVAYVMNf7Vvg71ARBrDXmxo86CeLnpXCxBv3epyKz0oglYJGZBvvtbzLQJLwuX1sIfmXF2Gk0ePrCwOPmu6Os8GCnM6aCYZzIaHMgW4vPLXU9w8LUXX2uE0LbZfeh7nEqVqFDtNAJ1wPsibzzlNXcgLhwtmRJSbFpxfegNTr5q+fIzavJER3SwElrr1pHtYKZDnsQ7FvGz4leA788lfjafpbWKscwy8XKFcMkZnWjL/iPuhkwxr64zz0J7s7toMGQ4tqWD9dh+AmTWZi0pyM1ytaM52E4V7LnL7UzpaO1uNLfQb3nkuw1cwQyHTQobqZd+ICkW7g0YGGwospFq5aDFgyZvRFz1mmZXKagnVZzU9m3Z+KC1EkHWK+Tlz8uiRhnde8XupS5EL0qbgt3k8pjKGGZcjBaag5HmhjtkYQ6USDfZZrEHI/4J6sqBFGIRrZ/9hgA9W/dMWBTguevhBIc9cp933EhvFJagmxP/0cXoVvThoxNZk6k+e+AHv84izR+hVTIbcryTMHz/iiLN0MOLWWefwFArTA75ODVxA7CnC4S3EhvcN0gteaZkEp7j5B07e1gg7VOWN9Q7OXE6RF9btZ1bNkaQ3/uOLrWrwZEqwLAJ2oD2TVrlrXZ5noZlkcHK10P1lt+nnTZ7iGKF5/GMUAacfdC2qlAWC9HEbEPJi1jWkAenu9ZAUKfp/9dPEKG8pRobPnE+6WVRO5UghYqv+8Sg0=
`pragma protect end_data_block
`pragma protect digest_block
104f666a82098a37445ba247a6a9b97425f85d0ba7ec0d9fd5d38097336f8f39
`pragma protect end_digest_block
`pragma protect end_protected
