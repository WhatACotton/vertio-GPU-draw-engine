`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
HEewWruckcHJ7XZGk/kko2G0SzxO5HgfIN52Es37FWpSL3ZIL/jyUHFp0eayzDZi3Lw9CFGJtTV/O90aqWHc/t+fEZGgkeRJ7vzjxgBB1wqgeQ+W/hk3tv0DlSpMj/Q95yAqcqQTw5HayULOQ1r64MZk4xtGhBN8gsuGH2mOgvnDNYPm8dZ4vYO5U+3w5BdfEynuVJgkVmvL7ytMcYCdLP6RTmvDi66iczQw810qGen/IBlKYTElh/FvmVoR89scr8CMeTX467CRJ8R4/Rz/F7ZXxXETu8YTaPO2NrkH5mdebH0u27CrJTx1z2OgVnzQrvhg9wZUSvWgYv/TxP3/ID8wtVJSlxy3UIEbZrsffYaLhCXIO+b/Mh6a3TuU77CknPbKsJ2ajZl4Smrpzt/kwB7yO3IYYCXzqFolQDdBXrlFzgF7isQZpZCZtM2K41kkO6yn4KOLacwnuHohZumWZchW5s1c6j11N+sRgbdeXR976EzaZDf8LtIPCgyCfeoPNqqdXGnYlbYwn+JXzxLQNks40UR5TlWat263GYGvp9hJmom+rYJ1ohHiUqzGznYiYVUbZ+JGgHU730OX9CPqvg71en1dMrvGOye6bMO4ZwoM/mJEJdrWw9uK95WG/DQCJTwm+FwUzr9Vm44GCi4g4QDhuUFduCEZZd+PHw9oBxNqIjjt+g4FgJMjcy5DbRyAngGqQNN8116F5yM25dOcgS/UpoPJeyeDFld3OS6qmaQbKOIKgRhe9yLPNGRLauE1zSGcl2jWU6zPrP9hDLW0otX6S+JQAHPrePv2KFrIPQ0xp2TFl09OmZ2VROXfOVwYh9rx+N76cWViOmeKRWrMXX3cBio8RDnajNvC8xPhd81LEXF2VobSPj8NhVvp0+IWLV3Y0FJv5Do03vBPGhpw0gRl7eOWlgAXGNvzWiISzfLbHd6q8Bt5E4h67rHS2Dj3kXEQZmsoB7lrl7J0sjnaXOiyNNgfSlX9JlcE/GOJJEA77Nm7N8oodvBAOfCpeyTzfc+Ti8bxpYEYCs1pLyrDiWZZ899W0xarXrtA9r9XIErfHw1CZF5NrX6tie8GObuBRKEYseJxMJ9oRxAbLEHb7KOyJ98Ww+3ncN1m4HehMEpZzPyYdh/uLGM53DbiBCn9QDf+AmVaaKHGle3NGPO4JMLxjhRT0jijUlSgxoovgUkOYE5Br38b2zVdZ/tvMjQjZ3DVGYf7Z/mscvhv80Hz6DSI8a+Z0f2+sbqYb1vGGfmv7gQ0e8N5fopLGEnl8XaeQP+UlVZcO5s7woeHbG2AQkQf/JpuigUNxC1zD1OrP26fuenzaAMA8iDDz5HUsY+NNbBW/aXYSTG/3eP9vXfIR3vnBp5NhjWQGBhhy/xv679b+QpWRQEKzl9nmDXOZm0F6dtXrUq7oT04UlHeyPiKuUthK3ntxw4AJdFGd465TZraUreBARBMmfUeRkV2t8j7SRWw1aSpvQpOp3v9mA2NBT3T4Ba/Pd5uXDD5ZNlVRKHeBAtsOhazeOOxq7IkvSiBBHa0J1j7DTtL3CteqyU3v/olbS1AOt1qTITAl0TbJVUNMevP6QeJ/x9KxnG67GtLt2GqR1Ml1GIQDWk8bXsLoBZ8AU965/jhhxg+MXNlPAvwJMZ2s4NbxFfeoGx7N/WGhsI47XfmpQXxxAdttLOvRzMKEobWvcq/EMv65CzBWMugb0BybnL7mmmtnHgQh+DZ4xS7Vrpb9m2oWcKjCUq68HiQvPTg+f3JKvrMP/jLG2mVccaTLgxXF6z+gaDgyR20xUP+85y1Jm3Sa3GzULfz+OBL+SyME+4ojS6Y3cIaHVQwsjOQPmRm5OJmBkb2Hi7bXsHfh/UwpEm236Vd0VzKniDQRDxmko9kki/mH6Uzn/dZxGAWtKbBqjq78guPShGP9nsHE8PjTJSoOff3sUB9k0TUaTPoOWoPcZVSA5A62Bg7J3RVVtHd8xZNor+fa3jKg2k/BxfHjzLeNxk0URAsc2lSQyE0AJiSSsz2g45wTZG0/GW34zg/qXKf/azhDkQgt392FctVdenkkumRwvuzy2Ww0Cb66O7RxycD0dalyaUqgij79eEx8TUyJ0r/E6UX9jvUC6jLic6ZycpJXOHfKicSll9uiEP0r5FNz9UuvN2gt4hwtg8aN5+ebjl3k9YmabRhjS5AH0ELiq4G6qOQgwIj4BtdSVzD4aIUt7E6SuNClDlPslATjkz5DTnG7QIkZmS3RZkWsM2CZSykJ0vzmQf4OFtGkJ9LV1lAQIhdMQnr47gjngluGGuKDlu11Fmy/Sy/w+uC1DRhrv+HFn3YAne3n567Z39tabyZyhr8UbdbDv8ckJWQ7Osh6C++DNCbWMF/Kx1cCzFalE9FCxpe9iqjmXVPXFd/oHXqavHhw7c71EJFJtOiPCznyEFo0flz44h+fT/BgahC6rrDxKzIj6uzWUqAVec50jwkaIs9e2m93gDxHA/h6COIDNAnjzX49tbA0D/QjbQvMI3q1xmUE4BqJxQ/LoLym1mYBdieKoyPNzYipt/Fz0SPkjyKgALK/DbJwNkyTIz8JvP9nQNPRGllnM9AEaIIkmKOQl7+8NBoD7rcZXDWd8hqKYi/Qrlynh5faT6CI35TJi3gT5OQu3SPEgzX9mde+nuemjyXx+T/tToG7UcfBja9Sq8w6AgIeCWlSBUxANjuALQDHnSUMIc4DmZNLh2VecU1/nIAzKhq75EXiXu1UjUnFTTzLAAJVvZcOHH0qbrCVceoKcB+ytSeskyD76NlSlS7Od0vX1h9fPBufA9pS0o0l0BZeOfkVi62kPWc2G/DWK4vKd5AFXkh1B8tOmlLveZ1m/1iu28RzPZGdLKYRPGKRBh+jzNCrggi4IFo815IgI+DI7mkI8kRooozZy92Wcw37AdQBt2F9t+djBHzT1Zh0Q8EXsMuRekpkGh5YHkOqUwe9QBKE7vDNVyFMNJtf+NPqB5+9NBisvkPJDQuH7CyYxYwHile7j94/MN8et99fF90tz/CWdbuue1RtethXvFQ3G1Q7zaO7pP+9IRsFn3fIbNu5EYYOqdN1/R2m9Bh3pLLex25k52gXTD6gHTwG9dOUZ7jHgNESC5EXlzXanV8OWJBwWGo2rvLy395mmRNxgQfvAHV1UVuI7DepfjnsYnjfe71U5ynKV5QV2DseLsp8dfGPpyJmmBiUdM/CRSQT7B7gJtJ+KyilmDTU/jqFL0gq31MEMmkwsoHnxt2HZVzN9wsSGrPSEEmzVTZlFjCXPpT1qVH3is9pFkjO3Gk7jN9nQ91K7SwKA/24Fmi2HxKmHXrxlg1wLvbRP/PwOAAJUXOUQoQn2klZfWNH2gD5p1xetjgt5dp9wmdmKQQYjvd+dIAzsFJIg8zzLc0cwzVKfrenTIRWLrcZV8hksbvsEvziulhQ1ieJZkBmoQKnVYqs8gVK3ktRj1SgtxFfZzF4gt0vQwQEe1GRLeei0LOYNq6MmhL/CWVtO6b6ppri6QJgLmB6mgL0TzrImM25e6rvhVcoFbBjsgn3ZQoZvzc20kZfmq9P/dVtQZwZje8ssvDVmZ8HNpHTNVe3Bg7lFxv1ouc9Caq4Kqt3fTBCW0MPxzwFYAAuzBEplYSi0pk1SKXSRJGAIM56YsHtxOwwnUowgAuxQsjH4PfgRAbJIYgxDXZyU1O4vgbDKHKU76HaR/zr1iYRKWD1I6HKXGi0pqZV6kwrH+8VI1er6Fc6PRbBf/OhcsAUwVHwyHx0+B+1SYug0F4Q1dqQyzrI+qHIfp3mFA0VEexg5wSxxKmYlWfuvwE//FGA/tMOwW0tWQJHRQNcATlleum7gRyVeXIe7mzKewydI3qpKgAYHni74LDmxMJezkGybcjvP5OHkeoU1vFNCHXQ6PnXH1hj7caLIV7hVnUgElWMmDt4tFvg9SDuuq2VC//+BF6B1TLuxJqrQv+XNBxl1prWoiDubZmftw5Js90cA5E7vpML+8gl6BULUMBxwJZ6pimMxcebh/gioVn/ZbLVH5XJzFfAB2ztDtbk1MJET5iQSeNuR9nN5MRPQKxZpbA0CA7LY74UYtzVjuuZzKF9+X8T2nzNoeKIBrKncmAuoVfjQIrM6T0/cOj6eHWydO+AUUc+Ocy+aOAbrErKH9dlfhWNYGgOyDvDoZcIrT+ubydRVoRn3SkHxUX+5yk0Ai+493ncUZsUEpMZJcqBeQnlgZn+DS6caZlX76zMsxoWvKPzE4HWhn+X/U65nt2sRUndDwkUWZ8jhtyuv4XTLfkIHTV4tSEUVgRr6ezCpENGd2/sKdEjVNruyV+H03rX13r+XrfRJly6YT38VBnkJt83Oub+WNR6BR+FTOwfhMX6v/I5siqpXcGwZ0tQUoIgB775kc5Pngy+4cRADjXS+XuvTgTvX3mn+X2Gpa3rVoaGfoM1AFwIA8M8W815UHsjbRk+mHXLyZsRA72XIo/skO/1dDU/T/BT5vpG3ybbruMsYKBx5MJPb4y3HcRdbBne6iIEUpyhvfwFA+G9hrtyRLntOI6JOe+VIPYl6Ujqxx9d+okLDJcCblXCOI0QI7v5I0RtlEFhwwhFECp83VNW2GsPiQCjZIRksKskUinMB0p8l2rHmbgwHb2aDBBkiHLmTsfEu1U3cJTWUkTtLagKb8IoKC8ynzOPfqPy4MJMdrkZxS78gZE9DTWCttkYYZVJs32hFjrQgcvPnH6pN7kahBAJy2pDpm0wPz1JMuwVzt0FswnoZYfbo6vOiYdppW1yri0veDfczRnlVWIa5XPTV5X5obDnJAAYf67fDwOY8yl58IcJ1HCiR0aHybHxvNEB7dKk4bWOEl9zM6x2r5ymwe7y9HxqujUdH9OemUDWepTkHyLdRZIQybJLLaB6xoUn5b60TtBeCebFHsSTGWq585I9llD6MaNaMlZY18gH0iRyzllcekRIo5Kr6KaFk6dIPkn+illYVbxKjL7LHNZW63jjMDLSXxBvNWshGzrSwCFXVbPg2uwFHLjsPJavmYkcoM/X33gbC7+TL64+0a+mG/tjLD1w9fH4teSTI55oJO+uGqL/6LEulp0cKrZzo1idvUFXabP+bdx5a5jd58v1Xb58WVBAJxJqT7WR+NeqIWXwPKRhjwsyaoV/VBhdnhbOiL+1I5ptZHTnHxgz6OO2NuiqFoPQ0dthtuccJB2YOx8ArQHEU4+i3BZW/OQbkho0SuokzAGa8eEruzDE9SCBTbodG6z799BaT768UjTCVAWOdAnCEsVJLyVPq89d/z19j08tY3S/EKbE7eJRb8usR4YLdydVV2Aj5ZndttJvECXL7GffWQcEba4HABeXhYLutt1GXMQUBd4MEgdmg2CNQ2mJ5wAwjdoVU8sVsaDXqzm1INObJ/tHlcmixcqu3Q9H4lKierS/Gi/Bx3Xowiq/ZgQ0bZbaN+A4yNq2wRKyvyhXGdEnfiIIrtEOrLwY+Uit7D9bi0eEsY3GNiMc+F4ThhU3E3QrAsJykuhP/3MSjdyqIRr8pi3tiq4u29/fRqP5bdVPd85jkp+n+xyV+e6e+tytZ/dcJLjVteM8dh9I7hykwPDPS7iHpjtPO+y602zOsBPhj8zs3RYYXVmrRyCqt6wJqv2j2kXJZ8OlMZCkuvcOdhBGjN7yaeYc4tzh1YLh7fDuf4wxNxfg7T2Jt5ds2XK2luiBcPRDnWMknkLJNBUHmTi49z0FSK+n7mgtDN+srkjR1sZwQMjlD34ei/EKaMy64HxmmjLkuVVBlvZPivFjBVZVfZqzpuMwCa0HD3ANTI6P31TotwdBKuRwW0PSfbEu25ywRWfRmtr34kOdxsfcEjCHNbpPy8gsN+XJN/AUyF3dT0pLSFlzUFoRTSoXRhcSUqTOSdHK6eptw8J3Pf5nEgA86JjTKcxAmsTy7Tlq6YN6kO1SOWN/B4m4y1Kg57LnNdbyeE6GmopybNzPJYxJzNU4CHccRtWB4zVoJA+EZOdtY6/Ek7pVTPiQ8skSTt8FGwMCMPH7u6DRnO5Bl7Kbigfxx0IeHK8UMX64ZXWuhSGvSIwKh77CetieMIH+1jnpgTY9u20P3mFvWOb0njsLqPbQk9CrHl5BX8pSOi/Vxq/98W4RWBZwT8jR708jYAWoJ6QGnHz1cbCky8eXCWAo1endOXSxh2pS6NIjz2D2gfMZCWamBPPTMkPYrFzYCABe+8m9vVxfBKiBVJosnoTDgWNoIGt/4lCldupfmfyBZA+naNwrIHUIgyqStB9r6NdjmYT+W3JbBB49WolPsgzCKnY2wi6MdNUDZp0GRTyqqz+/HR0EZDpYZdngym9Zlcwwn1O3jfrMKSV72pWoIYumAdlf2YENx6sLaQOFnLtI/gias8mTp4TOg+ihJmmhQQNh/3AVC7tzQ7ZlRLmjcCb4wyeGleOPY+kXGphK0yejLCdjl2FfvnmUM7x5RpyUBCsGUeKdkznFU2s89XC229ucbgegVlWPEBH9W6rSpR/BCzzJkVKbQ2moeIr4mZb7Jd1lBWxgFllW5N+f4XvMo7irANF3Dh2RsPqSVZDCLk4QVXOKqDpoX7cTThnUx6y84HoBHxhHaP+czqBz2lJ5ng5d1eYmICZU0P7o4MLJgdb2P9FNT4x1O9v5jRgbWo2Q6CAmiAOl9ZeE4OxDHztqVBvbhe9oeerW8bL9JofA54ZaIHv8/Dx45ZG47/EpHHooNpzWRPgr83iBoFkDeu6hyMl5NLZkafuhNljCbh5SB0jdA65yXrGYlF22Z14ZSrid8iUMK7RgSzjE+r16IZg8sNZdEm72CLRVxGJjSepG7UN/qhCojE2Y96/8r2xX2KL+siENQ1K2EkYPE7jcfsVdAevDIXn1kCGHf7RSHPF3g6RkV/YSU8x5IYvRVjNCmWSbqD+OuoXjMdRNvw0mOLbpBbT83gME8MoeyPwT7reEYdcN+LZx/RaILJ3/KnboZTtXSEZ2M2DHlZUOSQgTWrmTX19EdHjSD7x1s16oXxJMRlhzwdtAcK/Up2/W8+t3i+xdwI8Jjm0z0GCKnTPg173Ou7wt7zLOVaLqUVhzT5ZFbR0XyGmLAJA38EE1Gntw5k1691f1perRXf8Of1dXYjw86ZkzrG+OS5UnkQ+OVyGIHLOAMJSKY0+SnMJj+iM+lH5D4fPKLNiK4Mgw6aWuYfvefqUgq+LW04T7P+mN4w6qHyBtJXHhAJPXlptm+5ruFpI4ubipXUlb+BruRrwMAKCXNSxvWeE8JH0ca+wi1kRqE+tXFNGKZpAqdn8CuqIn2UELjJg9L++3KJmZu/CDKUvw6HjjewDYd++8kQibRWyX210x20f8BPGDnyHZvRXpCcDB8vNjKdRDaAYKzzLv/Rv5UPjRXosXbvAsXlsRqDIhB5s6yxK9R0DGs/pdqlX6kgmusS0HKjqWp9b9vAenueF0rmZnP+tcC2qYAkMHcZpbA4RpFmRyiHg8iKW4niEqps6pa2vjCdMxHpRTf9ZlHM/JT//57cV/YT89MeCgYGpOAZFDi0A1KgXR/mUgc/LIhySGQUcoGyJR5Xr1NBXfpct3dMG4lHezQU9wHgugTZ8938Jl34eCiMffRZeOpbKpd6ARD+T255oP3RWa97InTzHKXwPyRAnhtXeUAV8NmC4Gettch4dN2tUEMecb+jAhZqsa8zMBI9nD642ByzQAAIHsasthNhE6fouWP9uDFihcjndxpSiECX6qGIqJhW2cfl2oYTVs+P1/Ixp0msFb9mhyFAqvJ2T/Ls6cosyXT7qjLWNUAIaVcx6QS6xCB4hLVnYxqLYNZKFZ6D5OkGKbe6OtExdYsHOE0KBLmtAEIpGX+Ti83gucOp0YCxC/R7G1niqYcn4pC6Fq/UZo7zA9Ta9Yb5zWQ1cqaACzhPwaCQvhk/o/Ta9hzg9w9pA6QK8Y2NbRmqNaSCO4LlUVbrT6f+hRE5mjCe8xjmtizHphY8eeEM6IRZZLgiUceZXLMEPYIt867rPaLkT7B0rduHKg6Cd8H0qet/DL3wZ17QA2YXs3tGs5sz6IrIwmDPFmXtN8QBaGJw270yqIoIH9kP7pLzNouBnPTy+bCDUIRpJ1J0ZdPbbcCs3S+08dEF4vCbe6vxolLWrqr/OXgvPj6OynPw+RHgog19lCtvT8ZHunXGD5smUofe9xxF54qF5OqT4XinTCeBrifP0YGM1L/R7fxvgsiD46SYjO8V75G0Tod0xqYRGD6jpxwHjuheiSZGckzB/Wj0V6AkNq/Hux1zdmOGqtj0ZAg1LSfYP2WGAqYHsaFllxqMKlLeVWXloFu+fkPdL44IZ57JOtYmoJMqgMqBF42mXUA34skZ8iQcA2yn5yJ2ZrCv40O5i8kr+UF4BsWAWeq7652ksS8CZtkUpd+OiIww0o9Knhjxq9KVeI4I994Fcl4c4CH7/02Z7dPHad6EoOpawgTrl3PjWUi/lCBrDtBMMd5DC9MvrPxXRG+momY4cLC1Np3Pdbse8HDT7SJCQ/aa22xUunCMLpqwPH+kC92fPCa2QAZaw/kbmHhYC+kg5yzqVHWyYVCTx7YOYNhUfTof/1RQbQ17288MNygo/oVk1SL2yDr7Ej7ZZ9Xx0CYZRhvJK+QbEmdaZ1T+IpONybA3VRgQZMEoirAysD6Xg7yd1DxxzmMjK2yA3UDdoHyjpGOFq04nkDipmvYD4CYj7aprIAhBBQIqAyK3Li/7RV4EjPVK415wPgKstg8jW0JEBcryXxArNzsjGc4c7kAairbHq1fl8QU3ypiD6OScaZ0q2AYZFe7rT1B3bJAPcwFqgP1myzvTtCdNjKn1EkmhnZXM+iY3tIvz6i9B0bJI+v6Pt7PnbyjbpUg2plWSLUHAOTHNObFvRpT2HmffS2xSnau8bMfGCrXtLk0TWGRsZHtfAB+9jnLoeC+JaP74JLOiyRCRRrD8ipKT1jOA9YdWnhKZXnAMyO66ZlhVmdAc3zhvoGg23y9x/AWzQs+izay8XCsgRQN/9FwX4s3TCdDYTLfuqosNYRVwcJyRqmlc0BP8ehyt3PoAZq1GImMFdRGyGAMCeWum1FtFrmdu26LjXiaNRC3w3O5vHyybOtDWjXYmoNqy/yCsi9ZySIoaHhdQTFR+YJi3c5BP4l22HvwWTWCN2VGM8867iSidjRobq8uzTfenwfUSEIy+44akDettyRY9802wFBUJDWJHx9qXToe8MNwS4AHDaxBjjW+ttU+76zFxGdYLNraTDoJVl4osGzc6VOqf55+D8F7sXYdJ7IfosQsSbS2HPHCPYNiHbICKHOv1DBBhXKcQf2IQ1YmBHNAozHn/RH3Vb+6BIlN5/tqNY5xj2T9BPm27z+He9Dt599mG+BbYr+HVoVsvisAWZWsoBg7XOxFwEBNxX0uMcVVDztwQIwvzg0gdCAva84qW6w9O5VoeNmTSkbj2+ZkHS88wWFHWUVLUP2uByORQ0ESR0Y0s7jMZKy8z+3Osq1/iRmzzEwGJh/Xmsyunq0bhja8zDLMZl4yvI4JKtbQ1eXKFeqBEALlJwvzydGfB9BZC+HCmsih23IHTy6RHrckZ49BrwTvMqyUbZSFkSd6SaiX5TfLIsWgcayubLRSwAO01tNS3FcyFCAgt3eVWX1Nd2mBh15R2me1a4g/jwKxdYs2T8tK85bGyjE2KgkGBx1nsjiRfwLySuXSRhwie5jZdhK8sUk5pCphiLhgH5I2OXY7fPR2/jJVUFJNIl/V3WU3N/I93pSFVS6YAALiB5tllVi890Mgw7DssqL9ZIu1+3CTm0O0OeSBFVB0HR2dCMtarDYYX1IVw8i0KaTBB5uyCdvtQUkUMmPN8JcRtWuDpgFOHymxKTdZ+MKIHnbioFOGzDvWMpFX5/qJN/PUO9lLDTZqqL6KsdgoT92Qxf+dJ4JEtaN88bm8G4pQiOjtfDwr1LwG1jG/wb3K2Nza2Rco6t3opmH7CSzJtFRmSkMg28GbyM0HOr6AYPDm48e2Bj3clc9ALXKwSBbXqg6stFhnllvtdQjh3hU+oFOWLTL8vz78TDiDUBmtLuO53giB9b2qk4WjliNZQRZL7mLb7btxQ3filv1ayGbV1jyL14MB8SF8fbP4ZchyIouU8usEXHWDHWnQdFzO/PyvA9nYpu3WPlBNIv2cDHsV62WoanH1YmLXI4ViST0MAmKvt9gYHIxF9IGY6Tc/+EWxV1xU91mq9dw9QSKufmmvJjJN4cvNsre/JC87F7m3rWmrt3Z5YymnmHcLgFc0nkLj8DcLO7YuTSjHZc6Zp7wAvYv2ghzJKlbiDwa1Gzx16CQ3Az8K8KxJaYM86kX7bvZ3H3WGqpLXRlPo2NukIKNlnuGuFcRnmydmFCQUIIFcBbUIPCKFi6qx5t1Egj75lsP0eFeXax7jX3nFpdVnVIrp7sO7yusojCEGJxfLA9RXgSQvsayRzKZT8wqf0An683teNWPbBRYLezMdOSPrYQPDGB1DD8mmfUwbZKHW1ywxbOAUVSB9LAKG580hiBgvLjKCVsquo3FPWoiCIu3AubgF6pDz6N+6dvVD+aDymVqhkqJ1LMkaIYK/Undz7Sk0yphJBdAQjORTRZpWTnJUJ6zGDWrFssMkIxlHQsfVo2L8xMGzwjEdVnG4+YiDdsmtXhfid0eDSnESwHttf3bQKizWwgOPCkpMw2MWjSpw1leqs43dq+LjQ1rTCOMGBiCUTf9Y2vn2jrDAh802xSEKDh7VlECoSsqifJmIqWFcdY4Jg0uRoHW9Um42Pglz99eOsomTPRFWogjZt2riKwpwMxbCMgGbSvCPg4AXfR7d5e0ww+5mN4P1dOAK92lCquS+4h9oPC1GGgUvt0AkSeteB82CeAQkH8hT1J8hMaA3+UyXLQNvlIXwa3zBA19NevnmIjWTFme6lmtpq0Wj/mVjRGk2SzKM9EXdkufwkXmtH5U9r0791gKCi/yMTWXXjSYUeTvp4bNIrVZ+ZrDBQJQE2553Zk2FZfCJkMOkDG7lajwN4Zps1rOQAhv4oKdIl8oUu/di86ggsAb9RfxjKeo70/hhcqPIRixbbyCafRQz2mXZgia8rGDsfRgCBLgbHuzd25kFkng9mSVohjUT2egRsQIgqYNLeqDPJKdhuDWeVTmerkWyW0cRS6ZhqiUnpM9T+6NbV3yGSQHGH/+RTV8/ONAZ2LKI8g3pG97PVxXfW+HJOahE1WvAYU0p6vNcItfdtQfOGNTbN1WVRsAl0fTmBEnWndvm4Jmlq4Zaam9KZPg9TazLpjMB/zP0ZsaPaVAxFk0RKFTFL7DW8CSnpnT/dVsIRIVP5UFTjLHHgXEwMHCNkfNQkfH+FL683Fvlr/tIbJBylR9C7tLR2j+dpSXD0SYNwbfJ2jdGqZU84heBEobON19fCQAFoaDrgiqlfJtWR7Ojy3gYVmRhL0ubJ2jSPA0NGpVFieOh//1ASrEfan0XGmsD4Xw8zoiOPb5vY92qK1eL9EzkpPYW5fFjiTNfuzyqllExkYjV2Wr946qjyxu5Hk7XFoO2sakkMgzdyWZ+SFSgpKxaJoLOe3SGTZ4Fzqvg+p/pPBPu4rKBDmKXCdTRdoSjpudGOWpCggfm8LdZ+AhB0O1+YGppeXhJc7AEAw9jhhJKDSuoLvaAbnRhOOjl8XxDnzTMqnS1bfk/71UdW6M5kNNyFqIjTTqQPSObP7D/eEiJO1LyqWtn8dlm9goFLmse4r1glavM0BL+hrepuqBLlwq2MdxUX416poYXSEPwq9KnOaEY/0NaKYE50+muJtVNgp1h9ECu9LL1PvdXiAPyJHRJypmEkS3462cdAVIoeAnvX5p1mZIJ7aKkcE8gBcPSC81HlzhqG20iFUT7GMqEtCQSilDUcO7A8/k9kRr0gS9OzUdGlvmOogrHfZ+sOa40gNjVrbIyEQeaenlRibeIVLMCywuuQzKy2UnxAKyv58EzipT1nmxH37Svrg9+sUb5HJORqddyUiVhaqd6LUXT/GUm6BhOiYtTrRUgMWKmMlhmpqkE2dPKX3r7mP3pBnI+L//RtPvsahy915q2OVtf7dj30IB21uFAHJv9Cr8GA+jm/TDHXqPuOnbVrPsbg+ONOWfPk7Oxk09d0gUYdfDSmKreishurY4RwniCOYwuH4DdndefNEZ08x6HWA+ME6v7jyyHyu9xLsxI+87HKB9AyT47kGl5kFJSSb+nQdB4KVt/nRz6BJ35bkz3ztLuXCqnaWpgHpAXuxzoUMaVSKb/jBO4Qs/Apj1ZZZwmnQyfQQcm0WXoWPVFZsMAEzYisbm7MXadvr7muAwM6K4s/x3+LXluuZcQucdgEmPE6gZFtoLV6RVyq5KlakgByi2cm5QZ0Qdkm09Yn5ppPrUnuYnhd2YlZg6LCrsNzpEmcV27E5xOPAyX/FdxIIkcbCBfpr2dkEiv1fkyPNGk41yEd3notLAeeXFDGMFWTBbnjj88don7R19YLJAXmrqeGrVDgr/JoQ1yJeoyNigQ5b//zhcVe0+XH+welrPb5XKzHaXR5kxGEDOWFjpmp/G5OFOZYL5cb13x04MHJYPifUktW8l3Fyqkr8KDMkYXr0Tv37MzKW9xaICOfhYcGgQ6k4pt4ogQBhY6cV5f+aCjc+deL+m8KwKierz/TI5/j1uKfQC0tF7Pde8aoqmWWWYYjuCONV8S6DnxYAOCwBfGvL3uAvwx1GY3PeDe/azNxMbTN4V7Lhli0Xy7NyKSNmKzJIHGxRmRoBWocO0k4n70vbzLNAmnUxCxfICgMfc8xrCBcgLCI9g0oWKmNtKEgktiQSyg8U61A7n7CngDc4E9OOWMtZlSsnma5kHkhjZFETCLAGKKS6Z0kJ6W6NXlfjCxb2JrIMyOahTLxx/lwtmW+E5BqAou4XcE5MTmdC8fcbV8i0e9q/HLZ/lWKeU8b6p3QjA73aR6e207vQw7o8FOUC9AC3BK+nsnsb0XjEgvnatRMPBYycwHX1gkjJAW3W9mtrYEHppyVqpyARjOycn/W9q7JScvZzZNB0DyfMvPjCkB3YIsnCcAcDLM+7Omn1GNxzRqikf7xUpHTmwOgOFv/BxcqS/zUM9H5hmxFxnPw0oHKYDrNW/QBpxU400V0eA6OWJLeWvhIP5hLvkJK/kdYJ/N0DUL14I4zMJf7nwGiIxRt4yXK4zs1MwTLu5XkSPeTXsso0iYc+v+XFW480zMPHe1Yj7/9kYNNkbltxqwoFP33k0bvphFZ/yLeY92l0ZQeQEyWO242OIWmX3UMsfeYfqad4UJ2+IEW1NO7nwJv6JvtMTOnA8cGg91MKw+4sAoXrFerjLXA8MXGt34XI1i5p7zU3erJkbQq6pvD2vDg2fvzY6ju2An2kvTU63+f9AZZWlvuV16rfoqkhp7XVHcTndknt4Ozv6sAqGM7XQhEtI7hyV1okGJAmlYSDSh6PnwMmb1vY7GaWams0sdA5QffoRlZcAsAndzCxMupDC979/VI8sViEd6RVs1eMQoD63HSWVRmtZfr65O0VhnqBkJc6dg0kCuPcC31tGaHycowgjw8hyvJI64Cho0GtHbbiPDGunEQNd7RsfD7IGeJEptBImeadY1+761/F69Q1swZTJ8POm7/wqBbeosxuVMkYu2IAQfzu3TLe1xyAEkvo8NYuHW4LwtfUEF+jWi1z8Rtkl6/EkCP1ku7ciHbL5ReQtsoFggExOnltKyFtNgvm9GHBHqjGNbKv8AEvpJ/g8Q0fuFC/aatScPB+svJORV3EQIVo6Q6M2GiBVDiAsBlVF5JIJMn1PWir8iqPzLUwuaaGWwyiqu/63ArCZZOctZkEU+IW9HNEY8qWe00oXoZjgIL/CFsvUCnutvIQ3H8VVdrTh/9ulkfW1MFrqsPoR4sxdO8bXiF9VTdeh9YXwBtHdbdivwSOjpJ8qpHPM2ib75+5bPEUUAK5piSHb0Y7kGbhgAf66YVThiZQVLkB6AjkKT/H6nQV27M1d80RHMJRadZFDSJPEIfvXy2JlheAQznGkJgSKNQVMAijgcGKRPvuupM3m5knaaklyLMpUzlrl/weL0bg9KhHydTohlLldBlmmS7LgA4Y08U8GCBfnf/W9QiAH1s9gzWMfMUvx88FSCQP+vAKEUVWu1r0Rc3L3lF3O1HN5gV7HWu7BfwPlQmmoyrzRyo3BvVDKIJngbvob5INgW/EkuEg7n/RgKqKzfOksJW3trlXHb+Cuhvu/5JW09s5CdLAn0wYdp6IbcGwNvXShPFR8gpckY5g3urjg7wfwBfkMJIHSESn2G59K7DvGd1Cku6zwySV+rth3ktJ/jqxgNZedcEnQfbp0KhjKCeQbxt2SPdGIMh+LgMsRUhkUSZdX6v1hbOhnQ1q6Uounno0VwBep8LEW7+5aCxGo/4HkA2JM9t9xHMEBbDWZ2WsqbY9YrzlSgJLndaF/+rK8upFYpvllqQLF4qr5bmRnf/ATFHOmWB4s/k7eewWDjtO5+20igPM4eOPseGto12zJFcmh46tws0giJR9ihGJyow4PVbtTArFQJPEEvvgi2gZAWvg88f0TlAeY3X6gDlmeZddW5NtPTm02vPDUqrjHCCV00ymUgEaOqc56uehgaC9c/BYBBgyTRSfYlaL0VGETXXE/ZgyxyyE375Do9oOQZKwrAnwSMrahn6DafbuYRHKhc8tAjpdtixcXR+HMPUxPlqlUY85zFRMGoNHGBUzm5Ft1ZyIVSDzj+q3p/+tgB4lM6S2Y7eEA2Iuc2Qr8+SraopQhlWLZ8LBQNzM8ML1COEa/wCRNlKKzH7D9i/lZ7E8KlR7WTxq/mV1VtsByzRnGGD5fKSsH3CV8QQ88D3UN53LFMbeTAFije++YAYzV0B0piSfkwPOnjoGvMy62gFO4qOush/XGRRbx/HLNRUnGPKemfw1DxhDO4bBN4qi1qm7uKZZam4fYj5Bm6BYGg3S3q3lDjY0YkmQXlMPavK3f8KuRC4G1OJWgnf4CO0mwMVwajCzQzGmrIiDbGO8vc0zInunEiuBemSYUZiNp8Eem4QszRA/7P4NChF3AojYh0iFsu2fkQguLoAb57A532yTG6LC5Hlh1XYfW9ugU9ZHZDnN1MlSpdLL0fP3mk7d4+AwBC7TxXduu84ccb9b6PkppSYsK0j9AcvhH19xLjJe7uGVRFaRs+K8q2hJvif3VBF0HzPSdka8NPeaMIVyuVToeRyzzK8JImlus1gszGTV8hEttj2eiGwiP6E7PO8OHdCWbzVS58Xvi+ZyRnyIxIcMh33kBlq3T/VdG7vK2xQ5S9w2vUl82xAPj+qZWuhQrz81soK+plxafftl6JtliB+GYGxVDYckPXoc4MCCJE++cmpdrokAiN/nsmIPkBp68QQXoxnsjP4VeUkQgxrRkZ5VhZHgNtct7gkaz8HM70I231B+oQ7KCpB5VA4EVMyzGqdYK4m4yl5F0sKoUTLu8wcGwAS1ls0lap/QXe1RGzxTJEU5ywvOmDeSXFeTNDMipf84nWG+5yTAWqN5r/C3MxrnVYtJkH8uiA+eGvO8o+WrnrQy6KVZxAmDWl8bWnoIQb+g1zsDLHemNXO+ZWwS8Hz0TtmnljOkpSSH5gtAz/gqXvpJ92xH7z+M9VEQeF2ZEKzimBHlKL6keeF79h+vGvx/zURUdhmdre8I+wJ6Gp4UORs3sLxW+FDZgIYPlYjCEJVGT/tiN34XF41NMCG9fnjV//My5YMfSGD9P3ZzgRaJgmdkEB+M6GeuLDB7jhWEPXzj5jBporyhGHK/9TvmTfbVy0COn6RQtyaCLI/oUAq3eCp07asUOixsWxH8Py7mMv3AE6gK+has0ter3t3f0sFpelOWoBcuoQfhytBuuTNS/Yv1dHSV3y9GVSHBVtd0N2vJt7YqnaIylpmWO5cMvcLpdoaUo1WUuUM7nAThYnBpu8BC5aiF5rLwscwmSoKXovWBX55gyQ4gkemVwrbSJn12UEQkxgTmKJRHYx35VcsDRAoYUpYnpZKaR9Vowpf1ChnfWvOqOvrRqELyMtTe1VOKZ3I8Ez3mHy/Nf4M1emtlM5bYEwhGJlIXlWFc2Ik/q0eKk9JltB9liXBMwmP04taxP/hzAMSLCY1QKtvPQLLiZto5fbls2Fp3doYStiYJCu09KjtrdANJyfp8WeyGZJhVa51+IPRJ8/zVOkcxe49hJIL/QIvr/l9nwKDirM+cWPPXMNfV5XGukAvIPleB2mSpTk/4Zb58+1IYQEnaBcOS9VISF/ewOIbhW1LWNYTyEnX9I5zvUTX16h+IeAcxozcjxcjl5cnz6NX7osdZIk3d13ZBu93m1HyPMBl2ZNIz0zuxr/8/pYO9NzzEu1+vL1BXky6LQoyVploUktf5eMfEukCm6z2pIeg+bPplw1K7Cj48397O21SnE6ivjCK8zJ+UhpazSujxFZjo8Yloz9jQ9uMrTjOg6mpORtCetm3DlxPXohf8qIf5xN8kbQOlbTNlKAoKhVcuXoKr3uhu9wvGicu78POMGtkKQXy3RDeYstbtIEGGcQTaRAgks64Gp0NZykfAqkcvHrq8DLyDDEZ2h4rwnD+VR6C+KjrkEPgqOxGr4s63t1f96MymwimKH+i95xrNKhPMp5qBvXYjVOUSKFTAfzhPhdbkYLU/TWN2BjyitUa2pMbYstCiUdbM9KA5Ue/NKAvHLBOAixALpnD3Z+X7x0OgNVNbuGWbJh4me0FfFsgqD4h+dU8Lxyln7YjAqMMJbWcxd59j0E8jQL7H/fyQ/x5GPLT2srDpVH/xAHdLENcp3QI9Ae/Cpi9kFe8+sQJFrc3dFAQzRSt/2Z9/ZzTea9fEl4qJG06RMZJRElC1cLUWPBLi6Lqs0BYb8Ck/W23R/MfUHV8n+Ky7UYkrJGSDC97pPRUqeg3rCiw9DKYyZ6dykqJTjpK/gxTnu680hA7CsY4fKaGkqEGq0Vd7I2uHrV2lzbx53t8/SnuRRtG62nPmTcRAFrGhhXBONbdKSF8I81y67GWBZATw/Io+wl6IYaAPhTDJLJCTFMz0WIEJHGfvRzYNdyl5RjZ94AFDBE1SbzwYjeFVIx3lpCE33B8A9Fwr3y0QqICBetU9q/mhRCE7cAHkLUe7VkfhFagQK/YbWc9FeUIx/DumwC0QCnG4Qop3jXz8asleFZz5ajxoH9lpkqTn6ExQSEfyfYU6gdPaNFkvDkrid05kSSCiSLXJAvQhSWawXXg3DqhmyTw2BehEjOnZrAbtvCYwyBVfFtRaNZ4VyygXwAi6p14mBdP2xeX7j+kQxz0h7uAVLgSkar1KvH0F068Cf/4mvy0GuBg0sP8AUB9O64WYzuplzo20mvvrBCrudrIl5k59gRSO2Av/cJ6N5xGGn6a9WcuA/G77m4tkP14uKMrC0IaTB5HO0lQHje3VSbuIIs5Q8CZIQa8xVVJkxN30Rf9zOUTMvxY+FX+ki1pvj1NEm8QD6w78AgkKAFf3EQtkHR0p6Mbv4bQ0ZNoEs+pWnHkqwfNUpMoKgni7k0vcUvlp10veXxIYlQhd7/dK7utTSYq/1eNdJgYFd6EFIwzm2j+gmihDKGv4vTOFafRxwj/M2+hcXXgJQbYsEEdlxpTJHXtFbTLewKMA13WYjexh8jsaeGh0rkMe+usBS0zqRswS0dtHPT4SrPlCMmISAnmOAqdbhZf2RdRO4CJBQJvdQg0WchrtNYR42UxeA9hKZDUWmGu+yBezWXICQ3ZRfbjpP1t9n9lWBLeTvBBAWzxA+ii1TmHVEX4obH+tXuMJQHfOOkADaGZ6DOFq3Qhiw01lLOk+DmWh/49YNKMRr15u9zlHcUKsKcH5N5k/O4m5BSkyBQSC545lb6TB2COrJe631jVEHF95DoT8NkjrtRWO5GMw38mUIvn1cl1iPW3rDh1IdeDP9Y/FP3ijyFqx0cp+lW58gkONmTjVgXlby/G9t8iw+7awpVt4IfQXPLpJyR687G63ccOKAd4KX7fo+QipXj3lXMhXgoi9ZUsAUUN2B9tQAiKdQK9hF6Vou1rokzuWTwdLLQO2Xy1S3lMfCnZIUuaMeOV4317olrAl8YUcPE6xnSTC341sRIlCJqsiZkPLjQ8d6rFs0iAu2xmTIYYkU4XNrCeaAbY6ak4aEHxHWTGyO4OGtE9IunZK3CEcA73cG9JeWTRvoJa6Kq0typ3MGRGzOaPM2NWH0HaZGlgvneu7UoYmVqdQxT5BKDTXV6TJzLpGnPiWzF6JtyYMcUHip7LDCNCvRQMHOF3MtjhYWDXV23Orjn6YsNh3GPq+2CxOGeWfvsBo7Aab2oKbUjL3+LEBxETAUcbYluD/wAQ1ajmAw4sMlLxvmvqWV6VaXMFARNtBFVbPiaC59UJJ1Lxt1MJTnEw4Ul+dlFNnv5QmHvasXw9XZmeRSyC341+GBNi4O2dxg2Jv1TC0B+SKRr50fT/tV1ByAUf4HZPKvbxUihXZvWQyL1QEj6aomrHRhXWxgIHNPn+DNj9KKxKmpa4qa5PSnjYIsNUZZGvdZN88a7SNJisx6gmatGv+M4ddeSfgXRN4AXnFv7cp/I/QjF7Dw1ob3mO3LTZueUit9TjPhA71V+utdOUqZ8ptd9SLf5TdzwSiURc+k7hIya8q9EpTH+58Ll6TyPV+XWoNioqlHYojKWaW8zYp3gLAMuqojTroBRNMllLY8ucNTuX0zp33BBnIIvtwo142yHrFTWhrObUZDio4MN5o57Ly7BgCeMb+apIpnuTBBIitKoydLkD37AP9hXl4jAVsFqU3iw1JM9NnqgdFHXgwkBLrdWKK6t2JJXMPsWPDN96upMJVv4rHMbtCxmG6Xn7OF7Vt4gjyiyKliT66rQ4yeRNnRGnMijbGItlN5/xM+bXmSmazz+h6Ux9KPykLRQb17GaRipTJDBTJFQNUgG0JQgzpV8c93Fjby+7xCMwhFbSbsZxwMSBeVY6/lyo48h12CVg3Yi4/UTt+Q1rz7tv86t4pfhoBySsCRpNQ8qGhdls+v+PJauT6ptFFVgKc2pY/YShVrHW9teavgA8rPurRWv+hc9cK01CGvyRbYTHCHBZ6JKpz3ndT6Xgum0AxSHdc4WSIbkJwMLHQYaQTL+ZsjeuhkQBnITsoblaGY2ky4PgG6jVtPaKNMIZehUX82Jrxcs8g6+kNuyCRdb0OLPP/4eSl+WdffGIl9aUY6kkWI/AMRG2/qq6uSOrrFRIS2XKD/psJ0EDULMnIWh8iYWVh4o6pwvD0cImSwmUkb90s9FZIBLHzL6VsjAIYadTkdGE1rkfk6y4cL14T5sO6ljCh51cNbRFOHQdgz8aQNR1/CFiMJjgTptEt6ImVSX+QAzdY906U5Q2FbfQjwcPlGkSqThH+kgdcRCkmq+xeAcBS4DSbdWWmURYnPtc4x/z/raa9sp3EfyUoR/DaVOx9E5Hr6l5hEednjLxPGehPhxZdjnIObEV82Si4obx0mbBM5wJe0onfKUIwfRVes3/lf24KLi4pymiM7crO0Rb7j4ZuCOzMMhai0q8EKtWfZSYaiAVuHCD6Jkuh92RnbRxyK3jR4Z7omGicF1ezW5xg6Uat/CHobahgjvq2tmnmiUevxrhs23CcSYwjKuZYrSNa4ccvH30Ej+7pLnMI4Nb6reA5AjzzhBljXZlcxXeS7q5/mwZSxMFIu8+GdBop4VEGfHGQ4ctl3RS/6rM6MGJoy+WfzLuLwgBughmF+Uz0NYO+Q7yTMoMfjYvdgGxz8dpZuIeI5LGUa0wRogemRWGUKE69hQqVdvGCX8x5EEkuRcnkQJVMO9tJpRkkCwgoenxvU3SVoLkSVfw6rpVTOdE+ndVEW+ZRGc4FeBfTxP10/iD8x+JRF7Qc9KXW5J4AOKt0fsXir62/2bUpjglMc9Nj+KepjynsNxeI5NVDcEWjlpj2HPPH9UGuQ3wY/GHpSuzWldZnVpN5xb8Ov0Jf+RSlKInZKUjKn7JLfujFbfwtS/aT9ZhHLpXSgh+gTXw8xzXY3l4Gd3VcT9UM5Nf5QzUPgeId9+pGsQ+zIMsA3Iipr2c5OELeeuILqLeEoikwFvnCLw8Fd6f6638F92ZuAiXDx1I1Kk1i0Msequz++Ocd4rFHWZaH9d183ycrujslRhNAI4okfcSLjj5wD3Mf6B5t/2R9E3LvQk5LQqKDAHMDSw/tf7L9ysFV2/Ah+CoOc/Gj27dC00WJeWwpM0aS2Typb6HP/aqDanBrsW8KZqQpjzrbNeDtvS62ab+gU20DAndm/Xi0q8qHe54POR9EYYR0+3CashJp3MUN0YIWI+G9sGqmvc4mZF8ph34xt5Ib185K8ZVCu8DPhy/wDsETfMQxUDrvE+dyfoTbnMlIqlNGbJM4lwPAhIci0wCTnNpzMsJKRIXyeIE0Y3fTUviakikK3QoLkMxtVB/qZOcAisarrf3II5rbpFE3TCae0L7r5FwW16ZjY4eiMyIliN/dOT2iNELV93jRGj1NvyuKlehax2R6CdU9RedZoZdAH5dAySSn0eeT8/SGa8ayBamFMCV+QS09a8qO6AXezdCJ56oS2D1eiO1s5LQGna9u/19A5ZccrHx1t2mbEiDw2Q9VG3jSd3Z/YP4Ret+uJz9qnBPKJ/0IAauZH0hjBuaR/jfXY6xiG7gCC1/3UNwOp7Epv72MA4E1IAFESi6AqZDVOQoud6vNroAdEE3piQL0Fm5+TV6fE+MBfagHHOncW5PYYFgtpUtoNJd84GjlJZu2R1ZUHH79m/IRMXrHntXobe/oZhlJFY8Ymc5Z0hGpehr5s0VZPU6Hq4uzeHaXtemIHOMK2ktK6SuX4lwkCmG66P9rApLs2EIn6qygsotODNA8UuhEU3lW8MCmd6VAGXm4bKhngMncZTaE2B9yuJVhpYp2f0OiteSqmncyGxviGuMfrZ6Gp5uHojDc1N5xx8blfbYfdd2Fc+oSxJ9K8WvCSG391sdktTkxJDhZgPD6mvBEpbtXGxmG4yKmwAg9+fy1YKTNsHXZmkJ/Mbq3d0VGr3XGvLHjSNpO3AqbgA4MDUWk4A42d34Jb4ZpV1PHn2SKR8IDQwwKgTokVwdZbfSpjZyB4ie8Qri+sgl8yte0Ttfyi3LjvKybCar/RS8PbXbGlh6KEYLzyKsmXP6h4MIMmf+8dAYiUuZKcO0UXWUr5tjLhFaz73GSy/hCBjgA3xj0tbMssnIOny+1N5cXnI4TAq+h/wFbHR1IsaWrsQV/ln7RaxHy2wCewRLJI4vWhKKUawnctGeCfhxe7fVER/PPJzLdBXCgYjHJ/fGIv8I/U4J3nZxGof/AbkPQ7LkmhUfjB8tTPsHgBER89Vn71WA5xZmcSTCeH+RycmDkuccb5TBDX4BbL7qlypQ+72iD18pMFJRr+2JINkt0hfPUCnHloIrzWvoUYSlGZmZSIC+j+ua6xplPdVwFfNe3H03+rQa9eu9YP0suqraHFKkXP1etJPJRJ5R1B2f+7zQMahckjstWIRQEwDq3qMp6zbTqIJnvA2HEK9RQIhHHrzswY+Cqh80iOyDJ5fDChfatP9FnP7J0ewhN0qiY2g89aMWdf8cs/BnNq9UYJoxyJQYTrh8pgm3YSnQTm6t0IhtLPjZKMcZ4Qx1o+D2Qy5HgFzp6rjllnJtgW51nrHPEhGSRGZYXkxmynh7ht7Rc+lrA3Wahd5tjEtkCKWXw6K1iRFW5NBmZC4r7NysFPdksTHX5nj326vzA81WdPkvSKf4bf1UwktDsPI/6w7qYer1eHirgGi6AbvykcDFRRBedYf0jyqdPveC+LPXDe+mdg76MWCQgx6AFfKifDh+I0bfuxHKyF6Q19uE6SfJJ25MqKJE0OOrc3byKtM/6+tOzQaYfcVLDcjAQDbzAQkXxZQ1MzWxIrd5Ah5PSWZt6uH7XXQIyxDC/mP3xCEfNSn55+0guUkfgg+n9lRNmgOt/cviW7A8OZlAmPmfiL1RKXEhMgAofZvn2vbHUiaYyo5p5HJ4IafPchBTJaw0Wrk7SJBoTF9K46prJyroIKNZVNxSJx69/nW96mOUwl4kbt6LBehtVrYp8bO/LxMQrmEbr+HcaUR3abPebQSfhuo57aJeucJ1RrHpuX3lSfJ2c70Ntb/RWck8qLoqH1EuPBPV05p8LQaGNE2qLwTeaU/neU4HpbdVdiOOSQ+NHqikgcShH+fM70AGrLcSAzd3ErKZ+n4fdmtjd6efTHU1hJ+qZ/OpWudFtD39YMDegL76Q6Qhb+rPk3iQ5IwxcytRYpSEU5frDo/UCrOg1xrwNUnzjeQhNTshJ2ouS/jtstDuC6W7wxCJOgW/jGtCAIOvej8Ld8DwGW4LGtA9XvENGlb3rk3PE0sjetlDrVDlHv2814v/LH2D1Je2IEizvUshI9yGdcWrpB111bL2oYrhRKVSP3v6Iew9mDB1AXzH/r4jBQ75eTcfeKbxFioPAOTvtRiF82UrFXpXgYq8gNyqJSK9YyATtWmDddc4muUJ322f9kMRshIJuAGhg7yzZJhygRvTyGQ3D2bXtNmML1In5pwWDX1W8q85OgTOUFB4+8LvNGIfY3FttgAPrJVYYItox3dfBoDaH8EUpo8FAorS9veAmfWXqSzRYiwD5jSIiLGrOv8Go4IxDyH1PDZT0n0KxyXWh6JFLbGJuaAsRJcIiPTMNqqwRxGgoOb6MJhAIvVuxxkOEOj0hLXxJpgbMyk1ulglrpEqVSmqEPM3gxhlPkV01JR42oYxCDGrYDe00DtIDETRVOX/UADn8no6gUjU7rzRPUDYhKVMP2JKGMBgNAGx6XZ6QbIu+3HHocYFOo+5qhaVDM1caN7I4QMkjk9WhtPIUFa76zYaOqKHePidqER9wKCDN3/NZ3ev4mj8kFeZVVg1EA6FEwJj3zR5gtWy+BiLtL/pwurp48Ix04NnZZly9xXuD5DxWxxrDNQD513pTMfYtb40X3aRuqaWZnMsW/zpN3do42+P1K55BKIH1yFAYdfWSN2m5M+IyXHSaP0qBrSNAbDYwPiKMLCd2rRzHLUozbsyZVSKIX4K8X0pPUHCkAu2iPpG5MOdCeTxO7sAak4qH8l0IKE/cMgSBrY+3NllXKo3N8SpoQtMMTH4prTkCYxK69B9e8b5l3loh1CjhyA00bdnZmLcYgA9NuFFsc+QXOChKvieHvqD2wHJX9J1Mg/TNhG+jQ2eZKDeep87QfIArv4LpShNL52rNtQHE3r9qHuh8nTnjgRwCL6J6jznOcExCflrc/rPzHvTejDq2p8bL41LRfNoLYFrxNNyg2osBHcMjaigWwRfVigvgkr93hQNInxbPy6EggJ8UTRUpSiRXktfTghiFy8f4/5NkJR4SGm0i6wCBInbSJpoPRoekDiqA5dNSJeKv/00R/+u155Op3kglFik8ywgVfllTYtcHKQXgiswv50KNcqH6N1hjAC9/jG4J6HPq1Ezclsr/Nl87TLkFjLOrRiBO6HkEBBeVht+hjG+e5C8JRA6eSE+r/KJoCP2Pw4suPb81NLzV6f4KuhIKM1/77kEBCUlaeEzx5CU+bTfnQxBiXCE7fK1oanLn/2/y2VlqLRnrpRPxsdm2fIAv3QbYCYqXBn8KGdtMxlx2grbhYTtm+bAd3xIhyQ0ppbxqFoHUE3RLRdXE4ic12d7iOfm3/bcFtRWZTecx92xX2jEUUDuX8PFHh60ncXlmqjJQdQVu6DOakXlX5VbXsUfbWvYecQ5r6XQeo3m+pfuqpit351cK6qVyGUzRKJtFlKAQEWM6wLZc26ala0fw+C5hhUsHR5jIWShcF+ZjSL5XNH88mHLXOoZTMhGAgxR9SMdXgYvBCkVx90CFEO9MOxF+g8zclpZRSZIbZHVmSLUA6lbu8xfasIip/4H2G17gp0qH4t9yPMMmZkC2Wls1ohin4X0n5BWlaBb/D54r2+iDQHYajAvx+7eZteU107pW2P+vXfhCB7+2a2/g6gmHQrp853Zdi6tUY8FbfHUT/3jwhl07zemAOj271AFwhQt/tMg3AGwAX+6no1KnUNh5wt2l/StNsp0ad4GwO7jUhdYsa8ao0hvc+KG4/srfPY5V1yYmfqkdiIoR3agHuZtsjHKw9joQSs+V3dYGKELjQpG1nNgLgWA4e74it5Rg479LDF//+3Jql1+p7KxpG1kWO0eUogsq93AQqeBq/r3B133F3IBaWUp3b0E6kZOBuddVGQeBIUSztTfyNz5ajsm4jrlxrMeVXu8NoI65FBGNrzlm5hK7RPoln2T7oN3R4piO1+VNj2J0SObWa450uXJMY1QpYCjZtBgvouqnTeEM7oeLNJdWXXXGkm4eGp7v+4G0NS1S95CXmVwg/5xi0HtpuqVf0O2C9hnAL2Udgbc/PUI3tKBcNYE8rQ8rr+1KJ81EpbJEJklBVGIfqRofePMEZD500MsK4AGKHKQXB8GyncaHRU3ITXHC3FxBu8IH5MauGVOSNm9dWUkLzT09ibcAxLpddy/onoxL3W7R7Q2ZlQFYl4VyLsuhgf7xK1j3vuEmwcvgOxFY7xXQbU+J9FhRMIYiadC2oU3u/B+7EaRaTua8k1KH93qqy/F2WeCg3A7u9eoaYVuP9hx+kl/0O/lfhiuktnlJrZJbMqODUUus2zTghTBK9QttnzUJmeGOl8GmWY8OnHDHH9AeD9fzWZVSuzrj8gI6HYpC/+uDeyTpexF91sg/pTaFrbhhxgt2+B2+TUDeAV5ih0KJDZlI0wEvcsFuVD//0L5lXYcqqcerlvm6u/ku6IE6G75YbqYlBqWkzIOQO57DpImIbwIleU0I8WmTy2vIeg+cS0BifynAJa9uPBe8jWaclFVtkBLrDickHEHIIcnNfJQM9SkhhM4Y/rlI2JjqKB8SLbhSLb6ImwAJQFEGXjSyc36VXQBZ30F23OrqGhMqyzXwIvZEWLny105M+AhcdB3H9L3KPiAsjbbIBHu45jXB3dh3r01oNzP972v62TwJ26FgHvrwjo0j4v6vKo0GYGjyg4WDx8ZNWXOqz5at0xVbumdjCr7Gimfc/Y6bNL/sHQGt5pNJyNCiBSLKB+6xv9wrmeDBGqKuKKdqhSjOpV4yogmFYfWIC4b9rqCRHo7lbIIbiSACK1EnW60xcoa7m/SO0vSdSd4vpgjKs9Uch+Jvcc8gK8B8n2lismyy3/1wMj1mqoXVR9iIYUYvNS3w696CIw+iLU3BpPcP9R1oSADm45h1Febl1e6ZTCBM9JLkiJ9kuyMhdQ3jIixBE5H19VhpC1JjPeJ9KMIs6h7NO1hy1yqfVNi6ADt2JrA/SBtsA8WQcCXUmOiMEKEjNbOS4MPrim4Wyd66zYm/v9YgKmBOV9wKlfiCdMlM3Ub+CL/4DF5Ft29+4neJBZn8gau+TfQnHWbrO2DWHcmsUCc6FKHeSP9OswRmPED7gIjZtLx6WcAsaru0vACsYC96J5hYskk+LsUSwHhJlZgeUlPY76x4/tUDxncY9IIMvWk7K84pZ8sEpYi3qNaWIPsVRGEHaPUEoP7JsbS/BsDwBlo56sRZnWw7jypCaUS1xWL0NU/YJc5dtDtVJ96i5c880Uzno545kyQeF20mLtyAPovrrLY2Kofkqb2WSuIc8haVWsAXwz9pGyj6S2tj1xMq4MmrhCZJKOBoxf2JPqozyv9pssYUB4PjcDVSA+yw4ZGvrOtwSOc9eo3xXGnGKvleJPBLL/IYc3Mnz5DEFHWyEv6HyUP6s53D99mrVp7U+oYNiEUJFIoi2rC5kDNIcoRzUHNT3W/Uz3SdrXiaNGTpkUiK+LfGsJVqWBannHakq5md/sWTyhCEJPPssMMtDEt5JpMKVlcNsz4nmrUub/iL/tHB1ilQ5H8PfHai5QiYelHzxt/PSWzwN/OZCLX1G6knu2A3DxaSBzyHGhtq0Q+ciSKEuzUSJV1UGPOI6WUFCBvyH34vVJlFCpX66Ja2rU0a3cSMyD9xxCLVtmPLEGG5AO6C0xlF/lOWPjlX73Y5LC3zbnTh0jKbjypxZOa/QbBHQnfAW3gRTirsAS3N2rOJn26q7aDMa4mvYez1SYDUm5VcLChkZflMdZwJBLpz0atJtX+6AiH+X81qS0+ZL8zRzEJ4DzENjJWOsZM+Ofilvu/Ic15zsujBEKcjhJeFfnsgEQA7DGHx0TdwPCawNsBktXQsBthBOTf6Mk1jJiyk8omac7n992r/XbRvQasuAMAAj2kf2YduTOj3FD1ZOha0gAp9tH6k1RgexiA6nJjcTOc/uFgi7jjZoDsEFbovdW2T4timevxuZcY2TXsJRzV/iqzc8f7qWamiaG8euPEp+hnTTy/yi8GqJueFMpJqPeNQAaSVmBKo9oj3cP4qGLOTwwKmqzBl1QatptF1KSK81XHBoY7S1bZJPVQ2SLllj46tXN/zw3+n4iuIupJ808jRNXw8vsRzWcmx7/OkU4UPmzC/4kxsF0ZNL56Qt6Ct9YrmW9jiFvp+hGKqAfYF68s/re0zk74N099CzpIopqvtbHvShWp3bBA/EeW0aeAdCHHKczPi+mi+vbEJPamR/NPoqUQeuEAkKw8Hq5L2kskICzCZtThhQ2EN8tU2zkeqMiow9ZPxZp48AfmwuxxgHmF+eRKUk/tKe0DmXr8qbQWZD2uXdlSsz6cTKRyZEuFS9UgsoeIEMGfAHXNJbASqrtPKPOZXQIe40adtp2+JVYxVVixwYE4R5N1BkFr/bK/eQd89q7N4pIL6K2kPF+0lXZGFX+19nqliRHGrBstJU8xqT8U4vU6vb1SxyE+5ANRP8//OcIZzPuA3Vakq6AWO5DiMvhoK6Lt2j4d804VPn04i3U5cmFKA+SH6U4VAE4RrNhrpe0AunZYXLQRRpa8zaLQ/LCo6s24GawFVg1IlezSv7OIzYgspbeG1hLDFyuOENEJ71x65IsI1Sbd/3vHanulew7pJHSX625cKPrT3/Ow3uW7b+otyAjXIw5j27ccr3gCynZTrThOSKu3wOTstGULYqvVeyIMq8EFwInWnQyyF1kzh97Qioa/XHDOntzKjRMqYIladeeLZmDfzmBuxCCiBpbzOObHe8o8C3C7sDeSIQj2kUOgv9ygdTvEhF+y17hC3ViiHApxKnXdapM59hdvJSpjQIvMc8ZDnlJIwWOU7e3W2qyvzXBD5tv3wSxmyS0IpoBnydrFwkcOimCkv+4VnR/m/r7DIW/g4xX34EilQ8JKmBgS4GOIEIOS7W/tptGd5Ok5gLCe2bEdLXsaSMRsuWgrw3iiR1k1W9uai6JKLey1XuSGh9AcGcunObahnjJH+j6r4HMQ0hNTdMeXYcc7srBLS7oopnTplXmfM1insLezyv2WRSU8EMb18WdzJZvf7kNP2A4FFMYiz3/J0iESVIrF7ADoWtODPi/d0dut9RBkz36LGBHwSMEZIDMNbJswuq+SjPIViTNxs13u+3HOsmyjE8D+X5vfCYP57B/qDwBlw92/Ozw4Mux2O+PHs/CZGYtEneXsNeFi9/kw0fE/P14zh9CVdkQOOzYjRGpZK3T636+1vAnckf3jRD1gZ8drD0bykBVajjRmu3UEjDqKysOLSSSWNsSoaTw7JJ/fFD3GcqiJP7n7CsKxo3OWwD6XYRUgs8VPhvzs1HNU6eiKbh8zekJgynlXtqSlwEdXLl0tTvqg9ksnEOQWmFWqhwpENYOaTMyLFLyBrBnTyqx0XE3Pg8muTUcC/wAtCWWP16JLig51lakCeU62wQU1ymMGNuK4xETm6zgB4QUlIEXyx7oCxk0N3R+Y/cRQTN/fMZHpbdpBCdsVNTCuADf2SxwLNiDmLUiPN/BNRKGxG/F8L5mOolwT80DxNAoBtum6ZM42Vnu0tgedmmj3UB9T3JD8NTUrh8I5Y1su+HudxFrwGZJkk1HG1YkyTXB0ASamze0A+YCV/ZBbyiayrjp1076Y4RRU+o01tN5/oQztj3orzqaBdQMko5I17F0i+mXLszVWwCg67KtmhKAF9WOWRZelh61Xdxo3t3h06HODGMX8CK/QHWMfru7o8afJlD0hZW0/xn0Cn9omzEa+1TvOGZFwvRQMl43cqXqfsFh+ROQEYkvZI4pStQ3a2n32UrcfMwkRfSYz1dn1j8Hg7WSdX12SSaqI5OO7rBc6qrSqNUHBRpMC6v7WcDGZ4PV4p1OnUE8i3jzDo5BKT7O17e6i4QNPWOboNtCf1dIrAYGi1r1ZJgVtnl9Tezm8Giycn4cmnnjPERjRVue4LHkWdda5LqE39LBh2g1RasJLJ1nqOPA/82D68Wwijd/zHNp80pcdAv+Laa6HPzdmRRSG5eTg1pbgo5Qo+xF3qtd2z7VDSc+yKlZh4gYRykwYU+nCrKyoqRASZAwcBdlinYMoYCYZnkupzWq1E5cqLP1T0PsxycdP8TEhLA8nNhRR9mJuQScBtYQlNfbsPJZwGK255c+tez6QMhQg48Mp37YcKaHmusXKDtjwUf1UogHGjg/OdeXFHfVJo2g+QmScL+kzvaJGf6hoX2ZalcW+EyAEOzlNtzFZL5jPsRhMw/toHK1W83zKY8uiAU/LkolRJjwLpTeVoC98imUVoZE2cv8sPd676zQ+T7cXYZgS8xkrcoTYEuG+FTai8QNIVyFNv5TAf9kHXBVbrMykSjjtIiG+WewUFjC8eeg11jWh3QNySVeUzHhE1ybUANNYt3VzBtrXeqgAKrLN++1gFDoDgZtVT2QsOL3cxYiOAfCJjOQsexetiS0ZJ05CtdmFnWUM/J2gxaslvRIwPimpPkJiuZZJmNqOR8r02F4VoCvZoEH9SOF2SQ7nWkb8jG63BVMrsIY/hkpLwdRf3VNE0XOhG0YrIBzw7ESpyH9kOQrGq9jE2/LyL0TvsaN7XKw55MTiIfcnPTziLGHjFzsDUiUQB6XGJ2O8AxGhZJ+Eo4dGVFiy1Ww5yRMuMS/LT0fIObBs3PoOT8wUMpYQkCEnhme5wbAKrVBCt6Bo8NWDhcXCPcAmB3WKjLmJzQ53FnPV3E1NfWx5v2wPdrp5L/yNzhxwOxy9yD2dJOR7zJOHl9AyTcYgxq8jstQhJBnFZCstKKs0P/Ujz+s7rDuCTCrjWHZKk1JdZcGVj9oF+flVLrXAPzSlgcCQK2eX8AGvUBr/Oa/gm6hwxwdSyw+se7tTpEWYpsND5nrzf1lybBdYjijBG8BCgyOtutAvEiyHuizmHebRZm5KADZn0r7fygDDCEtKIQF7FlAVzlMa4TKG2KSetmjk9ihHVtioxCQz/9I+OCb1VtHiptonWMfFLKutwWUVSksVbvs9UvuFuKP1gspaJE21e4I/zLhHe3PSvqcB97FEp3MH+zGJShgNKJfAyJwVuMdYifDmYt8K7OTxXpUaI9bf2rmSWyk1mfCZNfxclL4+OGKpVAAnl9zX9uUYVdSfnS4oP/sN+Lscly0kYPaKs4AWz7HLav9p1MxP+pLTe36yq8kgczxmP+z30WK7P2/mjaD6cjiEaPSRYoKUewsSYcYZwZVHvxnP2Chpqgw3fFyqXTV53ag3q14AZ02r7CtE+RN2caQJY446c8Fn070svwZpVzA3bzNmc4wHD8HZtirRrY5o1J3O337hfP9fFtXNxq/p+1c41rgLYrzmGvDn/5zGZDRqWR1FHL7K2sfYgo+8mSkiSGX6wNqjCQzR+BdJZ+vIwPwuLtKDZ4H9tEZKhh4mO+7bW+kwrwBGMLyGCK1kzj/6yUGFYVtTZMvf+ojJE02ZFuKBJwtebWysroJM/3uS9x+g4qlCnytdXm30TgM9NuJKLTaazZhEvKkntH4tj2FDbdJ6NVJhH5kyvkBP2kJiupwqwmEjYwm+46krQCle5su90iGkFVGb/hWwWOIR1CR5DIvYKZA9uU6JNfinC8WFwCCh7Ws1wYnENdr6BGfGLuCT8018lUkMXl/QnSXGL4an72n+f1MZcP4PhhySyNeg7g5frW3ZO+Pb0BKqrSyQXJl1QTH6RBaxDST+FblF5EBObM3rIhQg3CJP4o3YiRcSgl/M51JutJYkglb1S95PJq7+U0LE985jyg2rs/lqLKRH3Gdje4r1/KBysu4rIVrb+VObh3mkCdNPzPI9WJmgcQ6CeGWy0y74LET9tqaq2dFQbE7xjst0LSXZ5rs4Yd/bVU3CZdlIA+bhwly+VwKkdbPnu9QbiInpq1r37qRCR+Bcl7TInb41iTPKg0T8VyLFmwrSweHRJ+t5jEGoSu83hBXCZcyTj/RQerpDq6QRZKWokqTcXS16CMKHWpliunh6rkPJAiym9kdAjGoFWQiLWVDsaA3A2NatQ64B3FufAO+FP/CTq0Ty5twEuBXuzD8q+qlMvL8aanMWvc9JOJ/EBBtN5KsCqp8IX4PjohNQBwLsm/zQ7d0B7kl+eFTqjN7sFRPve/w82tghGgRNFyz5Edc2N5LCM6hf47k4SlRo2Ly7W/UwSGq7U52XDQ9EMunx1CREkhfo6iQ5PrKlQyKXH12j9TxUzZrcO7qKPRbfZ6GrnCkMNTCoLeHzlxGX3k8G5QjbK90AEHroGehEdajlHZB5GM6E1n70kAlVPiJiE+c6TmcXoh7TnrBPVVRmVygEIl9TYZDxNugB+r5AhblB8/kHQxHbveSFUETPVxf3vpzifFbZJUcLuViAGyKb8nXnnTtlNw1Gj9czJowm5OMXiF2EvYXHA0F2CnBxNQzlTMabdSaA5LrS2vEPfa/Nym4Wl50kemLQqJN3E4dxRFx6qwWHEuoMSRle2HmwA9HoBKsu9/9llakNAyStCnaFvG6QCIb6t1udOgCvSxGfzdNMQJ81qdoCNQKpz27yzGQNQSPvlntjo8DqcRdp7rN3rg5sFek8Vk+KfCKIZXp9/4VMCbCAvvnJ7l3lDWzAzDEl5k7xZEly17n1FcYhA4t4uSzv1xmVdx83lkeVg2VffZIcKO6cLmmSMvjvdFr8nK8AhHqiLuO+KqO/yxN3XAQ6tlmb3VtbuqHbSUfDeposBtPzwq+5e3VtrTgOVW5fQ5UioRJKMe3K+ak+1S0fIQ8lNOj4U++WsfDBxJ5V560wKRr7KKLLKHE3zmNxeaZk1/kpTp2DxIKauIxFsCqjtZGBIx61ZHhqmhrbR6etkDQhOXEQVIFfEYStPkG2F47/OxYY9pL3qGV6VxPrax/1ZoByV7TqMBmPim7Ve1UI00GSyBCmeXMqeQjp3o8C3cS9ADCSnAnltHt/UGYbOhXbxonz5SfY0i+bChGuI8GEWn8mLaOnl3aziqYt/aOUz2aIIKNAi+5ERdldSaRzo6ckOQdAOhBN8nMd6YyKoUtfblobdvQfLhg+quxoJK20VfTkzrmRyTYhZ7dCDzo2ZUftn+RrasCFUVrT8Jw5SoWSd+CUD++z7w0oMwT9jM9vWRxUvx3R5VId+shJpznpukYyg9zM7K1xVGOy+yiQ9crrGAqTK9js0HOfj8b5H85KHLukIkNjWu4JyMA0SEuWj+zQ7cr0GhPcBubEfkF65+p4AaZ0d2jFoPDSLxYV33kAGZfxk/9fg+D8Hf9zIpDErKhqFJ0tbzXw6SBCLEayP0MrK73XgegI9Y04tPyV3uc6k8+ANIpc0W+4xOOfW0VOOJ6tzR/Xqdene/8JrYNJEDeHAhnL9vmf+b9AlJ3K/HSbfhpWaU/vSGQf//BJfePmOs2jVZVUtn17nqVDvC8PazV+4oyNK4pozMztPaLIaYdEZ0jIsIGLAIgrmagJspRkemKn7PVMZZ/c3Z5XTiycZ55XtdCVsAktQd6vxl6TVyjH1V+BOpfLCS4e0wAUPC85YGUBOiaTGSe3jL7HYDLRnc83lFfmEDP2kb797lEX5En/+/dj5BF2hCTOTxpbvAFrdkLwSTzg0Rk8SHFq7r/a+OMYdvMv2mYs4Cscw2Z4Z7EGh6mpHHJjgAGvUKnq4cSywGwir2aE6tLIWfKXDf+Yj51LkJ7/hv47I2ZpXvfVocZ93APXsciMiY0pKXj7wrJcPrO6SHLc8ZqtxepUoYz6OyYOPcQpPFW9zpdQmekOdRdmIqtnoabzDJXuQ1n6iPTlyaWaeRRV7plszdLGJPvbdsAYI3Z+NrAxrIvjvcFnBApOGpokmlvjeLd+9R+mym7WC3FtkCQA2zMgkumkS30zMvgaivtpKUGKysnDnnixB9dNCvElPKvAatHND1y16FX1ZJ/swskunDZEECgCN83zY/BkmIwqcjarf27aa1OGpgBzz7GnuOswdeZcy7Gk8cpjj/r1NL0pC/gYzCcXQCoaa9TxuLjyQCKO+JfjMb/LzzAAqSaGEBpu02RuO1b0Zc6pxHumx6nd9egJFi7LtwAxV6ZShbsPhbKz4AF2C+ep0T3ivpDNDIm/7LcoDxeaVS6MFFKtABEPczDG8tNVjwrrmnyD8T0+nQPmfjjVtIMvoNhKN7Kljmxcduz7bFrNw9/7+WGE/mnZMyoa6I+S8FSdzCRNo6VRCptX7j8m+TIkR/lfsHOG3tlm0KqXdpn4BW0FVyEllD3PLiVQUGHactk4PE5Q739CPYh6I8QUUawcjzZa3aOKGgX0U0FDkOGKT2CES85jWVFKWgpniTyHhuwhE300P8dUM9G1E7F5BaLIuR8MMLEGHOLY3wauNZ7Uy87P6CfSNJu3h3g2QS8dq1qUtCFVE1JUsmoDkIu9TtEXkcPu7NCGXAZs9UK88dWX/W7ReUnZZVsXGvtfUJNp6SJDQcADXzVgIENLcY/5cMrPgwuf8qi8a8wZPLoP/Zs2P5griKwhsQpJCYUZmi1jr6M49Z+ygvx4OC6KfhdUrBOkkyrZTKVCu/bYI1NAqDKFClJh/muauZR+SjkjkWQRaisg23Bx7PfX1RrcCpLUMH8Day0Mt6s+30stU12qWJJc+/kWvOeruye8CB9ID+7x+0nbTE6x8eZHB2K7darEyT7txrcYFQnr/flfQPTlKXuHAijDRtKvvQU8lK7enMaaGllzTXFBAhfFww9IxFhLcIyfdvUr4HeanUX5GqA4eCGXXoD2PP1OdUPiuJrz3zQDW6nRmcV3CGAo0pOiKFld23kIV4u3CQ7NOizUjUv39Od+2ne0FiKpHlJx5VTHuH8G1PQu3AxmNGLGYJcm0GPGlX8qgY8Ize5+h/MPt2U/WANJYxO/myT5k42wYkg5agRED8zxX7ARxmmQ/3I625aNK3/aFtBgtyXuUm5VvnUZLDMyPyv7vQdVW/5SB431+Eho3x/WFKdAiQYfmqvU7l/PbEqTBk33le8KbC9oqvrbV2VhM9WdotBPnUIycj/Nvosr+zvk3k3NCN1evyTfacXRzIxt1YVGxWDrWizWIU7/o/LvvfGy6k3dXk4M3h33eoXFR5GnKoEwzyLSUw0TTTD4CHTKAQKTe0ojMNvCcAF5FMnJgPY1DvcTSRaHhj6C6tnpBwscj4wXg1YC7+dUyCzkUur6Qm29uioR3mLvhj8WijRIbgLJjsYgLoYb8toX09WQTpXJKqtmfU78+xXs1c/DxEsn4KqqqMre6Kyf6Uxg/iz1lFEL95f7gT8gcXxfiCguIm6b4F/x7fMQleSpksaC6TCV/VG8ZW9AOmrQKHO6itq6sqQsdKTXRiRFfNPc4paXrLwIvdPFLdg+40YKxCzbyoO6bTV8VQQVoWpdLYnIQiN56JO0wBqP1+1g+cAaQn3K9pJLBCVpWV3Xj0mH3nXpjR5YOLBOgrGAQalWkVH2gJsZmxxxJqHEMihcqyECW4EB6J27tR8MsvAKntbEoZgbQxneJLS1f/jyBsI4W0JAFz6oYaRNlxrgGVFEM9USnC+5w4Tih/QeHZyMggy53Qqd87pYzfFYKMcZz1/ticLH6r3eueWKiFg+e1B8nDg3yeM+OPZhlZSUm5onz5i5t+v2gtN7QbNpe+mtH0m89pVeSiPcBGexS3NIUYHYlfnPJ9Z9v8UXn1GBv+dTK/DazcBLv8HqlekmawQkOGjZisXaUK1556i0g6kt4sSIy3yedB8pF8kJJp0TVyYqjwiJXMMcopn7EBfjI9yoMNco+PhmX+6BNqHJEj3S2CA5soWaYTbHE6K9ubS79uo2xZqVNBqn1ZXdK5L459Ylx+As5jwBtmcRbqNHWR7Bt6I5IJaXKXyn7h1u4K/6Mvt3FZIvubUm24ezLCXU4kP+E1Uz6P+HJaVh4NrX7rGt2+p9kKa+ldfFCSVDowBk1OWHkguQ9j1VeYPNXhpeVu7kXWArgMrMcfe8H/awYNWyTJ2tGEZ4wLf/YWsfcADWEBva3ctIzzlnLY8m/luCcsZoqbrZdgAdf4WPCzsDujtDSXRM90zzD1zzkycwa8Aly2TcDr6sFBXFusOHknjnqjV1EO0n7k2o8y+/JhO7qB8pdW+e4a3W4e9pDqkTEgkYAJfpDaX2r9x4hZuuLcfOaxZBOF2sjOthD8k6NdFL1koKFjePG4LtjrSRitMPNMN6sx7TgWm9dw3HS1h+w5ra593adxZLeBQQMxDArblBi4DFkiVHMOFzD4OAU44wIWewkegHscUk40j3SYgG4gaBSOGn/QRqhOwMq1w4KXde9VslavrLC27jXiGx70Oq5oi/KVs6O8HG5B0TlS9ccdn+IQdlt8bALRQfpuB3nrSlLcJjfHy+aQIQ4jeZIjsUdFGVbh73M5B2L/8kYpnSAla1jP+j7siLyIPX+/BfHXR0pfovw/qNO4WgevAD5loY3G8zpkUwNj878uMpNjlxun6oDUsdUYNMK5+BHyBJ5UqWSq/Aj9lPGZyOQhioLpvX3FvPhpI4HVsj7YzwHzzkQ/WTQq4L/ikb28DLVX2TYV9Fd+nsrjeW0XQ5H1pLzQQbOlkt/5qprkHYU/GCFN8Z+pS1eWR7ih4ZwrvZNypyx4xzf65C9LMKtkbUiWU/WQvdDGrzQiAcif3jT3x7j0nrTfC/ljN2sBNDxYnQxfhCoD4ySZFXhUNYy0n2PZu1ik2TAopzbSik5L98kVyldfZUbKyMhMxSms8WuRjsGop6iqESPOXoW4K4uW3suK36Nta0d3rkzoLy8X9bMYrjvYx55Q8yM+6foMyHo1RVRmtxrm0gmvLt7F/qKfF1kKMpHW0wcaktXoV2RNVfSvcAG9xNoC1/w8kRK+wJniCBP2+7/S1FwpaZVNbBx9jYooeHGN1P0VcBkl2pBM0p1aDKYbwBkkNjd9xsxvE0vJS4H+9eXjsOzoYN4TwYPEB0koyb4oAuFgrRNcuNZSURcf8Ui8oyYyW75tqr2KPIX/5QflUSUN+KqdlvZOgc+tjiDLb86inrtm+srZEktpIwqyHIGgQSDKCpvZ4P95C9vpOREY+9XEXReSYssBy5sDRuvRTSmuAQpQDwBwyz2Y/f2hiXvekmVCmmjQMc4h5MfMW0Ma+6/dKwalY6eGEmqzhBCchtAo23+DhoO0TKKpMpKeNqnkPLOC0dTJTzXtW8U9cmNAZBkD6P2FnA2qe2uh+r3TWl7eeT+DmopObet6licmVe/C2QAuigAAjsPQllT64m9mpFYHD9GoSlQmmZ7S+l4CDdCOzckZMvQKSwyWWaUE0AmKkqmQ6ZCajGSILeftW1/jQrA7CMzdbG4WTRbq021d1ALrLTq125qYWpU+aYokdw7XFJVEYbc4XT5gDb8lZTNuoLUXD7Hw5Tt31HE2pa/387afcq8SJRcEjW6ss/14PVOenDYB99rjCeU4rpmYm2PbhkCyCU0QLUhiC+ZdEkTkNvMiPrVcmpKPgIhaDxsz2aVCWCHxLmbqjh0S5QxiNzKIuj5z8xGcL+KDwihc3VoE6XOTipfwe121NtHTJBRL4xVnR3nHicLy6tJJU6aVCYVHDUYVYzbUyrm3XcLCWGbSqIRLm0V/BVvb+t2EwCI66vjxx2TdOlsDqFwHL//0UOFHJWQeIETUe0KVaN5yZ8dFLW/6kHfud73z5G26k4yNMjwttcVV1y4aFX5YOfsE9LdThin9Rhp0BXCeLe+N7jpk5EPvC/tr9LFqMh4BGz2XDj14guZ0ptvWyxdSlABH1dLEIZGH2u3c+s93LhzHAMQD6YnDjlHE1ORHchxHJG5qDUHUQGn4lFzLfK5M8tyiHEdl6rcR9YxRIKUX6ctokz+ReQe54FsqzAvSipbXYjXQuAC1dBMPgCKyVL8rNVdu9Lh64WAuYE1mDkh9J5bU/hVvW5ZAqMrmuGqRFA1kMbmJ14IHFqBAtrkcmS2yJr7DhaSs8ehtiQ/QB/hRa4HhPpbdDcfXDMtJnotymU1++yeLYkqOrxwC1p6YkpVcAxCxnpTVaHK25+urSbHoZOON4DX6GT+vBnQRgOpDc2LPJNjJdhCklWgSnRV4IU2FtndC4IGbksR10w4DCGvcZ2pSKEdZWfvTDPr184pBF2VaUZmb0zmSrZtujCIt9cwhAX4N7qhq6Xpm42/4SJ70Phxips5CRHhN9LA1MPahMwjoXweesFER1le7dKjdr9+jDDDipRxUF0Hm2yO3jvMgLK3Bgvlkxq2cngHGm8n12mxl0yOTpy83Mk/BV0gQAOi2YbO57f2LCdCsQWTofSf5lczquOEq0EwLI5zTCKcdG00qoR8euY1ApIY2k1fGlwkZzdsX3lNL5OZ+l2uDGzZVw4wM0RN2Oz/0y8gzMwEWRUVY520f/2O+9sdYU/X1qN3FyDJn5OvPjZLYlIdMCafBKh29GBv7YesEHMqzmfW6jlWUvMPMp6V0L2XdJ3TTUS5/GNYOz0DACNlUbtA5BAURW70z4ufCK1xMm3fY9tSIRtnIj0gKUeSJaTG6c0qk4hEVDwQwzmu/9AyZojdBs+fcpjOPuQrR9KC6FuozelQI7K+6DYahdwXuaK7qqtJLnl5fQnh2roU4vBjZC7jCVUL/eLauUJAJbi1MoMnpSauSl9JSJGFjbJhVtCJh3RqSgMfB+DcqhMADg70unlILKW0kkbsgHB+6ztqpq/r8vDjwXZ8T/bDEnYG/qZxmO/TJt21YGUmHoO+DaN1p66Y450v+Nb7uJGQibsHde6VjWk3plqLW0LJQ5jgqy7pTybidEt2AFrAggPjKy+x0VNtMZ/kuB8/W9KAftI+RdBKOi4caVAUAO8J/TnQ8vAlw286x79Wek6q6oBMuZnn50As3XsruCHfIfwvv0ZWoXlb6vFdshhl2SBZSv3ZM2qeDKOYYSZllysJjrWwpzPSbmbBYyp6peHibEE6eAZH1obqyiNvmH7YRUAcpKWt6+2PticmFk+0nZm582kO6W2rHifbUTVEAv4uhiZoGK2AKlREpMQOAK8fcHbf2+G59T2VRDoclbuD/1yRtiJs3qxbqrTUJhyJrRYlC1F525cZsXde7DGY6tujuM4Z+yc3SrRWOcG8Kv8mQpNNjBvD18OvOP6Sk53jUAz9qxgpJXrYVpDROZd7aNv9dQI2f6wInyD/2Nyx/X+lmb35vSNlNxlllpDj8ucDoevzmUfUD6lHQltvktg6HFMeEsNtSzBbuOPJEKmqnnkhp0FLtqPrDekos8wN7DzzwnjtdKt1XOxdmcqmv8Vbkc4Ue9l6jqZeM871kr/AK7Ch9nnagY3iwpCRiwTDSiQpGyPdTxn1znEB5O5yZhawtPh2Wu/0cq7wYr1LhzYJHyu6YszZGfzpn5PdTGA6DreE3uhYPM5+BEsAMiNdQge42O3Abs3d6zkpPzO69S3HlRE72lHzi3FkoMsImwii2kkm7rxQGmvf0kJ1D/zmTk/gIqxPgIWoUP5UNeLFE1bwdxNfE77+Xi/I+z5+GSsBLXMXUaljLQ3DYr7BjEG0N3D1CY+9fvmLs1r/XNgfpmaxJleyoJ0EiXvjsJQj4Y0mnQtaR/N/tKux3yk4FSIdgGbynrXE35X+vyhgQMbLgtD6DATP8A2wjipQhZ5aad0J2iNcNMiIKEa3QbwNzdRZZfKHpfv9n9TwZuZXOFmlmV5wTVZ4Pkz4V5m4oETEVK20X0UT+ylhTRnGwvfhBHMx9lH7mcglsR6XxfputvMtb/MhU0Cfkkyrl2P0QC8H5YSvVn0g7ExykbdzoOu77vu0B7hkxcrHcBDLazCfZ8iKRVHnOLXVWRZXFTuuRqK6KUNIWYvbX3GFIiea8cNSwOkrcxwg4kx2s6sZ7e08Mmv1tTa6r2O92uwEpomaa44+6eKO8L8z9ykFvEsaOP32llPNYVgW7nxRCqj2xbshemXKHiGD9sr+uZiIjBAIPoJBMpv9TjI6v6L8wsvsiyY8g29Z624sUGdkDHw6u/qLgOB+UylAePDv2ujm12Gctfc30bVzhKhpFXdY2kvZ2Z/do2R5eL9ujODwsWnWyCpl3eA8e5zX4KdiQR+NBUzJ+vVRhaJFBzQR2hAvcwDXcCM7TO7EcEMXm6sjrfuBMD/bqxLmGLtzwvUTyKxZLYWAS3lz7wyXQj7RB977RMz/SQV+D616tIUvlQfvGNM4BJLQWmQCnGXiv4bBsTTH66tXv3EtkZRqG1spvUbc8N4xPfpj7tkACYDk4oTdC3xtWWg1qbCG5XRTajA2Myavy3gm1n0fIA77R5M3KAHThqYujH5q40YDxlKG5XWbfYXq7r67tH/xcwIVz5Ulaje+SH0zQQFchG16u4mdonGn1NMkDKH7DLR9l3Wx3nW0mO+eFCCfpanYPBhDJmnqB/nMDC7QcBrDsWfdMuNcSaffD5OcdYx5XwvyTV6w4YM8g03BYkHJ7cKFs6jr8VFTDUSOTjFXnuFEpPrQ/k9xitfvJTWO8Y4uy6RBH1VfErOsjDjnBjevrfAeHNSBSlDsOtva8c27gp6LmxblrerywAL1fULwvmebHW117bt+e1Zc4B4nIga9sQiViIT5WAWSsk4b4rrMfaGArHwifnIPMPgQrgP42NpnqWhnegV8pjnbZ4kqibJzIrvZgNvttOaKm0J/4yYKIEedhJUq63bOomJw9xLBW/97DKL4Gx/gHwly9tVqy2fE19Gc0hWTxp0n0BLgniVH/STWuUy0x6LKZbB8FGDvyjsOy1kTh9vDXmKwNwrMjoihT+h/ZPf3Ab5V5Z3ubJsUUHuf1NtWvQFf2hG3/FeqQ0PGNQud59d33znd7n+3lsQqsVStfXvrvKP/H1QE4CF07omazdearRrOkQus9B7/wxuohUEcdHUdHzgbNNK60xIfS1wWX227VxNjTHolesqVejpwbCjN7uEcBY1M11mr2M9zf3OMBt5FBPhUcbhUJyCLcYY+ZusP7M0T4E42/bImxrbVrJJVRQVU53+oRwE1bZi1QhoM8bMXK2PwK8tE+s6VxzGIhtieHcWA94gkZx4Cst8KvZggqWxuce5NjKjYL+aqiJpJSA9vFRZJodzUA2YfFXGoOqi2Q+nV2U5eUzLKFsbtTP4rTV025LQU33gF9Y6B5Q7aHVLjGKbzNUy6s64VYahUZSg8lCPqiD9I3BPRCjKSu5qcynpSsm8CYKuZ5N+EqUftjx5eGA0FcwMZvzY0xwuMVWEbnjVaed/2gVlMTXhCWe5kBujb6sn5LeeiekKFJqPKd0K+eLxjJ10aScsMJ3aYaFym8fP8cscMrA6y6/Rlr8Jy2MAm4N+Vxr9vxGQy+A2Zc4tE7yM0gD2IyzG3Pb/QnJSf6986wN53JwxCHy1ese/jik84MqYwWvCdAv/ObUJps+535/jEo/xGFYpsQdRMDBuYrTX7BrCSfC3sRHaestx4Kol5zc/cQyFcSfaSFHW9EPle4Q6Pg0LQ9dVmJpS4pg+vuu2Yfn3/E/S5fDNGdfTWkL9uYbhcEXV90ENzFqudcVY/8pYRIlw0mVD2Z8LLOC+AO8rTSWfC5elaWi1msrO3a8v2L8hcriZMV2Ipof4VZnuZKYMNt5SNJdODcnLxzwHib/GJ7XpTJvwlVgKAxAPiV7P63Qf5gQHPR6Qw/4YHq+Ra4mdb9hiW9Ucx/t8rkXlSJOtVlkR+SKYGfhXCFCKOo3ucIbFEtRunG1nEbAnBHgtav8wKTjvsImJfoXDLE/U0jdKnxBN6ZTVeHK+eZ6DHcO5xX8nT6kEZYdmi3/Nj5ITdGvRPdZKSh7DJiE3HU8dO2v1RpeY/mxX61DHRMhKrYLTWURKoEuo511zUd5B0bQUjyz63gmOCO56ishwwlxfrGf0+1bxx6tBbEY021Kc3iGUX41kiRSPwh/9h7EYoYgxuIDzo6aKwbuTtII7QVnT0YaQXmksOa6XmBBGWKvR72TAgA+p8X5YIHTwSWqqy+q9ZVKw/DkuyiVTQUa5GXg8kXqSbeLFlVfs8qzPZ0gt9izhpLNZNDCVORjBnigpeyLHxBe7tDeULAK8gpsCuF1CQjnJn07g+c128TlwhPVU2d1QDtH6KTPkc66tZVeRjSNPUhPFyTtubWDEpRqVG/+dFLJmyal8Gf2Ycns1g6nx38HMx4bbB8pAuYXJ5JI3dgd0pMdhavSETu0x82f5w0V21FrW1Va+RGA99KgfTu+aNYXLh/ORYuBnNzXHkk9ux6BLYo7BMBOMnRrDGc7y4X8N1mpsyxUJ62DwtzyXF/gAK1laulADh+F8XRsGkYYibX9+6Yll3869Y/lspS0AKmEy4oj2VIowT788oT3spWckj7XmIG+UqJRjCtOqpcqA546QyNgxo/BwO8b6LZyOoe3bn6JeVYkW1hNrm3upvMm8JOyaaUrtbiz10sGNcNxyK0xUd4U3AumE4hBon+fSJ3SE=
`pragma protect end_data_block
`pragma protect digest_block
15649ddbaa08db67c4031f6a5c73c05e9083fdfcc81996620c275ee3ffba6267
`pragma protect end_digest_block
`pragma protect end_protected
