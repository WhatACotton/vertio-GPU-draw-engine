`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
1AjH/5CFBUim9EErY57CcSg85tYymyw5mbyaRDJtxnjs4pxV1tF68tsxd7ANWCui8TjssYRxByGuJGWSuMg+3mJgv299K9o6s4DuYCeYfr7tvhxerlrdwaUWVeYdD//6EtLgescYnApb7sAbgCGCS6ylEpvgDqEj32JOgX0Jxguh+B6ejM5dUBZ+ScVFeK/twpGIwbbdD0Ic2PJsQNJM9H9eBsHintGVtbpdYDejcVsNmT3s4fz2Xw26zSeVCj+17Uz7/+gFRkPisclA5d20jC98FT3eG3u2Ysi6zpEPTv4zCKQbzf7hybUy3Xsu2nb0X3QBLSL/GNumZCnZTUTnYlYbJh94udzTzZmajkzRKuUdpsfxmi1L1YwkIrKzU7Zr9vj8b0Zdcd06EW2Kyw/RDKPEnml9RUilJgdQCkwzHFmA0QCS+BRk/5uXQP32ZLWzYIrgGuLM1+aEYBNhhnYYD1Epvk2DAcB1K3q8tGJPE7s41vbLGgivDsugjW00kcpAn+pYi/A64x2MXKoFA6W7DwWTNRrIblgJTmcCyTydFkMjL0twJkuKE2wgrodzufK55V0aGK3MjqBybW+tfMn70Y/WmkUpXnC8hacEwFpS1kGp4Ym/AwVm+T/qochffQ0sXyGupNiSE4VVn4cadcQ4zGrPRMHojnQGKNcklwptzXMkCUbCeInZA8VJUQRyAbsv1kaYS3trOs49mCh7ic/POqvtgTfP/+3fKFKjjzeQT6/hqiwp7GSTgWg15UKbhZ9C/lBjWW2NNP8Dik1XaaZYvgxo5lj0zx7YPk6oG9viGR8whgxfV2FJ+gQRbSV0CsxEDUnI6YKP3IL6/gwNsP/gvXQSL+WOhapJ9S3GlegHnoWHeTlc2Re47dleZyBhwRWoUBfqEupySd21JAM/9ug6d27d1jhU5RhP41gkZXM9FOUbXkCgcHt6Rjl6yId5WP6GymGekT0+/hjLcv4q+sWK7973fG/1AHWSH+k2p74KD/5qpoIhITDl6Cqvb1sbSG4CemXdlu/Lj5XdkaPnrbdcC0Dl5gejorFlV8zKG4rnIJdDEwh65egBgYIwHMwbV4VhSmBtI6pbigsusR4ImQL3QxIrwCCcTK1n8t4JwxLTS0K9RLRLxaTalKywO9IzfR8haVmMUNPph9UZC5u6mql3uuC4bcO/ZzK9+gZ4DsVw1aKjCmCthe4IH/Q/LAIdciJyqGdcjxXfRxqN1Q8EiJ4/F9tCDY4Zl/mpWlqmmsLQBIc+g2vsbHxARIM97WXqlgZgWYcYhtg/MdubNkRH9Ku3mt9jLkTFuk0gF1eH6uZkL+18k7z8U/5/62hwmTN1pYHxNKGVOGNCSqBk+jcKF0LVcQnlM1IiNBH+GKrUCNmGi53elSVcqlPObngLnBPxSy5HAcSD30hCZcMPAZOdV6wDizdwtSTz0wKFe4fweqzd6Tbt3jV7BAp0NCYP3Jo5PNHC1laos4XRbEOrXzZ6vvEqmPMUuyQvOy6It6ltgg3ppV78BHEYcwxnMxtI47R+cTBUtC2RUie79nBeYVWIZ15WDPv63F9Tg49xkjLY4nNLwlEyO3H6xc00eMR4ahGb6JHH+HiFp1EK9bishskXAQwTPLC7PuYODeN9t8NZx0BWHAcOmh9susdU/x9FYskcone/OmOPBr5I9FwQAlB18DkKyCbwc3KpEmvfPRhMwSH4AsYfyU+ZMGNhep1gffJ2oIaYORTNJ2F4iatOuj/f3eI2PzfGerD4e/7FCTlxW51vz+N5kF8btKt4Sm6MrLqu5PtMX7Pyb9tuhwwsngmUe3S9DNiHHL71h6xa0Und/Mf7JMn6YfAYqRv7GTOLkxFldn1pQqoY35bYEOW4uwuvLmfu3ZFxbUTyjxtALJXNm9ZNpwwDsiWhQbGSCrhB4KWEFemrxcUW3wGZk0WITZGdzLYVKFR+j57GEoa4t/nW29h2R9Aq/m6E7PuuOB0Zqn8zHsGoLw5pO0gLq+qdZ8YU8+g9ymvRg5xIvg5idQvXKV8MxrqD21pS2Ovoa4kgaWDcHNQP/6/wuMZxco6lGzaf5I+LvgVa1c+6fxLS7MyjqwWspHXhT+A4N4uZyMnahxAjW6p7+FR3NMLPjTw+Uszel7dB1MSVbPGwA5LPek/Lh81BCa5t3iMJhDvezuZ31e/hbVUkyqn1l3Tjf3AOe7QiFRi2+vi4DwJ20EdI+RuxuW5EdsB7AR7UrqI+cihYTq16xSbNmTRYnWp4/odSpVEmP707ZJwciXk04iwrznbeGe1fEk3TizKKXH4OTAaFwN/LnfoRJczJ5MsdC4Aa7hkeGgH8falDkSS1zW3Nt/Y3XK+PEVjtv5fQVLArN+boTBywjlVG35m6w+agDBrsu1Hz/AsxRKCBAU5kUjUrsAlstSprtdxXSvE9ZmFNGrslP0XCsarzppqNu7iw0X8O81Wy71nxfD6rvCmFCL80y/YYM70xivPlxYcsdEmRFqlk4JtBAN+3Lv/n+9Ux+sVAdkeX5kbkHI+Tu7uyly7f5j4lj3o491IMT5GXlylci6hFRqdm2ai+c+MVTftAIEIwIaMkLyWD/jSzi64Uf+eU1vEKkte8C3qsuWIFIw+fLwknJrx8mPKw/LxOhRSSs3kogxJaI5N9cWfmfaAT8MDrillwLvHPxhdafWM0WQlmcatKaqnGMFfbZ8Sx0AQrR3bXkmgdkVLwtYp4jqrVVSdHFgx5gCc3ljWFHAF1lQLKG2fIe2eAgnAQQjmUeqDIOOBWAA6bUag5JphO0oVoxKy3g7UJ6m7gmJDTyYZF/mXWRMJ8YKajrhsYu79vUFTkj6ZGexO1V4HGqYy/Ibqvprc+uB9ejaacQsryUBEVPAVXeFUKFr42vFU68XETT+R6z/QBWI+1Q0KzNRmB2vj3fP5GUgdxEtKeas9KSeKpGoQEnSAgPZtXmo3uck+VCVCNBWZJIdKWUFYldRA2bTahFkJFTFWlFVdvePxBhgBZdDi8BO41r2Ql0pggAXnyJB1xFD2HpDcbJAhl8TJt8S59RYQ5WWB8iD8fQFi3mTpTolwlxve+DP7N0DGQfj5kKcpcUSvOuB4HR7uqkceBq1PddnLmTpCOsJjGeg4Btvlm9IENzdt8asvwJBa45VsejX3svMX5JDIFcsRoJii7UMJXmmgH/MuT1owMUH1wQGP6KJqWJNf3ABD0Zf88a+czbmvKbXCNG0bJxPcMCUHgso1+6ULr4ypz7YEdXHHQ2aRuxTVkLqE6FHveML6YbhDVGSjfJNSJ1JxghvNWZGo/f1wO/XIKrxef3pp64hx/n7f9HXj0/Z2HYgujG0FvtPKUasScrExMIic9JHGaV3xgysQN4guJxkIiDitf/wOFsFcgIcnXovk/eyWs2nWTEdkopBMDIEtWV94tmNqu0YFkPAcPXD/7g9ICt+UHKTEqX5dQBnToWWQrk0C0BhIlb1TveNacb+IJv+VaOnSIe0wHCd25m5EkZt62jy10fiiDzHqZmP2i0swYXhDLjzKg2c2XrjPPueesZD4QC2yQ+znS+J3O69/p3o4PUueNdmo8N2SSrrWOY5XoQVmO4IIPRS+IgfZeskNc+BTgaW+jYiI99012gm0Ow1n6oBoihP0y6OXHk3qRsSmU1SW1LiZ+xM4zhOmJOYmhgvJDRknBIv7E4HhhEd+QtUF53a5wtfD6sG2c83RYtJJBaxQLNLG60K7AzBasnWz9Bx+eMOLqsZ7qEJ70d4mGHKe2EoNU9iESi9aJ4H9bkIUXq3eIYdaDnHYwQnPQ3XThFLnCsB/8drU8E1nLFCQ6YUthJ+/mbaeIPelQpySScFv6c9ZO4VrehsSiCE3XDu/x3ZpPyTBjwSRoNigcxgH1gM/o/2AeT1rClJGWJKKUpL7bVbZEMdUBpIEBd3AiKGMF5J4zYM1oAgiqhBX+9ioHnh1ZSJOlWEyZTdQXjQlbAtMwpS+riCdXXK3M1mAmETzvRU8Yjs48WhvZy1Mi7lNzyFnTGzcKCUC+sbdmbKk4X0okwzf/757EszRTPIu35JC3bYtxJntYnVT9Xn5acsLxfS/pqqcSZXhN0Xw/BN1dpi4hv1L+veFBXpzD422JPDbAgDtqIsbp0KQauJB4R4RqhIk+tv+UP10/ofDbz4yGkwCgUZAxl0FbNGivdjmlkDhYl7uOxYDBxM/bTqqyqhGv7ptg837OGXtM4d/vXOcYRLebQECru1ZG7BDJd9XySfoDJhW+U/jZmzjoFmVGfFvZ5t0qVYl1Vz8pDicRuruAzksN9lyNKoVIBe1GleBsF0QcfKtwqgZGPFSpriV0C2flmbnHjFD4dyydiVYoQQMAI29q1XqgL+nThlVv7BR+vxrjnYV9TGg/BEoKaV2Qk4fCznSL3J4faFcTkVC+oMdwD8bcIS5fp2fVGuyUJH3HL6iDbVQdGe8oJMPKyc30NtJOR3aH4REa5yNANiLwsu0HYCr8Gs4AFhTf88qcReFbHSblXXRjEfkej9f+p1Jw/GbBokPGqDyqlxeAqzsMgYiODGvl2NHl7Tb267ylGYrGAvWJPkjMhOmlz00QmBhBm1wqV7ttccHQN1N/kSOytzVs5Cnve3BUMYQXiA6b9nW2JeX74O9KMXKtkn3oM/z67BZalqVfu4+zyH5q5/l+tkoIDwSq7cd9kevNc2ZrjK2Gc7SnolTg2DKX0cXmRvD/n9YfWql0NAKY23EfVIPL2gmzIRAyhUeIxAU3lB+gIktbilTFC7NnB3VLiWBQRd3cX0sE5Nge8j0mFHG3gZ+n1t4I+AbvGYI3W3GGsO99id6W1yBVli8WCmHFdQM48wShGxKMT7ioawsR+EE+URY7U7yyHXkmq/llg1KF1OWivNNdjSY3hZMrVYjH4ALFnS1958r6nixP2v2PCTB1Zsb3Q5JGjYs1UzzkE+edG9xNMTEa2VBmQedJJAh7fJFLJCaD2dijLUMj/UZfVoEkMVX4nS9kcFpKmnzK9XcoAe8AgUlQYy/4mUY47R3bJ+/j3yvPhqoMGU3MJk6iyddmLsaiNL/M/GZ3zTtpvCMRoviVvfOfoJFqHhYRKR1+ZU2p46pIG0mBAda6VbLIkc8KM7/bL5k3xtv3fqeUf0lGU9s8eUvgEQjoeoZiS9/LXn1KY+3390eW8sSfYjk5ou4830oFqp51YNPhtanHRVYvDz1b/onVyPP86uR66EHPILmvyCXa1SL7ywGJRWdlsgpD8F+LosFcMEo/mkcqYKgFWkHZXpLMNf8px8NzMJbkbOWl7LxzMkiwnUsy4GOxESr+Nr/AldozxwkG9dl4TBw6OB08IR7HT/r2aPFgFEAm4qQQ/hsErKO66RFEQkxdxLdAbvp1eIjPR4IS7CXsh+vsTHlPxKymHRbKwJIOp+VfrrtVm36oLhlorT0j3ei6FKMMKqejFel9VgOSSRMFRVGnAEM7vSoVKF9rGGpNykbB6wIiDmbI2AiRPOq1J0pfRHgm2uVWkKU61NJGycLaHvZsre+GTF+ZFlGzUZMAocgin66qq05R5kAOSvl6hoHBAfCteJj5DLJEUqP+2LntZNVpNdHaZ69Hk8e1jaf6HoN4Gh/9EbBshDNR6YUmAeeD3sj7lPTFyQjlOT/I2bOeBJANS9RHSnciuAC4hYhVTsx91fF2uiCQ+megV4RFnVeO9tJ3T5gbCRyyysYswWdHYNC+2EIIL2GMgzp7cVLOWP9ur6HlMLfp3fBJ3pPeEhXx2f2ReZYXDQRAYbH7mEGyy7q88ZiWUc0b9hq1T423pFFyiQKkksTeVRlDZNBjVkyJYzhZbEglRPmg2XUd3bJNENtuUpiY2TMQsCQQ1Wc3N+FaIgpUGltjxCWzNNEAChCMGA10DL3CB0yt0V4uCJVcNQKGoRfcQuJ4dhic3O+sIPbdqgKJGzlFCwyW18u2ZWusyYiWHrZEAkfN4U5xd/CpkRQKhni6UrkJ0jrsgxkE0DMausGq1JG9HUeY1qV1qDnxkqtlSqoXuanEq6ivTr4gAtUDJN41PtSXFRzbDSQ6ILEg9KUZLg7pfWYoRJkreJSziZUX+DiSNA7ukIHHhFXelTaedC7O21QgaeXARSRQh1vU+7SM3x/V91AzrQkCv4qUjO9JsRanYZ5UjNCJtdp42xFsNyPWfF9xyNPYzec60xfR8T8wJKzWUGq1Dn7r6S8regUrdcKDVf0gPNlWLMonoa51nR7MfAyqCvaS8/fuUnCaKxEWu9MYSnVPPeVCbOvbROjM1Jwr1eYjCVbcfuKsLl9dyMMTVrer4FD5AbN8mWVQxN04mM5UM2XwqaNErHLVzv74rFYZK71NsNy5kN+EdcWowDztD/aC+Czzzn/TDekmfpv3nMcBbpAH9s+tDjN+zlhaS6ZO37dp8+rXLZebpeds9/aicT9k3QMRuTn1bFpcH0lArNRRE+hSnyxwd5y9VO0xOsBkQqxg7WBjPYY55WFCQjrmlTVz2wNU8h2eWZk/abOWrt3dmMV6FFL1Igzbk4usGYobBetzYPyJIruncl0JinrdjM4Mj51A4pNcS4H1F0xA+lVP48lfk2HSIiItUvLPDSAknlH8Trl6IOGXwmrKMdj3PsanREDu1AtBNxUW0axT/aYHKjvOkMQjHjj2143HbBED3sEN48atjvYAXoUOQll0wCPwYIAYlMJPVR0LA1WBFNnYWKLRUSflKjYWiGKtubyYPCxpP79eGAgdlVidVKe7y6arBpxx9f0bT9q3RSc/frB/pCXpKAxFHGsIBSlnzzqQO7dFKOmCiSxDttqGaX4Uz5lSbzKWwCDM5D96pT/3D9+WM8hMIl8BVxyj9MhdeurDb6hpMoMSS0PyHG9wa1lpu6r7Dh5MbagqozNVmE519BFHCm/zYabVhFoAoYknHO73X3NXhDid4fpp+6pDsFKKHCn1fNFPdCzIupb/7nZULB10k5hhzUkLyaM/FHk0HajIffN+Pa9AHrrxEweFs7g1iJINeJr5mNRjpdZsbokxrosAAD/AwBJI5aZPfdoyd5EOheF+AgmEKpLc2azO7ESwDRnTmuctME/m96ERY9o4J2QeZPvqDsormP8NZ6twmGGHjSZRFPg9DEPB+/g/AlKA4+Wq0RiDSjPCMkYt0ncUgY0kWOTDhl/GK9rBGiIo2836d/DzkvXAg4N0DVrTSI6j9IsjVIb9JJ+e4MM12eG8EOQ9MGJrA3QEmCrCzRCKxb/1OdxguRASGcGHgjDudWmlwgWu581H8XJAJ5AeDQjtLx+WkIpm6Fdc9E5Xrjo+8nXmdAMqx3UBAsnuV6fXfqAAdL2BiDOLACURCFFyegwG1eYTZ4YZbQ/vN+BTyI/IFjkRVC2Hrz5jpU8b4zx+Y0NmOyK5GwgvvFXtY1JRk6arxPI3I/nuTKlvHd1MDQvv0PW7P20EcCZT/2Hh17ZyoRkEsg/Mg2SmywRhfMYkAgkSwnK89fjjuf5GeAECAdc8MWBL85G4M11lbQ+C4Hy+br1ZaGmxJeOssdFFHUxnY804jp/2vQQZ6E3xeSBu1dOes4I0Y1UzU/eVDkbuw6UbDOzsjJTTRvXduze26XKbKXFiP2XD3wB5GI7RUAxs/rynM7F2+bNf19J1BNubMmEtpCGiJqzVpRDUJvuPtwKgbyLo8wuccundecdoHSSkGIUOV17x1Hd5IUW/4bvPsIQ3pEoUQhI7UzdEoDds/+ml1Z3Fw5+aH1GR0ceTatumbfiObQBtX3sHSc0rTfEndvaYmehrfnEupuUBTT+we/rQFYf7TTzNWpUgsXfbE+vdqBtmuL7Q00ClAODmpKRIBchhGvpaHSQchKWRViO+KCb5GNoKfT0Fp6rXmu2GgmM/kAuA9h2lVqpqzXKV6HSlwEkkr8iaf+UfmCr2G3hLL7wFqb+dyoUA0W9Z80BEmfuWcVAASlst6axa61xO1jGJ6UCIedWWDPEay+sbBm63Exla4y5ohH5Ir2bVixDqhE23jdIUGH8QG1P5tdEsoSml8IujhfvsI1b/QH3FIp1f0jMR13O/zcMGb1gPOCVOz6JSyu1auTlm1xcLVJYXamuwsWfjac71dRw57FMH2pMw0JTY/tehUnITg7eiW9AFnpCO2lAv/t/rSSSLHsXd/EAu+7bwmaHRmI9vcbsvmikmuxYzprT4zLPX/ZLIpoVWOI0g/a0AJOSIi9CoztehI5r9gyFrKzo9pfk2pCtgWhHw9G/zENiEO+/NHUpEgF18n8gmzjAOB/1z03sOSF6MijeGXcAD5V25Z9eDwEtRHmZT7Az+0nau7sKcHJb6JHfvsdhkY9WqvrMvLat4f2HBVjoi0M+Fl+YT8Gwx4q2OaABbEim7p7KPZKKLvQilpCBJPisSxzgAdettXQAk40aE7U4R9xKNGlfZIai8g47Jei2n1IAomlxguLp/QboyiN7G3pWs94HWO3dEey4WM9CyxOemJa/wi7z88oSttmVhy1BBA3AipOSUW0H87dLHJt10nKMxMsVp1+LCxEFQ4/1f7rUthSeSt9lqr7jdmtFyGt70MLc5ZTMtVDLQG8Z48QbDSMggc/oUi8CJqs8KwD20U8AIftH0qvqxJiMoTSXGHFkmhMP4jbDj14+quQlLxGHN9TgZwda+LTYhEMf9wqWTbbQbUWA2LipX6GeZvvr0I5AigcLsSTILyKIq3cf1p/XiCA7k4VRDA3s9PMbIYLHmo8lWdNeZJSv/ywG0YMPfRwe5KPos/KIqHYk1UUsATvUwagUIYa3DlaFdLWJSt+Z/ybSdqNEX9vKMluOC0ZtK3JoL9VVpofc12759tClv6Dqhw3/mZKe+lY8wpUXpirS1nF6G4ds773z/Ps6G+SQ/mBh/aqB/pD2BjzK+oJdwT9MRqFKAos+7BesY4uvzNznPaZN+k35pWrxSiF0ul64I5EHamZVb0axKv4A5+OQGIk5gQFhgbmYOZUq0vnuXb/WSgRn9KOjnfl5FqDvZvafdnKtwnjRAzrcPYGSPFEzJMY/QqWocUeIz/bMpEQ3w/v19LyVXOyp0pUtP1kNj0lGws+YkeGOXtM93Zq/g8u2p8iGzVa6uwkHcIfyKs1S/pIGzPGg171aqJile+FgFSvf91/6Wat4iKwkpyE5d+bP2E0+/acUbAWFgFbK08kv0MaHlbB3AF5p92o2/Q969UCQO8uFCAT6YfmVMbz3fdMC3ZiaRIZAz3A2ZTTgitYZ654Q67m8V+61gAqc95R2g9gqzJLdeIMDPWOanB2EeunPu9uw+uu2HiJLMpBaqhvDJx0CbsqzKotekXRn4bakvvWfCiaVrhQq8orPBSA4nbrJ2fVp2Sz7BI1OsI8f15VHP+iE1a2T8tQSv0YqSp+Xmj4TKaVmqCVL8biNjmNPA/gA33bZNYqrGQJUlr5v+s4i2LWnWtuz/JuarsfnFu8x5v8ga6hd+sjumQ7aepDTjfZSVBcXIfY48c/Ou+G90o/M/M7u5WDlD8xGe33TmKtTbi76gvUeEfSnQpKMrEOEpR3q8SYIaP4rDbXJQq0CCTM+Tu9ooWRdDVt3sYCc6jwdcyPYxjUVukd5+MBy2PuzSe7PltfVJXmvpETG56dceKOet37R2/mj+Ci7aHxmgKT8EMMW1nIbugxkhvSE8+Yr+aKsN233PTqopkEi7fBCjh6FoE4k/foJ8qPfORFtdnVIhr7VsE+mI4jczmLvgQbxgFHbCn5UC6IBaJ7A/ZviydaLv1Mz5qUkJomWdGxsjsFu3HJKZ9ScI0IGvQGXJlUe7OZqUpgpFJnA57rVzJJ4lZxal1J7iaWTFhNgMft8ldkmGNNaYN6XPw/8vrvFltll81woDdWR9m1kfGdw4oN4OJuNHycnxOF+jfNTEcpPuiArYEGlesfgU5Pfx/MHi1Jeh8NidQfjKl1GV97r0XOJwOvN3II9eCW+NTatcNyoJ0K86nipsbVhLqWA36uiWgII23S3Tpvc6ExhpKss/Kh1iz2zfm8jVjCF3RchzJNearI0jPb22ECjC1UkSg10g464LcaRytX77bund/cNgz+YSwgaJaNdntqjCuHOugmlP6fHIEe352jLrX/qgKz8+dHCVS+JZ4C8zPFrwHDn5VBXxJ6ZiP3luACVHfrdFZxKeXQCkENMFdgRLrCIQ+lIwxyur/oj5HP5W5JrpKcraCZKNgFHyLP9KwldqQDoC1I0LGYTHzF77pY3J8MGIboqvc4hoExUj2HvkEzfe+98pRcsFq1e8vjkZ9oBJrgZgEx+RjYwskzAeF+DCWisfnEmPBC8/42kLc7xNLwTegF5LVXOyIF6sHYZHazvPZGagfre/+j7K16aX6QKe6LPSF4lmNiqdUJYv3hVmI+iXwnLFgVF3cAwOHsdm+kCk4H6LInHd+v7JWtY4S5eaoLha2Vq1pZwu5wGLPjG5EvX1h5KMLbYMc6XcoP9L0U38WMtiPgBuyALZx7pCTAqc8wmYFmxqwTZriIZ+TRyquUV1WvIuWI5waD399RT+JchcJeaoYbDQSrYbM78DtyFTI3jrakvFT9VJV48UwFwyKJamDk1y2c0zh61ppkG0Ku2WftiuYvVgciFAbjdXVcTfVnVutfIRv+G2gPfvJwEsrRU8dJZmQa5kJo5kuKGpLNwlvjZM3K+L/81w1UPMHsisX5LuF6NPA267pZn4YXzCrImJgUtYGM3GIN+6zbxgu5mrd8YFwPUBZrhbGmC1Qdi40FnaulPFhc8JfDfSaTFfa61mpI7xsRCcsz4N7wHpO95phYEUVNjfz/MKrtEEhMxwswF9k7YeegHKga808WBKwziExK3IheN3XbaSaAw2SKhA+jhIJypVB9vprn4GkdxvAj8IHUysRZ0o3s1vVPwh+YBalinCLqMpBjVRnvJiYS+/RwTxyp/nPkkofkzVbjLU+Y+r3EoFzcIZyggB1v9tXrfirDB899LS/L7Wsb2MdsSNodnHLtHxQa3oYRviNDcbkDqin+NFdd0b8rzBdoLmVit+gPmlKQOqcChdXjRbusDBL6h01iYmkWCEvasFRKIQvwQW0jt72UDnpPQlGJJu4xE4OHkD5DKpP2V7NRAXJapqLQU5p0Ucrg8D4GHFfLFORzdw7MY7qZnavi75NeH1ePI5XTPzPcthmPC2rauYX8esM8eEReJx7GzGwtJo6I/W1qFZF+onPKwSzH4eKJh9IFjzAAM8H6TZi9w+Hds48JuXArHqgbT0VF1J8Ti9Ctm+fTKee3AF0N0uDfGo/8OtHI+A67JXObPFpmhs/BxL+eR+abujlVOFLPBlkDsB/G7BaebLu0C8E/i/z1IEQiQKqlQG1l6t97WQkvJL6TuPSU70RsL/T3BE0zV8/gbQfYlqJ2zhPm4OQFd+VIyMwzzGtalP0Rw8cR2lY7UiRJ1HJRsQLhFPvBT0COPBLi9RnAxH31/6dsl4Y9+7ETe7wocWOWDbuP77pDS3F0zTKlBzmnj5Per7r9PblZi439VcnVFj0vWScBDaW6sn6uo4RgzfXKn98tHUmWDq/+a3MLI0W3Oyef8wkCxyTxjo5C3mGwSzemhCGw0xrtu3H2ZzOAXlqqzTFVyHkas+3YM8Muezhd9Tot+Yr94hKtqbEU70hKDKbKk2+MZ67gSK/UKJfQl5x3ZxsusowHInh8aUGjjfKNHLc0XUrJUJqNw3uEciwD9NX96FLNMQdI0gRSCJjajkV+qwVhsrVjPOsbzzACnTOLkN9ID5r+Q79cX8ZVyKFwA1U3vUo+zOK9Z571iN9PgGpJQBebSj2cVeXfsKsE1HKgu6yjb5Dfg8oKK6xdQKVFpjt4uV5iF4da/JrC0N9Jch9VnSPzsO9Nx27PfgErfJEBnIPYs6cxU51L3LvNdWL6XOzFsnHlxqR5xWjL4H/xi5iMvMmHl7GsOCylm0+BH31hYE1Qa23XHK/JMrPqCh4QUmiM9BUMoa749UZOzE5X9EqOQVgGI6Y0EN6eKpqpYB+aEuTmVsIHQQIGkeKA/hj5jaYbpBZjnYe5YjUysdyBfrnyrM4T4FSCB5/H7DQv8eSSFi6N6+naxGtGldHUESerRl5zKApNCQ5EEwL2mYIa73J15Cp5F2BHCJRpYxNcl/Orsbkxn6gRREp2iNje4arV3AIwll/gHIveShdxEiuC07WXWKfwGXAKbhBCzxob0uAMeqQU3wuM+erGfTzHzjcOEfVpQVY5x1+nyGCgf6uyF9AjXNyX1pfZlrflGl/Dlj09rLzwDIv1gzkrEG1tlyk3AUqcZXqWQNEHRAzxhY2tHmMQhSMlNpFsstFLVYl+dQePxtpF6XoNbl/OutOkxYwxVRUXO9JzutANKAthhwR8g+yjDjDF95TSOox+WP3WFwdm3Fq+SyA4geVrDo6UKLiAmStm+DC41q8EMHkCSETqzJM3TaGaS9EtvRfq1uTxNCYF8UKnaQRlmYBzkafCdVyuJUApEYNTcJR5aIIQEEZCpSH5neo92y9gPn7jXF6FZbeUfUsjzdPmyPQ4eADfabVzYZbXIo9gIVCiXolVSPj/VG4PaMQq7RZ38c3q323Z5F3BwS6esybzpKwnmKukQID4RPeCXOsmS5L2cywWY68xC/qmrcpIDOzAgqPCssVoc0MnHdpXmzqLuj2pKCsZrqMRP8bFw3eAKrJmj6/hWetR753sgnT36NGm7zbnR9Zu30SnzJOGgAh3+krMFl8hBt8MY74frX2Z3bOSD5YdH5Vop2qRSus+n9DMqOfzqy4O1Of+nYbIlLdAudeFPMTJNR+UZ5PA86PJgk/7PGhGAPAmqfYklCcgd+9faCSAOb1rpazVXE+vEZes9H4LxqA+1yeePMRaswWkWo1peB9hX/tabA3VReOwII8XS7cnzL2x9vetx2lP0LWOLPCX0uoWOmhR3ftyr4fehSOjVgfa05A2/3+i/FC0XhxEKRi0dxj9x6ZvE55N/3C/ZDJrawubC+kYSvQZ2BgRsVNajKJVAkGIcYCf4kb5MgZaxdvTx1RsEjFgr0QU23yaYHduuB6rRqV2jsTMvXqdIvgm1K92Id6SwqNaSaJlorcTCHRIVrqr+1/nWOj3pk/nUwzOUvLP9YNkrLOEo9RulSHNsLoYQnyo9r/gGl9a27l5MAXffwSe5ms0lPozXWAFVuS4jTQBWGlKDDKeb83fzpImTxyhsVTT7EG/JYQwz5M3bT0kYiMMKhiDiGSO+LD9tKLLKAVNq1R7N1AIpRpixX3ODQAitQL+ENBOJ+9uGztYOatR4cbOrdmNSVw6BpDZBvSyKPCdCnm60vCB+ahUuREzU+K3IvhMeZrT0UbiSoaQb2881BKLtgXvARRzvd4deBhuq2V1mP1/ntX+wbntpwdmS9Oa46xxfc+gOVBcRURdAo3TmO12TXXbidSeREB9GomQPl73mJW2pyKrlF+e0BSBx+arwsjXbCGoTdw38C08dhwsL93xN0NDUKTJPhR6Yl0R4/qqrlIw18jFTXNNlAVE16Fq6PtvkPbwI+YpBQQAbKLxBYsXIDbDW57hTYRB3mYwB4i6PlXXMiHz+RPI0aEdp4E4UmUPBQFoElExb+5SKOeNnLbbQE8kf0i9b+6T+OrPlFNd2g6BsohOF5H7N/mrYBFUpf15V+K6EYUVus6RqYYvwK2keEacouL2YIp5sv6Osn+Ld9OQD9f9AxtvKAxs4V9GynS7WyU/fe8IlsYVLmcUkZSkHRDnHkQvAfpVHe9qWdBIVVa4XWGXUxXpwnXFPL8JWyDee5gzyLzuwLiJC/kfLzg/zLj/WkKJi9H2R5UlSz/p8Vvk4tuv/Di3wu5uhRpSAv6MUIxhhW7mkEeWA9cd3ljW7PvfAPXth6YMSsshJbM97VWdcMv3V6NhIdw44kqhYTlmMQckcaf+Z+OUwsgIBuYahQypatMU2x3W4SpGmaTAv7YPPQdignNUjJzFzFWeIlSt01EcmAoqvWzOROlNVK4c6JmFyNIAxPQCe2UcSdyR7AMVgLVzD97HfcLoMz0LdPjmw9wIMtyP6y5fHy1DORYmW9zSUWOZk7fa5/x1KXMM9vSIP9Vg2ChIejyiw1jkngpVVXPpuF5V3IGkHlJ0DRul1LH62Fe2NsATb015JkhkMHSgBFSF8PdhMSkyCWkjHpd8GULrEKJkc0WbPQuq9DnzN45JIYPuAEXoK5tDOzFKsR2WiogaLKN1zXeIbornh+vqYafJ2Bilt3Gmc1KNdr6fpSCBDPJG1nEs/Ly00bMVILrjb24slVMoDaQBcA0JGjQvMDyh/LRVNTN/LEnpRoe/D+lNRPAAZ8klivCWhUZk9eUw/DT+VDiC90r5LMSU+lI1rPp3+B/XFKTgHg1iUCpyQbd65EGa29+WAM9AHeE5AzklRWZYhgyQ7hoMxzQiKFSGIRUyUza3b76iOZSwDJL932J5VmMppcsmBfQB3/Aekq7lHQ8PTgkxO6+IDDgw47yhq+4JFzb2snXSUMGmtSLV+byhKRLqX8+fAqSjhP+eL7yE2lNvu/42KTPqvSDJhxZ8iQPv63VL4B3WZ3woYBkQw30ppBqOeMRKm9bY6kgXWm8qHUKHH9sjmsJ9Frh+4vgTxRpruuffC6grhiueZFjC0m+sqvINgBkVqEbLZLlsyNYRquNnOAHurmcEbylYSEYDNSBbd7cn+G3qol9MJqUxrNEOiUiTHdcdng1tr61Rh+hwSTKkZd4QL0y+sFC/Qh54w015EYqVFqzuosyP6E3AmrkD8a0BscAi/d6iGF7aMA6GPBMB/ZR5mphz99RJ/8o0mjUzzHRbQqrD+MtNRpJLSuucebr4G9+SefZij77HPmtePSjpXy5gVlQ0O4PHmni18IavAcE5/F4T9wx6RbrPamDjMY9JqdaQbFhELbSEjHA6IpzdnZ0CLdvq2dQ0JYUJvC0DUYkTba4Eq/KgmOXKwHCR92altwTsufaVopVnaZW0ITgw5LxVSt6cOOuorgFo5PX+e2v1xc/IYuiZGn68xU4t0eI9RMhyoHTekS5S4rc1oqDuScneskYJj5zfxaBrY9iXrJTQiJ4QzOXJ+6U2PTg1UzWbgCPo2I87e5DWJI3JuU/d0BPPkW+oSqFuHKfoOxy2xt4yIT2SGUPigazqw9OBmdS8bVtGjQAaCDoAr8Jkep9qGp9etubKDp2wT01AGOHBsaRYIvWqMuCEKM4awuMjPDvAMonFcrin336eN6giOScWe5bvM1pEnshdsOhWPF5n6qWjDnjPLfI88dB6dbGfoQwd+1d0+mZLWEVFd8eWl9eKcq6pch4/J4nZOFtYpKYUsmMyZJSJzu8Sip9mXlO5M87NY4l7xBurzotrfaxTlgJWWBhGhU8UqP7MuMpssYd+gsOxRIjQQTeS21/N7xlY3bG6nUBfa+dL25j63SXczhZ+UCajLgptQF3ZEpeLGp/pfKHrff3G7APxjEvloASjC4KmCJBqbntOBlXPGnZK8htxBjcFh1pEEI9MSC717VnaG0y5tqMoqaloLT3FW/E55jj22i+bu16clnmQJRadS9q/nnQBxJeMS7M/wKn0nj9TM6yHVioOBCg1wgVAUgCkKBSkGGETAeEZvqltkE2c9doi59G4DdtHkyKt5PApQUdTVfuzzOhLhh8nP2cloxPNTRKoBvfQqQIMLAGJbpz2gzaQKmhtnBCfStqplYtMm6Rr8OE7fGTd5oEsc3MA8EmQ4Ko7ROw+hfUS4N6ce60OLHubJQWPdL98ZUZP8s3/Z3vA6//OSkciADckBf3KyC+5c7bfb39ug44hZwOLhsWRaTqhAzBMRvdTpzhSM/81l4G3H09LTDBG7jX1gTNIcbr+dYRiIAbowCq2ywVa7vl6S8tn3qqh6rOjmaogt23VB6uLsn8Zsxp+WmkfRqHsK6+rtvBN99sblQR3T8Gm0rlFohUEXb04KKkcvjQyTtzCLlzs7lBut8Zjhr17v5TFLLIVHk/pEDFYG4BQgPqChPYeZtv9uzgO2HhypnlRn2kczwaUkbfHY1kAHAL24L7T2gcIvKM+nawAKFB62WB8RpWNk+Ciiwh0v8FfAOI/fWXicfuo3FhLB2jdNbxUc8JBHmH2MGQOx5evqnZBdPIxURi+Tfxc2a9PNiX+c1r8t/mg1emBDJOw1kPV0V554fRa1/l/xwpnivgfQpghiMBVy3XGgQUvjFnWI9PTXoq0Aw2b9p2UnbQdqbX2YIU699rgQ6Jz88Ekk8YTlyEs3IDsF+DkMlFUUDWBKZap01Kc37HTsQ1rpHvQWsju3JeMi1jDbEosklYH+6QzSj2wHFf5ZUWrnUKcRtT3GCVNIpumpAn97T9uviinhzKBpaKL1wQoAQHmGzFyjNfZq3415Wph2ISKxN7yLJUseRMW769EUcgaLwadmDrNT7UsK0gVD/2FYeMcZvtEhjL0/j+GDm9HowU62rv4B+pi4pQ15PCQk/IuXHq060YwdGI64nqXBTDFG7J7KaKbh76dmxFzK1peQGMw6XMeVZN+PEFM6aRJzhIZCy/9CXEC+xk43HmV1TffzVj2OZ0/A+wAkMujusNlyKE1uAEELHGrySSkQvBTjoZxvPmripPSd5iJMCByZnoDMraPk42kfP/FWAIhQm6IKj2O8y5qFukRWbMmF4Y8GWiHod9f8NQbvL8gMQKBFeInqOqsOpdJcgm6szhCSfgbagjIib8fhYHLs2mFttdrGVzJfFYA5VCfCE62C/QeazThOKaZbjuxgl0bl9nRsJAQjDSsNpPX5HfUD9zC9ZR/rl46YUVQvFpK+eovgyEEwpyTJpT0rWUIUTgtpDgJkL87yKla0/AhmjiQc7f3BFYWb5JoXKBJSOsiLRfgCipzFtMbf/c9XgLW6R4GYCm2bM/8d/M4bmUVamRv/IKXNyfIjYCOEBnNLkYxG0Q1N3S0Wr8onoMkZohLZRXmOA6rD2grbM+ubo3FY2aQkidZ1vAWEObsl+xU3SmoI6Vn1mw/RpdJ0PyOLAtSswhJOrixVz9afmFrYOlqgIDhirzpwzwwr/ywk7IUTv3GYJ1zI8zvtSMsXzgypI4axskE0HPULoqvuuZnc7t0iK+1TCfj5eq1D8Qs/hO+lR44aiPsDzTW2L3hfi3x+SLVyCGzlPLe9XbmfzDrHJu2sIIxrMb91huyurItNms9qQ70/U/n4+TrSHwE0bdSW7CnohMnu5digLMp2fZwr9+25sNjwfOTot3vUJEjK/pe4ixLGYBmqbTKD0kcXaGPc/se2XDLq/Y5hL14g5dSKfJSTCET2bc3U6u0WAVbWEySpoLYaeCn08erNSI5yURe+81ztWXmpYGCzIMv++iJNi3DQaudUPDyLgr2VAIIu6pIa08rxSuNJPC4n0IsQs1Yq6J8BXE+eILHo5+S0YYEA8Rk8riF3z26DlwUkzwmAU4vF6bMJRJftcpuivz3DyZgFGfwP9Jg3UhKiE6w97D313KG6xZFXUnMc3uiVo652Oti3DXQRD2FzGbtKMfITROxK0bfP2rgyjSG3PJYnfmjP1vsjDDIqPKaggy88JZFPEY19uU+KXvo+FyrfNKyjdceUrG+2DDnzTc82U9QC9Y0dUgL/IL4MdyS4yofZVC4CDZjflytxGSoSpe8fWrHu568eTT3fEjA8Bu78qijsgIbH3QDMaum4oXZ40vbT/d2Rx5JHqrJYNaGmHSbESevNfTnSzqovtH1JBdQS+l/6ORxmwGy+N+60TvYzOmGpEw1bldU5QhKD57dh5g/sG+UaL6gbo8T+fdacssKngl9XwBD2siZv9d1NT5pUHNXlbS1hi+LkXeq1y9pTnoZTJT32x/XWI173g7/dahYgHghOgN97EnaXw4Ok/2ZT0Y9QrbAcZm9bLip3V1FG/dQL7iE3Z+YjRwLXS1k5qpz5vHYcuIZvZQ2rt0LBsdZ9o9yeH1spcyV4p+qG2FSitbF1H8USaR/gdFrob7LnRmUZIZ9Gp52mt/lTPVoLSv1btBrBwt3vxnEMan9lEryfZ3U5kb7EK2SSAUQnZ4FYlbSkmc6p6r27K/2Ghkk/ntC63+Ge07pyO+173J4aI/2juWSa0pC/furEBCeRizqWasSRJ+PZuKhk0+cdB3zix1EAv6Q3pwF7oJUDpmUub2kbZFBUisPYNF/PL0LbFhkc11Bz9pkZedFHmlvfgciNueKQ7GbR4lg7yEW7wLKkUY2DSASrgQeztpiaCCQWpRgTYG3Auo1d5HeWo9xEhZ00mPRXgbYawBjWPd6/XDsgoLIhAAw6yiIYr0jNuIXTEX3P5y6ZK5Fa5FnnZBsHvRle9bVD0+jTww5sQ/gNFKi1CQM9UtNYGR0upCBJSv1KKm8eo+4WMaN7BCcPuo4+SyxxL/WxYYr8A0v+jOvNp5WjcWEqzt8jZ/tKLgc5g6NIuTbuWGZUb6tGOGcpI4qXIqdKwoivkpcUv23BzGZmuHWLT01WS9MAeu86ES4l752bzC6qm6kWkQRADa/dGrzQZJ6BVpJB63dVodhDq4u/gxY6ydVGKhE7eNqtGcSIGwk1ZDaNC3CnVsY/BcdT4Xl9B1ozOWUjpUV1iGpv0oi3N6ETzPQfYFZCVLGm45l5TsHlQ9e0oBLerxuIoMLhf944WwUnneJueX4xp0LZJxzCESCeaUYKNa5LabdhOIADKFT5Pg14U2amhBYl/WsxzpzeTxV5hgBRU3iLX5qXZVlUXw9K5M8NE8LpujYDsPKEiVjJFxZkXe/akUbFtHqwIOu3oAEZsUWX9HNABnIuG5Tioa50crDy/yUq65hCWq1ZB7oUgh+n4Y2dauA/1cGNV+JL+EdDOKXSvqzgkQLvKpnDHZv2/u88uo5fmPWZ5Hd8I6WGNFJ5SZQKwRHD5QfQ1N6WNP5EhrTam8sgkHM7RqDsFs6kYf8MWMzPKLgiX6BHEaLCzRI6pHh8i83Z/qF7BH6jUgMQ8Kvewrzqzxs4GtsjruNk91GhDIffPMurcRfyrgSFOiXMc6x6Wl+I1WSfhm8hMxDLQ6cmQkMJKJSvcZ9uMgDcwVAhTFHXjZRo8wNKaUoaLWV2rIyY3xmcl2ygRsFio5JVHAeZ+uoeKejZrCQf/EUu6aJ+3okMCgEtqxWNyrWeRNQRjIj9uvBcSwazPdPyi37iAWgmaYvxw45KjpNoDjJevBZFhPwhYpJA1W6ifL0050x36bfizXt7QyGEe+LGUMytZn/vbvuGpRElrWtRU9lkJH5xD6Uhy/CXBP1PjkR2KSaQWL7Yr2bvnCKRLiL95BBiNW2OTZQHpcfpwk/6RR0NQNmlACU4BSLz76zi+Hm5Q7jjjY3ZWcWB9XbH2sLWmqznhxjqWATsEviciL7bgVuoUHT0zk7opLuuvCfMNV8J+xcUymGmbNFZ/G+lp/e5FBDcDwfHcFExs/sNdBdhm+SswpsqJ7k5EAWtm4HOSNBtPrXArLBpd1jmNrkFvx8i0hq9SV1cyyA1WkYOWTZaAGbNuJiQDiThfDdp4hqqWOx5CSObxodNE+0eLdge/kxyXFhOp6ZLKttpLxtaQMLB1s0hd0c639cmysH2fxpuxZgDbdPufb6v2W7DHQWYxzM+FoWiX88cdPLufXOUKnmhXAcF2tMfvozYZZnqlj4yLfV+9UnEuNrFyyywfI9LUZgGx5uHxPcRFNo0gS7m/L8n7bRaeCdFeUSURY4EereouD1KSVhETggFapW1hPI0sUQm+9ZbRoaYQtJnX1PUbAJdxiwipxtQHxCjOvBXsZjx6FdFmNk4uQMe54ntsHN+RWa9Wi99ADs5omDgQPywXszfPTJ8MGA0T0ulIAPG3iijKiSQ18vygdaEys7vkkEZsu5g8E/fBFDmOjGHpS1UIsq6OynzBXalIgDuw4fnIkXY4v/azezSt7K5I2nk1Ny19tc9DogXnxn47dUU+4s9hbrq3aSVeg3HF/NjdWq5jmlt0CiiX08VUGhaP+eIi6XEeBP4QBqUU22gka8hQzKvsqX23CzeaQar/rO1bvLBUSlE0AofxtOGrh8bqhpAJ1q0g8+DWXn2h5ulZZQaPyet3UWEyonJeYtMHPxZ899ZuQWroIk/Z0aHT7GVd+GRLCyNPwjZNoPOiKKX3ienTkiQpQ5q1o8xt+/yEUmH0tGYh4UczdhvnpMxmpwIbV8oLb4rSIsgUPUZKU+ocBNaJKuwzg/QexHir79q4ZGYrzKeGfc9qgx4efhNo708rWioBUmQVaHmzeLX9oztE4xhKG6DeWaUS+XtEvVeFegu/IJeQyb6ttLqp8PpMZ8CuojRRy9kH3V+XC38nfcdVe0A7V747uEeqw3nVq1rUA2L8v92dHVfdOVdk9FmfC3j7akaJ6yDUEhuMAR7HucCp3DWn1Wm7DidRkPaIpEUTmNVPVzMp5/2dfi1TLj80WZM1sgUbE+dtHxWLsxxUGCuujEwiJ42xCpJj3hBg+JNHCjsyL1LBMGfZG+ixw97YwP/iNETAvQhJPzHMttTl2qIXT5oEgRgpU6qGbnkq4JokAwP11Ghia/DyfJZPontf+Xbd2JZaDuTu6k+63ufYUypYr2XdZEKJ58R1fp4NOQWnYsM2zda1QnqY6YUOWKuJJ/n0ArIlbAdqKLVzoX/jHfQEnOEEKaD1E2xPguA8kvXTLFdbqt1ctBDnTnto/QQGIuvde3+bEAJy1U/2tk17TROwylnJ2ZyTUwAXWL/uVC7pXqEL/qJzKe8f6GpAox+SvMqc0PEeBnutC6lAKr7Jk0q5anzKUiEG9j3WX6ICyTaNZDWQ7b7fqK74S1kiXRg3o7s/G7AKGwF+RiUwfTGlpi9e+hKBlfLFnJTClbbhajEMCb/xBNR+dGXVQNkEjFRtIQ+IWPvF6/fSjdwRnGqadx77N2HTJ9FkSWSA7I69I+u6mcKLooiLbnwffzmrqLe7V/6ehNEg6FmYL4w7uaZbAJ2QAabGSjh1FFIiSe7kQEOd0nbppawfv2J+tcb/+TpB40dkaBEgUdXzgckJqWehK9KjUnsIQsrXgw1N/qW9xrTxkQBX11N7iAhr/wit20Zp53veFPqrAgqlEIQTzC2sXQQDmSG2OyrKX2g0Zd889bADlDXkI7QgkLcVQL9++j4CIu5J2AHKHZn6bcBn4b1FfoJISl72ehWwb5zR+Re1sLbUYpFKUt5qIfP8RH56BExhA2IsG7BuYWNNpWpcmgNHJxVLPCztBIqjmUGj+FwylLaVGrM/Y5cmVJIe088YbLYpmD2pS8my++jVN8J/EpYcqWsDe4COI1M+hEm7EzT1Wy6zuq++67Bkf8U/QFVYP69XQjlXjQys8gvBoyCwwSKRin7z3VnTJyqJN3KLzq4DMwC6mUaCqWtwIfuZE5ZWv0PKIiE1+T3x0SEEZMG1IDG+NtM8pFbcW+DqYE5LBWEPH3+H+uCvXtRa8iAbzaH3RYZPvhIbgDBR8nkeHxzaqneq1wIP3XphMSJ75QiabhNhUmHfwxMKgdB2k/D/ebkPTl7snW4K0xupzEOY872L8nPcY/mlBvaLON2O8+DTE0Ecko0Zrh3HEfOBvuE4OLeB/6MwHJYsZdatmJpJwumZ6Ip8uWu8k8wDu2cpKcIk3yNJCmwftFm3wfHIP6POdpU587pabu8XBHO9nAjYvc0hpgz8ZQZygX5W1bvX6aFhndquHvvaX0gtbfiAVG8PaJEXTaYw97i59/gO+OPNpJ8R245nUy8i6fWHLfZCSKhS0RWkLAfdM237mSGtHbeAQIA9B6fjZ4CKctI1FB/QkJK/SoAfpqyjCP4ENhJzFeIFUjP/K868rb7W5e4DFURYACeW0xm6T0+QlJWvJkDkUx+xxg8OYiUL4dWQtFPcOP/spy0Ua/HWlaRPzxToGzsZS5fLKhjxKf6vSOXHZ297G+hlWPAfb8I3xpZIcWbJk088ZRi/dfMFRAV+xyhrarnipg6fxUt/5bdd6IVk7ZartqKFpZ7QVvJmXD52tOdqH7ardxo+ShXjZDuXhjvjBlb3/tdRM66PTH2ItOIqQYXbB/6LPX3PYAfiuYxUbqH/od8RlaJo66h/p/R0YE3GMhEyvlanjAWeNK2GbsqrL6IsoxwFlXePwFP3cJkWs/5hvIKWjPkrZqlQOQc0g3G9Lc5SWxiOXYFGz4WaPsLdnlkqTSm/5en1r/RNdROCOC3F+3aOJOJPP+L9M5Asb1sJDpdjveZym+elvgDinDZfm/yVpqy4Y32CwpgFMsMeyhb0qKtNxSFiu7KgGDanfj3O84I91bIv1Wy2IiNJU8kEiZEdsi/L1LzF8KLPFAwsrBRVHPgEqAO0D44e/NFimI2/8jfOxBxKu8JZynqa7X3sF6MaIRYyseHHhSLpE0QqZpr/9VuzeirbJjVvWiB1LENp09MJUT8sDdatnK7cIWuDHzHzXVe9sDSjmmG1G/dFaVPmx2vrfnw1DudY/hlC6sR003CeMvW3RGFStz1rv+BlJaLR9UKraAvmXuO9PqcYt2Sn6m7kydCyCOrXI5MBWEOf4/+u1PFhmcEqz39GvoQQuvd+jR0g2E5yGf1QyTb2RrkxdcMPqYlivun6z6ux/DIvosyovrY0OBAYguZUKMmf2JN0NF9mp0D1GmzOACxkLJrzz00vS8hBQQm2OugtOvrUrFCBYTxkBeLKesaJuIk5Ty6molI3XejjvfX3g464ymTBolkzGTuksUMcxo7dN79rvpwRMx0Xan+SuK33ArEZ5NPU4DrzoaM67QzsV43stBF1e9Fz/4iPp7b9cco20HwQZg1XPjDMD4QnRMEmn+7TC+sgkmNdwhGEpgWfwaStva14B+/aMIFyjmaJdsTBIunimMTrUOwOFXDQK4rSq6OeZv8+rKeG/MzUSNrVdxqPsbfgiBaBprm+2XbuGjCFOpHHwE9DZQnSj9rUDIF9EaDt4a3SU680jgjdIyOuYRKpuiezdO5knKLyethii4qFEXiiQ0ovg8I+NCiKjbGUS7bK1/LUjVTHVkussFS6j+91hv7X8JNbc3ONUW8n0PjSjTwCvoXs9hU9iEWzfaxc+kZQN1cwbF9FZUu5/ZCRdzxvtmUL74nn9X3oVmDTaYMzGuoI4tKxYvxXU1ewId7WviJpPk9tSmIk+6sP5kKbkSHhPlMMYOe0e39tcuZOz567eyeOZ1rxRigvUZFb9IAtJkTivSaVLUsqrjoLSMm2fFw2MpObDgFbRtf3Ci8PFhT3e010afzxN1PhZkFSiIsZi3yl9CKGKuAHQjcQtUFa6I3XXVzP3yuy3FWdZQvDp5BONobIkMBfDCavacpeto7Fk8kPBesyC36Ot3pfsvkiqLxKyZfXF9iRxnrLuZR4+ckLE9BmlPpszhANKhuZNnmBLEntwKOFymHaMtk473oRpcu5kMr+DOaPy/cfvm0s70EORxxGi4XEv13IIXyQnlRbZuy9BvPEeIIrXwmZOL4422DEdoHlgCDQtQbnddBHN+lA8aO2Xr6dRjF+hP6fEQBs1keyyupS9cmnjGLJ2fwUHA8Wb0k4l3ZXbOYxiUsldV/xOtJHBCuT4uMfX7BkOka4e2lz37iA3BZIDNAlXDgGkradtXuive86LAfX2rN19Dl3kYp6csRHSl8FkW8yzvPys0j7LVirbb7Xl3kW0CljNc/o11Mq/l0Ymh2Bwxo/DaXAY+oPAyiwXpsbE5EMEmdb0K3suiRx4d+7m/KCyc/+7MuNCF3ToNNmbbRa1c7kjpIW7tWXApQL2t0kIhCWNIlML8rvo9oy9JMaINLKdOpEDwpDdJKQw3wK/eQ=
`pragma protect end_data_block
`pragma protect digest_block
e1e263e850999ed4ef54e306644f777b3105a1a34f97f500067ad750b2d1fbc4
`pragma protect end_digest_block
`pragma protect end_protected
