`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
MQ37D/dwe5OaLMPNOHGpvcJwyW0otpOU09S2WaZXbohoITg3g3RFiFW0jZmOjcjBXdq+UL58E48E2H0eRJNA3OZ7kRCQdEDaLH9SmtbtsJaDPbPZWIgW4ou3R9ZYguGvFlZQ1EYuvL4nn6mHokk/OQZwmKqxawfbfjtQpSB9hgf+CF+SnDdAC7PJhBKi8mWZ/1iBkcKw+Na/+HcYLr6cQTQxJMZOmRpNfnKm/qa+eVypWUp8oMEDYNPsIhql2s/gpYSC7fadEBC2bD+diLYCRa2Sjj9VXfmtZoXw6O7ccvGY52Rm1US6jnbW2gZFuj3rXOHegqn7w7Vca830375m85Siem6Et3V7KbWkhFkFANz8RdmHpq26eS7sTccM5SXbk0uS5ZLlUxDrdYKdeuXp1oVDgvRNizUJKILYcyk5gAEc7Q1pWn5Na7uq4PPyG+WZYGS8COgKUMHvWb0WW/Npm6R7FEtxDZv0jSkXoSXmRgBLDfoSGQ0A+dutxt3woWEmZFsAJv4oWYSZRUaGAq6nAlgNKJI3IrJ2Rh41TUjSUrY851R4jdFdhD0mYEvKX3WJlCaq4hcexIDbJaQUDj9l6yqg2EX3Ek1vkJRsoAP6Ilq8UyXfdOMXf3A8kkq6jAUmip9eFcln0rweCxGGqKQHItvDY1Ic7xeeOzGr72QQ47r6uMuBKwtf3dEXjgqfUcNZgQghlN2hNBgIuMGzz0GyBYOt+ltZ39ZwYiWsrZ4b0F31gPmzO27Rh4MOwPK0o5aeeUF03PU4GnNbX6fDYgjVNpUBThGWU4oY9zsk09PyqNR/+2SJILg1+PFJf7dIwmuQUWXuLb/i4iV+M9oP9IlwBZTCZwT7fDjCWkYV48Nnh3eh+/AroLAQw87L61/CnYZAOfM98lP73XU86rYfZyzAqaqEhaJf5rHJyfssvNY1+E6ycnUlCtGeZptwGIzE9yVzRuyzyIFd8v8v0mVie+GQWHiA12bykWq1nKcCzEAK5qnMbwyOGOpbAjis3XFpw5lkOWjuFyqUP1mBmidIqb7M63T7VNU5QoA/qln7GuVpAzqfWEO1BGIpnspAW+waXsn5JNtOQ/AunXyKlUXR85UD4KA89v5ejKw85sgFQ3wuE63f4ZFuV5ZhiiUcAmw3WRAtzWXJuYu2uEAr1EyU1AB2FuFr8g67x47opj93cKBEtnfjxvAO+w5KzYVQUGbKwJNIcyQ9Up5R+VN5LlR9TuuBhiIqa2vfLdLkPRYWGWjdcJ62Snjb/u0bi4Rxf58f+9cHRVvWdajcEKcuUurXNsGJCz3BeN1tEuR1fpdDUJrEzgQJ3Y66B+0H4l1gGnnaVrrfUrxxmghXh2Io1d/Dg8ZvRnyzFC/AZvYH9TJzTIybUlSloYp2fyZ6uG3o1iLYj6/49UJ9Kshg10pgs4Qqw6hvjT+qx8TV1r2QxNVsGBHCU1w9Bhjw1d5gLQ6uowkwbkXegNqDkmvURW6iKhqiOrAnd9z42sN+RLdLpOkmkUHEq7h8hWmDxk/MNpYmf7NSbMZEiQiutCmp5ohofVEGyLDxfPwIDqgD186EIITzHa4+GxdhHTMbmunilvU2h65CcdaXza4g+GdHRMpTgVv9u6R83ycJLmZXEXVHbIzPf9B37peJECHjosHs5q9PGtNKW3b5MdwxEjcaGR02e2dAEpQvIvH8K5DM73cgLwX40oqD1FRGasGtG8TWUpdVu8Ao7V8ix8MVra/jKYKO+HbZStIXGqZuK0ChoX7Ek4gvxHRq10DYecbChSLpAL5SQ470HC96Q6tB8vNlx6/DWUZkZEz7uGRC6cpD+sGT9iJkOx2j9ULBZUQiyR+6fQhUHGzQMt/e2lWtX1/b6F/1fGhaowP4T3Tvfvv6UIZ3o2R6VaQTY9ybgMUlzAgeNuJHMB5o1NC2SPU+4xDY6lae9hGlAJNJoFmzz8Yy4Xjrgu5fa7RmzkbZBK45sqRoC4zLrGf+qAaCSeUpyEe2cXp+fIRBgJYeP4Vro3c0fW06ZGdwRKtsUs66wbrF+yT3aOkE+D5UUgUxOAS4QSYFYtNGSIa/vFa4LwQofjZuRh4iCkBFrom83WZwewtn00+2BZcC49msRp1rMAnWRutnAFMZIs9GR+w2yoCC0/NquLey7NpIs0a1mdTsalf4FBWk/8zF9WooI3jHlvfAP1+lvrVE/BZfYTePL6Qgddl4z4S6Zembg3yKZUVjQg1uWnoLTxelKzEFw/ZS0y+hbooLQ/OkwOtJWvMe+3ZZ3u/r15b6KXH5KWl4PvVbJVA2+EfxNZkZ7zvFrUCzrkCJJk4DGbxJv8aJx2TsTOqrNTCEzb8jpRcrom0qYFfLvnSFjv+fYDmQLLyP2B+gyT5gjRLAtSX9E7a9R2mjREWLoV0i3+8tMXFe787wC7OKueqI5ETakLnj8POtfA/xjQlrycZfyQxVCEpR9zj1n8FFzFTS2LNljMDuKExVSGurtpAAF8q9zjBnlfiEaXU38D7IM8q49q7bYMFq7aO/UImsqmQmjIrvRvzN/fgYcRIVIBlbOQj+RMzonMHx47BUt9b9ydYQBEH7jaV8YuHsm2RqiP6jKh4N6yaZe0D2igHHbwW3kfp2adep24/8jB+RwK2hmCVWadgG3jlNTbdS05y/8FgJVMtVvL7TLGjw22LCOOG1wvj/Gfg/MPRrobXS5QB7h+7A4AEiVHi7jTXc+NUENnkDkDl2+IJz+xGBL5Lggj6tqfwhQfKzhPgUDZTi/4FoY080HBRcWcRnTY3OATZUy+whzANPuOy5+qcNr06Ixevg3zq44iEz8lHMKV4ar7+7pEqY5Wy+KpD+7w9ScpRSn+kzEp7ODLB+YnCuwwsuDptjPiwiyXlF7X0vBkzGI6Vrj3rrNp2veR+lbEgYug7qMYy3mpOod4AIpHT93RBZyQ5Asr3ckOCnlR32hhL4jR3JfTFZK0HGSA6wDVfvKWrI8gCKysMam0wgh3GRjnqpekirhN6BiERoYWbkBTvHu+arWZFcDcC1e3urIOPydC/hjBC/5OYZU0MS0MCFqW8/5tRjRswluJs1yBlpS9Q89kf2dhJWAExHrOd4qlfANqDF+5b9459/FaD5Nn9IzDF20xSo7YHcTMqmb96gHzXuX19hBUA/F8v9h91cdtjoFW69PugmyrYIKX30PLcMpEAMHBsc24+wvEscptoDmVoKsMoTBMl/Z1Ezwnr1Zq9KGOLdo7iNR+AT0RTOHDg5XynKDzyz4CvlxjEgnOmdOGSsRyOT/V4ciGWyKLbxDUXfmrz67cZxg61ybJk7X9i0FH4dMNo7lfPIfh7NLumxS3k1riI2XtfTAiMAUp+NMGG85/F83znZIFiucduiGOZhOCraga/irASZABtd2ACVnZrcP7UPuXIvIAqU3B+z1TpqJH24jO160NqB3UdGb3xz7Z/8e66D8G33EVzJsXOttMhdzghIK78g10rfaU+AP2/VvtdKD5Hwn4XUoSqL9vZEP4rdY8rovkQi06c0jU3CwQoNLbQCUl7Ia1aodgZ/ht4bGvcTRpgQC4Fmm2vlocVwdUYywGARGaH18OnXvhtPj7wN9NAEkLahzVqDiWltqg1rhI8+2rIi6rqPyLxJUtVs4nK4qico3Oy6yOQPkUVMMzSwfBs38fD1DHCSkwZITvBwK4AZprJD25w0RL3CkckrK3rVmebcuBiS7dtrpqSjBMTb5dUY6Davhd87dDhbvuSVoyCS+yYLBu4+ckemG04OZ5/3wSqnTu1y+mmJqm3PNX+zFZEzDsB7JkG/WhzVVBXW+Sdm8dbThgtbnjI3tXax9TlNLMU4tppXiGvh9ZIdiAxL8Wp7mNQZv9IRzIPR0Y7xe6gRFYQf1/XBliqkI9tz8k7/sQWwLWI5gribvreySkmQbthh/zjqKDAd2vFFt/6gnyZ1eM5I7vaD26rbUEy41E7yxdKg3Nnk1tf4SR9hmW2O1XPBi4Jm51lLjCO8Bdy5JEciU4bIg1jOwppQUAWkuc/1xTNzXqHuwwa6lljsxIG3Cvxrpq3KCQ7WcyU7PN8S9l9e1yD5QrJwJxpiZrLCRTy/qIkv4IkunT8d4cU7tyxG2C8riunUvSet1zAoqaAy8TGILi6DdtLuiX++wFTmYzs0ZqwajaCksrJAQd+8pnYcMjehEWl1CFRCw6NiHI7ilYnvGkm3ics4591nM8Xg+YRf2May61ke3xCnd3IB5TPz0smCDfvKSzcTquhbvDzRfTjAmmJX3J0sm0XjtaNUgfG3zkWITO0ZZFagjdcEQLlbk7i3Dw65YTgzIGsFjLthUbYcOMPSVV9UwfmiXs0YUlsoZrfUkqpWXl03z5nWSFUCi4ypvpJ6MwTlvrfyRLsNbehDUx4yqOObCuSUPs5G3kUh1AvnN1j5csZ/6ALel5DQ4hg6QEy8UV1TrUAHBirgpzMqG1CU7eSnAbZU38C5Ss6/aJKco2umkVLi1bqiW9uDzeGyTwtiRzytIVFNZI8OWELRmOjWn9h88TO2a7UReBwTBUE4dG7YUo4wf2AYekLSCKwf1aulKx5vzSuzD3SY2RfkOAPoa3DvpsOW/bIV5x1ot4X9XWHOUyi7kRlsR6Z/2PyWmB+4t2OQX/e8OviPO49mh+wG3UZDecAMYpJZt70gsePF42YZBaMEltF2DSIV3/X/wPlMNL6KpsDGbRGbujOnduL6UjtwsjWPPnSKVP7DKukXZsbTXUOzFOYyPscCEGyIcf3UqqiRcYXnrWmol5UrsygIS1fSYojerylX9sFBzfslHgKR10dXgQkPir5Hg1l5WA152jwKSBQEimg5na9SYyjEnkXjKvNBF76s/1PUC9SONmbugOzEPrI1Ym+sAyf8kSR+v/nbiVzVcn7TEsXUO+pD29/QJ11Fx0mz0ywrtGmw/0EJ/rsw1DFQ4RDnoT5mZrTvpEIffGcfm1sfndUeP/f1ZuVzP6OAYNrur2qrtYc21qZ232+myaFmNUmbdJBh56fVCx1vPVgvEpyi2Yhm8yRRwyfs2EeKZ7gZ1RCeLeQPJsIFdvUMdQYUEMGdQnkX+4oDDIVesGJ+LK7Wa2dAZgsB+K6642JO+V7rf3g+PLXqNRU2ZA01PhaE9D4zuayd2pRfjr1u+3AJuSEXMCnv4rmJ1nn+OYsbr+U1eRY/eGH/CqoI1rrNAkBje/KDmOWhrk/hvOCaJjNnGPmGB4tCZWBHoZ7I/Y3eaGmO5gtbWHBS+ggvs7XXKyXy5gjnm6uJVO+IvTnuo99REQ6Ck1HA1FDhE2eJADYozjgd3Nk0EHVwG2dVKXfL8yIBOf7g+AAuz9nc7o5X5ETmnqTfiX+3TqZxltc8m+31u98eLiDZAbVUidHMYiz3kUGwILJFY1H+b/5L4P/ZEWEcMXwLdAwfv8bGzdsPFJcAR7pLyOJxWuAIYb2v5C0MVI3JUYxocK15qVAkkbdL2Nmx7tzq797JwDMgbaLofgBzfXFAna9n8P3S1DXEhKssBertIuNG1Xwzhbk3SmA8z+iPfkJNIp9nY7YJRlUJ/uVtGKTnoZofm/j33hChrKUY+bQeuurxhyM+0jFrXe0b7IE77czXMzZVCzyaWGMeF1KkNU0uNBVeTnkvnTUg7FMHIfjRWu45CH1YdpyIBw2X8hJaFiJvJwEJq5PtC7RSuuw84ljA66vb+qtcAfdyzR9Zdky5+VI+8tRrB4yzSIgfGP7e1zESuKk9O6YZ0d4Zc/aMktmh6sfguvDQ1E24KrlxcnA43dr9MjEvb1vixrCPVwduvYSNdfLmMClzMH9wv/5lu0fbEZvFRy1SmATQ9xdd3eixS64T8kknyYTx71Lgr5cDhIpAyIC4SubYjOKS1vYdaXqZufMC2/+PQMLsp4NT5oRbHykPOfa1SGsnEJtXVtlhU0bP1rXy14oCHp6Dp9K2RNCkX0sZwBBGqICi4Xn5Prx081pOVhy632aQCoOrKRBWXWxhGQcyLuOGcz1/6dVsUSW6gCeNXt4r1js1k15al6SsQSwlLJh3UDz1KrNxLBePmni7AmDC42U3qrhMYWyK5zg4qYqAA0ZlPpqIf1COD3oyfksNsTgP8PU/c42bRaE/SeLbY+nJiofDkZD3rqjgqJlcvwYDQzu1j7EL01riFDmiKWwk8K0VNtwuyKFnrG8IBF+N0gSyoNj3fsG9vLxXu3Wlz1n5f/jnf0BcK+wi8hn8Cvuyk5gvChK2YsMTQD2mlxxaGs6gOgL7rUC65cCvb3z/yO46dO37f12ypYVUylBTKtGIvekYxRhIKTDRVEen6hKoiEdwLiTLjPy5Z7yfNgQV9UwTOI4sWkMRpp8vgh07sJtRPUmgbzv9x6sPa1apnnYOQMXGp2vkAE7dAPNfNCs85cjfDrxq4NLUh220sV5WgDh7QS7o3Qk3AAwuAxm4Ap3/zb8arKmZm/P3UPzetrySMNAP30XCGu2GWGMDU7oZ6P3XDgg3CCFbMkqO46txnd7kRfrGfLTFqQ4Yawd9MFnwVZt4HvVnsMQA8QVef2H++Q2nCWQ3h/b9aZh02m5LdKridMjAAJcanEe/fz2r8YIazuiN9cYyqMCySP1MYUModSdvG1riYG/uR+NTy+qzd2+aI8hpJeNDI5wwZr1pLp58qJnnu44/oYkCzupJujDbjXYxa4pwcJZ/0IO8WszofBpvo9PbHDDnQEJ4AUy5tmWrE4CSATqhOOMdaZZ0Nmj/nYzlwqJOD3fukz6bO4t2KIW7K+aYhvcEN694OuR6SeE8Q4FW4hfsY6jODhoR04s36I/MzeYX6F2oT961M8O7ppewsJfCy6JRQlRcrS/6gxjbw0kgnGkEqv89DnJrxn1C+ow5VrmMlQXzycB9CzfAJiyAXFs8ZkiFuaUKQlJdmzKcBMKWQebgoYkY5Wn93NuSc5JQK3ljPJzxBCV+hflPNBu2BgBIWm6rykAJ7jO/8MPvMvGSVjELWDn5ItDks1ghNpsx6nstjXX3yT0jjTA2bly2BHeroTz74OJaL795z/eAUr1N16oxHttiYeU95l/26pg2UvjXmlXVsItadJ9DnGqaV+1lM5ZrfStzhvTAqx5HYdgvI0Q10kkW5fuOV8mlnt4YiTdWKaZJqlFaaSLI6btSMC8u6rGX6TzjsnQmMDVZej2PeqJNubzSVysSY0fnlLc2ArUw03XZRKJG3XWQeiroZSbVukKLWsEkrgQBF7r1WDu+pLvhAA1B0YEwq3v+aKVX7a0lCsU/J1BoutxZkHFcGKUoduF/5RGY2Z+PhH8e3NsaSi0ve09hwvep7EkYTnLrTJMEMBgN/fVBgTVDkUJ+zCTLBCWPpCzN4qg6U+RRTx4ZMX/vVxi3BMIcezOhayxnyXeXI7ULvGRfOdVp8jRftaJzXIhHa1p6FDT19f/G6Q5p0A1uSLX+0JSnEAFiYLG6sz0z354BICXRL/YDfqqvnpQ4MVtrrWg0Isg7+UbIdNhfjBPimBgTK1F4b2/EFnbE0EIo7vTGvUIfAsQOfP/m/GU92xKlV1LDvUGfSUS6t0vVU8uTA6dXf7+uLhUM0R9+6YDZ1bdU0POwFCyTw916yi2lousoueXiEFaNtharoJssQXSyySa8veGrjRId1SYa/gNi9nJ7ojeQTzXBXCgobtLBlEFfUqxjHzleiUk+ptaZi3GBUif/d48WUhJDKBVILGP3RTSTuUy2lDE+dFtHP/4Mmz7uu+aB/2/xvyADEOFP0bK/8dfKk3Rn8ZNUsDDIv5835uW6DiUKR5RG0R1skHG+iSen0zoDIstr7LMN0jr8WhEIazWji0lJz3W4NHzV+Iv8uqA9cojovENTS/qlLaa/4xFlpccdKQFpSamPaStUEqL/Cl2ycsZcNhzu+taNn458RssCQrwBk/r5apJ3m5CAED3X0wpGnQwZoRGjXXRizgSKd4q22ZNtMD5Qjt/lBNzBhhfv1kbAetO8KOXPmqQQlcECkKVqfEK70hOdpj+72srmSDiWXqfA3SDGYsA71Wv6v2i9oKRdfpSdOtBRpis45lCWdkHlTCaGFmYng7BBJPgJK4eGKd9b8qTKb6cxN6IdOBS3yvbOv5x6G5//o/j7pGVWS+kNs/szRE5u4j9iPsJrYldl/xDtA2q3NH302+Mo7uH3HqcbYRZxcQvY846iqsMyaD9n0WMeDI3wpPBeKuJ7nlyobhf6mVZpkpyl3WTjv5S1rwcC/B/euxy//kmsNfritISspXkVhHtbPZz5D0vIXMAdSgpsWkshJSFnMlqNcsv2CG7d6zLJ8XevGbBTa8txrb49s76dhW4vgcjv7/KGEMdP5IeMHxhbIKQExV853QzCkliktgkJrOf1gR6wigCG52uM36qxCV6AuEjrrsW/K+D5eAcnl1meY8FWosVxcIbZnhcI94nqA3PiuY+7gW7LtXqBU5gWP9gqHLfQ3D3+wVfTXjdMQpJAEYrZ5gQm0qSiro1padvNNmo/VdgIV6hnnNTm9Uxf70huKtSiV9HS/vwYnlhGXl3mFl9gQ2Sp1LkLnH+V+7iLpomrE6TxXQmEbmh6byP7S50ZWBfciOP1ApAhk9s5yWDO7fPX8wySP9OZyBMeaGUCWhQkG2ZEVMLjOOIgLt+Bj6o7QOgVtSz/Kt3NH0QZ0mYzwAoKWuGM00tSMutP4HBkHXrRop6TKGVj7QZNOQr2F54R42vK6SmKsROKRnP6Gc4W1klYzLKT3QHn3imP96cBY5HbXYJIb+f0mXDlsKDWgBIr7e+xSb0/Sk9H4eC7QGtnoWBIynj2GjwE+IstJLip108zdfd7H6Mf6UI0vUwPedczNzcBoB9BtHS+CPbMeI0hV9wnqHfIPNBcoOwstRR+QyvV7TlG0E6INeJf+vH1OrPz6kIeA8kX5rWv0+cBN8f9HvztWmIRoakxzHIFFfWH9A2rImzs3uRbrBtUmYKvTApiYevjkbHvrXnNX5R2+luLQfDe+74MH/7JBY8SlzI14HbDdxNX/BXUyzEKRq7dTXZHXbzBlp8xcD91Ad5pWozDqgpMtOa8wF8gFlew3S1pAoTWsYAc7lYUyqv8ltxt+7emyqKznwXA4Jn2bc2fAAmYPqlnf3MShqoyWa6Zu+ZeiZJLenqf87iITjpBmE4vGxtpziNp2AF1Cd9Yc+vikxSeVdMqOR8xJP/jCcx6LI9WhOisqRnSTo+jAIK1YmqBk0y+XqDM3xs8oY9zwCU/cMs2BF38k99q15v6q19LoueiGSSr3V2uJwcZvCvtDbRP2TSzAH3kKQEzZvHH2NtsVOlqw1U4DqPd8obAoVsGl9xqmrFBCm2VYEBnSawHV4BOdTvyvCuAVBvMWY0q6sDviwuYbgUo7UWIN0szxX4yn+JrTLHbRsQTfcTxkiDCJPw3BdE6V/zDSBIFkUjB74GkEVvlu8Q10cJ3DUt+wlgOLwzzldgpzyX1CwLdCg2X8MuTlnf1I//QRhAk/q3bzhrusYPRsPdg68g11pzhzh9ZAj3ZFg3+EawhvkFuz39SSnN4ghEtJU3ZZwKB9GuxSazr15dhIkGYu3pLpUSQ6YJ4REeRxzCr7zMQDDHUW/lHV4iICjs2P1T+10RtDygvkic8WgroCntX2g49y3wvmzlcrlqoQSIqw9Rsc97Hq6LlaZ/PxsJbNN8w8gD1vdc1xodUCdDZEwW3YZ1xUvBogB1ZrGxQUtdZ01G5jpelM85CMgCL5HzsRaOAHeBmGKg55OAWYNEJRws2cw1nIR+8CxHc/IJvWKYd14pxyty8VNB+ozABp9JJXaQSuwANv8loqnzX4xVksGuO+uG9IOQCfmXTgO1ShR86ATz8yXPLSPs8JKy1XUqQADsWAlx8bNIJy9Uym++lrsPJFK5ZL8xNc4SZCvOBDtYpty6seB7gS34E1xY1prGjHPj2rTOvOrYVGgWa0uQe/vKCOIxkCD3dBdSeCoEcHhwhNXkqjiJT9abBOg6KWmMJpcocbY+pQNKm5zMMJa1AYevhFdZcBsaJFuw2w6JRjxIPOTgt1kFQen5D2SUO2OTH5QhkA4boR4Ayu7UFjFmM+O+DBuUvpR0Ja31rbXi2hb/ANhvdxkEvQ55wkfERecFYYSiaoH9lsmO/TjPnHfFLWCZOnng9sfphzpL8fcxDdgaoiVeK5bDgGvHsFneYV/zKi0dapTxN4u0stP0Wf3a/yq9WnMWU4FDfcr+w1wSwqZ0B5CiA1uwkpV4Thpu2+et7rroHRlM9tTcLEXivNEJFcJ1elcsAFI2iI5BrLuK/IGQyMpouKwPxzeB9W/KvlxotP8WFAfRSOtIWEzNRbhiFxtkOU2FykQw01caX+2GWr2GhG7Gy+aAgar6Q2JU3I82A21GV77opEh/G20HhW1Ihz8VY2sQrKLUZYuwdc5lrWfqWXAGfVscjjbXqSwsbKcnxKDEkmw80oKA1alpRHwpfAToQ468dgSUTptCmEh02rymkW0VdicXuPsU8laPk4WnTKHLMOTkUf2X6DcvxCMPe6VJG5eJvFePJDJbGpEN4MXMAlXhrmDEE0AR3J5PaogAqneJcaaDMxni+Mt+ZuSK5GDJKFzzA5Ct0e83jNo4PkthfWelshJ8gDl5md90wqi7iZkzRLe+nOZsaMGc7q9UdOcTfMFO9yRfix0XkGFQdW13690NxpBRbtidUlR2YfpDqxVJezvt30XDB4HCetcO1X3UQSIEU6XR6uwMLl3RSqhqwisBtoAck8WaOlcX9hlJkI2HRF5vpr6ynJMF5NIvWNFXlXmV9Wt76IY8MvLsdn2rwyp2WPNR/cgoAraBoW/+CQ6KilLUXxaG0P4WzMqKErxAbIcA/pBPatpwnpdG3aEY78qFNKmUfNfg2F+l8zUSPv3HjZQo1A3ulXkiNMOyF3M7ZarUJo77sZXWbDj+ewjn9jlnIxaLkQT4x7W/KDlXjglSadES78wc0YkVu+n/mhbl0kya8REXI5orV/RKNTVtG4S3fDfqomKAz42vWIkz/IuiH+DAfcXdRHGW4FzncBVxjWCxxls7rz4wY9Oc6/CAtTPvecqZRumlTL5zLpcq/LMQA3yCiu3Rp3/4NmWzMPgPzmgxojDvC+5NGNrI1fj9/wcoPREdQ/slbcEXAPpQIw+QgQYQFe40nuMU2ARVNJ+B10kn0HtSjggSeOSNpr8ccGy65TRs0QIE/uFLbo7EyqojBBSWXDcb49OFc47w82HfwopDIbY+T+TTMS0DWcyEiUmaz0BofSQucjkHozBkvDq93jTV6rLIV/HbUk8vrbjwQOop2a03253u5CG2U9Ub22FQozkjx7Mw/Kh8Ne3l2XzTMgimvD9fg+2jNB16MTzSVBmncdZLu+iS1xZeyN22eEQ8n84m4/sBHZfsU3TOiQEkl0GwErMABRT8WBGDHNAmktn2bcr6JqgGCFDxVZZtrADo64NXfEYajBwjKu7OSZMWZDF0kJ+LkvfNq1lP7LYjaU3ibOAQ4Uw8l0yPTgwbOxTMuehkBjZMnmMocQXOEqtLzDdo6b6X5wF5+Q5Jc7jxT9tcIZS00RjOW5uq/aXdlPS44tmrawVyF12KKaGKE6eNiNlQzJ8+XcfZAQKhpJoJ/CoBPduf4hTYv+ljRy9i4m7U0DYNSBViBtrrW5HqwcHVHzSQtMEBWJSLzkRfDWdHeJGbUnB9vWmBvwyVBhHj8N1ZoNVAncHYlsE+J1/XwLdStW4sXEcQRnA44PaheXlPAGb3J0/6PE6AUA03x2tqHhZw3tvuPhh4g/AncuYE4L2JmzD8oqr4TAfcRHjcfuzIRT708NQmnMIl5TSqpBioaNVLq0ZQoqJSndtBLcNusx9g=
`pragma protect end_data_block
`pragma protect digest_block
9e554990da3e56fa85da0b3b4d904532ce60907921de2129c6ac7fb90774023a
`pragma protect end_digest_block
`pragma protect end_protected
