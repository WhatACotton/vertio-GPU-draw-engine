`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
H9DE8vSj8SCzBV0sYkRtV6jKeNng3OeaIRqstCsvolU/qcrQQGwnXlygMfMGZIrYnG4I7bbB/8a4Y3OpxLO7KB9HvxC/Dd3J9OGgiGsqkHwYrh1zB2/z0fLASYl+X7JBXg/2mhIRm8ZwSKNciQNY2lzPy5Xvcvj9/IlCQLzS1IZ/k2RYKSSxX1iAzjUS2W1ePMQoxWsicQyxNrLXuZZVhuGWvgpzgRj3kgN0sscQoCfRWkKO7x8QGDupoTJu/YdwIySyJARasHGuUpyF7f5CdHSpyxqBezY/RjrET+wCvS9I3HXFzJPyTD6MVYJW4IbRKwZDVImzs8k/Hha5MDNR7WaUJb3+bSjcZqgcGTBEIj7Xlp+x9r4KoBHZS54PNN26woNYRvSZT+TANWl26naNMzBCBQQGGnvTrdiIyABxkpFvaQtHZzhkaY5Tv+s47e0BxlPs4BjDhyYmNJsCQlDbYzaW7Bsd3khJBewiKdqYU/a42CAnDSvvTU3d5wCv25RMmS9lVV1cYY40++TxU9uIG5HjeqNs7IkgcLdnXHrab2xmPT5ahEcIszLadMtcbHAjtcTlJFG4nq+E0uL7x4c1t+kMYZupdsY8zj+EcfLNOiUMWsfDW93C3ZceXF7mQXUqR/7UfyVyMCXhP+3kulqg2O9ZhRpOo4Zn942a5WzyL/7rH7utgfB9NPJeRhHHANCzNk/oM+V402WhJjkbakHpcUMOoKPxRTzN9EWkAwWW0YLyB10ua83FWYVBnF2IGtySYCd8bVHf4ZSCsjf3RJ8poUHfly0Ke3l9oGgB4RVkL+icoeawSxkSM4OYAihs0lDCRI3PUhFepwntOKGmDnqx7qIBuWU+6CDHTSLBGpdAJniXneW6TIEe6A+R1lfhh/y9o10JXi76XcuFJ8kchcSsFllln+e7VqzOoVyIVox1G4saothiTgUM95rOZJWzTrTCf44xnpQGO2rGtF1mzCiRYFyet/1YYWWSDOQiEma61wJTA2HbrhwA50FwdgqNRVDtVzYL+UtXzGZ9a+fWSuw4Al/82y/S+TVQkc2m6y+zenlJsFfoU4jxRSAIcfY27soZB8k8glqhL5zmLBwmjg3b9/852mg/8d+7VWQh2DbqfLJeWQZudrVH0FMex48mx1Ibc+UEEZUg5JwspKkEOWkqvdUVsI5P0OCklOG75lzh2IoPL8rdNmDgtVfx5x7KDq5HUfZMFSrwTYhbZcKzmU10EjJQoMgfX/GcfKpZ1m2Osq0r7NrjefVpIJf8r3OlwT27+dQdg+jagTiLmvqUN3plzRn5ON+CWYRGQoo4A1L7PbcXjOI85zfUzSn26H7VSOCKKSl9sW99ATjpdMK1aoaZVBLy0aBzPAKRwVFpZLQi/SC8iqHmD+WEXRYjYfs2zOGgecA8DrAW8of35q65zdYUreN840uA1CQDnbB275hTbV35hPVuJR4IxN5V9hQ+XaIBXbpmjTl23AYiq9BDHVEGG3LldxMR6nqIAO/0tH/URHdNIhjxe4s+3ve/xBuI4obLCv6YszU/KHfMy8EB4+ABzlkResPlPnE6B9kELT0oacWRNhDHPDKTLB4ujFHyswDehbF4goB8JXZei6cqgfRbVYXIOUhrvWJW6sr0rhCTBdc79rTFHDPbxP+L7x6tSEuxXGcexWO3K6It/tCoAFfEzfGl3Pq+Ud1uX4GLzbjTvd8I8d75grNHcmUqsTBpOE2G2igg0PMMtAuE9LJiRZaqe3HU+zrO+5tGfxpuweKnbYwQMpTa4/Nd7bz5WYRIYEDWoeDkWo9RGlxfWcz+FTm7Wb6CI63+M4i6S5PwkqeK86NIYnObO1HGCLZ82EL3TCgkb37ajQ+fzUHGTEgYDxMK26zkNmS/qWiVUJ5OMbNuIXSgV2vo4OQtG+/tCvdipWpFxGutcrUlhtKJ+9Y7eS8Nzv+WXT9eXzGnzgmWk1iOhZDHutXPA1RQ4lXeyRnPv0/EiXHAAQdGMr8VZG4ZY4cqODBiNdXnrBbxXOCqR2eaf8BQ6Gzg+wUI6b2qYUNzgFM7onaeHTzGgr3284NsApxoL7LZFutPz+4a5W82g6cl29cLXNatSZPO49qRKkyz6Vx055vRMoa63ZcpeXDHYWaeEMkYkZZ34ZPGVECE+B8gqWIqKNpLUiq0TcHTQ9V9TqiNwL+pBK1lYtEyOl6xcUzXRPwdhEvP/3hGIZNZfHmCUjIwFBLO+Y5Jm3IRg2W+kRYhFqyjeEQYr1oXJb9e91P3EQkM5+iW6szr/1X1zvYRMIt9mcet5CKnC0p4KAkLBBxMCupKd2AiziMKx+W/ndFXZQyOczNNJgiEOI7jZChyQRc4+/nyNlf1daNe52FSiKsE27j/qjG276c7mlD3k7t/hRHSjD2776rJoRRTaJ74IOTpfSxcfLSl+oA+CB19SqI78UBMJclEdyJ+IVkN9X1krpLkaRA88XPkb8tiW2Md4lLl5AQnevegTvpTYCKK/2+DW7PQpb7lcILLcq0tPsTsPfAMbvXb1KJkLPXWEDXMlIo6Sy62KKyYixyFqcurhQUlJVCqLVK70L3mTkDXmwVHi33iKMzVLJcfILimSZaAbhyTjSuaBgpcbSIl+rLidrTBhDYJCZdjuVkcOox/S2zL/oNxl69ylLs6t2N4xa8PtQAbJVOcWFmREC7jH+b7TZk+OCr9XhVTmwc0Cj7M1Ec2jtcUzy61asytAx43a1X8vmRubCXXMYe99x9wLTIXSBfobn+CKJANI9lyXx11FrOq+ObW6GldH4cdoEDzmosOX3KsGj9rXrXCJJLXhsm7fPSMMaEIFO4MfZ128mjncJ2tUP1OVNuaMhmCJ5EWpqaYFkvDg/nUGWOpaTWBPx0A66I4JP9xl0FJC0upcSxb3uulGNin7I3bOr88eYPwUi4SUF5TaWSLBnm5qidecZt+eVljzPsM98RS3tKCvWve59TEW/iuaQo6IyyF3PPHBgcawVSki/3XO4FWLl+/d5tmjhu0mozCippEr17lHGzBn44jnaQEKg1fazipioxdTU9bowN8hGEzU+2/k6jw1mxYafD4BbrXJgwNVguTjxsIpFCTgvCILrt5+Krd0GnwSe/qMGVeMGWzqzLu/xV3Wbb4aLC6psrNFBHSx/ci5ka55xE8+cjuIM2E0jH40y9Z5qbgphup5kowEFCCoIMNkjfea/BoR9RVBpNRZak4q1i9hzoqAfh9LWyZZA1JgAVchDOmc4MRSVnt3+3nu2qZkoRIQ+lAeDbeMmyRyy2WjEfGeUlT6IPfNxX58NLZRnXBYXXPuMfghCddpBf9ayUKTHmlWm43/Nsn7DwGOAEFab7Lpn36st+QHSnhay3T6WOiF2zBsra+Y+sfa1WOfwruZm/zVUZC7QKk8BkxYoTZ0eS8tW7lQTiFojd9C/Hw1kyAjQC2wa4I8RDIbAh/4zzUvN8EheN+FFg9yQ1AwFeVzoIkBuhhLnp1MH5CzQdO4MxpTsYA0cV3WOAcUaIdZ/OW6mxolv98lLNH61RDN4TQAn7/sSkZt4WiCSI8HTv3q7mIRmHyHC61sx8wbhrG0AE1ihzFF9eBqaBwe+eJ98oCjgoL3B5q7Z/Kvw6zQS+PUExbdkBEg2Qx6HVwYmmrCIZ+j3Q2fT3MooL3P9YKGqUd5xQGw6diYRlvtdhxROHdCiTkqJIoeHdHWdcostzoicGFiyKTx74WnHhLW7vqnECsyl2ZTYAfqnTMzNrXIfGYNz+AWn1noWoNNGcZJJ6K6fd5ZIvqle0EjK94toFisJHfu1GxxKaaGZV1gAyIFdoPtdXMZcjHeLUMJW5sFVdxLyyBJPHrxMRolP1qNc54+4Yef/25W29hU4QnDVOJxFhvbF2pgPWQcouBjW4OugH+i2JDb5OmusKBeQqW3kviM32Ovj5c9FptjcG5xrIcbyk1poeb53cCpcN6h4+qT6v5KVCiUhZZ1wYvX2+tM3uJ3T5HGCOGNlj3bNBa0ZB71pK/kYe+fBgOFfYMpYIObrGzO/0TCqp26bimsYM9NJ179DeebGjUmixHXb/mMAZx6A+YtvQMDM3vktPXmkYod1UEls0mUV0qQvyPTgPaU5yaCjBKDkeRjx++7lxSpsdJNrtan8LL5d0p2G1SgcJZLE6ZQYw/D1w3mMoEW9z9RF+jbVj+XL6dfodvhtkuhkwpNVvxBR0FeQGHsCdC35zpQ64uF3wO+pIGL4VPDDJsLPpVZcYjobmYj+3WybB9kAJuopaRg9g2o4vTg4s4LoHcyNG2Dy1m864hDLkgT4wYKX3FFHgEz9NXEgcYphksUD4OULT7ijuMLJy3GtCol7kHpZnitXA632KpxQlRy2sB3hY/E6hGahZ8K+XKMapvMPrJS2OevmOSCyhDz+SiylYH74H5Rwej7Sy6wI78NcnZxYYhFwS8E4MITXNFSb0L4AF2lGm4QkwVEi+/Ajqu4noR4vHhiJtg+SwG4dY1VU2CDXoB2NRRDC0oxHmKmfOSkmr/oKy7J1J0uATDx8ZnkiOKQrjM9S/6WM0x82faQzvXqX0myeutaIImtcRdClbzA9PkwD+JSqIhLGAxCaBjLH9ya5mldls6ymRBJQFFBSNcLv9d3eeejoh93F/4blQWDPmMhV2n8Pw5e6ArelsYsKpOQcgmRVsSULpb+/Eu9YkJfv10EhfokzuRuMk4N7eCXVdhUbg651xHMbBtjXen5g53zlIq05NTjCxjTCpHfsBfyX1l1gR8XSZMnJuFWF+xIdUKVRGx7O+KCehqehtBhCgXoOeRMOQZ78R2OBReYhqtjQykviVtlx21mT8wUOCnLs3p6yWD2pEDJRMYUou2/vZe48Ny0KGxogz+UThUhsFty2hMU/Gkh5+98S1vTcalNoH1q/vFm1K6RFUDmGUBf1XN/Y90HLzw7kygIcatGt/ciwCwjerSYg7CQw9NU/qSFftQoOA+vKwHgFqzUd6QYl9CXDnX6o/6C18d2SDmc2+rbViTalrUTu3hD9i2W7QzbpDHCVvlMoHa6VPKSbyJSKr4lVd2xBKs2mtMwXu4wHoSIXv4b2hlAYPmR2VXcrLFfkdXUGTG+ohfRgxn9Jptq6ciSHL3py2VPX75hslnEeBL7NULNsiAd3s0eoK/Kkt4vd+BpGLtwLBFJri4HpiGwHYL1i11YcZ/tQvv6SNZHjQ04sBo4brF1qKyuCjs01Y1y+S72Xa391ioUYXHevZVZfcoxjFnnOvkRrVsIiJwOUeIOnqMnMr0rC63TyWJUriJwO7RAbvrYRGh0LlBsAGYz0CFMgtN1pBbSx0Y1WWdUj4UXwcsP/xWaR6lGI2cARK4YWIr+vnJ6VqVvB889yxIgwN3riWYKYThq5+gmX4ZuklPlgCfpWXhmXOtzAOzsQTCpdfZ8dq7PgwP7dbAzHScItLB4VhItMMAxKM0AzYF86rSrBC7UHU+FE/SHVWUdq1oTBpZ6SJXH8XdOYfS0qR+cSHVrvPKnRjm19em1wSrI0bEWrwUpvMLt1/IMVqM+9P+lvta9nMTZaVC/n5HLjbmv+g2uDQ0MoqHKm/7LHx9Ui2SvD0XkvpAvHgFlj+zO8psCfV9Qe3dV8Xm/qfai9O9sqbxVmBRsN0Egc8UIK6dF/tpmz/SYKzNN9i9Ws6fNmH/PlMi0qZtc8LBQYkJIhrkC23QmJz+vJ8UB8gBxN0dMDPx4yS1Klh0kUjAbeLFLR1HrJqPQklwGH2ksIqMje/SNNGrkmqqt85QHG9GwpFdIBXfxvPvplVrjjAkGfg34Y8bFqPgiZ6HvX/mWsvEQehZaeLDYRsADKejzv5dyv2AjOhSdVn+2Hq2/oSS91a8pXytrZoEgp1a1y9TQdkbEOL5J5sMTuxbCBb4zuU7Q0LguPu4a51E5yD+lTMbRtWZSHnUfa1DM2INks/TlR1QRqn8m2ZqnVlxSMCHLRCTdRX29l6o+6fZd41GF1ig9QKytYvxaDVONHjwLmvUh7KhrJhCQsYqgJpNP9fRUfsxisfIAVS6yg6+Luq/JRRLyMI7JNtUa3YDXRrPM4QruhoacV4wbWUGjpmuHnr9HvaWy0HLCb+VRSHKi8C+04Y6ioBcJyzCrpNFg1cAIQtXzep0z8WJ6a6m1dqKWzCjzqB3Iy/t2Jyy2VHI0LA/cSufvM+0hv4T7JCZp8+EBbMDwMpLTQqk2D6eNlq+DjX5Hc0vf0ggmQm6tKmwXtoFm9jOgN0MBxlCSmZTHaHwhauVYWbzC8NNot4A6Y63Z/gMIgO0hGLNSoOvcvye0NBGFP/CuJrIu9ylugAmUq0U+f12cQXEpuZMStW0J5KAfC88qvNcJ39/BwuEvEh2B65i5WvaBfv+rm5gkiXVS6JJtTyLmDuovvnazaMX0qiLqvkpQSOnNK6/r0zN/98XxUbfQHLXLJ05YUojtYX2o1aLBsBgptvGcJlKPRcVGw3Ob8XF1hDfrM858PlHnKBZp1ugoEgSWpDO4E0R6TjXFfrDaZIOlDt4JIAKRH8FOAWjB9J22KZaRWSnFja6+OX/bI3Y0mcdzWkxIJh0/DnjJO8q1qvZQzedMAR18OCgRYDXkPwa4agaTzbAgMtsRJUDGe6UcmQ4w3TAyy7wG9wlIdKZXB5/2c2CoeEpN1fsf+pdfUA62fKdF8ABkoUse1m+AMmNQLeEYu8u2nwq2nJLiiuixHVz2K4HgfvHIKSHKp85CA1FWvz7bDahyFuLsVqjb8edRGJ3NM2kVuaYP/1hBmkCRC53b9OqKtbcrMZ5c0BY9rqVb4dbBYGLydqoEkHMaM11fscof374rnurHPRstv43Y/rGafgY7W+2ilasHsXziZPlZBOzQ9OdbzqXKV/qKR7q17m/DKYXEbbXebNf+qgjEeK2u9t4jEw8+NpU/LIKhCDC7UnUk2UcF1/MtRL93kc5pquXKwHi9ytDVFE5CWVlmeFmOdR30wkseN6sEeWBrWV/PlemK3qT2Q8pi2XToGTm2LyKG16J3R8Xfe35oRhmeoSaUrQkCbPFhNQf0B27DHcyACw2LBsS4BKfAtOKKkC5tKO8uXPSAosw8+bNcJln2HAgjgrQkHOa7dscg3uNGmUn9N9ilY5d6mA+j/8oxSwZRC2kqTa5pLXEJ1cSeQyKyAlfTUVFvTqDC36N6LNp/pPYvWYGh97O1YdKcuwjmz0x708FnIoGaaCPLLCUxhM+s+bOH3QgJxoLCTgmKuQE8mTlBy3y6D7VtgbI8N5u9fd7Sp1k/2lme8Vc/0ur5m2EWW1PNbF+tURXnlTBpUHlPFcvyjs5/iht1lPHXOvAMhVAHCkkeTw929FJs8/b/mjTvZDMNleE2p2guAURHOR1RWDXnjmCxYkBER0LJHrZqAkN0h9iI+QL9fPiCLQecAcwnDDuXZI64NZkxCO3LHg5/bzF6mg6uKyigwXZtJAkDc+bh2sn6ZHpfnaezmbCnDdu5DzKBJ4rfZFfF/cgO33dr7fX6pGwqqy0PiT9s4Kc/Xlnc//Fi1W63XOjiiIRIVaNfiPn6wXuHJ95/KtcNKmdaQuWmakUYwYyIE1Hx2VpLoCHWAoxnD6qbYimeGLikkXUD+Ujenm/QEsX9D3G20sX9XRiNz6xydgpFhJzK6y5if0vvTBVmd3m1ts3S/i7sXytkqDzAyBvl2efFbEEmx/FnQogLV1lXCRfGYWL/5VqhCPkkn8usIncmYzk6nFDzhWxdJm7fHFWM8tnanKeTZw2ykJn14lL6OsZC/28Dy+vYInPffpLUCsHRGfz++gix3WXI0lHsoPH/qp/BI9TNUVseyuW1P9iT0h2o1Fc3MzzWOGgxVnA3o0fnd2Os65PG/ArMn3hIAgvqFv465zT0+x+tPd275Pjhv49AocYYcP751vzOX6SA9adgfkvmA7h5v2fbjv0H8K3tZwdtXjyGOWRouJHCSh2Jzv/5qq6fhow3ee5dFhblCwBAl3qO9SiH68NjHOV90W4MT8X6bmhKxMm2SQ3Wr3MVQL+VGc8D8n2+nrnP0ysfzytl5dPNsQee7056U1xzCgGYGRP72fFfAGzV0XbyPIEI90kVOt8cwJaOrQXWFbajyvGpyVLRHbiTH8skUAjJU/SpytA73Rm9gPmrbRnog/iw0OWKx/137Z/jVxqR+NsSSsCeDifJfGRNv3/NLOnOVlO0MkaG9UCtZQz4mKznTa417vybDUL1+51hZZiCOPBi8f3qrBS+fsO0NflWZPKr+WYHvVbC94uNEkatAzFglIwOBd7iinz0KiEmRM7noGCbCbq7mYUVgiaQz/Y/5oqd8uTYAP81946jqWjyA1ZcoXExJGcl9CB3ffqFTVYqE2Z9t8AcBIIMY1YZ8wSKUOHG9FhYygpQp4QmW1/Z6994bzP0JEVbw0Z3KweaEwxxJ0EGzF+6fNPQxBYYyZO4LQ2Ze3C4/VQGlX0dPToekh6HQ4oN/D7xElPa8nRgNAqXAMYH2piuCmy41zAl5ND9aecwlf1e1nzzlr+4Xn/L8hTwfwhtacYrNnPdidycCSoCVFOyt3liDIAHHrQgzo1dd6ac3Ia0VMEldYhbnyDwOGNixUJsFzYZALOLLpjzAsLhB66uCeuHK/6ihNObUL5Qf38ekoBkkZEKS6So6YePqg6g6TZqATsfriLQmFo3w4E71opCHcL53jiOulNtnLqdnuqg5uVNUacXEExR5TdW2t4U1vMUSVUfzSPnvMubBV3ARU3cH88nS2NtVKhXpnK2mYw/IjZ+ocIei3FuCkesPFnB42g/3ar+YnhKi2W1Zv9E9/h3CndDO+gDgp1naQq2wapotxYeeV3Ovou1PeHrnwPI/2R/hpyQ/KEXP3USJno6KnWKpFUvLaUmrh42Ta2NEN30IgU8j66SrWDZhq30PfhXnHOER2ZfX4LPr7CqDs2M00+Zecf+/lFok0VIbmRi1IshEVe1+LKXEucfTh5pPUIZ5qT4Rnclp2Jvwt3XwawmrfaAu4m7AqqwfycQ5ZrDxT/+/tQdaAi69QbYeRTO5aHaJ0tHcmFBzMYEnc1mGxrrYmD8PeRkU1DnZq7wODnb+Vfp1MI7IyvfjgHEvdduyx05cGJBTCok7aTbIClsre6QvfcjNBLubTzRayFWB0mv7/7kOq0728ZnroDliup6D3vy7lVR1S+93vHfUqCQYm5RXc3hwZjkfZoHqvULZSHDUJxrYEW6NRXDoXFVAXe5gU56KJlKUOU3AAQfWISMeanJulE/5Wys6thpa2sR6KUOFCmVSTb+4Sy5PAwXIAapiC/K2ENpdnt2NK/XI7oGvsbnjg0+T+IJQ1ds+jNYyWC3QxS4ka3ZbrR984VpaiolqXbYA0pbRT0Z3lc+uQhaz93DBqt6orFPFyjRYHcQoMN7XGNgLs1BDUVs140lpGFZsqrx3u9owRzT3yUsLAg18SkXKn63Yt0a5IaL3USH7tuODrmJ/hvPumsiJTIySJyzvTlp1gNznwy7CA7rSov2n9HzrF1JBecKerCmf1mgN3ppA906/unwEotSTvh/2sWIFdICrowvN7IhlMOuYR0VdH0XTZMBkY8Io2Q8Xq9tg54g++RlNiIsAjg7EN5rvb5lV0h3ZrIj685HlbGaVVWvuzJX3tSaQFb5sO6o6on1W0cYNjrmm5FGi6yce9XFxKVa/AIRbGVVr/CxTTY/ioyfvRZkqt3mQE3/CluaqAWL9g/Q5xu0K9xlINL/cLsgIDidipO6NcCtsEiCoax65qlr0Y65Om6WYtzaoERsABjVcowu6warLjDnAJc1ZUsUYHSqnAyaJXmKYSoBRwBfRrmd3QJKTL9q8/mdbYxIv/VcJIauLIcn2TGXfBSfi/ylZM0gimJyeXqDm5I49tXk4Muy1s4b/8ihX49davDkk+AWIVijloSRaWFrNlf4nFFEoemlh61qVyZ4KGX8rBLLG0Z5H+ruH6BhVqFenm9H9yW6swe4uPJvg8o75Q4gt9ICn1K7HAtmOCIlY/q44p72TEeF5bjqezHNShlkICfktPKg5CLwvPk74iAJRzmNTan2HRMTHxjMTCo1Pvcok4QZXxLEeUUBIALVc8641oN/fqIMrZQhwggyZ+rPjf3BdD4CfS32jOShrrU+Jqux4rMGz67oy6+xvT0DeThBy00RaHv+ufs13vjGKcagC9V52Q2beBvyhn+5ZU6nBUoy6X7H8isXrSsBV2NEuxGc+/SFrViMkH++B60I68sLbRZIDqgUtCYXR4PYSt1qcy3Ow+QI1OEwmpEMy5oyft8Zs5dQb7hoLzEXgHmd0cMv7MWO0/GO+K130f0DePDtiuSPS37RSmpZPwOJDXQXQWKBGGQgYYDOFK8sk9Zh0EdanPjhkyEryXEwNC87LznaopDPsuAUZqfL1MiTm6pMbWzNM4uw1GqCeTP609vqBFRSGUrjx5Q8gXo7s+LS/Fe8UeJvEU7u8iDcrh+GLaW7oleEiP3m1X6pEQNxEJn+z9zKpq87S2eBnK5e3idyC7aEgdkOTggbmJdCzlFZxzKI+YvUO7JrWV3RekdZjJcd/jRqya1VRwi9urQDSb+R8VdWJG6QlOZkoMCROYCnhS51kHkauzRPVOg5ftmpa9oZG+LtVhQMQavf87hqagLaRMPuwqfIcs8uYd29xk0xybqXHX0QGp7LHosMJ+XmEVAd7yJdpU4BjueoFkl2VUeQ8ofussLmHEFpln3wY4sEj4Ju4VHWPtfPpIgJNzFKIEir/vrU7d/JQ4I0O6u7Zk6oSAdkYJH/2BpY+E7LPGpz8wP1wP7gJ2xiME3S1pwTuad71Cv3uZsrLsnf6gFi8tWs1ZCvOWrm7Yc9nK4rehozg0yK7X7TDDvpOk3xX1w1+N27kKUIAle/tB4TNA82n42MuW8l8QkxBxbgsVB02MMmg02wa1USwCVOoEHh2Gyi1iHT2NPx6XrBbDmPiCpsHqqeSbBsz9LlmLCqEwIprWwyQQXkn7RRKsSQOxzJFc9zKWt7m8zmJAyovQcR9JtrYFw4cWP3DKS4l855aHMq5NqDz3poY96bjljrOw1NN9dgy7uc/EVFIWswtSRQz5rFrxdILRoXbmcMM6dzITyd2z+vurvWdM+H7LkQww3khebDXEqvS2FqNzNBRmYeOHj5/TRDnYpeCWwBC0IaNPpIqEcl05Dv8JuYtx3WmwCL0rjCY7vtz0VFDsPdPX0BsPr4nYaxOdui0lp6j5Rzf6GxbghDfu5oFKjx+QuuAKsO/68oOBOYepSZxa2Y4XIxwwxEHHC/03Gm2QjtHwG6ePWOzJdwsMy5NcpVMQo8KafPcMgqgLH2TAhUrh2nSgZ+5iFqAr+PrZqg6qdw1/qUpYL8DXXQuHsXiytyPu1IZjGBvWTVroLr6HCjFmgWm8mOYn3NNRhuKITdkdCt6MocFsYxnnqYTGO9tj8jp7w+40OXW11URvd4Wz0sOIO334++lV3FP00tW8jzD6m5K6kmuFCSQwTDmN36jmyIL7e5DJRXGlieh25TmKIWt+Yqop6GllnvHebisVOIeN1t+DLv9yYm11nUJiZKw4AE3wh//8XqA/6NwXKSnVHT/cW21ohtU44Cx+IzLwEcuZ59JOS8qBcGA8Fgqym5wElAWFKSneb8CBi9EJjx71c8Y8cTqgSYhGFlYV9fFAfAHnLYXKgLUKU0UnFKcaHS0Xs2RT8SzoqG1vFgQ0mkZs5AGSWtCn5685Mf6QPPV3mGPd+SKc9Uf2NuKjd261tv0wKc2h4B6cvpQBlgQYbHqVUIuUcoiI/2XT8epr8fe2gaKtJZwPIcUDTfvEGmsYLsr5iQfSUHKlk78nGW8nVtRS01H8rQ3/zsyCwNG8VdeIgFN0vP4GVnlJbiQtcA0Rz81AqB5KYVQKPoDfTENVNRMgNZbRirqt1neFuHcSbfK0ee5vZefP4OQXPmirPlwZjpDZNZkADtvZmo9YvJzC5FlmuLOe/iI2kMJMTnIKqtd/E5wMWgbWn2GQyyCqnygaA3P4l4lGhDP4Qb3YcHMawnzYn06LtAe+NNr/4sEaDTqSdsqku+kIItAn82AkwUjM5PfmZf1/+tmMUdlGYC6HQxMwCX56TSWPpqtb4WIydNYDzjCyquU1rb3oWcl+rGhrD8/M5XWRr/ZBfbCVGNydxw83ehD9V4O3VARzKeVl0VL+qqUVlN1I/qFQMAQ/HGaB+0bHCbcmwu14z6oVsv9ZUnsp471qFfj1snoo6VA2gCFo2JODCA7PRA1VA7e2K9h7do6KeoKp23cM0pqHNoGXqyLMzQlXIHYnan0bbOJaL+4FmbEI2RRNRZ7SYTvCuViUuzORbl4x/NnirCXiuW4qzHXH3V81kEcuF4siIcaovE2ttBHG9HMWtKOaFg1196+I48euvybUmuvKwFbrVwckZfX6Sy2f+vBpmkr8J0iHGXSLpIYTXXiHY68G59XiYRmDtLJZjwjtxO4YRVDNmsfwf0aKDJL6RQW1rpRkrro7zaAgJLb9V817kvTDsK2U73tZ7RrPbazcWtjEzWPP/Y1ubjbTFy0qg8vx6IEagymxWckiJ0R/b/uNSOb9r9hNShWfILZrbT8BuYfgo6yL6mDp4dxXIETrJewuemaa5ECgyMeCR7LaWLMAXVTvQ9aF++2ymchVZ1eGAMhUn1SldIAV1Qdg9leP/RtNP9wNjNDpL7mqTKYpFYROE881sn+MXbQEdpQKBNZNC64f28N96plVJZAxIGOyNIwOeeMUhlAaESiHKDmaICB0g5xHW+76BppXHDGR6LubHVGxipJKa4FazCiBKASDOYJzS6ifEWaD63YsaK0UeTbUCZ/p8gdcWoNfQ9al8cx9uv43Zg/lRKq4+Kzci/wpUOBeCAg+y9G4wxAJaoSuooH0VuBGMR71gS9kawrSMMwlzp6hEsg3WVV0UZ0hK+YAEqXXCitKkzZUkVzam2pNLAq5tP5vIsjU8P+4RGUXqDH4IQ9lz3IzWu7zi0Vc/wnOv2Z8wljN8XzXUSexIpscLFaM5OqU4nnJCJrnLOjTIcyhaib6+moTPniV08kRo6aWZOq7OBoMuZKRKN3DqAymc6nHY6Rgb5RYeIMSKp1yhAAVrjmrnjx9llkWdPUgTcxFJ5ciG4Kl3nYzpu2V8Xko6cdvgr0PhDsd8gCsKuSLzPd6SLYjEM4/5g212ly2f1UIx5CmWJqB54iqHYpfA2HXc1BtzMiP9zCfJwjJ6xenY1vzkJGGZ7EPN1GK4z/DsbSK9JMr3Ba7YeXO+Omx1y8j5gZzY+QLU1Z9pI3uDZWYv48jvYAqBPd3rU1HCZipRyDaQdjX23fvNkV09hywkJcY6El6KfXFU73V5CIgmmSY9qJt3b0W8bqg6pDOqm0vqW8O7MnYL3Upxfn7O3U3QxLV8bqqnhrXbv7aaHDp2y8Vde6AjhuvcBwwGcdlwnxDcGgnwNuhE/WgkUmN9Q9IcISX2TJQJA5p/4CZupGfDPJt24WX7QBir5Ne/wM+dUzWrE3hNS4FblyGWF0GQUuztVWZtApkMuvY6uL8fNrSs8crfxWFGjeznVHxgZFwxcEJ9JzvMH+53Lb8xMTfx85KS2fdXXKtO/2cVb7QIP7M8Ruil0PsqaCbfjTTRnF/cpKXHFVrG3PcCKmCLDh7+mX3KTdh8UDNSmeWayoiw2y1DIjZyI3aLJJePGD+g7ZVg/QnHiogLy+KqI6AC9s+LRE0dsOtajWdp4PB5PWq0si004xs6tE234QKq1w8g5FJY86jEkJ9JYR0VG3gRZ9GlX9O4lyqj56DxSeoDX6Fs94c3gsgRF+VYOY+NZPe60XY8UtRAskbMsMtt0l2CTvQSBdZ335MDR/T5jFUWXUHhra3mA3T7KBhUE+yZojX3DtZdI1ck1x9myjTz4CYomGJpETHZAC6vefS8Attuj9BBjcqClifeXa0urpvIRwTITWvBv5ECC6chiczJ8nNtPUihX1Bc0xMf0Xgmq5M6HYFDibEtg8i6X2jJ2IsKE4O3Tyj4XXGTUem2UYdg0Pw8VvSoyhhMjf0yD2GVx3ZbUF7m3nB+NPyDd0AM8QaCCWokWl9h+LbUKRul7YU40dhRdYuCG3qrCX0LudO1wh87c5jH+zgXJWZ3BSd6tL9LcD+p+tnN8HWaVRqEIPP+JnbJhr56vOTQOjdrTg2PSd/R+E0RGI6+QJGIP1ZLIhGo0wGPMixxuYToYGEjXX+Hq/OUBNK2UzIPv15UmjSsO6dv5mrXETFJ9rQzyGLSKA+NOG8Sv3GY4o6E3Otoadh8FcXeRsGWmMXUVyBdhiz8JXDsZLTqVkeqv6Hpolh293fbM5gpVObaGOb5BZ/QIX2aJOASwEVq7HdGiXnUtKHcIHF/FOlqHI/97or+H2VF2vfoKs+bRvKWLx36GiMMkgmHHlKNSPExuDEo0RNOUPKc8fXuXsNEIINp0AuSfMKa0L2huNIXcVm2/soyQjfnjURvBzcTNKO0Tso1oVmGeu73P7tUau6nyTcJEx4m3YDEfJWy0aW63O6TUE6PcfgO8R8rAJV38PMBzHoFAItt5+6540ArILmYa2NiVWlJEvJ+PBIi1XgPlRoWBiIIRAAITo1SLBtL+AaM9NrNYsNBEtV5aUuA9LszEZOVjq77jHVh9F+2VMFntwDkbDhpmeG8TVcfiaIH/Qhrty64uQPSSEm8/jtrUid4DB9DUwmtDdAOfEyydBhI5/y2i5TGo7Akftby2aCwykygc89RTE36UZ3F2qm7eFBtZH9Ng2z02DzgEkIXlOgQNfu2xedo7IS1IczVRP3Z9xAup3muBV68W9QogdyeZ/gUdku6J1aaFrewcNM7Ieygxuh1R3v88bshnZz0K4kxN2mZVoO1BF6jzhmXIaUapuFVcsmXGwcCuyN9xepF52p0kslzUAeN7MPF49Jxnm6ixH0u1KsC4t5DgNoMox/YRyNnEf49KAzXP8RVW7vwF6TQ6MEXTXJGYG9Y6jQCO7UE6vuyBKzaFzGfEKY4jbt4b3FtT+wJssRsqzbZ0XoDLCCGTuqVV8QdSa3PmCRh9jmLqJ0QVJiqNV0iRrgRu7TMVTPC0zevy8BZePT+HYuMzNkQN9ySKEH0M/WjhKM7/5YmP6OSxtNHU+VM3J7VtqHpyisAbOpukYdwNpciUJYm/a1afLeMjU9clCmxk+E0vnbYfxNb8cc06T3LwcnIHBWLtSIXFw1l/o9/70508OycNXNMGnkSf+hq5R0Dbka0iJjU/LO3FSYm38wklYIpNPp02Ne6fTRLBF63rxTy3uasA/iOT96xXrbNLw1ZZDVmZzScAoCdvlpMEujIhlGjQW5M4rlV+diL0qXHfX9BHIkLcRZauWd+wCB49zIvw4y6tZj/+WjfumkKN65rLKEwR4Q7WK4ed0vmBVcTVnrNUg8wff65R63eTjyEiK5CFiAgz70GPU62o0jzuKYdTRa2Bk7zJcans6aTSmOlwJmQDIe7Ftwqm2wo+Er8xbeKwhJV2NSzSCbkY6dAvMK2qUCI2oxB8r1e1M4bmAp7uZb7SrwRPiwAy3bSVAAOzBTOi0we1obi3BSPmYIEwB6u9zN3QQjPLuObcG1fRCCrcEDHTLUgBVQFK5ZafngTSWufh8tmspGW+Mx1DhoCoyD5XUz4+kQueL8hRvtHuoxFU3rbd2vGlFKUoC/PG89y9IS7Z0AFQczb5vo6qFzhNFQyjPYNl+40fprFc217pIUtooKf6Y1HSxzcFhh/Nm8lrI7FaeduubctqtV0C2xh187XKCVHsb4PkiWgWVdeGMwMboXUy2j01MscwTuVjUbHABa0c1puCew1G8ZOq1hK1BshZxcFUB2eDZsdvGmxDRrTNk7gdzOzuKsvvdI8qrg7oXOo5mmCh3bIMUrpTq77ORJhaUeKHM9Cw7RvzZOB+2+Rv1jV9EQ37/Fkb3kGo0J4Z8xXiDt2T4/Bg5MFzvti8WUaM3qqhUnsd64pZGj32ir//ruD18lvrCFntCDwijNoBsvnr3IdW6Nl8XiP+pH+nwIPD/3Mtfy2ITh3xzSG02FyGqajcqwptJblqjmVfnAeqqv0X6gMBIksbczwV8KFzwOpLtNks8VTIrRJOgPliqNOvXW73azm0R+naxcO0BX+tpFcK4vsIu3uNHx5pGumu58N/4f2ahkEzx0rOjZsIUvSVytQOMTBrxT/DnBVzakNyqdlZKmogE+fJvsCGZDieM5INv4oCnnQZxNgadxbklLsJS3Z+yLKjN1H0djvBu7+VGLZ43bgTgKl7L9O44NXS15ETRqXRCUf8Zx7O5Du+12QqgfebnvNzjhqk6y0m1WYT73bmSnZL4k39HFIIuoOl1fmuemEM/YM6jGqq0UNZNUloo+s4mvIabpGnQe3irVwPwOjzrIeWH7nB+Rl4WMEY1xc8lwNAcc8clKpo/bpUgedxyTzecHZtj9uVvE7Qgek7aUTyW5UIG49eCuU9oB8wsxs5G0fx9XF4vgZF4wBDYBfP93IT/U39bVCMJuR1pCUhlgT86XZ+xWHpLckUBTY/iIFDXgVwkCyJerx1CCZ4z3wVqhnLxOkTqOiYZZ/m7kkuFAGTtSqJGcswb+LIBKnFWNL23P4Xo296Z/YxOTYRCVquTPAUnQ8/porXZWHBFznQz6x0VyKRmaQFEjrVo+2fWtMQghU+0dHr5P85F/2I60/PVW3CAqR/d1moL7IBOs05u2134K4wgQCWQFin/HrUhSW5GXgvewaWJFhkO7Ocb5fUvsO2+J2za3fLG4Rl6v7Gu/W0L7grd/jTgpnv2YVNDtDqFqo7tD4vynMHMFrE1NVtGV6P4HJZlz1auVf0QVp3RkGt56vR9iVawwSXeXEeCDunc4rMAdcfWFqWcTFD+4r6rzezBqBPEXcVAvNSceE0wDzBEFYSeis1jKotZtQogphW9BYh7UvqlCudaUIlKtYcRZwFVNuOOj85y48V++v7njrTmyEqyCtT8nXCZxxBUp+Mgx4sRTkdpgB4hgmaCivK6dzuS+RakgApJZ0H4qKtstleDUkWOQiygDDYC/5LSi+vMYRUUa0LstaWrAhGxU1juHO4/di/LUh3NfdfPGYW2ZcoML6xpu+v9R4/Or38eOso+VqObzmshaEuzpVFdxHupvE3rXLrHTWlpqTEqgZIW+Mh4UPVnVWUNwlXufzOHd0TPEQ9gsOkC5u2+lnPqsGCtQOy6dR1/iLABUazrPCVW48emmId2xAUXkLwkGQ2A9sCgRxLNHKl5Q5KFNB0o0o1W+JNASjcasLLdzkbxXKfdeBVGNvZBst73c++OWHPYfs2k4KAZ1fluLnidlTnl+HXcs5cGFByEn4Kn7KNwnDttzTQGp38rBjPUtcLJf2sWxJ/wPAc/vCpUtTsiNiXdwrs2iO1A0jZL+bxm1N1n7k6owu3bZwCfh2aTg6SL80Gyl6//YaLRdMaClj7poTquBr4ic1Q1y2/pXR/wKhr1edAU4+m9sUkzixAMEPQ7IMV7nArCEkAFD9Z+e9zVSKJwamV/f8nOx2PhHDgqKqjy3BcOpUUKgKXmM0ADtq8BUOTieTTgzijpnEDdPRbIegGM+FJV4tZmdEAnJ1yv9AV4vrgXDiMi1PbsYEnsdvPBF8HCcNn2PNTnZvHe8DUeGXqZ6Ev1yo1ExKPTrsr61z90P6o3Nq5BSkz2cBh1SnvJDmIeAoc8K6K5lqpks9cQ3DA60COWPlib1M+JYQc9Acb1zbXTlLaHh9UG6T7xtcedSL4LnPzWot9FyTCLpG3bGZsu9ir45L+zbo7rcXB0MIlcd038FCWtH1fbI4+APkm6aS6t3AFBDVm9IJWla4nmgQJa5RNO5c/npx5HeC1TRbswDGync3+8q/CgU+KRMml2JYNMbJuQTipHNL76ygo+yflamAMv+ce0VcMGjwJjVnTLG71NWmuALJz5T8ZuNLMZoMGtzNEodAJ0vlLV2zQb03feS9DWGQqfh6NMcndUiHk0f8l2qObGYH4hI1bsdibmS/3t+6bsZiIwR+TRWXNYdVAhXlUVqJqzUCVcO589pZegqp2DO/tdvo1CmTn3cKYyOWAFV7TLg/0nRA6aITIC8RD/DeZr45Cc8QAKdIdmd27HjJ9cvosxckSEyB01TXbNhwC5drpWuG9e8/AcbS5ItDoFopk6+E7DYNx3lZLeS1c4Hd4IrqL9vWkg1mq2LHFYN2vlR3N1lM0Dv1s/WuclEhIb4c2hs0agpB7iFil9IgZ6cGntt3eEREk7AAaLnYDBDvCjlrBy/zBcseg30mI74blosIobMOZE1wJNd4Qv59wiEKhj+7yLdiiqdxuZWw79jPbIxRbM5R1wKpxH62TRRb4/6Lf+sS3gDbQ452u9Uec75FknApBNF4Ra72smZCsdR9kaJsfPKNO2tbSmnt4o0RCrNlrF9cbiZAVM1p0gculuvTBww32QSglDjyOZWO80ccv7oSoRfR+NkTXdSiqs5dca5k6w/YXf4N3nlCHXJ6weQyW4JBFIFc/ncPJEg3q1nIxb/rkAtj1TsKRPMjyVr2tAe0QJfmh50/X/vyu9CwiDO1MaRzu4/DDPZBquOIqZ/IxM46lbe9ob3SKrQrRLfvFGgAozXi0qLbFt6s5SFXnsyJ4pDIO1+btYP2TpvQxKZRruscNuxnDx9l7pRClbD4y4HmLo/hqUJPknvE4I1gLhxxwo58Hgi9asE5UOGDwnPVySOxCRB8Rr51sNQJ4ARfYVeZAMUNzuPA55Du0QfGJa20MYL4jCmDqKa0eql1C45K/EBYoRrDFTyR0N9wszrD0TvGlJHzL2vziE9bV0ov4gFMWr7JwljtndJ9N37FMu5wYvs+zlEn0O8o5gwf/jw0D6hkA1o7OhNDGXqWpRJiTyPCri/lZEn86yU/D2gxUIl15lB/Y9WdX/V7tEHATIsiXg0ZGOyORNOidMOw8wI9GJ4brSqZkEVudLlKDwvjxUl0N/8hg3xpIi+Tb/wDfRTAwTx/ASfCh+E/E6KZPNyydcZeVW2kOpP3OK+YoatE/qfWCOCk5dI8rF7QQeZuyJoSyvZ7E/wOujiHByGoMucGazEl6b4CEhKUvkRnga9utHAxFjXzFT2Qlx7MsiW6Kd4RwP+43FGeigU3x5keEoVHsYrYfQ73vHho74bSOubBs6xhCzo/Ty8VJfAei5DqOHuR3zN/VTK2mOI/SVyoIyMEYJxhZg3N9tEsdB5kQ5SfS+oihJy7yus6Vq12fFBcH2bUqlD+oXvs1HkMXMqJbiOafz5Zja0MU+FTvbioBiviqvNU10mskZ4pYmXESuOWTqBzHXKPHvjX/qOqGNj6GggOrr49CWlHYZChYFSAvMhzViCvD5ep5X3SXrLHLEIwts8OLdFl8rVtqAZGzqthOu/Vl/7dvcj9Gh3DDCCVkWCKJwFovl0gRXquj4f0kKcyms5l6l9qo1y3BjiK3hwP47k2tzeAey+HFI/3fesumWY+PIVgTM6vdbPvi847Q2J7WVkW2cKtjTU13itsMgXzDKDzJkRbHeofY6zGcVdDuMBAN84b6p09KMDk5cJMrwwf/BEkvrwgkf0iUXFRr/SY//uShOiCuuqRP0rQ25xQke4I59Je0Bm7QQP5JKeB7KznlUTSZVDlI6/Xv/YwqME8d5ZtXlYW218mnSE3qBDvSqf1GpLUviQYGcpt50aBXHJVgz3stntXU49OYTerM45Ezi1ZP4ksXggibiswpbZGv7Bb/bAGYNBSBfv+O2dotE9Lezpg9vyLjMx3c8hcxRCaYh8XSsA4RnOnOhJgeZyZQ5jA+udxJsKpRoNSHGyI/DVIAJN8l0hbRO/2YpYFQztyb3cFPGwVl0OguZiWu9DOFVdsHSCXZeQemYBokh453BCxQwIArBlHxtbot6/Gjs5xE0CFk9OjJViFVg6688HUvbO2lY5W6YWZgodLCC6HR6rDcPgEPZI/mKgsnad9jYgfC+W0eOXxmBYPGVwG7W6jhuZY1WCCdyW8Rc9JJMn9cx8UmSrE4KfoprlO7MRPAKyTJu8qF0EjdOtgqRGpA4oLQHDWvbW38spG1rQpgOpq1JtJdygGGMBCzkEtirKtWu0xT3bkuqgwZfS9dEPIkH443Cbl/gSkLMWynxu8eYw8lPKCWmYtEkly+N/QyebcLcJMGJKYG8/aPCK/24UD+r7kEdaAthdbmgzOMu7+75dxRtDYFEOTosLzBz9uPKfZT56K/gdI6raxbZeGKRvRV2/TXX1J20lmwvat4pA+vR+ku9ir9GfsyHQZLa5i4G8lDcSIWsVyexzRD+uJXRbzdOgKzdutqfjp5Ra47GRc6AMXQ8XHIZVDxG/nlmOH5ApN3vLB/JZM76DHGicpdmoTXVsjUVlbetzDFxCGBX+zJLiau3Xi+JP3nYyZRw6aOYjfIp5210dKIVNXTclBkcs0hzt3WAq7PjOkOHyCWFQpZONEk52rhR/lTj48S8O2cOk1HpB8qQcvxeoxKgwe8Y/lYm3MpX61R9p38GfKz3+Ac7HjgvtLCQyNdhrF5atOXwUVzdc437PXHpKjQhZXkqLP41i1SC1N6kwLtWWsLTO51HqC+k064i6I5VTDoDgWcCTPsI+3QIAqhH4gGEA=
`pragma protect end_data_block
`pragma protect digest_block
1c22d08bc4c36762a0a49e9f6e4a773d38f5268c33c4a7d54fff2a4732517e01
`pragma protect end_digest_block
`pragma protect end_protected
