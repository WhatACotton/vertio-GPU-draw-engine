`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
uTH/kavPdyR2WY0mWOQYrbdWQ0nOILPuavYkYY/MNXGEUTbJGQUrD0nBQUztUNlIL2oWi60D+7A/1xLyshDqilJv6Q/rgpGp7NkxGkoHbi9fr1GsZWJybsaAAKQ1oXieQs6YHymA/Xoelb3WaGhshZ7yj/5xB6ys2U2+oeyhLZioGGO+chdo/x62AoUG5FC0h6EXr3og+O/zUH55nAVOGd3UrVDooh6sAEis/NCtgYaex4fI6S52k3Qgu1ct3L0jmlgajaXP+Odl/Rr/YWZKGMEUd0gmiqy7XOp613KNwGvvbHnilxw+SPx4/abWQwFQGlzEtYrOCdLGgcVcA91Q5lfXoCSNN17jYy1aFLwCnwo6vptqI2ONKSs7155PUVoddHxIVjAjcaW3ls0YV44B12+/WGsAglyCOOs7oAcs9ZQBf+7EP/cxMMaA4D0zJdbqb5Bv2/+jF81drnd4twiaNDDTCHKm3agl2S9dr8+81v56Xjntf+CFC3kzla7b2CVI6GdTyICXXRXX5qHpKu5dQkU83HLBqXMPa1fPIWtPMj4T+luj1qjpHC6pi9WT/i80pFMsKZwaLLhVkivfYe7wBb16D8ns2uE1qDqqMO/g5paKg3vr2eyd/aHitP/PHnBTpnnNXE1j98vcUaMgJu1YET6tGiXYMAxOFCjzAFdKs7nd/OPT+cdUlNfANMov+JcAcQXiJME/NmwIWUS1pjGXan4Ee1hRtXEpMnF+e5qMQuxRjU/UjjadVNx110+kvojnw2X8yru2jGKbE7YbQv296ZTmiq2A9MfZnPfz4rHzGxnUe+Pr9WUNKQ3CCLEpEkdbYhVech5vi0mYMi8nahcW7JXV+fgzCNHA2deWx6btv6BVMDF6C8c4K5q2WAMZwkDmBYALx37szqzJ39d6ql8u3BuVv+J3pPvs/F+iulN+yuEHtesTgmhh+NhSGTsg6F1ZWD8hFlhrBHEWcxvGad9btxYu2aYg+1v5L5IkM7EqjlZroynMpmQ2sWaRSC2t5LaeGMlCKXztihMEgu9ugqb9qgzzo5zt84tzQWevCrPEnRP0jvzz/RmZtW5iThhOHwCeg8C+m2qBHPeu0KEyiz5wj4tQ8rH+1ANt1TYo+1CPci8si8yLH4AlNmA5LQ6HL8qYkpnoz3Bbq4Epa2Iu6Vq8XVUWBfNdT2B0v/bFT07fuRXmCmVmLi7NI2DRJWTiSGwqI3qihl89Dow7LCP5kN2EqSMWNqoVd+6zVHmksmf6jGB6yej4BglE0/gy4H0TNoC5Wkb6lq/MCnY0nl3OcOQpMr8cvMymFnj9wyl/DL596qT1Akc9cGICPeORttlEIkWYvhVphVwI2obIZrDNepwyDTUoFrUDuHNy0XQUsBSP44KUM6pvBQmEdM7aV0iUT9GN10gZNmCfd5EB29V39iRRAxGkvySLm7ETDmq8dFHvDiGsXQ54+BZ65QW+sDYMxzFvT6JfWxhp5Bi+JBuJdAkpke6O7fF3zLoxQcj6sgnSFVDOJdVE7Ebkm0GTEbegvmGWXs0JLZzNdswQ2D3rE8MLw3zrfxZnNWVPYQfCj/iWUYRxcEOgGsrB6i/DWd6isAxrYD5TYho84w8CF7eBZCtE0bVR0mC4l40+q2zyQC0Uf/cr9xaxvDeORJHk61wger3C2ICBDcICry+LvDaS4CrorXUaIdo6NNmX2h9H9OlaLGuTLFchXAEFeRX5G09jWgHAWkyJoqrB+nWU0v+oKRga6mWa2/CzQrLPu+cGCDCoBQqca6AYiTtd1Nk7wsOz0B1pygaRG69NZl7KVdqLQXMkxCdd5r3dESnOzQBJEv/Wqbg7qNwBagoIRMVGJuRFlakKO63xUBFot9tcUHCcAXbmEs+yQRtiiTltBtpmTPWq+y2KThQYSKWmLicaBDiQFJOtyjco7NgievLTYwQFrLDy1AvsAhiaGPDNDWWAeSD2gLyi9yrZm5X4SFlMo1Z4F2gUPOHxvj/kbvIyWDTao+Fa/busLsDG8E5xVopBd7qOoCSVyC6DSa11txipnk4Uxa+v7bvKBuL20bV5xzni7JWIZc8fNeTSayMqSyrOtRBZ4SXRTZC0YNRIHJXsqQcQemsMokymlGbHoPp16WKAGoK1fbnE3cJ3JyF/1bUCCruuPLGxW3se04WcG/cQKWcZ3/7qJe9A7E/YBNn8S08FvBcJKHiLJWpe3qiE2TKPlr59voAPc14yZYq+HNZ1+fZyij5YFbECRdQ/xrVTWVPIKZyRr4LTu/v89D8fv/0Q7w5noYaTTPN1c7wO3HRcbJfBgockQdG3+FFUuc7QUCwBQXPhgxrToV3L4twc2zJiFS8NbU4GE5wPSs3ThlLfs+lC+kn2BEvrouSyv2T5TnYqR38mwv1Wjv7DE3ShccBDl41qdCIlxZVcabgFOuQCUYC/xhXAAvy4Bkjj1r+aDYhr0KNCRJfytmGxM8i06rPDxG8qzlOWYyVFk7ySlsey/P5qbZGUNuaWdBmE5zbpR5rACEyX0iElNW0H82ESdWpdlTjik5wes5/cbnxP8Um5bdaEFAF+yWHCg+jOYvEHUhb2SGd1dqK5KeY+SZpvtroO5fGzRpdecle8w1PXUuvgcn10V+ZFkmmWNf5GA74nQecNJ7V8pkMhkjonfrpY7N6kv3jgXNLYDLfZKPMI2A3q5NSKj1dHzScB17mtf35nxfsSqac8zOvPuuppnvP9ravVjoEdwS/qGr3csa6gid+x8gwmY3qw1PeaPFUIknau5My3noMHaV7YlYgRJXaaSiYOZLlCoZHWiGZh6BhlNx8NCokKXxovOh40UZtbW4bYMv4fnNo8MY1lCIEZPzAhXlGzMDV8yBxUPlcT6Qrib0OHDYt5yCNTeYupzQqR7tzlQwN35WgjZaznulIms5dcBx77vi6Er8FkQE+t4kKx4Hn58Kosgxxwf6Nkeedee7XArxxXZo/f5w0EmopXr1RaVuAloJUDyG/wiFq/BCkBXe8779ibFmRSMgtwR+altyPk8W16WOJNjLc+Z7IcXSjayiSgK+FwMV5nE/kyi2W6yNqaJDDYerhXU7NF4GccbLtqDK7by2lvrD5zg/fI+lQkMzSQWSVIXJjR8v37XSljuxZCl3GAzGrtpF7i7pHkX1G0izMhKh69+FocAzU299NO8CEmrL+T3/nE/QaX7ThYvK7B1n2Ls7tZvjgOp3Z7+Kz4XZx2wLs+8vpO6g2H0V3SOU6EY4YiMFDstcwGh1ga2+ZWSkH0N1zN+wzjgVsG4JD40cFsLR2oDskAsE+y7Btk774ID15Qqu8S1ZPFaYuFecKhQcj7x3ZmVTqRGG20LZTLNmx15Jrn2hggAQt2c77Nj2nQggiIU0u/Y3CXtJAR8IZS7CSLSiLrwopUvOCeGoBbPElrzvXLSYF5bNJJ1RUb2W8OO7NnFqRUmfp9ICXGbrCxl9i+dYkKlPkLha3LnpBXf9s94G54vGNn2ERY/0h4aW1RbQUxYps=
`pragma protect end_data_block
`pragma protect digest_block
48cc3b6015769d4972bae4f7cc3758583133ba968eeab49b16cb87bee4014660
`pragma protect end_digest_block
`pragma protect end_protected
