`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
XtllpfAhmII1n/Qsk5QjwJna4ZRbWYKc9UJ8EFJIfQ1FhBeyNiXfo0vznAHvCbBBA2XPMF5eQU9Fh+Uz56N555ST/bNq3NrjMqGEIIrWos5JGniU4BVsFg2J0la+hxRLdSHgV/wWha+nO4p/JkHZCNPOeqr97OCwL4n1ZYWzyQNRyGsJwxpkc3DXRkOZC8HWaV26HXJK+QuD+UITen0wAyk7BnOjg0YuGkAcwQSKOTeMhXFYWcYzxCxgXfqlVzrHJD0VCyie9k69ZatzqvPvUMVl9+i0KHR73NSooag68LVyNyshP36OZpnBDCekp3rwomBhBxtSTTCMfg+Z3p/M32ds7aBk8tnjlMVhXnkP/NWYHrlD+qbhQqeFP7bN/Sb06NVF6oQMcbRKtD+Ry2WFoOmpuaIQzvMwJ6JNAxZ6EmisDsNMe0QREZhhNZfSubsIK1CNcTaM8MGxo6cYWpmvifuVsv5WnpCXeQKL0B/fLK/LgTbZLdwgQ1GwqLZtW9rH0nd2bd98ERekEeKU6EMmU+qF1lDev6fzYy9AasTOw5761hSKVmZRx/THUP8ZHHlHIsd6cnP9BRAXpsw+o9J2eKPBM2m7gvhgdt3MmkO1BvL1H/uVjwSmQoNSG/J2MkUj3S9S6GvB9VWX0fWl0XE+SNzhO9sBwATagGL/e64IdDovIvDSU7sHkKZ2UOoXTo21N1m+JEw7bwswmezL2uihKeSVZYIhYuJvGl594DR9i9ASJlyz8tUF9k4XfyHk1CsUVI4z0q14LVlsFD2Zr0wmYnA55xJ0Xe5wpVeEIcEmtdAeIIHCxDeV8tfIo2G62Vrla2/vQO7Y9s7NCENZTzq3GcuktTDtcX3Ur1f63mrvLxk8nUV3t/TYOtavjLZjdXiBLy+G9TTRVGMsU+LCrWF2+U4dNFf6VKLslJIp1O5bRhpa6CC12Wsc8TXYeGqwrZpH28kGs2/0G9YQlRiRIJV9cekabVJemSQfRDbBWjNTn8Jk0Hf2dun5OXfB9lg0vOE0FtSMJIdD40Gjtl9mqRBsyrOCCrVHDy1bEkKGrjTug3jtLiC77UaSN3GSJL7j/1GgQv93Hi7QRXmhmOP1w9zWIAUwKjSyAYvO8VrhZ0Oyh95eqsamOdm6+VUq0TzOM9HO+KzoweW4WoYW2w7c3Nav1IB0OMjdMspms8MPON86+Fi0bGPjxVGp+NXK822MLASohxyMSTOtBifNITIGyRzKNYFvUBOEJrlEGd7xdBO13h4/Mccq8E1knGf9LCzEWiQKS60CsEuabzJjAryZ7IKgBCsnZEOsm1PF/WjqmH/XxIVNRzm6VUHQekxpSj+873IOVDDO7qpqFlMs2gjEqYni9yohOAoVSAC7L3X73AbSKwnasm380LyxPaSTm9C7/IYKAFGViiVrS0WEmsS9fek/d7Hpq2uWOn4w1MkWKmrLrIlgONDT9dxbyTS/L5bjO8UUYCcaGvsqLchkdoCG5uDpXThs5UVLXRPP1L9DiT/nOl7ulbEMbHN8kTWS4Dz7LXbzVR/y6t390M89zKeEjzCg/wGX264w7CmPw/GfkaE/G2bfnmv/XJ05/4F+GRUSea42OIOvdQCBWoV+aKSTogrUCQeKK7lkpARaMfisvkfYtJC4MshHSJpCYt7asYCtTOC+Vt7+nbYjt8kZfVwKugPdxBm9Q7QHRLGkaAN4qXQb2m7Xf8Hek0sn+xtoXlfDNqCv2aXdo0Cq1lDcZZqUMYdqBCqaQtAHa06FXFWUzu7YOvHTmGis2qck9n07CeKUMFqn8Pqm7sWx5v4cgRY63wkwrXETLeJnCJULdQ70UjvydfF1aNkkl6pTwKxhHY+U6L6nUvJnjPlmpbqUUq48j+qIsflOuS6JvJKxNe6iD5QccwN0rbMidjOAvSk/sP8dRw/0v1mqNGDEWTThHX7R1pIbRJoP2+rCwBUkt23LXFksf6RknbNkX3afSRiJUrT+GmeeaXR8vH1L2moHX5y42qcc4NSw89Qlbcz8NBH8ODuWWA2ZstyBHRu9qFoBOkabH0Z90UrlWN3kl2i0gBdIkm6p9fit/P7kKbDFJeTjRoiEo45iGDkoxCP7xTuHZCtRX3FJEPkdhIChDNwr2C9ZJRrkSIdlfEx5Tnba1/9BtsiQv2A1xud6paxU3SlXEi3chw1I1CNwCsOQgqoc9+QrBvsoqGKAESQnDL9dwvXNgCtr5WWxw1AnN6DQSimOBkFOqgzfzTSbg4nT0HOZnGW9CnXg3wFY9QUfA5gKED0qzqdjomk20Cel4TmwcCUbDHJdbQ4FTkxd07kGuxN4xCN/6DX8fF4BA/Pp8kFMqmsRRpaBHM3tBr3GnOEprqqvX0Ue6xbQ0nMtxhuVdFhkWmENUcs/m0Lv77nFVDS4TNTeH8OupWUrvF7l+BoCUqOqQL5VXXJaQbcl/DjhKzV7Wsa2Ca23CR7zTNowpLyf+5e7SlRrAOf/TeJ4EZSnjkIHaSdYNJOVWuXjcC42S3cvGqV1lwFyDGGtpcmhSimwGFvm0GibUvoc2PhUFX8SywQYoWFlayvwbWkZigGvuBrqDbI4pz6lNczXNhvPujCk6yxNj+pBCJfR4rJCT+zm8MGKfar4qzANhLgVoUG1QZRz6lVqjYHDoClzYwMv5aoPkh+dOYaYp5pGYzQEB8JTsTponeW0zI25W34Jr0w/OsEQOaFghx1hTaWCtxteC8FK1zGPzaib0WP/C01lGMtpdvdKwmPTAE2eB3ZolGJqXpF5qZ3b21CQlOtSU1qriI0SbL3FMUXgFvlKDpGnRKFDF/mie9luWFr4BQM4BZ6NGLrKjQ1TmZ9uAeB+9oRhtKKWu7JVXpH/+JusiWhfs7feZtqD4h7NmP3CabvraAFb3JiPrg1+BXo7vvd0h6+VACSq8dHoGr+h0WXTk1Yc5Kn/iqusu/vPA/jNlnyESQu3HlOoYM6bDgcEeilahNMLN56CtoOSHQE664/vTV8k9b7R9T3T6sk7f9uSPWwLQRZGg7Mh3QXahIiC9wXJSEv73ZKyUbes+ROTsBj0oK310ar6Tm3g7DBGg6qAczLlodclJjknczzmP7EpSVpNnLtDVVWThGfXQGwzVM87yO5tmI090HzGrhrh3abtHyEVD6UROFGyI1wl79YSaOWIo4udlx6++pRddGJSxCQnVH3gOOxUQIe2p54O5KEaUNwid7k+7KbA7t4MdcWqdA72rf3cq3ArdosJZh/8K7LNoMJOvO5sKVVo7Oouu32KOcL4Y6DPujJxNuAkFLajMqYR/DWhYdrw94/bN3KECOAZMzbLcWW1DxaYbqNeKN4ciGJUfv4w67JcjzY9vyzSeW4T02BV5mZ/VtWa5+s9qEwaxc9SvgmJ00y7JNvGJJDKrua40gxJSO2pXEejz/aFNTSiHYcBPOHoF2M7gipDVowBPTdbY2f8F46mFEaBoLeiQjdXb5sAxsLJrCdfnR/Zz/DSTCCrU9p6qe4fs6HNsLbFbsglz8SrwZVV1sXI4JqSV2rQHxG0mTSlQT5OycXfTZN/PbCCIXm0Fjb4HnqjFeB7ODmCAxoo77Kc1WZxWDx/JFQOiTIWJ/rls65m4GYb+QIwhHE9GIQjirKR45ZhfY0Axdft4haiInzLxgtsVAqATGROzpyLgbKpLbWAj80bjTKedmffYhgWM0qG4RmvlJgdptUBgNST5nanXzRysk3JH9HB9SHZt5Db1yZxgsGK5zZpM5laOJW6DdFvByy9bq4NPAFkpLdS5x+roo23s5BdUxiEjQBNelOWzwe+7x6Wr2LPVwzFKxMCmw9SmyWlKdrFmcnpgXKAS7Nt3bR3EeN8QypFJBFyyeCtKHH3GMZ0nR9RGcuQr+O7v49iBWJORKK8V56jXuvW41ceFFMq6mUzjYzgSj/fkwanQyq8vBujDW+CcdrdoMxjfnexFx3D9ghkI6OgIoc+iQNeFJdGMwjMRuKbuIyWfTR33w7AQnnRB/zyigGjNp4V8ZYeg+L/OPtrw5YHJXcYK20Z8xCB+BNslPle1P/gPJA3CmAJi0u+BYY5Lz+c+iq/xliz+G3YChSxbdNc4GSXUqe//P9HYEs/tuXi+dMkUl9/lukj5Zdpl8HUi6uPaqRzqA1KczgXdl6g/voToSiWFnabrV+YTftUGtCwjMnc51UVCDnCi9uKcamcSNACL3l93kDblKXxxcTrOBKWU642Ve+VKlxp/PsmWJFgOAF/wYod9a8ZDgOhiajZp6CBNZixArVvHwl9iWU53nAY0eHelL6NZbaZh5xJE7qjympw7fEev16STlThGim6ziwnh4YXwukXC/ga2c1v03krf7mTACXunN9313KGSWfR68jequXpGEAObN9KOCU8BEntLMhyO3exM//dZZrkgb8e73Cb7Cqyrru/d2zOYKgf3tfBK1BLznWLvN+rHrMxQuSpHP5ate/9896IWIZOTGuZYZwhEm8kOAZGGCSPTi4Qd2E46BraJEQwgpyMaoSOQ4nrCxyvAAhWOWGjD8Fh7qzDkOOvqnBGivkzrMieq4ExUDTCTl3iGVZM5G7TPXo5zCS7cWJrUbohW1/GSLm7yjVxBMWokwBQFqCvCHRwo2aqrqG8fz8zQ1UWcrxg3oPKkyi3U+QPJqOFEXCqKdmcWO+PaVw4amUnsM9bvOanG22GpAWGDeIC/i4Lfb5Fq2meTw68tNPVryaMTVzwvobGHxuAuBYUfg0osU8woDFxgEZOBAnXS1Y9d47/SSjZJEMav7BeONxFp3hq7oXK2k9YFYUfKoYoK379A73IUhlCKZ6tnHdg706K44sDNYbLuDVVQLMX3f9pOQ+IbkNEi6m0iBFqqWjCQ4gQRfYzD0QkAlbIwcr7uS06xzaZrnTQESGwb4EKiLxkNSXd9WzaDCPW+sx6+EFLCD0WxlWDSfTCTLv4MO0L8QDM+t33r2Bbg9ddxiZ8gUat4aaSBW7fZ7QPdzi45UWXLi12dnO5vpuzPn+6cgq983caQkIoxD4B1JnvuAXDIsKB+1Vl6PZV48ZcspuNagvVmz6SaH02s7tsiAvThyqiEmuDoACLyWhHCQXAi8AIjw1O6KOsBH2ojUdr36TnRyTJ0cGi/u+8e9bvBPefCIpUv0HVryP8wyaGcT57JromBVlUZQI/AGZRwjibHvpl60AEN8JcuW/R2qLA6sAOtsSaHOayEfv1L9AebIyWgDV01s72EfIUXrBguPPl+ns0bPvvZ/K0fzMnW386q3/e69GPq/428Cy3nYDDEGybhflqCPlAE2kSHxcp2TqCN2fO1XrqPRxKNnsdV1zOYGTDPR35KuzcLxuWVLr238VGyVtl4iDqmfJF4cZsQPzpAHQhAdvs5HKfne3aQhgE3j3KfvEu1LF3ASr4pZtjS2FMUDTBXCqUhuHvbT4rnccsQPUvtsfhu0jNEItpcsFjMOQD4kX5OuXwuE1TsDKjR1flNdhUHgDJSRqMbdaqY7Nz8pGpHPAJGlVlCFrYFFECOQMaSdEROE0bvhmUXS6SX2tFozmXAY7VwkGwd+Pi5JeGnTgvcuoqEfspzbU/ZGf9oQ7A52NGGe/phrmW/rbWdw0RctFgOJKE9SKVoRdOmTJK7Wi/HQMMNON2XKbhufzokh8n3iu879YS602Nzm2pX2eCtBUNm1vPhmNdKiTbQldroK2mSqqSTC+Iu4oDQuFervt6EsAlkjaOrKOTTCZ6QUQhXYn086lbDCgOWghs6nqbrgvrSytnxOOl2pPohoyqbdum3zX4sg3gtQBlnENWgswW2SYRnwi9AKIMwLnUZsDjJ2fXtXzE/6fTqTTED7+6FeiU/EUGC/DIL1ps1iQm98havzmRSQFU9RVr2AhEFOhz6hkWNGALllsrzMNShmD2RnWcd/zfHr/p9U8T+Ljp5ffN2wYekbi9GdarAtgF+sHxVVA4b8ZIc67sSNw2+eC95sgnQnkv//ATRDUvAXgK3rwyTFFWrIYbM2YHXOooHiPHX3wof0HJfkhaWwKsd1FhxZ+UnyrHXQ3tl8r/tI+iEWwlFo2rQonUX/HfkPKx6Delz4wIC8Nzx9e/qvdEy9YCVjPFJrOHRlUt87OnTB/qnolilbcROGAdohHSdB0lAKGAbHskC+3beqaCh6ltK0ByCInmwWMQ70IeEZNU3upY1MUsFvIOx7kiS/QO6gTFyEq3XAQ/pWxOdFe6nOQDtpQu5FFx3xolDGatC+3RO2b+9/jurBPkOcKPfqTf4PmRSmOrhqpbyYp7vHk+edRnua/Vc79G6CDyKUpzId21YECxqypbhDeUCpMUzaSKzb7+2oewYavKZlb7pJyVeSzMN3t/iHBDQdoxypPGhr/+tmBsj7Nnio6WBf+qiwk+HufmUGIARyDJA9xLyhAwqpZ0faoPTU+L4pXzEXlPmkErjsOlUWZ267Etmw2GYARR/s7H6eo0+8wmeCFexp3wDvO3hGQX/pcXRH11UjJ2UGRw73UvfesY6p0Ud+lNsSWe4sHZx0F0FQOHX+vi1U+cASLwtwCfuLece4gJmE0TCyE5YNMtNTQkiozDAWAF5ojejp+ZSyGflYK3e5lHiALlf5AV7u3oZX3UDLU9rX6lfoOUTQqVfCbjBOfd5fe68s4q3OODT0UdvT/3FemD6uEqg2KqzM1AIcGWuUYgQMsDe0xFuzBzGZ64B4eLKdfxpiTfMPQIhR6lmJthZax117zWihN2LpFeGbvpJIT4ygPScWw3TJOOjrUVMiz81dEKj9MnURPucR+ppgIE7v6oVem8MJ5yOo/caQX0qBEH+71hky8vFdHtjYpbE8cKa8GDZnUBgX7CFlMt3FTfkj3AhKakqng02ycfLyZhK6SWVFdemh1jcaKKKNf4fTJIUbPIdRjFSm8Cjjlp0w59LP+8jmonSUq6Rk0C8oBeWNmsDzxaEBo7i4O03aeABZHKPv8tBm7zJMDEAOdS5CWqiztsmyzFMVdGifR31dTrvEMthMsWPCyXBfVf+axc/WtQdjmRLsxzdUrAQtpNqA/GLszF/rMR0WZBiGYDzkDBCYiF2PT03tlScZ0Cna9SgLLUkbYL2Wz3qRv8zbT3Qfiotwy3OFMJT14WMKgyw4zkqnRuENVwee+6SyLnibC1HcVK4bYC/e1IcB2i6B4/mXP2vGuqXiCmSgnKLWVy+TfEC31X16/T/vRB0gjBxmBporW86CkoTQfkg5XGTb9u0aqhJEFG25eNIWVbiNzeCT/YSuQWxPBssMC2uTvfvrb4eMpbRizoFxiCysYg+Brp2PLqo/rIJT1GbTzaTr29Zwfig0ZK/WzeKQfmtIvimlWfIexsA1pmrKnCT/T0A0OrHENCthTfazcqnDhdtXDgigcs85OSW7LcR8FCb1tfx7HpgEpJAemL4VygAK0XlswVlrsDRpNY5/mC/rS8vc9KTukPeu2GPyjCjEvMOe08jFHbJwaxeezpvM8q3Q5QcwDLnjJCz352NY0NcVCWoFV1pFaInDpbxDuN42rYBBh580hftVCvEVBa1Mr+1xw15pli3oc/VaxcUL4s69i/O/xQSme5gaoHFFXdOjNZMi9VECv4L4UkR+cjWD9f0+3f5S5ruGXZSKQ07squ6gvgCBILmkZ6OhbWLfsYGB8gUUb4T+NXzpEJFsA+ZuPDveaiYDnOtInHNpjRAqWeYgHQKMBOcFnO2cuRBd6dfr4VSp4w39EJNQUVzEi8w80v2EjkjxwdbPsIxdnbGZ8BTuaPPaKPjHtADKnlEUUPuDa9A1Ht1CY6sdckfgj00XbUlJe3Ay8gUsSkytolD1vUqWTpd0WFFQrwEsL+y96/7J01Tl3MZ1L/wQGmdCHvuM9ai/ucPO1HlC6lqsGT7Hj05/ZpBybVvcNgwOW6gqXU91HCT/gPAlZAbB6Ajqm51jK9FtfT7wiLIlOSZWbjJkKZX59BM37eibL0jhcWp9rfLOtaHkhBFYFdOsL0LNEWmA3Nu1sKSGlpIiwDEBj2I85CrpMBPPl5PV7pE587lzE2ghb2kY27mFYd8TQC/z34F3AnQMAp4NY85sgD9DKFdU6LUqZ4ZrlVeNg2xtz/mqDQMwjT670xGT7yG1JG3JwKYSJK1qflpLfj///F2K86QBlPETosVrymL1FlJPGTiTP0yr54KFLi0uu9911gzSa69BE+T9qBTe7jzW3ZWrDZHp+n/sUI1tkBtr5Xrjd0YGBnH02W3XRtdlSGQXKaQLYYoVKvvuEKz9aJr683BjG+QNUHgVCLIPsxPKCSs3YR9jt1Uvz7I/huIKgvaB2QS+BrV/kCl3ZeobIFYEFlvXAp0Mxqm24IdSNngxZPgpSK+J7H/0sDdQmRPNzLxy94vPt3eU6oNfYMR6u0N4fLB/X8ggmS65xKYh7TZ7tTvo43aFtKyurudRydBXeHGYiJOf/4pJIgNGh/Af/3J6RkzeDkeELDqGgizse4wP4teHRR7DYBnB68K5dgWeHukFmbDl3CmU+L0BZ2ryK3xq83s4EGwdbxKKTtC/azd92buRfQ9Hfm37if12rVyC9iN8LGz69NgzZYu7uXEfJod19LC5npFxX66rqfsmJB1CcKwwACL2PQRhlf++Je2oB4mKAmBzSLqa2nkh9XQh9nIg9soyLT9sRFByjZlF6PlzqZrFZdbTt8CoegCwnwHpPX0nbAfGPOJjbu11lEx5UOTxAUK8hNjSleeumCiwhcfo8kH1JOak1GstknxIOQM1ADlHFfoMjwielaXhkJY9ePH6nfFEe1j+y51KKvCdfmlnpOVvzHhrnO3yS0CyiFUR7Iqh/cbt1YWd4PfcctrUyI5qBTks6WfYXvPSVlmJRnL3Vxas92T+zu2KFlwFht5QdKipIfHmyNSsYvtM7verx4/WuNk0Fk+i2eznFw5W8f4kvm+ElA2v71Px4TgiTz8WCL+HP2GK1LBuQbcl0JuBK/99quHewWXp7GCeVPilQpvEbS4Ck9VlPvObqIBZ1SsEmoxLE9uFfCrV3JEVqVJpfhP9VnhLI9Qvs7ud5UipjH9Az3SU2+rXUd73t8iynb+3ynl2qSDN3IezYK71J07RYTdYv0YOT9Te0Y0GPF3Tt4UfFPsvBa5wGcADyAQ2tF2YXpLMm8ciciGH2AeUEGYEioY2WEFmwpnJgzAf7pEIerfwiNKeHyBDp43IJDAOlXat2pSvHMKZJRoWjbioCcwCDqMr8qP9qUVh5Q1ETTv5/j/XP97MhaPFb+YypTpBbdDvh4OSEftmG9JNZFh15UPLRvmf3w0C2POhyHoMPlqQfUYoAx6l5QiZt6g5zUA7u6qJsci2XYa704yrtyllepyW7r9cweBtzb/O0RuO1+vg/KKGay4286QwlOtjWWo6ZDhMlGPayRehk+FVHBFjO5z+8FBFE3ZIz68BPVCeYbjYpcs0dCaUe8PlYSJFS7YgNfBDVDXrWO7d+AUVzixB0C2AkYTyygGyuo4YMxi04ufw63tube1KTTCSHoj4mwnOZIXajvBWr4uqnt0702pHhLxc1Ge5LOEDsJAk/2d5POv+r6FKFMjSe5Df1LNF/zMcwzhxEYcL/eWG/4FZONbrB0LFxi8V1tTiwE598HKkUIQXbvqrehLDKZ4X+iwI/qIgavbGPFv6IJsb//ryt7KG9iQ+3P6X/GvVE5pnNb8VL/SqtEzKfvb8FEZn+4FNV8gMAxAyac91aenBEiGWms5gedqYo9KiOdu4P/EI5LSPN9HVfki78+z2jg0FuUik5KiCnP8SMff6ATjQOTAHJjPKEJ0+8ZN9TEd63Fi5r4QOmW3qisggEOsD77H6PZ162miMbs6myk86v4TtILC26LEk2T9ibqUllBB9UPLuOOk0wsQS36ybj1DH7WD86FHGn4pc/v2fjr48I9ZBpBGc+py4bySmqdLYE86iXv23I2+mxyI1vz223cbJLj5uPtSmYuBuE40zgDnqgvJKVYokpfc190LI/9Vj+PvhnQUHwK7RrUieW8VIXjXnE469i27dIjlXyauECO6BGDJ9ftoiQVKIBZ6frUmDp0pgDkRt62cuWCOB4GW9MoQrV/SL3YrxdRdaBntdSi0CjYXtjUQM0n/X99MBLfNeNTy+puNzETpTRSOEb7xa4XNaN/4Zo1GsLTT+Edw5i5GPfKgNm6m1IzKXL6BXh6O8tYBlt8eROwoVkkblppMOiNRttPP9i+Pl3h2UmPE6qs2ncezUcZygOgYexLBDvjMZINC1IgzueU2wUcN16p8msWhjLWQkpeNiP/nbDo6hVDbNORSaCDBOYvMDYnkfMQkqom8T486YWLt1sth3l+D7XlUMp+UJBcppHBY86JyDgcf4QSPLndO1WENC7sStETwvVDofLn3eckScY0RQqIq2y/flRLDZMmYfgyRjmb29/gXCxosMLi4IH0VDxxpp0TxDsWDAGOW0cAgsSRoeamQCU0Jjw2VFZHHCW8eRL/VIpRku/087ONzgDnEi+jz1TUmW8+JEbrGpQ5uDWojzA+2oDqpcmyH+voexQcEwiXeJZBLRd47oQqnFjgdT9HbR2XrH/uNwT5kTGVlT3LPJV37D1NnYF32YgtyoT0rCgZ/NUIDXjbXfFOo6BQXm2uyr05GTXWW97g+MOyosoq6ZhaKGACelTKdkKG/mBiM1qIv7H4jnITDO01JA8N2II4Xv5P37+948RwgMyc3wIudo/Z9Uit5t0MZEW5Wyn/1eUGbdcty+vYfa0NNHwaU1PcKPQHUWh8OpwwO8J+6oTgDT5ZzeWTs9CDXrkbWcPJJMU6lmQRJxRDQ7v+5T2L6o2lYT3XVwx2iWgH08hoyn0E3pV6uD4oHLfSz5BPuUJelE5bD6FaSkTJ8V3FsuSh1WftmWUcTyWw/y8BzCCQ76HmKBZ30Fk4ijQXr4vaHxll0qHdiJYlrQl963ByqMRwmJlTvGfkkM/ZaqrovjyQqc0AlYp1DI6K7OIoRZJBVuGQlQuiN176BgvS8016TZ5qR8IrNhwnkOl6ZRdHocV5HNo1+q4Wx+h5uP2211lMcgOD8BkA6VL6mw5JKX07le6tSe7QEtXslBgQwP6Y5XksJZQDqw1XHdvY8XpR36QN/8LvdHuOwk3iXZlJAknWuRysCcgOuqu5MF2z8/skd7gzHONB3ly6v5+1cK0e5NyelYt7ODNLax4Z6Vw0a+/tCG+85pu5qgDuLHhQLifIUBvsdQt+SywUHP2jq1+giTd3LWIoVgqQTUGYVuKrNfgLEpzodUHv8UV6i/DvQl3oqMWWEMo2jrQWHb+dcTXQpRwhqbrTlT07w0whVzYRr7k7A8exmpphg6u0i176hIDSMeN20wYvFc2ELIVNYomiFAoyhBMAs6nDkFUhtk/QKupV9vyYnM/oj1CTB7vcJVQpCLqftsyXywj9d11i6j/a6sI3OsHHmzNwC0qdwDIqGH5OjIJ4H3a9UYPq2OFHEN8aa2VpK0mykvEdcY+i0g6cuZkOYrG2aOsaL+CoZKjmlIzeSs1JjVdigP7oaympATDJAKLi/4HA47oC3u/LGEKh1oeURDunNpvQR/TqsTtLxdXdpZrcFea+4dAfSqP3uv4mVNfZN0pw9vRHbI/yWSx02bOrf0fb7ebh4Am2v/JT/qC1A4CccOaN2ZS/Hs+Kd9QqeLLrge/UQ/XsCSdum7j/7DbIIHfZWRhK9dZ1++7pPboANJywngaVcFo3AXTOgp2/JL0X38gZWmVZvpWqInIInsNXUWeAG9mJrCZ8gPS94bvlGR/KrbgM7/DBIvqfO31Ar8yFgSL4bePeeBSyDb0PFhRGWcZFY6t9Q0GBsNFZzrAN2E6cEQ7MO+Qe5oEJwCOwHSTex/DRLecgKk5dEPUxcZEJssnFcqfJ7sMkaOW4POCVR4m2p8lWlYkD/o6NKPWp13KWmohg4s8psc+vWvKha5a+RHO4l6LDRM+2v9DIc/XTTa69mAMIgyoUjGiIMg5DB5/o3KU6Jb4KFT9oW8YtZ56AHynK7m2T7eznBQwR6p15z0Oa1Y3cQxMaYEWc3BXvGP1mE66dLdy6FUpPJh6/5FTtUMKYsWdIuxT1McFiMzLJdY3mHtZ0dvC4PSobV9aoTaRB1DluaLz5StKYGGxLV1f5vkvdXwbxy8cQ05lIeXHGZJILS24tKq21Tqt0kSz6iMdPL2DvFdXqufWRd1wCBt3lpfixJxxIJS0cT+KgadeGgnnztF836SbbUVi/17OXFuvqGNsl7X1GxRwECTMshnqc1kO/uSRvhPK0NVY3g+8vtR8OvR8uLoN+Z3CnbuRCLEq1I2sGF3YiA9RpCTncf7tozNZqm3DiNMsfriWgvtr7gIOQ6nwu7UV2el4Nx0IE98I2q05OD97fHsG8vZeTmY0RSpZifk/tA5YP8nzWIy3TmIDlpp+5vh9OY6gz8PS66re1tIwajbNSrq+0pN86T8T9k7GJ4txPWLL8xHm0gIi4lJFpdeU4WtErQkZAbuje/f0lIX7M6pqNTwt5D8pYz6SVlY7RI6oVb0NaRZTRG0SvWdyXP5vC3HRdA+VEt4mHcd7eL2l0P56ccGz++K4FbKWvbtRpVL9sl4TSnKOxQL+FnmRgZtzLfyYMFsifR+KLo4S3ST7CxH7DgqZuKRA7254lOSYosAZKEDIXV09eaqHKUQzAbGM2cNqMKsNvY6k/kYxxES8qwlOFWLpWIM7AxTVKzCIn9Bk47BavuKjs6C97Ngsm/pWgDUvIf4wBceD1fZS4qYGybLIiEG2hnr+9qYjm5tGxRWv9kstJf5W2qtDgPs+CtAXWaMclYud+iYm9/hSnePmjNoTl7LjDW6rtt61tfy9/XE+pVhvf96xMfwPHC81OGfBduh6GQiQOudnX84AxqwKpQDKurJyqIRMySO9PXOLCE0dmAB6eVd+K8SEJ6Iv7TYazTGqYs9zlafxb0AGTuh+idNWuJ+PNWrBw0WcdgV3NjCd7Vrz08JQ+HRtLox3U4+ar/KBkjy41TxvR0Iim2qcwrHo81DZjyK2iWKEJR/cxSHVVjjuC6C3ihNE9sht7d705aVs1W0apY7+mAtaqjySM1kypVbTv/ZyLZrfCP62VHrGqbT0asRh6WEhpuSlzm4vARyXQknb7r/eL7HVc9OrmcQZHO2QNsdzP7kND5b5P0k6E3dn/O87PzJVdav+uTXa0gZzevjwoOWbgn8tBYXbIfXsV29SMYHNhP85vCQQ02ve8ailKR9x1dW6pmbfPJja7x3ULg63bk9ZGn5Ls+OOgS1WPR9WHlvF9rqUE9ur1swOANpgBYfzcSixW2c3z99IzwX/JtQfnNxFP7feQBPUVSpaYDRJk8j4NscIEq2Zt+Y9TFdxADvYcBazaWGWqevSgjQ/YkFNwmBXIpbTq+e2Mw96bR/hUGl7U6XeiHGXr2mAdglAa0/gLMsAF4X1FgpOZNLT0J04pOJL4Tuf7VNLTuo5jCqGNLVMSvLWYjeqpk7po8ybiAdAgNIYIXyQu0bV4KvxOcPxx4znnok2tfNXrW6dvl/uKqYNgwLd059yRtTPH6PkfbKA/3elM0ULdmX3CSwwQ0th8UO7cyKeJTrFMp2Iiq7Lyov8oY1cYULtL9WVRijkDhIM++SlCzvjo5ah2kpf6smxXzex+i92mE4LV2XJEIp6toDMqeqOTZWExyosRJleoPtaeB+uaO83FjHfwlxyRKlDqg6kNOAVnoi6JzeKqDcudY+gAzzr/3Ou5o+mz3cZp0aew3NKNpZqXqnW/d44mGxYjQKCqCyRkpds9T8UizTVG4JF3Mf6UkDEQbrwQLP2R4d47QQEQL7kAVPtLz+qd6yoS6EXEfhwuPnlI/pqEyb6+LCpQQ/HPnRqpujtlt6NeR5pf8N3fmHz4lS/IiZ7n5cgG/maZAV5Btsqi+Ah16FCLr6B2XQ32RkAqGBx+YLDmMVRJzZOOodmqYKnZH0f/dOeBYTy2LyoMVWxeeHxEWLf2xMRD4tyUsogM3pFJHaj7Gqg51V3IU+RlayCJswMH3FKUQ5A29tGCbklhNl6uKgLrGw33hQKi89q381wuK+FI8TyMteb7Mr4/2D+DoNdGB6vmSM2hMUgAbWqg4sZlNu8xCQGfGTfIvqh2uVegmesJgZb3T9obpzondfptoOxCWmqFxunv1PIejF0mAzn5UNh8CYFncQiP3EzKpjveKWXcRRT//L8GH2hwndXX/CM=
`pragma protect end_data_block
`pragma protect digest_block
3a951e740e2b8e4ead1882b5a87701b6cd105003719662662f5a2d7ea5fa9820
`pragma protect end_digest_block
`pragma protect end_protected
