`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
ILjCU1MTIjW97VI2kGE4OCnBGD652fR+r4PgnbPtWbVfZVgEHLPMMYf7dS/lE5m93MGJIfz+eERfjnd8TL2LU6ptje8evv7e3wILa1Ju/ELMk9SDfHTIAnJRQ6JJ7Jruxb0TjIvgCjyF0C5vkTdUSWhEopkfC9tz1Z5tQjExMODddgIMqIvUSbcMaU0wZJ6QiZNqC0CZ4lG2Hb2ghbOd2QVGpzlP0ctOvQZDKKe2FEUA0w/5QUcx1NI5KbR+x/Oc1ELJyvEAjRksJGryDYlslTOxa/0rE36pR0eI7ichgqtTI6O49i/7XlLeJB+aqkILrVS50wvi36eev3YNLQNp8Zx9XXscfcRM8QTZwMM/NTX+37iTKnc1CwwWLK4N+NE71P5HhsbYN/8o3O9SXMN7t3Z2twcKl/FUIVoTmw4n7FWxf51IQYkKVTW3OHDub9xxCB/HYd08DQMUqyGi1uZ+jG0BgUXIyojV+2ibp+Hlq7BIqkqT6qRFhFGna/1QWNRF2OshpKq+GlZyYJZcxGsGCYlkF0e2RJSFrB6UBID8yFd+/yMD9wMZoLDWrMM6MpDhnOSLmSejiEntfuYW4CGI8KrXtrwvatL5jZd4cy1trF2aDHn5bag3qOBEjItdw7qLn4VjTM9CrsK2Zypa0em3o9mb68t98JwUiqFRALKI81hAfRj+8G3yyoWtyZnziO2foKQZ7l/4+E0V4XTLQtSPhj/TWgZ/+yaZKVlrry/jZPeI9P7CT6PYaJbaNTtmpt9Jj06nLUkEqR2SaChTT0kbdjENpUmNxifY1i0XfrecYmX6hqACyX9y38XBwRPWQBrx/Nru7e+bvjG/yeO3uX2YTbZg1uX0fJj6DmjASVOCt//hKIH60xCDOFjfaF6hl62jJt2QtgdaRbOCzwHW6+J1dpqdtQ15eNjJGUGKnGIbShJsnC/gXVKkX9My0EjVm/3tuQ5WSPE0sPahhxIOYiVc30qauEaXiiMG5aiPaX6k9Ir8kj0AMMlerzVfmegWusD7NNsX1MljEeokivU2Xa5Y+ebBETh4xE6rHixoWdVgSDkRyFq94RjqG+vclDphy5s1eBXZBFEBkvBKFESQoXL+dGzIgbFtViOVdETYVSPfEBx8eL7BytOKZjDyH5Que/Ldv+iXIK4pyDG12mKghwJ8M9kR3S8aZqn1DYi8aYFd2ZJu/Qi7DyqIhrUmt7MgW42WNCZkTfTUfwBMX0xjKjRNmWTFo54u3tFu6tLoYsazLsXu2ie0UmFhHQQ3dXb6xGJn7BA1hzeIpHamP91zICsS4r9FxIp987P27kjQllXh4uzXJCKo1I32X35yO6ytQryujvSFKCsRg6eIWFzS0Qjm8rhfDoIz+oIsPMagMcINBsUnLO+MfduN338GtoESkZncqSNCF8v0eFCAFQB6sBuA8ABdP8N6bi5TLiLCD9YS+nk=
`pragma protect end_data_block
`pragma protect digest_block
19a41ce667a71a6d15f4848570a07067e70bcfafe6a818b365f2e41d789012f1
`pragma protect end_digest_block
`pragma protect end_protected
