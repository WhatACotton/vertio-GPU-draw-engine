`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
2P9s/9h39n/RY4MP9iKbawsOWI+8TA19U6BEneKcpuWowpUUbHWFN2UJC+LLKi/p0MAtrv2ucigEY7+1orqZeOy8eHr3I3oFZyRpiLOA1uGDAXyJRK+JN/46EphqvRwJLGLtc65YQneSE6OXlwuKzAYPpGjsQQ8TNBvfAwZuz6NgKroUea1kUew6bh5Ok451pywZ+VIr7pVUreG63Z6EeQzWH/kag5nK9CX5d3X36/Tr/lnuGDmnIIEH70NGql+cD4JoLfFs8oQfNKtzZg7WGqrNCzVRq5wsieJ7QdX0uTo01kVFlO87c550+AqvFhortdBHwVU8dGP0kvvHqQK1libfnU3b71H2g4QmFPA7msGScXVbOGwNAGBiSge8zUzICMx9HMT5X07iP4RwSf4sZJ8iEGBZM9zvBLBLOz28xrz8VMyoyPEDPwPwLQPgO07Zo1Sphz3D5o+93kw5XtCAypjz55hcoj/T3MrkUb/b2rM7DWAPZWlqj96qteot3t7t5J+JVujyE3M4ydMhlJwWx6gukz1TyxnvkW5Sxs/hR7bRqlO0V2mmrS1dYF860cPo8yayK2IgN6/f+kNMF5kR7r+HQRkE0JgpyZVOfArqWcDGikm8V6d03gJQv43dNpRaJPRBOGIIJDe8vegsfCcAYCOxxTcp9rx8ft2bws46FvBXnWGqa23dologR060ACzl8kjBrz8TudUVN4hhnlW1AaTT5xozhGiQDEmKyj3veKD9w7ccdKoSmqoaJXCDvVg2ig4wOnk2SzDlaVCq4NMFIa6fXQz55GC4reBB4cduYmPSFP7KQq8A6AYU0D7QebSnAVJdsiKDrH2DgeFOWFeyKBjXdhuqTJhEmx1oRlQV/jmxuLOAlyDPJrKIrMNGGMgyMN5toeXcX+PttV7X73VbF59fktHfuXO9J7CYpl5gAqUBOJLdVkbq3YTd6U0TuYfKgJJAv45zLZ8JO6liE3Qzs8i43DDzyewlX+L0K67mgQYTLrkXZmVo6WVx3lhY3IAb0TZvMlOpB7iZ9SuPwy8pqTaRpGkXQktSKcbGxiCSQAxRMRqrVqCIQGiAlZhRxsTBCk2EOV1xK/SwUUVgVjGvVW60VTMKyKtBWWvJE81Eq9LZgtKNWDOzzl2efFvSdOMufT+haQZiqC02kwPUqwMxe2cxFhnqKO3T3k7TEeD7WIf52qX6k0Yp7ZUMMWJih5nhR3GPXlN418ogP7xB2Jv8UmDOwpwC3sNOgolDtBY9XzZtOtzVCcLDiATjarWg4+eoZa+pbnFhowb9rJ4oMR1oX5115yJshrStkanzptTZxInOlQ2VdG0+j07cLg0bQ+LoS5cDdChY9GMCRDa3Xw5XsRVR6n51RDDKey+iq5dqqQbg70ZuCeH9YXx7i6bj5SQEdu8Q78ZvWexhS0icSgL/zXi4c2IG2VsVmxqfBrobdXx7V22WjC4tXMrWFwf08+HImrwKMGG1UjCAy3gPQV1UN9DQD/mS19gmW9WEmG0rhj+3gCncOl7EC7RQyZ6GjK+wwWVaVd23S5G7jLoKyk5gQSfFGplskMO2VfSNdcJX8LiJm1ETuvb/inWA+1t68xYC57LbX2F3HmLqfj8mtvykL1pwfoACG/CO9dH18T3JH/Um2QBGWTXYtm557n9Hl1wiYUwdo0q08bD+v8HGLDhd30sbiXXoug6Pi/QmH9gx7X43CegCFF2RjBeJVpldId3wqnjQAgf12/UApWcMGUg+gBNv6FhJAPivf0aW16hBLeLrL7Juk80HnkdscmVFIrFsWIPQeUoJZa1lHum8xPFOCw==
`pragma protect end_data_block
`pragma protect digest_block
49dbfff3208ebb1bb847d1f37e89d519c85e530efc0e81e8d37c7dc945391dbd
`pragma protect end_digest_block
`pragma protect end_protected
