`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
0ZH6IiQFFR4Wrt/6+JSyd3jwhwiq6rzKi8dHxxZAebnx8dYlN8Z5uxqx0QrKHGKlxnOSu6aAiCEk/IvrG8Ec59QLDa2ceuZ1olOx1/ZlVSqfBvNKcepXPx4E4c6iecYtqJdcZroA7ElBMlyOKx74J3j9x1ScpkUW2Ympl55xRItYD5PftwCHOIQZzfckAz4mLwweq6ZEr32//Pp0+0QCNUhYe9jTjv8jV5rRKxJWkRqNwMMwOgCEP6dNYWeU/I54e7XutGUjpWue75oIZLjYiBkkcYik+AIr5ljctLT37fPOz4EtmLcFPha18VhUpoFJVWQYBlhbRTzrvtmDM5laXkc1cukjoV3byt2HHwPj7cdw9YYlG+g+DWNR0PRJs4P4zhKyMU3A5Q9N6iZUtobx0yQ2RfF9OSjGav6nA+qqklNFTkCENEVgyXWQstJoWa/M9squusoX7uXJ3anAPhZUo3JNgrvDkfjFN2Vo1DCsrv5RfV3csOnwtNL8nsqTSRpf0ltS7v5HINrgqn3apoZHkVYaMDpFm2otPTK+QOj5488qPez+zSaKiRRG7lpZe/pQl5NdbTprqG9fGdzp+sSuzd365q4O1UiJBi3Ru2CwOryUyRVyKnsHmoEY4MgqdY+tsu9P4UH0gPHhU9PQDnuQmQWf8KV3D/+gXI12VWNiJh6i1hNb+BaUXSVUm6+2t8LVauGti6YnMMnEHvkCI9RXNUqTU8JRCB6he2SxjOmdr8yO+oOZEXRBG9PCNq73WxDkW8fsBn9KldB+RMerotP9NuM2rjtvOdfFGgFmWZrPSOY7IQz+f3FMyfuzJZtscwfnScahJGkpIylWX5cFEHfi7VsZyN6VnqYS4lOA7y21YGXNpy9dgDPs19ORUQ6uywK4vAiM23dx/IFN/LATJUZ5MGF/qyzlGa/8pO3pFcTdoZJYRb4evoZVICQQQ05aY/WOHgGyPuujGl+UhJPASJVMNhqfYbUDTRi4JdqCF3Jnv4cp58r2R/Jq2NC86wDiyLKNy1SXUDqa6IfiJhc87U+3xBXU73vz0Arrd+59BwdJuQ5S7tmg468OFlnzoV128N6dko0ZGfUcEq6Hdy9zhkZ0BvZAxR0+vvca3g1NrOxqn0wugrnmkrVzRVsMBrbjNe3pbND3ASB4XeI3pvZEvfpS5sgDt4Lq5Oc2LvnGS/VtFnHUB9581uOL0WHajiTUWnatqvwHSjM6lfnNmn4AWxWgOGtzqcwXI1jZEaZFSo/acfly9dzyiRPOqcX+OwTSQTsGfJRCnoiIkK8qjmHuPXliWPkxSWB2CE4yX6MT7d6ZYDMFR5eSmQl+6eZIXK/JCOBJZDBT86yP4CiLLjL++9C+JiCBabjhQybM/WJBkJLcTnOA5qxNE/bPOMgOUVPk284jyz2lijWhR+cAcNix4J13YQohl0FCZp/kacpzmnde4x0=
`pragma protect end_data_block
`pragma protect digest_block
a12b223eab168b532256974cfe5b251ab33aeba2d2a4e6a0c45b4792f963ca32
`pragma protect end_digest_block
`pragma protect end_protected
