`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
msYD2hMZarYf3wJs4y4iEj03+l/MZ/IlTX4avmLcRG5R64LFuX9UcIPV2AyNxMmr2gxTf5BVmY6Uy6+D3SvYEdX/XtDm/KuaxuTkd+zsLLi2g8uNTFxaGwDXfvfk2wuVmR/LPvq/qjoB1c555KkUeC5QRSpjwqkTkY27Ee47vEVnvhjQYVCaZG7wm0t+QgqYcXZSkPmxZuuO7wLWCm3U3qlsCnWuNnBP11vCQTSZ2OkDAiKewQbaPfonvXedf9P0W1wLmkGOFFvElvsvnN1h5t5Pz2I2sfA6xBdN5s0JpYvHLOou1798FcxieQoDG2wcMsGAPQ+WryAfHA5M7ynH6gaueWs57llfQBwRweanup3uUZVDBPoEF50SIIyk75tXRbmoQVZ6M/qPpCD8gU2Jg8oia1Y3rA9iCZFPY9xKcC0exYoRwuCYhPG/yGR3dtLeaf0z3OP1Ou6ocYQNioNYlFr4W0fY8kXnIRXzOvJYUwBC315RNz0XStBG6r33Z8LM9zh481mCoAR9h5jk6b8h6P2M4/7CVGyo4cPJGq+Lz8ZpDVp2vTlZkk6S2kipQDezIr+rjk/1eQa2PJj9Jt5Ns3quCSnxUxNAlxqFcfk3ZCdl67/QHIOFvWxEKrb8fPf3wZxEq7fwgDNzxveSurNfmmTD8Chso9HfTN/NPGVBpy51slOxYtiDfKwHNwWen64YqyIFwuRN/OApa2mSAWQbpvIJr4Cl+KloGQy4GgPcearqpR+/3kJuy4FK8ni4eAkVjt3UoFh9iWt7AdfJ8VlsZmwk6oVpMwi3ov+KEKuFWxIS1WnG+kDDuwC1ZsXZfg+eNQ+IpIUEU4fjSKEsM6B2Bv612w3NQFNGArND4MT4JYq83Zh6UWOB6YhPWefFRB3rt41rugMoLso5VVluHVxtRYrwRR+rEE2JUc7CWRe1+2/Dy4Jjhe8/PcrlL+2fxgv2TiMx/zBapz/BE4Rg2a4CICzE7e+I7L7CdUrY1VDnh3RnrE4+xWv4ABVe92ZCrrTh/aURg5HzlDsC/GjjeOvKTmtromzGfJ/rnUuwdQoMmgzy9Ksrau4QAVJLARzAmq2NjEXYy6mwaZ3+gRQVsqvgE7DnfvSHHtZN4QC01OZ0lotoD2VGxRtkJEHbcq0ueMPpZziMV50f8rv7LOZin0AnOTTIN4/cjQcD5N4q7ukof1g52/pV5vs8VZFgLvSxiP8rtlLHSU4OgM8HW8ApmPaGQD9nvIACmUD+Zsu3gbIXGfwGlNvV7ZlVArSAKAol1zcJhyz0Z5OtQuYauu0sqBYLJJuiW8LseJ385RwwtIw9FRc0ziJEVdK3VRMd0huztKWysoT9BwQYPZBAaDuo23roS5KtM5aJlfqkA9OcfcakSia/QCC3JGCwy4GfvOFGo/2TRSjUWjI5/02PO+fSOAad7gg9dzhpSE6IVRa2ni9rfuOET7mkiIjv8rEYt3ihkC6nAAlwecO+jzpQoIHlbswrpnuP98i2oETTgjkp8RNMXTEPDbmlN0EQfkBfglj8QcbuAqLB4PwQKN+jSG/uYYD6ZaetFfzeMj9HwlMiVEfgplYiO4vog+GRWDTxARzTCoaLFER5N/KmQ1syeDOXuOmWAPchKo/sHVNDKuHfdviMrIeFvqEOHhyhDUiBWunWAJBFnaLXmLWd0YKbL0WFb17vwec7NZQX2pGNFCHOXGJp71Btba4kyyVhN66qkyzvQnKay7ceRmAo5IZfiUv69WwlD7DuJLiupnFCjOwsmUjR/vq/SnS2LEBNOjP6Es60QGoJdMOoFXGYplDTaO82bCfeAGchtYmsa8ARl/1Jdm4dK3DVKT+oxeITT7SoUFU2DlGGMHNIajGgjBwWJG8f4DOR4FeNCwRI0ZQo0yMvl+ykLTNlfIoP+j5sLPzO3rx7rZ5uZ22c/L/JI5lhMaeIbuY2IuKkcknqTepE+Dtu/iiAmVUfrTow02AH2d5rFdaj2StWmkzIACbZwXgOUnOPnUq+BJWX0l0qf5EGIzjscVHmlkU3R0V7i6IikNYeM3on+UZkkObj+Vks+TbjGAt1s9mPqTXaZKiqePXWLmpW27G9zLAxouTjSq+6oqwm/cVh3ghb4sB8Noz5i/w59ZI6LAjMi2o0wQ+J8EL6Lg1gLM3P9ycYa1N4mZWh3lzR8DIaTG6a1aEtoKUw4gb5UWNlCUr2Tcs1QTpWClNiEOEL/MRKw8pxLL6QgS9b/fH82DxpcHXBxvgiqV8EmDGbmpR3PF+Lr6faLzrjunIzlE3ehP0QoggI+clTBrivbfGAFfC+kpSztbm1P9qA390WBqj7j7MvqaOSnQqbfOSV1mOwcG43Tj6i1PNIv0iEydIBSzWYn023OARHGoR9emhTG0vGQgLqoVWzfEDKI0+VZnSzGrcvRxlxCIbwtIEzcxlg8gRtsSICjFeVYUs5dWk2DpnWoyIZvOuQNYo/mwB+0QcIekE1LjXI5tYVfG8v2KomxRMl10q3/Kq8mJdJgiA/sKxGTjCSBH/5SvOnwnlCwegspDrDUWa5Wmlgzb+m8VZdVsQbA7HK7AbRt6cpZw3mgIloDMc+Lz1cTL4ukV1MQoGNOLU5FBhd8y7ngpD3J9zk1lLo3hceR7atEihvYI3H8a7JtlSt8Iyqc/xGX/MRnJeaYdj31nVpCwgUG2nwovp2DycaINVHHxpItHkbQy1plWAkVy13Ej+tdvJNzLo8XPXJS+nhDg3DcFv3gKd6Sc3OZUFegBqi36R9tMKWpa/iqj7KsXR8f/08HAx3MxHhMGJ4Y91AKVWSP4P6Yp4k3MFTSd0/wBYiQYcVcCbVX6YtzbR1qZ8uMVHFlaKyP3gYTm7+brwN/gOsYi8u1JI44iHbRNNoyZtUvxFtdcyjfzR/uFI/1UcsZdDdRfa3LlTsWGMyoU6jn4Is9ZWaxFE3rmC6ijMBsvYLCUcn7GIQZUlAoYc6NI9ukLD8iTQyjjABMCVqpz4UvhdzYu6+590DfPJkP6l5UTTDx+Iz+iVKNqw3BL4uATYRDogKd2myLd4av5Rgbm6cKCGwb+r9ipektRSrWAXjnXkBk2exGowbaK9S/mIrsjkP3ev0G6E5XyUiEbNWGJZnJvztQ4rexqVYoIHZ9VDMpslKiqzP62muxVv7m0lC/vwmZIUowFkaVajOJi8mxnrAxJllhKZh8fd484ObnguFRORucpEbatcMbtWpm2cmXiDAsAd+6UXuADhU64v+pCc3m41bsbpmHjtweNHiLHGAeBNe3Wb36+TIt//IiTqIpcEqQPp/feLDw03Q4dYT2Pmb3DilPrLnbNAD4o8lYkDA6YQ6sHihC5irxEJdS1w0B1nPx3evVm1LSVqBLXoZRvtiBsKREAnTxFiDATj1FQnJr0sE15VdZ3SZUPohqgsxBfgGYLYmqil33UjQMu24/5X5M1rZ663QneA7lhBbEKAnXuzgGJ3XRtjypuBYrhH8LW6pAEPxN/Cfj2tIQVOZfgn2pUingdJKFLgSQwn4utDQwDxJKgoNdPG7Q5omaL2v5D5ga/3CfK7nQCpBYlmCRjgtv+SLjTTb8cIeC5C0Od5aQrpGL+rSB8yTdNO2beQvQjkleUP7ImReX4Lxp/6kHShYvAzYBqFdeqxDpya6n+x2gEMqXHj5KoivOMS32SptCWUZH7xjqDbRv5Cb/JwbkP1t+647XCClboTJidF0sl05e51uJAkZ4ef25PnAUizdPjYz9xt4aAA9ygJp70IJxjiO6YBUN1buWlQgRfVdhYzygMhgvElV231/PK6Dez4OzZoY5IQu04LgBqw7mZNP+6qxibwodjAN1hl5lnOy3iuoCjYtf7TLdbGITiaBLZbv0SY5kGefTZvP+mADaHwIy6gPLEUotPYSnZAgMZuzuNNgPWSNhMS7+TsjjtAo2DnRMbsMWFnObQ6Flm8ca6UGVD0Q2boCkw2IGdMv+s4UU9uk3YzzHVHJ9Sks+UQ/ppbxtdsZycRXNdS8IS9ffYwEai1k9pKPGbMeoGZsx6PFIiPy0PVHAZ5YhxzAeM9z0dbCQ4DZlWacOSzi4OBkrBVK3A4Q/mngWX9XuXgh6NbVJkfSYgJbh22J33OLJxD8nWsUt6d7Ix4fMpEPV4mQpKleGEusvDe7NlmUf7XfSbzukbKFJJ9VLcCEu+yG7cKNIU2jBLHZyAWvMC9ATrPHGst/s7cYGt0CwScnbGgYOlmHrDhewapD/54m3Y2xgeQXaGd3kkK/O0c8zdN1IinmK/iQRERQJPjpY29JwU4kG63UT4yFPcy/cuh9JI2joOCHFpQ/iDxOP8G6OMZ+3KqFahsLWz8Aj/HN6poqAxpm2S4KttFaJDCme2JQJ37Ghf5t1kHRe3pyUW3/saG29bDqXl53AeLqmsnZPn/qh08fiXG6iPJgmrvjuoOJeH7yXT2mDQj7uZwRpywpbyZzamjLcRub60sU3z7xSfLWEF3GdeGMhtrH5Ldqga8fWO5YYudPsiggW3513sBc+oWDlZVRlj7NfIS44K6DOpd4T1nwSqoGq19XUJPg+ycdrJNZG0H7gzIO7g3xpOBnbyCxEUlXzea0++GQprFiy+PCD50YqfMYuLo5H0p4JIAir31G2HDZRTO4jQiheMfR6bBxc9JiGF3PAIhd7tlZGbSaNtDvfhHsDRZsWafCSiukO2TlIEtBXELQH7Wds5YPt1iym3+lEen0f7aRj5UeusTkUF1cU6yemen8y1RGZ5q2nPX09kSeV13MWcOa+3nb1OPTYqx5xRZ+ZhH+rP04MDthFH+V5ThRo21SWGCvWUrbmOGdC403WjP4Hvmx/gXXofh/gFcw+ifAN32jm3N8kA9eVDVgPIh/lcTrL1o5lRWMsggGFb1uAL02OSriIiLxqdygfiymu9/3sbCdHOkqiaBlCIIEcFLSoUDjYuZyIayPAQeTzaWlwMCIveIGB+mgr+Zq+SR3XRqhFQOzZjMpto0MofMeKQxgzq83/6hWW0DVIHdC/fvxJG/ETApBMrmBgz+rBe7OmdvqdAyQT9bsgzWJyc8cqii24D10BFtwZT/RtaNaafK7pUo9hDv/hFJ0XgHqCvq7Pwb6OpIe4GgeXRCzKHLmCfQJwv5XMc/ZST+6oGJD9g9bSzd/4Ql1TnEV6hjGKug1u5Q3UPcJ1yb/MMmbB+qbmaW9vzH/cpqWfz/Z7pU0jEmq1RhhowT2vRd0Gby8+1A3YicwrHzQs9ecwtYbjLJiWFYbuKwZ7EFOARbcg8nXe1t4AbmASJe/3PieTxO8J/t9HZfErBTEpdy13Zbulu2O7vswrjjaQW3N8atWDKyqXto5HL9xVQr/U/F13CTGvciQLVu35xtLgq5FQQwU5doFE8Yh/LB9/mKd70zXdrtWtc1CsrElMwsQI7HtfpajCeEeKTO40gZD+aFsPmP56EbwXv0TqIZLwM21+xDzvxvvf4VS3m2rUxUI/qxs4ae4L9lWTOPxmV1FH9W6MkiMCXVkBxMq1b+tfdJy6hF6GsjqLZwQ7UlFK6NkfzyR7vlbdb6qi4avm4xEdodGJZt4HV4ssq9FXbsXLrN1HV7UWAJhQom3JvIi8K6upHlWYsEkU5Q8D3UEyxCh5YT8ktt0/e/KKxIsWeYgp8NRr3ZAWymZ3ohNhJHn7+ggW5LL4iVNzkmCGbeJn/XFbyc/DAwhZq6SMNtykPDHthCOK/l50LLExDhxDyVw/oQX9Bhsuh/2W6UYpnSvIKth21vVS3dP1SmLf9nllwKUbBZItv1SCjiC3lSQmQT4cojw3q6fQWL7Z3bjiy2mnCMlZd1uEOd9O6SdryOpH4e+Va2giTxhCUZzGVlIpP+DMdmyys6gxryAz8A1HMWGAI4leR37FUHAox2JiErGc2u3UOxme8Odsrez8OYvOridHxgZZ6eoymZAqh0hfAxAqL+Ll5MEcuxds72aK7Ucl1aO1uW2LwMVIeyGwRVqNtDxUJcPZ8QBpGPoK1Vg2dw87nkOCYBO+nDshAUvMkGcKn+P1Glcz5hjd5glIR6M9clpXvYcpiXdYEP6+R9Cuq0d9NIx5DyZ/tLWjQBsCweALhcsOnRE0VzMNd6bVmJENquoSh/k5RPaA2zFqhfwoMyYxRVqm6MVTaeZWldDnWABUgr65ncIURtT3sXBqz775QZwP3ExY3cL4JezilhDbmyudjsgt3SQTchXe0DW4ARl10xhfBp0LRbR+VCROUGogJpsrFoEDG8u6sKTWZd5fa4ajO522N6lDQg3xKpPrWCWCJ141czMG4l8TWz4NnC9M1cqT97+FBq3Ten7Dk6X2bJZqFEcbj9fYwHa5HoylZHNB55EUPv4xij5RQ1IkSvFUE+bGBzNDmSPGe9JSfhIiNK2wQYIHvYDkdS28vMQHaW/cDgoSaoVgETL0sm7/a498gZbyENS6xMeDqcUKOnfapit1+48EISCoz4QtiVfN5W3I2Z+SS05WmR4zUbDr4CYL4hEWb/InqT8Wan2rItSRpsoxpi0xeFlW3zaJnkIGmf/iATAWJdKyyoP40sEW1t/rax1keL/t5yDM8tWvgridi05A85z3G3Rc1TrdRhTGS+TKwFtwhsPk2YrSOK2u0NXZh6wU96pcokJwYM8FA9kycRmGtBbtT9VWE25exP6OP04mHxh8FyOETpB5fecVepgTi1LebLjD/fZVDD7HuZWxn6NfVv8k0QuOyHAjGtEV4FSmaBG+irLGTRfAOyXT9hi2BXby94aCQel6149JMaHiCrqXkJhfGCz4P1zsOTQHyLxIJIAxPcUQNH0GjIGlMo8C2vZLmbzwYKKvR5dILm0DIcT5+Fz2UIsHInCjo0MWE2kz+Kqq5fDrRfqzQe6qtNENKmkTnMBJwxbonMUsJjaOfs34/vnTmqPwp1+c/Ks4JiTIZLOXC3Q1x3E1Zl8t71MaHB0yFV+HcDZ3jGDUsz6VxKYGWk6hf4EwwwAGDz/PA4XDP0UeicpAZk1J0vXTGWj64aXnpxO8HaibmMpw2vyjng0L6lFCiLhIpI8E0CYxBqeHyUGul2b72LasBIxSTUAcOWOGMb3q8t0YoElyz2vXmxMYmqIj9jELJWXx1juJDiqTkTOj4YMjGSU4jk4H/CDkoKnsokxQ76YgcCellI6LRvozZL/dow4u3dLyXKUFTizuuRb2HD8MM++hrMTukQQq99Lb94Qv+s+W7dBN9AbTaGXpnlyukT3OaL0urnerArkOlBhtwrmJbejttjosa0RInqxo1u5P6tV+SAo1IyWQxW4uhQOdKLl1rcwP5wnfILMVptwhXtOvaSu5AJklvwL4JByWJl0CtNjyaVnZk8SVVKHy/Md7iqVvMotTP+yJiPR19e+jU9df6HLMXOcPZn+ub97VpvKFQn7CZZXEhDSivXxf9Ay3kpu7j/+5asEm0Fg1Z/T9qZxA1lrYGoFnfQ/fYSx3Jl4gFnB/DduBzFSaPE9b3ReiIndkwxY4RHwUTd3WBpbc1VbkVuoZ9QcFp7b1eZwWkPNhzrLV7gn6zanAymp9OyyBtrFrH+5298wruw+W4r+fd0JbA7lLP13j6vGBF7LOQRsIxH0fiRK9ldoTB9kLTs1ORswV6ncgZqegGlPb36fDH6FaA2z28d9IMMubn+rj7iG0VkTnUrPYYJ6JgJepugD0sCAtZm/k7DIq7cX+4doL6OCIb979CG+j3Ntm0r/nStTBFD9aHEtmViOmoGzvWtBXoxzzwQb4m1K/LPcGbajGdeYxNdLoRJxHWfR4GW+duf5EzQ4rWbpXWy029IDel3paGn9NfQao5WCHurXaxYx7TiBEBxMPQJMUpLefYX75+0WzD8uQ+fpKiX+mO0di9lR1JVyXNMLQOpIIRcU4tw7+05hiGYl2H5jSVaCzqv6I4EZevTGp82KTFLZIlly6rkB1duxbsvbrk8qtiOEbJePi86Fo6J3afICinRKaDAYjQPfcWtotEftIL/FWDmgpRe99wNudIxNt3QDNqcFjmc86lYijpwgzwiI5FVu4ElILe6SXj8tqNoNFBgWgqYzvPeZycPZpjTHzmB9Rr3v2DoJcPTj9114ttHPdpkvWWj+ILNLQwsfaocLwCqSMPlbshqYn4E3100fCs3Ybr2IB0rbIItlQJkHUwiMr7ybreyvgohYSuloT6N0iJQsUief2Jt/Ou7QXAPyxAdkwnX20Jl7Y7HxkV9vRTDzFBdElHc339qFtNKhdpwSAKwzwRH+LjtV4cjXSoqB4ISlYd3w9RNW+YvhNjhIt6+cfuMxgI4omjc4f+M2K1Q+g5w+Q0zbw0YJFE+8CkCEguz3h/hDTxBcmpYFmuwLhgI0JLx1IlxkAE5TMk9TboEOfEbeZWiKq4KHr43YdN4Y9blXqaYbHNECvVPoNmbNWkqAretjs5EREf9A4eqRSRnl+2u3Taz7/npFwSEHYUOEmtmOcpCrVkUIeCH0/sMReBn5Oc+gWHYcaUeYEeuocK1pX/XXc6D5cqWypGRPtkBCqOx7Tzp6KXiiM6/GwlCLD5gAT47CaxvCHPhVw4q9pk/rVshHkeZuQUiPYGYDQQBziSXlrNQfgMPFYdTLXabCfuydLO2hEjbeQePu242mczjWsvwS2e8uc2oFBOFXvLBjyj45fo8ZB/VMiQGPk+y0SLLj4mrKuknc8lPy42W0mlDzQUUHLN/LmlvIvC5ByCr5mrbyOmpemLERGm8ZSUVbA5JtDiwxjXrix74+DUj5ykDQcGpPoORsUL4xUOppeIfi1WfJaAUI6vABsTCBmMLLtE3EtKhtMIoLrZkP7eI7445fEAMYFb7knFJ+ceFkJTsUCAH1bNPMe5kdkFeAFkmKyiQsNM3ru2oJoWNH8qDPfcEtRkN3RjlSsw8VR5a+2s+aAZDOOrcYdTyXWD9XkVOjApDSJMQhCq0BUBIGNtljeXmH4wewA5rxENrzZvm7GG32ZD65BbLsctyASR2kIbEqQLpbQZ1v3pitG9Nfoaq2Seemp9/T9dt1NLQvD1UyUv8A43PacOYguACYzpOMm56VF5Bpdc3proMVVc+ZXp0dk/XLIJoVVh8Cl1jWZz0uvsu04uQVtkItT1aiM10iujvrh1FCOxaaZCZyRn4WNpxUFESrMGnTgroSfCRLOCYasfOGSz22931rU21Tn4sCobefZQEW9Dp3yV8HcseB1pdTZqKSgQ+r9uzZdIt6I2E0JbQVSKkW/pCv+GSShqzdoFnzOG+4E0MlD3dDrbInFjSvh9SAtUGGQpfrVg1uZPVwv/7h+hFcWZasq6Jz7hCunFIDi4tgWWnmKxsbu64yKk/+DhLOkcPi/G2MJ+K0Ndd5LMnlBxRmbFX4OdGJOoBOUR1U1cdMtD5S/CffT2gVNUC525JuE57uto0n0UwY5JtZUSLsI4QVhvP8jeJrHitKeJrX8v5bqnr80QAJ7gsupTxGK1m23xqBRNKfWlDCkU/D6W4J30KDlkQxjybav7FKIaxGU6NPh042M39oC2X06mN6BISE4JCno8lLRHKf56bY6Hm3HOL+NMQMTJGOPR0UTjVbZrPCgLF9CW/gS9Q89736C2febHUS36TujzAA/G6wgKNlB6Lcektva2/VoSCJUiAgk+oCyYQGdGPE90oKewEBV1mMNGSNjlSlfHNLURGz74wwbfBftxtcBSK+RKcHqvgvC1VCvAo201tG6ezQpfhQxiEJdYciEywM3IOsNLOxUqzBGRoWVR/oK5A9TH/CYrsCbwBUxF8s+P0ri9itknFMQi6++Nl5crucy3nhxo9J+bVvB9GAIkS8Dhz9ibfcgiyZVqEpRy2vtFLEvmAahZRp4NRnRAAEzq6wvJiHNFCzY46JYmcjCP4xACANlXrn/ISrkF9rCv5oukIBfLEx4F2+1D0x8pwZpCSZ8XPXjETDMYK3UTtDacMKUzceVnSpWa+poJDugJI7NWU6UwS1xeW4T3Fy33Cnm+P5X7nUuuOB31Hq0Lj3Mq2unMfgXZKNzziGdx0GPXFjWA92Vr3cSSmkLun1glvqRru88e13vCWC/tvVom0aefINSPVZzqWJ3NKu1vaxpI0Welvc3BpxPCdVf7/fcaAP6j1/g5IRTazTN9tw6jRqIXt6WHgnfN1atY+iyb2MFqNA2fg2JPcd+FOnYNERJQ6Y3AkzzcR2eyGcamK7Zp5NbyD52Wh56cdOpoHAoFTUHue+uTq6Iyigu2Mw9WyeS6Nt/hrPo9ZRT7BKGRdEocLIt9S5zaIhOmzpqXEKA8NWf7GWgghq68bpExPHT+ziMxT4VKIJyDkDsIi7Ewk9y50ee3jRhGsQRNzrkAwUGzAeuIgHo1sYSitrpzjq+DZ3OmZp6it0VRL3ItXgJUm69N5+ok7/ss+9Rk/C6ZcZWeZ9QKy2sDNBagbjWEIsVrjcxx2SFHoE/QUG7br5r1yXQKE9VhOkotgv4PZ5fEHqmyWkisPe45gc+1ERtiWOtJM8b3GCGnelEfgslWPBvyf2lP1cIjf0Hm+pAWG9wDsNxv/p3M547+sAlQEVGFktLyBHRpE5qTkFHgZWKSYcfgph9kfuRsjaUTAKqk+Zvq9VZTGoICi6b6dBWyzALzqXufv3madapLR6ZUz4emeXfDWvViZ2xcf1LTQFKXK2SBLQ/k6jW5Tu3MxFC88ZiRi79CAwLPLfvkRQW913O6iSbbr4ZwdaGvkd+82wLiqJ8eqK6NiIfJ6hQpyRbeJDtfOjbT/QLV13mj/Xh9Jxiom9W3K+ZLKuyz9RvQ4QSmrknSAHN0XIwuARFQDq7mWoxZobvGKVTAQoWlVLDNYfxPVwH9hgA7hJDPBfDH4pxEvDjYnKTYbHXjVMlqGsvvPC/wfkeNldOffOQk2e1m+RhPw/26M0ZzDuNqhpz39fRro8aKoNVkirZHnT2vyPfWvQx/GLqfCuTing5bBPr2ExvADSZTWWvIDnn2iSpiJrvaW1xIMrs1GrNAaEzXkrXxvUAdiRHuhy+q33FFp1wb54utZeSfLitrR60npFOg3YHp5L4u8lEJF9bu5w8gA+J0DXKxOIYQqAoN4WPIGGlX9QqXUZ2M9gh6iHG7SrLfLcIm3GyXxHITyw+2/8SmA/mKJslv3TQDLxdjdzKHhk3DuyQKh0ZAd4gfZwisrVs8Y+tO6jpR0XnkUD53Eo9eUoydRGC16Z/CwfdwVcCmRwN15lxTE+j+dg9HSsyL2BYnyBWoLkyTCbT7JRu4Te00hCMc0z4HkXf8H+hS3eqEoe67ypJJrdCTC3Kze/9BWKQeacjl1JN0zcu45I+oj0KskFsU/O5MEMTuFgPSHNXJjpMVeATcNRL0SdpQVyN8w9X6BKyqAGqu6TO7koshvuit4zsncrHo9D28YsKp0KxxTqKFG9o/cC2pEXo+MkNi+Ow5t6zdZtAJYrVOap7G1F7QxxrebXt0Px3HpU8jkf0UDSr/OQNvG0AskcFqFB+8x4D+Lmcwuu30kgmxrCKC145POWN2Mb45/bbyups7yZVwbaHVTtc+FREw4705Eod0i2WsdmqI7nvFP2xriILpT4c4uO36jEBtKljKXuvUqeLX3TdYggvv/cULa1FP1vXLsJgdoo1a7jNWIzvUQ5QGDyWCN0I5ckrdoLpU0Od9gRqPb02+h0m3RzvzHmnvTw8w5Mz7UuulMLAWo65rOhdBBBXBd/BwUYpOgPyz4vvDUfSPuwh/nX/FUbrGsiylSHUZ6mzexXFpr1/bbyW6N3GL0sZ9Ktera6aC701cVt12yvbGYxTG/peXg8uqesnjESiZPHQ2zT7cS2euDFkKnJ5pYwwDi6BlAY2YgGoVTY2JNGzKRCOQKcr5CcKnMflwTaN/glI8QMBYq12iUwTMooKmZNfMXb4z4/dfGNtT9n1B7Z/t+xZy+f5pUfp5Mp8F6n8qayCGpVEpRQC20v9LFcv83Np58k9W9yWtiSS27+s8Y54IKH6caQS1nlylADIRZ00hjMcSbYaYdv3EQKLM39YAHoxz892ZfMtTnOI7wTPnuAYLa4EqKEPpeccAbvAgqsY+BM8cJpjU99f74/qX3v6fsSVkRzeCJJDb0BvVAlG4KquneYxMF4GEAUwtUSIOPjcI1xsaQUQXkz/qfhd86+W0uI95aI4FboK9L6El7Fi/gP3pE6d1CMnw8S0ZhK3J58oyLWsKBMMCYqmFsQMdOQeKvEd8A+D/pJY+fV/8WHqGtCez2jQXCyU5+Bg/bvw9Q8ahmCNEK/UsWUgfSAXpPqfWa+uaoo/24oPiejeOkKxljIXfiTQsScyvKkrEL4CYKhHmV+Xx7wnD55tHu/8EmdmasFq5NsbEayTGNB5YNlqtDV/R1BGwxPiYGCNZVqupD8vxuQHS3mLYX7B9t90nlUUQnlUrI6LIVWjAkK44yfYLpNLlvYOBEjUQPZ00kQE9Cb0PL8wBnX+21Ahvq1Di4Ei5ve6WhcHWWCsreBvXZqV87laLMBKzs1HGkz1Smw5Yz9t9ACQfYExcuXIhUaFiPfm8Dfu50HI6Cd6TXGqfUmWSj39yDyTc6QE/GjcBoWn4nV4A/1YMZp8KayFiQJEV0sRGFG44fBJwUWxkUAyXnHc+vFDm6xu1M/TIbOC84CRSYryytBY1LXYnDwH9DGdeI1t4Zm5xciqbeaeV4BtaVEDN1pBRCkbWBaV+J4C7nAiZMWh6vVXq3RNFtq15SNS90AeTPQrM0ZHv1X5Wmu6UIdIjTaMw+ttLO2nZ7F8+r54oL7Yh1br1b2Qhi1vFFGvFIPsumHGuY57j6oZuowN2KYauCqPOenIUMaHf6itc0ag2GtWm9eoTsMnTYJxG/SC5JeYy8t/iyJu7CLib+6HAG/3sIBDmY+tGaW9yeTphPfG5ArkvzMZiSqUSLXsg9QQfF7eQLw8TbgpRmjn0slZGQKrNlRRLZolX0tr9pkw7b4d7GvH5qjFfr3XRbpSRqkwCtElKj/Rvsq4s1CaZDQmb52inGuSnZsNtdV1MvOVJ0iBS3DpO16ekWJBi625BnjZsMiX5QuF/v8iQ69AbTrPqqEMahnftDAbOjXjWXipf8TwYXHxqYBUNqJZXPUknOU0EswrC7iuYH3jnCUdKG9agXhFesK6ZpKdb73rxNR5opJnRJRagWv7VRc4xVZYa7F6SP3IOypmH5uD1LqM7lqPXxJRO854GR59Doh6fdKesblyHJXD1Aptlu0aMiW5rk1UfQh203I9QjSPrliZZTmFepsFFDUXJZvu/k27j2RNHp7b8IPiUoF2KiOVLMAX2foZVTQZ3KXl2AysL1fYu5LCRNJ34pow92avswfXjTVrWMsoiGk+1AznMUfq2kMb1+2IxY8CD7fo08p08KJ7Fgg+XiG7BNayMZUFT1LHsUmUx/8yhu83+W7SUgYQWrx8/2mqYWRCoxeaMKrILxZ2lg4WCosNoQmzrapSGMcbRdbTdzfyQIeqMuZyKIKeNpQe8aqhwOYsm+bJWV2J0p+EJJEmUHz8XIbh4oC98ZGerWjTAvfqeliUACtUGVeOae/oEQ8K6TIRGqJGYUr1vm4gxnaJcC2j0TGWlfSaFa1C0rO4045yNz2sVujw2B+uAEbeOgeorLoTwergXcEkftOAbj5PVP2OhKzDeYmImwj5lY5hDF6KWQvBoSADrZKic8eFMhvoxHyWSp784zbBDHWhNnHh1eaJNbe065hI1Spqwj2ScZIHyS4oSCgoRS1aS4i8fc/bRUQX3C2U14DY5XuWO/TLYr+6LkFFwI1GV1bmkj2JXafBcE+q20Em+DjpCmDwApBp8LhyEpCttr8w7CVBz29rI1FzVeluu5Yh06vHrWyYotAtI7yDb9pz4Pr/Gyd1K6JFnyjBQ34yF7cp+TlRUvWvuYVhiA6mfiX4frxfIyHntACSLeAYant1STtqOK1FcckDt5boOO0OqO5Dt7sATq8MMmlweA2BgG44HBIAXKcBhAaEoFuJ79b8nmaVbOq3oEl0SD/5husq8cIp+EAaiSHvX5RRTYL3TiTrfoDNHGY/SF39S9d0A+TOsQExD3WIXxAEESdYvgEyV0HYKgJhT+Q5vUU+hDgJLhvOGZ/g64UBpZUuyzEkXYBAyxZT40U4fbljqkq7ML9r1NqOXHGZhF8xrRvnWuNVpIAbFTOBcmfuUlm9sNSXSCz2RJ7/XzeUZO9DmTUPXgOO+FmHovKjlmUeIxavDfBhtRYrC+MWoi9K4umsvwYJAS9BumuUd1jUPlBXqRpg7pPv3benhkjcf6X+Xye5+6rsE0kKPd5smBV+Lwuvlubwo1bcw8HAlB+dmoWE9/fgW9V3nx5TPeuNlh0a2jwHpQyYVAFmOp4GpgZu7se4owXOXnhyyVJ+jSQ3MLaiJ9qEu5Z1VFkV4iw8bWcgBYedqJDI9YjaMqDOqCRYsKstANX3lkPzK7OyKS3TCDkKkdAM1IQD7ZEoC2Ns+v2NMJX66NBkQ6Xff4cxMpkKCUg9j6f6JtkEnhOv7j0d4aaCthmfj3N17CQPCGF7eovhYFvypkx0wQCjC27rB5q4Cp6I1MSsH9Ru/G+QRvT02k3UXilhxs00KA+h1JQCZeRjTHWcrF+Wyqdx16bcrsnb2DB1TbBS+FUm72iHm0BIy2je/cphK9n/UuhJzlYMyNYpAW1ZPD+l15ipuoM4iCQPM2r2p64JKydfejCwk2iOZa8fXdAG/BC258XUZDw7UBUMArGrXzaxC3NorxX45wIyy+XZW3IaihNZ+RiEAfId6wFNJAR1wYPCBiMyCyEJXTh1gclIPtN4lktCJjnkWYy8GNe+8uQR08K+U3uGxAqstzyyDmjqrV8XCCGGu2UdVr2uayFPI2dyj9AS0IpEBZbFTQnJYKsc8bN6dEuO87e0nO8DOXbbv8MxFAa2HuHJxfREprlj/P+UEj8gBVfcbs1PeCjIraICaMypiKbtQjxO1N4NWpuOuKmHH8DbRlyh8jxhCi3DBNmbORhR6AjmLh109jbi1Nbr1fJrQSYbzoPZmwOCF6FS08rQcEO6b9RCKYJcuMbonIU0zzvKbVWXftn66cCfZdu69bm+hdaBCPSPlcrDAR1Zuq8gQC5v+l9kJaCjRA3RRwHw7ijAWx9C/RNbgVB3LIKsWflwNIynBYfdkCKSeSLKkBOJw6hfCLTBHminTkpqNYymJv9hZWxXQm3iBqPauVEGxSY0w4f0vmUIHK9j0pnkKyXX3ssA9uOrHHthHN8+s012VzRnyWYI63BrNMaSx0u69H13CEe43uYyN2yGElqvS/VAI0PbmqMc1ALOIvLSKmqry1tobBERdm/8R6to21hzYgj47buD2BXgjXywO21ReKg741P9M5To4JYTFYzzbwf4c2LAfgn0wFyjrLv9yMqN9EnnPT0JuCZzxaZM4ieOnY6TXMA5Ju4MPKNshL1zaRe6llG5XbaEn4g8iYnvDX1Wmyi0+kuRggXuZs8T763anLAkfhEBL8d3es6QTRjsUwVNcrFplCyRp7xvMUH8gJ5PIuggO+s4dCg4MUed+Cp0WiDZhbSi5lXpvecYEqYLKTsxS43kODXlgZ8f5KtrSt3U3hxPq10O1oafOQ4Pbpfe6wVxDvTE3gQwzJxOkGXzhQKjXh4Z3FO3bfXsgoVnqP4NKeCAqvgk7ke7CGQchishRdFP/0OhEzNMz1joiqxZx6NdPis/yjVYd8HmMH2JfeWmGg5JjBRzY4zSgWjfoXH7aQTXTtCI1SbMUcG/+unsQZbHJGGXFBCWH8yZOrt6MtSnIGDxk/yVAg8uTUi0F0pFFgAJgYP+FTF8DIxAhgrQDoP+qV9qFuSAzpxxVZGlAjCTPuGLJUrULHkLeirv7f5IwLKtGvcfUkDlzsgmbJyhJkhr4FT55yYC6ER4ebOZ4P2jkuZsLFSMSHdKuDePmO5Kvl+5qg8xPya63tBFcaWniqxxRlFEjLWf2LqhPLbVGnfFIzQd7u1iJfgH9PwnuCYbRofzvwBCPSaQh27TNqNzIKrSyZdA+cH92OX8HGKzkcupM4M+BV1xRfDp1rWVhI1jqykfZX7Qw3IGAgqHHS030myYxDNGxzMwO+YZZspOK7akvd+N+7UIvlK5VN5hA7FFTAJw+X9y+sKtXRO/tMbBTJp5/wZRV8QOk8Rp7lHN0xyKcFGkj2lTaXIxK7KsCnVvTECYl5BhG9JGLFs17SaU2XyxCMXBweifqyXACfroKbfQXVryJydhumOeAMF5gNR6DiU3BNqp6KqIWs/PzfFPpAFzQOF3LQSIoW+GVqI1OcBqO5ZjB71GSlHuXPTVJSfb29ODDTZIlH+Zd+EBRlj9k5lsf7Z7XpftUEUHG6jGmZrd7iNghS15QjMudsBkLrWriLXaoCC+l0cvaA8nohCGOpPfdrSSAyV7OTe9d3JHSLel3Cx2Cf4cpKEXIZRIxIk8L0u/oBriCorRx4HytGSIB95KbVrI53GlMPKYlDChqPTF0CtatO7JyVRxl3PhZAT5tYp2v8cf/Q4jvtL9ny5PLnjsfzasiB74LU69sQFQ7iMZ5myA7zir0Z041kEt/B4ggHil3p6ZzwSPobDSB7QaHSQpDb44AqwyvfFOyjOJeM9C6tKJ8t3Cfr5zdggtcuZWbUoLxHfbGWhWJbIjBQcV56+zAhVpIwBvbkm8SlVOcpAdJ43Ht0+CYWQ2yMJvazH2zVEdinOxFaujTOzHCrgFCjSUb5SLcFaG5CromAow7Rhihdie9ysLChaRDryn4XJeGe7PzqgRfOe8hMhQi5t6w0ikm82zQo4Zy5hkTqcOhmuO8zTSTeZFy9hGj7wsFxYhWN9K7IJT13tIr0O0+o9x5VOR09iahrF/OGGXc9hOaSmhsD0kYlBhujbXxd+FV1fJuZ/hpSF0RrB6qhLWKjau6/eL6/svOUFDQMCGeWFh5yD+w6w1VSmNPUXMcIdlgnsQkGuNajUL9trgLoyZ/TpWkaNvvi1L18TQ9baRqeIVz0p1LzbN2wgp+nmaqTNVxAPeQy1BWw6asMT+82+cdvwLJFwBnV32KFBWaiRcvAwVC5Jry46zLn47FUE7NnrtOSbGMH6Xey6IUJOv8/3GKhilr2XlzD5LQXr6ZyC//fd7Q1IUSNL6P8b5tPOpjbaskr81EN4HdhAA+y9b4hFgJhyaqULG6uxbYtVzzXJ8jtF4o3qV9tuyQNa5OdVSxbJyVjRKWIyVVVNkvxfv7xAzASiRquFCEX//vDbOIFpMNxyqpCeNBu+EtOic+CDV7qb6gpVLrSbtYzpCD3F8jxnYjnb85Qz1vlQtINVdWwtChyJNWjb5yc+T5Wz4botnIgx4JoGyXR8JKauK6/UCfz9T2ePQsr/Ej72n8IHD0DQ+f+Y1t62zuVFhI+CnG7sb6M2i0g2Y/ZaDFPbpgMUqSqxtQnUz+I5xaSo8Z6E4JvuRW26w2MHXMylIwT7wlhDUBuQNoNSavVKPb+76kgQg6qAZiyakgo6jqb7S9NAQ3sb2piRuM2dtyraH4Q7i7ryXLPF9+L6gcgoCqfN/1pLlbclsd/qQk1hAZmxzOcT+OnNaKuDPXbl6qOpkPHu+fcilIlX1NGi39idqNWqBUSlp0O6srjmnun1olTQh5a7Il/2YWOnqJkC0yWBRE6sPXIBiG9ev7M12y0yPPAS12UncX8klZXpwoklJxaC11KsN7IS0mwf6Yy8X7vA9rTAFxOiKAh45D7luN7FEHkKkSNbGXAosgPqiwP3sClqt0G+TRC1cl/XKyBw8WFaHtg9EJzRZFMw3LHs3qrDm5gHl4V/lIPsOq2Oq72iLhpJE639M9BMRw7ZwkulsggNKFw2YKJYPZqGXDNP7xeh2c147o1MOG2HIGfBBsYnZDawSCM/rRQds0DKYlcb+O3+zzPmScFj+KoZpqCr5DBDFXGnjHqn+PgSSccxeUJSbYdnQR/ThWck8re/3TlEBiXLRSttToW5BofKk+38ecJ12m6WYEiH4jF3esacMEJVIJ+wK9S55iRBkI8NT0z8Qx8pVomrwk+hJuK5PqOLPocvTFAaPQ0MH/lzk0eCivRf+Xya/8YqQJH79rJNNFQorqZgCraVmZi6B463vw4tUgQuhVLoMjBshGaZgyHEUCHfGXCB5DaLFSSrxQvUVorPkbl7biA/jDQLh6crrSDq+lDJww7waqKpq7HEy8i431H2AKJIiH49V0W1apCuvBXW2INUeTpzVEbgQKjts+j3TG/DHP9CMNhopemPo4wi0EO7NDuOuh0WQV7SnxpvntuO0TrnW8fg6plvULjr4QUqeT9KenZp+lTVTRsgNBIRZ9A9lu3wz0luNQcrJo/9yax+kuy/ujVTTf8DkxgL7Lv3EcpO+QvXA8wrUS6a3E9pkL2JxsNPpjDqtBv+0E9mZ/NZbb1MYjc2wVxBbLau530bBGHc8wSWnmOqxLq9mW64xPybcJd8DKL+e2di8qdlBFnixrtRtk4eYcDNZTM2hf7h7UP8njg179n3mUHBPbs4MMLNllykb3ixVAk3oBJwxMdj+UI0JRyxaMXxhbU5yyRh/fI9bk0r1xZVPqsyk7xGfeosDLTncutpCbE1qGX5OgVT9R3Wa/d21fEuY7GCuML+aLyxuRPh68aplo9dQY/ZGXxbrBTIjsY8bS1mLAaVbT2486zfRTuI5TpcY9JFl+aYrjmOU8hE7BE1++VBt9yDFienLLj0JC6xXne+ZmF2QzuPkyJ2BaD1qAGBkjqTCVGftxQ8BD5m2d8+7/w8mCAGoh3BYfs2vvJ7An9B3PJntkwBNKv7N/Yx454JzJNRvBLNo2vPwgDDcetIy45HK103Ak7YY9k0chfnE9KXnYnrIY97x4t4s4LpAloZ3XZ4dLaFytHWe/QD6Gx/VFnwwJlJ1SOlJk4HNDGFs5lwhaWulki9Vg07qWtRrWRIxFaefZeNk5BTP6iyrdE8wn/6nxDD1w4ihzWHih8J49ECw3jVzAp2/Xkg9ejT/c1vxne64BlGxD084YRLY7A7a4yjE4tARQmPtwdaM2XACVxjpLu/mkRRHg7KY4jc9XJYPZiWhwxWI3HxH4s1p/SAaDQO4jY8I91bD4aaXwIcDnMN9/iohUH2MofakG24pbpglZZHbsV5OxCxbXdfCLSMxH8oIUf/bXhTtJ0+lykKRXFH+yd3RPXLLO2YgZj16v9jNi7G/d0k+mkbKeM8a9mUhnOnS3kUXgDftKj4Uvx1F2IrQoiNkTE4F2IhllX2TqhTzewGn0sk7liR/yiAtbbJZIwk+9MmBaKYxezai6bdnUem0yoXHhAbWCyQeBTJ/CBWAO7qH7RpKgR8UBJ2rq2jDDGEInNsxK60mep1gJLVG61abWg2ngh079yrJHkhnBbE1GzqNyEEkX+5jYZYUwHoM8p+/YTZb4bDAoBgjBStEXx4eHsir6XilXGqAz9ZrmPb1pm2IFSGCIt0HZ4sy9B5L/RRsJ+18z9lpxpEi0kM6MsiMl+c4uQRmu+mJxPGUxSnyL2AfhEyUy7E0dmGchXgMfSAB9BMVCvA6z+SRDc4PU/BJS8ZCIn4r7iPq3BefSRnMkLO86dTJE4ZaW4E9X826l7Q3n/IuhqywIEy3a8Bb4Q5/MclnNQdAFQgEEqkwICUXreME2ljrMp5q4sGG+wvh1qFzTuU62VFOBJ5lH/poR2ZPmct5WijaXIxHYrnK5S/6rxQz8zAjmuR3Rnm+UWchmMrsue7Ur/yxZ7273Bd7k85acD6thlafPmJAY7uBW0CWHeuhXSBwMCp4KUlEoiJ58riWeyjvO8+Tb1oMcMhFvQSXeQ5+sedUougt37diOVIrPPSgU/teytNPQTSx/ibDXCnH0QYx+9tW0SlbT11XnTRnQGNhAb2+JpQJbRxZyjYMjYTWMY1FhibdJrQ2il5LuFiVhKvXldWQdodCfCD3RODDHWTRTysks0KfrpMHdTnW0ZdLjDbWJxlaXXlDOUL3zPRmm4kQryLIIpFMy+BgrX4CNloW89GffEOLKN8SY8dUVC+I6ff87/gBqxtr7TRzqx4eFHW/9Ou/dNIZvzgcLfwQkfivRqZBY6XOfuQYdOY7QFNdrPLVW5I//3CDaMJhS3X698j0SnnXrLLU8znS3hI0jMQQ2yRUB+z3/FRTze8ikkUj2nZilofmmT7C6DT3j1LMe7n8LpGGNJ82Kg/V9D1/Iuc5r2oyALEmltR9DlHQTcb2BUZ53YQ0ekK1eEmdTKmoM4kl2DwqsjS2KOkP7S8Vhl6BkSYYGbjBnoOQErwUEVOohrzkihtU/kKoNdO0KlW4pBgrFqz+UDVQpQMTQfaDHhgeegUsrnr/kV4jxlUSWso4k8Y6jnUL+QcfDLN0jkWkeo0ExFw1fuGFFUPjAEAdhNfrqu0S+2XDlaIGILMrKzEyLSJw6XGmTtSTqNPWWVdIKaUNaQVvACOnpKbSN31mEqf86dP+Szy5cecdzgs39nGDlUlN593fHiCJNMqhh00tFIGBOzDVwc5u9erq7U4KVLtI/qy7oZCz/MDynHGZ8Dl5gsgpoeMJedC6jZ4AJnaKR8Byf/6SITxhJCKQ/bnX7JAaHWG2gecIzIB4CEzpzYRfeEv0K2slxNyEaLmeDXXTyc38apPLVrHp+G+7ko=
`pragma protect end_data_block
`pragma protect digest_block
e3d32260ca6a582acb4c8240212b438b5dca2fff09e4856826e50094440d5981
`pragma protect end_digest_block
`pragma protect end_protected
