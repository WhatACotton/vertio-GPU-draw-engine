`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
tZfDNCqyangfbGpNwY89mQ9bEgkGDehYMHvhxl8YQgoF3Xl/Pr8A406USq2K1V/6Vx6AaIRXayq8w1uj6W6ecMBUbTzpvjbQ2k955sGixjoKQ2/j4DUGLDmDIfD2oeVI66gFsyENqWinl/vClOUuUgHBQnBbXxYBAIkmEYUyw+YiQmMTUg942e8L4uGcOz7sSR3h8taMzLQ5DCmsWOhJxtIK3laE1T9Z2kPzu/fyt4zfumWlgb7cKQ5aV0IKtWK5O1Vh9nTN6FvKVAWkJY9G0cTBMXiWgNDQgYNNVXMYBuTz7Hj8aUGKYNVrEj+Vqagt4QsO1mxfbX+SBXFiqqi5clXF6+pplo0EJHu2lsrZXRhsMoycEi209wyRfGSC2H2PQv+5CdibO+8tYjaualAP9apOx9qkZ4rwhNJftjoWYzb4Au4Tc0FuDy7R+0xiOrXy60JJXkxG/j+VC2oDmM4ugh0AFlFR4WMknXnqFss9dxRjNrWd9KRTkqDSoZ/FDokyLVopPwiBhkkbKWWniKEYhZYa2QqzI2dXTt5GYdrOLtbfxiDpf5IeRQ0e9TszxF5EcVdLTYWYg12unTTgAhI3YjWTS2p9KYjRm/mhdGe/Dye9opqcFGiUeZxJi2YKQVpIMI0n+1BMKFZELEpM9NfkRdjmB9BBKlNWXa91wMfY3dfzxR6/DFUWzFwUkUe8EDMBAJTIQUFAcmiEt0mdebojMSvginiEYo/t+r50WurxDn2SCmRq9ontnVAx5AFoC5VbMMV/pI2+PC3uoqLUB+8tz4RJJhKRo+B9RIPpV6CFilFfpZjpJQ6LVM/xrEGB0YK/krAMvNatMybKXKOVV3++ts2thZO3LLn+D2sZXNbKKCB1XGEYjiiKQTbw5LlG6f4m4mstoTiyphwm3Veot6rcxleKzsh8zXgJubKV2f8DcaYKs0Oebgs7Q5OgDNX4Qo02RMvEKAWRns9tPSjN/aJ0trSTvpQ2Hqa50QBz0V/Mvxb3c34BZBBwFTeOkmniReIv4eFRzVJ8r45aA1xmgEZenul8y+ZCNEUzkvTYk4nASWTvLASGCvWe+oN/RdmoBbiqgBZ/160WjduYhABxoSirtKdyioTgYa3c2cmXLMREQ3rB7zD0APKv0f7j1RTt22wNrLbNIkoX8Y9YJ0k01/G5wHbNjfxzoLAaKkkuyVDwlQRfgRnT5hqQmgyPC/sH8bE4he/7OuZLEV9sDRpIfBqtrcq1sVzcKEUoWYHj2aL1IN8LIJJe7FY5wdYUJKRzEElckYaL6DSIZswlXIDU61XE6jfwx3LGPLokgwrmmLcYJaW5n9BP3u8cFt9Rb9oGgZGQuSCXIbtT2rSyWAzzQpo2Ym0CI2M1ajMLZMaut1x5XDQO6pO1DdSZC/La4UirMw+rgJwETGSWxXakCjaweF552nd8wfuii2vgalh+K4oxAoaAj07u70k2yXxz5QI1IOnnwRWSaiR73dCpoHCTb5xO+ljIAgRkuIFwEhQ8apJXSRREl8IzHWa4r2tHqjbFfhhhCpKeokyKWXxCp4cpjAxO9EsTihP7XW7omWQznuoZ6RYkdqzlpUsXPLUzAWbZL8189vPELHHSesj/co4W7SAGvkbgzqbaKR1OjV8QXvceQcpUANuYeOOrQnDJNW5Buwm55/e5ohiuJW4L7TDR1TwfmVqWEuHxtz/DHK4ucPlt5CnHgCioX/DIiCDxH2dfO9YBNMy/G1WruA0lI5bdtcYwYcDQWZ4Iz3pXLGFsaIKuBXc9sPx+Y/OtxJTUo2NCD+dPsrsLw2sJsmG6/Qg9RB0h4kELWqqYI3S/3MEtQUMUS25gXG0AT00hYJXz4/kcpdjdELL4r6hmptyavSug+3uCidCBpEyjON5p6Cloge9r7mEvqeeKxm/22qqq7RMGfemfpJZEa/1iOUzL6XXgyBhFc8DxhNdAsBIHB7cIEIteNv6XXjTD/XNxEJuJI05rkv5P0rM70uCtEQEL6C9GcGpJDvQvVzT5kqm0SFEZVxL+5onDR2+xYzZpQ3k3EbKVXe/ib+LnFvwBZzm7auCVaf7x1QhdqaAGBziQW3fCWaoYOvwsfftxlyALj7jI7HpXNbYxb0wvpR2TgSorTB/F1aLAPDdWT8ry/WG4bN5p6+/5yiWfj7kfiBvm4AkAtQKkJFdOVRAgQg9AGI3nROJfnyw2w6Fbtb904JQ0kmzujtOR2Y21Kle9vATNbOP/jcS5jJT7cyZeEboaXNr7gYn7LZfJ8CqVxndL5inQTOKgBpCOfvAvk1jSWiS4i3rAN7iaSD/gMIKBFvOymEshP7gpxoajDFjg6SfmWkKq1dgNpkiqUszPn3UstFO2NK4A952xVq2NCBy21dyPPgOwpYwVwCmd76Guh53jybk2DURzHn/i9JKf+c9miOzuZXRqJW/YhrZHxejC23Hb76FIrJksxNzO7mxx44M8bt5dr7w6vm2theoJ553p4nnmpR5BTkaBeFPS5JP6mJQYC8zP7t0Ja7LYPjR3Nd+hVEfssCAFzldiFK3mxm3UqazS16+PARCpZRdtFJoaE6kkJh+2wVpX0nYIPOIq3wKD82zFGmfG45AqCwVleOlTqjKdegbi1jVqnwGk6bAcndt+oY0/5FAcR2mPwZTDphMVeMD5zkj+sBDpxQNKVBrGZdJAHBE7n9SR6Os+rcwaFxZjCW3jhToR0rs6HUKmFPVMYM7SRXbylMvXQjZOmADuLqYnCgc4neoGjQ4ly/rt6B3dMT7zACbPj0UWWt7NJ4u/o77e19QYXrm4RNH6Yxsj5VxpMKaZlzBzRcaWgOHS/22fsxDaXez2azNt2LTfE+boBGFyYsPLXqBhLYQFHsXI6uHrRwPwJCvDA1/k47XN05P9XuaMdphjqjELRytBq4ZyiJwPag7iTUbXJV5ff3VGsiEjG0YuYiIvP1hf+YjofHf6Bina4lE0mjIFpBNg8gOPRnp2/RtrCFlIKNH7U0nmi0tJhwcmbafDSfBkho5du1vwExPkiJI5PkZ62GkZwLcsmx50gq2Y8awBgS1EtoUH5J6d1zjQMvrxbp5gsZ4grHg+IHoLHrX3wVDayQRZe5TZVLN2ra/UJPUlA/DNaOLLfeTRW44DXXTR/PZwJoscCCKzHgBY0asqq/mJT64EQsOWPmwjyv/DN2/my9jQgsQKNhG4eR7LzD6QhPJyCR5IS7LEF2WeXdakBLFGX0B7RoWsr2xKZNAQolpfbWCgd83aA1x3oTlJr91YBoe7vKh8ZUJWCRuP0trle0huwmA82QQCUOVV2nE+gaHyfe6bAkOkrvqRwLE5vNI7C+NdOw76eZzqH6rr38fAFMKJarB8l5K573SsyFSbMrcY/fk6TFEJmB4gRBccbfPHEwJ17+sGVbn2PqKuBiMeoTDGM6K6nDtR1nwSVKwQXteGefoVGyb1vlCw7bvUWYx2jR+hWeAR7QaLv4LX3vWVYCrhiJSnUARDIpZRHlh3pLYLp6EJt1SMBeIinj4d9sMbLLCwdku2eww3O3qVxz8SPeMGLRMIOiKP5sFpp112ox2UuoUl2y8U9mJo6LoQ4p9BZUlLvJtGe5rM5NKV3R+4MbB/ITlv/0A6jsyR0l8yA6et8HtyyAd/ib5CM4uJ3zHG5MrHcKupGmOR06o1fO5p8IEcVrKPZGF3SuWwnMr6AXL/jGlICHAs49Qtzny5IjEQi9Kr8wQwmPfeaXrxZt6tXKdXEXPvddQYubqBus2Bc/WittPbCdSpsuTxPxjLc9vg6NW9Qc9mltXOdPtUleAUaDTu2Dq++kO3l/FsBEZeDvytjMR61OQIjJ/2xbSZNteHdprWF1Rn1ovA8aWYThK9QG+gyN83dH+FGtCJ3hRVBCKTEuOOUjvmUcSHWVZQphEpTR7jl4v5b6i7iDMNYa16xp+Y3kiZz9u8FtXThgUg0IFxj4tKtOYq2AHE0HNvVmxIqQWYqYSMtFKAkOY2cjkVg6AwGnPU7vShfiU4rYttNAtdapM62iQHT6eKfhDi4BUOPGconthuStkHuF9SliLzX7zQvgYSS5EYw8+/H/+/j9EgQaQSggzS0DDYKpLrt+vf9Da3XqOzLSIUpjC2MVF12U+C/9i/zzxqReQXYD+ftTlZtdySwzXny6ew0urxw0Mp/JQwuynwv4UDLegXEfFztTjVmITfE+kJj0+N0HECq7tPboWgfV5Z9Ka4rLjqBDyI+qQ53r3VqqVCktDCKoIV3SwJGQ8tjbkxYGqDWk7T03Y0xz6i4pZRW4scndRjkWYzutFpcapzJyrxZ/Kru1y5GThxeU7TIqiiDToBKgi/AXaqmfSM1VExqbPWBJ57eda2ODjYC40VwV1vw07AaMF5qOSWe+5hDmAxf3oe9QbCBc5HSd5xEHFeSxrSupke4Mrh6Z7M8mG52/jfsZHC7Xwnp5sG/H9tsYId3jAxQ9kaM9Vr2T7sJbMFPaCb20qdd+IPkzX1qM1TnVCoWCHEX79EzPOLLM3Pr8/ry4nI+3Ry7CjXzEA33gR7U+oj4PE8Yke/hU+4jZXPabtn0/l9iAdoYy9LqGNAX84CW/UllEGVOsGmc3roh+kTESEhM6kYeY4ud9qx0v5yq/9JY9NNFnH4GD2C5SWq5CXUkKcNWglNc2AVFk8ETUTQZUZoebDVChRr/puVRKVHIT9EwKFVx50wC7dyEmxJDCMyT986LXCSbB90cgpB1979E9S9m5wS0g00wBNn49f9vrKEmtsFK9cUx8hlSlwRubIDUNwPB+zm2paSVxZxQc8drwFNA62Pt/XJSWR811Yk3aMFYCGAHBKmo0PA1yo397psCmOqwRsYZlk9B7dnFVNLpDui8C5z3POYc3nMC66s0aofAnwORrgMalUhFE7Os/pHnnVeM5FP3HDuwMVeFJHWipX/b52AP/CgI/Xo6eY8OVtZRJvBvoPrNJ4nzNxsFbwGCjxtkcZhDyfMk+l4h0sXIDc0TMU3bi7JW54AC+WY4CG++U3HfLn4XmfQ0cmhCpCI3MBQ5MZ6XJ0YKUHW7SafIcUpkBHSXvJFo+fHlZBQkurIZ7fnpQnToNPTz4hmc5YDq209VIEQN2Nev0FTxj3ywMFD/4Bks0yoHm5u/YBBEFNCrA0p4xy8ue7KbR/27RqM4wXrE2EN1UjucjSdSIEopXU+cY8I8lwusm9n5wAV6u57bKwaXMDAG0ixm3OleAksS5TDY0BDn5DmzVR4x8A9sOWK2dbmjeDFqH2ZdjQJIPQSeLJwI/1N/aSBod/uQSN4NWGRVlCjSnMpZm7Dg0Uc7KNBqD9BKXsiwVjt1GivSOuwVOW1B+VT409OQj4uDQ+rrs8Y69EA44/1Rxho+YDGgr+EA0ABy2tDyv7DpwpI1fMJzDGG5rYMss+ANjyaV9yGkVDLotA8ievDgfG/6rCxD4y7EFiLhRE9qAM1X6eCUIFf29+U1quK9P3sAQgv4as3ht1T6DFcB5ryujhOnWvXfogrrAV0JLAJjtC5epehSsiSd/49OBbWkQ3NwMbg9Ev0VSvh6RBcEmoRXEyP5gEIblREq6glxn5kDeE9BV+9GkQ4v8QaRoCBh9cgNdXGJqrYuoAO7VyxvHyi3Ba/AOAflRmSbgl4OMuxqH8mbCrzbt3/OSaD6knwzLE69uFKThZgLiEoA7guGm2kqjLQxQRVIuwJWNWruO+lIgXHaBjNg3kCtYr7vVQg+3ace0FOvgRcSCaU6d1I/xpiLgFwa0irdlkwBqMnzBq2Xw0Fl9EMEuHVWJ90bRy3G9Ug4dO6C8Qmmo9GRMVl88U6UUMDpZ83MvpGtk+2+a0eXDUvb8supwMQrEN6uhMMGNB22LjskhipmQ+iHlVIkzU4opFEgh5BPFUF0iJiWWPKl4A2T8eESh8jXMuXdfJeZP69f3sTeDocWWNWlETocQBnkj9e6Jq9hXnYvWBr79OILnulPa5kEslaXoa8gFHURqmx8DN1ZGOh6q5hz8UXdT5s8G1UyZG/rasNcrESK9LQhrn1EPpr31z4GjZdgRyz30zWcwCKis9mwKSGcK7T0s8C2SlmbklQGjK79m52jrf6NuY2vywsC1/cW7QLzYEPeUfh5i2VV6JxiPcEBU0vkW5Sqt0V3D4zvvJgRP7ehffUGlJGzwPwGydUF4CetExMUPFSBAxS1qAhAQvyLGYw5hY9gcwG4yzZ8ooLvP4HWUfX2myzCM/5GBGTzpXdtf30srrd9bVlslVdfzvm9ocbpLw08L/3LoyHjiPxGWv4I/rDuQd2UXKU/aJeGc7gpUE1cWDYiiSCcxGcLfjAc8BIb2fViyy9xjPapryNY2YQ5laGYB4FTXyyX5k10EmIeq6vdtab6e8w22KeXpkmMQTNfr7njJGKCz9OXX1wKFYllglTyTQLIqKoJA2yahOVxYCUNevWewxd2NYWEK0ue/w1Al20/MbkcaKP9ebUTSrpw/7RUpaRRJwlL5ClPJogquPZWYnwCmiMPLjf/L8+tFfrFU+bN64fYWSZAhPQ4MLZtq0PQbli6Rc3tFTD4zecRxz87qI2dXjdgzQ3o8wnlBI8W/ILuSrnsK184/iqW3yPndpIVuslht6bJadlahiZbdzvK7l3XPZI2Gi9TYvMZhAwXL31YuBiyPp+7AF0HQyDGi4u0sT/q1LuQwVPm/h3CNkLEZMwneq9fb3D9glpvxqe7xO3iJDL86FmLoLy43CYHXtOShTVgVHrKhHrXlIXjQ+saJyHlC1cjCouINO5SIPDEIH9blB/2kpIJvMB1hBbTFi8TJfwQXXMWDpvyN2G5NVN3/x2Po15FzJ99UOn7U6fmD4PJ1p2rsqtU5kUje4xO9f4y705fQavGB7bvAhrRBXg6EQdeN2DsfD1WsCMoA2t7xVqwqtdi//DcuGV+ODbd2Zr4knO1viAlI2V07DK59gaVv7SgT99f+Z1krsfQzDavTMv66KnmRSuKtv7egI5xi7INB8W3sAULpNpjrS+/PRe6u8MVJt1E8FFjXdRgLih0HNof2ioprpSjTj5OJbyDdKEukn3AgN5qO+Ki6G9+Dq608RXcG6M+HGqbAnT+Fsdgv0O4OJLvrBVLLUOH7A5/00BLG9WTfj977tJYTbZDGIr8m46Cjd5xjDqzbNewPTQDbpEBT30tp6B9btzdct43R9+6ZM42bb6j0ANUkxx+R6AYwgv9b/sm6zOYCKvWcwAum7ZW0YgxxXvKhMx6+AlSBAyM8YUrJRh7I2moz5bJaFKYEV5l1wwoeJinxQ2mJJ/RYMo8bjRhFrjnBdkuftn9MHHW0ioOsJ04f+lsCqxlYDVq9z4/6G+WUsZG0Oze+LourimY2XB7jUJj47EucPWUGhxOIGlsTKtapxRcxYSfmvU6pSNzc2PviiJ+PufK6ayTbWBxXeikq0XyeoE6I0kaFMaA/hB/MMOh4X0RuiYSab/hiAieMuVFRCuEPqJhTICrVmrBEXhAOuKJe+dqdiCSPdh0s9H1GHflOr766bYLmcP0xETLeyx8Qz/mHYGA+smULNljGD09rSE+7BQ0iMN0kUAH4ApNfYD4IS8xUNWhDkPKy8PI1MW+WiAi0iT+1dzqyCvW1j1Mw5kjtb7LsJT0xUr5rI6ggikq1Y0T8fl4xFSMxqqvQ9Iu7tZXws4vMIBFIetYliJUJHMLN2Xi86nPJZq/QnozNTx2XpFO0W5ZD2CZCW3B4sMM1WQ0GJbmk3og4GnSuEEFwfM1G5W8YGw/RWlcfmTKGFCo08YTZU+lYYxUI1Iy8U6t3q7sPeWnLbHwq3nX0XrWAd2V7wMotEo22CwjsZwcvq1DRG8gHRKzZIwJ6gTKY9ReiTuDXQYokDhXAmkgN3RTEfKoLZ2gJvYEpHRhA/sA10ocKEKhVxCi7eq3rrxKXyGiOvlKTRBLDY4MorqR6WJgVrD5u16qOnSO7GBWPV4QkxTYMjHN+TVM1pBTW5g2KLWKZxl5Nq3vz0SV7QsaaY5pDBLaWoQBMsW20nGMPtLTHdqiWZFk3JHs0DcPBIgktg6qFEyfypZAbm2sNNkxi5mgIqjbCbOEVcUgsx1K+8sNouy6KCeFx0n73lDtZojsuhr0sT0LDy0Bi0ul32LZczoC/5uQEeAv9wtzxAsjBEGMZJIJrEIQhg7n/D0TAIIP+6e5IqifVIr5cEvdfw5vIDpbPs3sqQI0l2LdfzhMg3CLVPZglUNI6Vb71bwgGtrr0FuG11KI0L4Hw5xlWemXFU2ZQbltKynbkR5kgPpWe+2c7XvTbOyrXzaZOhhTDbUh8XvpT4f5BOl15LXXikgbj/vrZCF2NmzvlYVjwl1hQiKWH1S/Sn6uxC4xsknq16UERMpxBfEnUcL9ZiUmu0sZ624nJnKMPpqB+BqLZPBgGsxQCuVcwk50krY9U/jLZ0jcn/amezOrn0xSXnxtsY86NNVqbA0UJsjqAL/ya9BRh/R5/5K4Qugl7zdVJWVu9mPdGZ5+GhPT3Ig98QsxaPHX7ywa85EYo8x9Zw8lLTbFR28ismns2WTmAL10z7tLoDoHqY3iLCS5vT5GsPc96WVt1Wdmr76emmz9gTRuKN/0871Oo29r0FmpDgyCBUgEbYxq0VCK6Po+j/ahTPmurNrze8mhNCatLB+2QJyp3C6WQFinpX3ZrxPBBCK+dQV6S2j/A/wobmCvM0Bc7drz9/fO685Y3P04+w4MHLbhjLCjrra/N2ZIFvegg0zEXm2YLZjSGbmZJStjN0FicJNS3Gj33vmSJaOLjKB7VIsD9D/Ssn2WsKhIwdyO2LJWroRNzR1Wr2xztVDrS9Hf33iopnoe0OxRCxH9iTeh+ySyECGuw7Pb6tOqhrDItHRfcZ9NmhG/z2ie7jC/6/21yjP3hZ4Ywkgyt8LU3MruVyWcr+/F2BuFzk9Rl4hOjVIFkKuAULvjFRxV9UBEkSyZEN93Oi4eDQQXJPfKfEZvr5u7eiKqJcl/X5Om6kxPloNilgNi8dR/4Z3cj4x3JZVXCyxFjLPPo9ePTRfnylYMXhGRnWJXly0uKNnI/98g1scTFSsfVMnUtOEsLJkJCnVoxj/9q2+SXOgjr+eZSnVhXhpFfe8ZpRl/oJnPHocUQMc+ZsODqT6qZspMaWayLsXsWJICJAe8e6lD05AKCFPLlV/tNcvopHsWcfknDEwRyX80ZBHH+Zm2C/oSmSihbC+ILYBZKdeF5R12pDCdoGFyO0NtGtDzflfffQ2bGRG8EB5mjne2Q05TvD7ci2Vl95gdB051vpyGxlFHPo9iCEZzxQxDPg7bzjuVJYyUnVjUwX9lGboPOLO8likdVeAbfN1+AItCRYaTCWi88IwPqymTtQmkZBmjrgo9IfiZtAo2ka4VXfBlM30T2BnKpZBrgmMMyP6KRHrcJ8MEEGppcRaECHWD58tLv3kf+a9rw9LU+WMyleuB5J+BX1OoTyaZkg8YG9swLnHWGgP9QgTdikgBsw81935lYdxPzoA9pl8vtT+Fg4Zatr2ggjM99z5ZJM2Wg8ApBNeukRaIIfFg6HwJZmHO4RehYWzQY2qeEGSO+QEXxhTVhjD/wR8wLTpWJz964+trcxFcl0T4tM6iVvUY8JzukuOvfvtujNP93IOHSeFCd+P5dOcYx69oj9kU867Sfln4LPt9JTdWRNEiLL0uVsU02jSvPvD0N/BNDGffLkSjpldycbglDsO9YOEstVCY15RlutR263w5hGMsYSQsJTRhuvAJuAbbZ7Tn9CT2V9oZtmgz09NLZe7fDw2xwvzlmJrOSVIyGPPEhlGi9XdjAu5QXyiH+JrNbVHb3PpXnZ/JTI4qXK724aZ6uEpcnHgWRhkV2lnJ3xozDz9toLbwP4vf/JdxtakzEWu0KLZe9hxaj00S68lx8hwbHyq4tyIGlyW1U3VA08iM6w7ZTxWqkga981vn9ZWx849sizsjL8diC7cHxXS9HVPV9jSR99eB+IuY1kkXQ4bVadab8siJV3yzqNHAUZFH1iTpphq+nEaMcZdbospjUfIudkF3cWFH1ZNQoa5vAVWMr9AB2+eMQ6iJCMzJc9EvpKb4Ouf04XklpJM8d6uyBxV4wqsQvDIBPJvKus7o2zlkxpVf7AqkBK+1XGVZallKXkR5Mj9h9Hgv99Jy0TMfNHNWyb1tKUjPx01Qsfl+pSxyyZgWETrDeOrUByOyl0etPKPjO6Mlztt9H3uTSDITKnLKuTlVy9WqEcs4h3s4gwdfkTVBlhM7RfwAJ1Mb9zqkyiutMOD4KtKvhooq9GILTKblm62m1JXVNzB41xU+OYxJ+RKLKi+Vmt+DGNEICj4LwsOLSHRlRucn4pIg+BjBAQadONxow0hTi0qt+m8QYrVKJGbGo1BbtfbSiM57FSs3aawWCLeyulrnkD3sXXrvIktcQapAlf25CWbqhGnDCkTpunMBMCR2RN9qcHsdtTnn9o61p0qH1gXcyNIVkJvGPY1q7M2bw/1ou3cszGIHyI11RfhxuR0neMB6B23g28bYbUy6HgzD1dRiG9noOJr0NVJ2LD3ZQ2wvBvCFlyk8WsYyU58tSlg2UwO/r2eoKmvs6Z+H1y+syvmUUb6vcdjN0dJAz+ehTuDytuP4cqggN+0aJzIsfseaqktfmtIX73KZK3GYuUZJ9/RdFpnl+auBJqZHiuTbOXEleAvVG9Ad7uUIV1wyQ3Y+IG0OpNQ7BFKts1oLdVlaD5HNGEVvRTWBRGuSZkfzBOPTmtMApfGKvZ+NU6CBI0qPL2qlCta2hAT14rz73RqA3MpopqSkll7JXwV+8BD34m5P667/xCS7o3u2n27m5X3o5EDJymt5/7X61fgJVyzNbEsDgAyhDaL7e0d02ILh7/yulmOYCO8qULRqXXC0eHkYYDwv7Wy9pJx1eBixFUBIKWYceqaylziSXynaZUnAUV6cdOjxDgvegw3EE9ujScrW/Oyiq1nwJ5REqeEh+yR4ToofpHjaZhGP1oaA6MmSXOW4yKXGHSNy3PYNHWArQyA4JJ1TLaPvKOQIyt/TH6VnL/kCrH/lwy6jHtFVyxp1gLaaDH66QkC8uI7Mn05HdgXzaFUYdGyw8NlGxzoo8JFC4rcVftgS/sInACAfltUoti/Y7RG7Rtg5UErMukPfKIUqJVX9WajEd4dfpzTVJWIp1J3WkiBk43kUUxFtlMjbHE7SDfhAaF+qrkttgKCoqjPROCtZjmEHw7ViIWdqFdpcwO1juXTxA7GU3XPbvzzo8t07CUq2aaBInAZ0ee+PZs1h7JHzODWTffGVz7xB5FiJ49GMnG7PqONOzUZUGCPLNMVee0f7Oq5BPz37awQrJrqjH7R5GdOzyo5bpd5hQxp44YV0n6RIkm6lEqoEam8NKbY7U+5nFsAJBImVCUKayu7buiSJZpu0p1GktMNIDzVYHChyCbdH0PF7wW14DHdRpwCqeDUt/vSqBkpPvWfhWjtuBxthGNKBAHPA0fWC96wMb+aPyHGgXSP+PyCAJsXfMf8M0/yOis8rj/C3GoAZb94zKbiNWzKxUb3IUdIAuSAwbBow/LS76QyhopOuim2/haAQeBYJGXE8oIp2IwVTdaMy/9GTAgFXS9HpDqXrdlGOSS2KjiDei7aGHQu+mCGmBbH90DYnXRjD2DxJyvEqP0BzQjzEXgBeCNJT/3BGKdsNHHf+izQh5AaIuTe/BN0EIK5Llsr7O6q7JdipVBktP+BJNHe/luHVkBeL2lJuxaTq/MB32Z7sC/hmNvrO5TyjkrK1ieuri1s/W8jdQigbnbjgTJ9yCh3yzFFgFxhTAM4Bn4p0HPal7WTtcT8Yo0D33sxf6Hx9kH6wew=
`pragma protect end_data_block
`pragma protect digest_block
816bc1f8d2cea1bd0a9c517d4da06457512efb095547767246e2181d93da1bb1
`pragma protect end_digest_block
`pragma protect end_protected
