`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
JYfHIInPKoZSnsdSDf1CygJJnSAg8i90olXEmH/4pf7Wd0A6XKnE+1Px8GJPNkNl38i265iAn0ym2RdiYVgZsiMWzWgmvs+bzBhj9v6RpDDdLVYcKKf/0RIZTNtx6yQoZa7zNXbR7XUj5rsLJBuZuRrsQ52w4uTfMr8FcJqD0NYvJgP/Vwy8O1Amx+Leg7fTwvtTw+K1TMJR18YFPOFxnDVfgt4JftcPpizYE1nu0Mtm6rtAfrRlkaZl1NSMS2KTPXJ9ndmHKHkY725mBlHHL1VpW/zyZztom952sIyobii7Y7votwi7KH9U28r4rAfZLeajoYfnJIwSZgi5au/lAGeJR7R5JjRwQzZQUaJh4QyGTjB/qeK1q5uemiT9Y+vB5RfJ2FQbR8q9SBelYIfsEwGX6ql4TOJIJihD15OHtVWXl53avVf6jDW1NVuhcC6yc7KSH+2nX3/iDzhR5OaITGFjdIfndRXXBvWmtWgZGBSZ4b0lmDUhS2QXOf7BExKIrEzuFn6gmgM+TKzA0UJXr4UuKeMqmXTnhxhU4htSPQKOfFrT3JURSQX8avNyCV2xyX0mbTbBTDcVcib3rspO6bHro6viYxi20EiJzoTaIrcRr7R3f0uSpAlMFA7UJmIess/VWAi8gOperYgGM22sx5+gTPJc04Jny6GSKs9C01VErVX0YSW6FWmFHZPX4U6lkiImwrOydKX+o3qRZisH+Z7icHGnk5cPeUkW/wTJ0/n3YqcmmIWv7v8DeFtkLyHRd942j83XofRLlCFU9PIL0TmRyMsZZqnfAb+k982YJ1sLF7yff0YEfHvqlzKcNld6u5Of4welUgtsDj7uTKFnRttj7k5DUMbWF5XwvBchixe11FEHH+HrxffVUN34WuhJqeC8Z68marKOGu4Dl1WnrVbHQkC+1qOsti5DtsWcEqklYUXnD97K+pDM+P7CDqq73+Au5spvaXXhwCmrkpHTWoCK+szD/6SHR0783SHKSC9OmXoEpqEryOYglyT2br8bUjD1E2v+i0BHUhK1egE7gj/UhYjS6nhpf3f+rw0rNGxdjEVK4Re1H/t7EqgJB2zpapLGcJJ/fE/YNBq6FabWuhC3M97Mge1MjG3LbgIooPVPHCb9d3/aRVi6kpBD0QfcXJKcss+31ibT5Fc/XHu5K7/P37nXcmrMWLzEDWu5wH1aKcxHmWPPcPgGTm1tPTMcMa6s+ZjiQ5IeZYFTrXClvMyGBhMWteEhuFXQbbJC8vB+VAjVGTxeepdtiDF6qmyj95hW4PS3XlrNgnm9b/0B6BJ2xajSrRZA8PYQjNT/jQM1kpzoUWCLeBsaqivHVf1ciEMpt0ZoEqTgMzhNJZmiqInaZRDP2ugN3jD1hxF7zAq6CoJXK+gDnIOubb/pSZLqzaDowAummhREv5LvivKziuvSDEU6e9F7k233m3OSPKhrPGEBANPm4bZ2AEvDSCLBs1EDvtDm7HmyIX+905MhHgjg5+JM8y/tTS7Zy2UqFRIwJvQF0et9z5G1uVStxMMaRdwY2QyBpuEiuf0CesUg2KZwXMB/C6X6fQy7v1155BZZTdWCzYhIWTlzeSXmvy4yBtjNm0NzRhg1VvYZ0sxmRtFTP0Y66LFqQYVNMwFFqADiSZALiguMvs6CJgme6oL6MzNPB6DNLURbLPkYalr8B7k3PZWRDbWxDhlV8MUo3zPiEOhMdXteR/OWlZL+0uskuMGZUIFXrpghVVtkNE3Lt0rcDaNuBinX9g+vaOu3Arnh9E8jUApxx70fYQJP/ejww4p4ZJabcKnES0r/DVo7ziqXo+vz7LcwtQKJco1SG6d2jHdDSN0zNr0QnrAjB4aklDJ/ikTy0HFypJI29yFa6GfSnI0X8L0N+7//dcJ9ueu8kkAcwORyrsEJZo7rAcrgDIGrCHHB+frUAkNy4I57FAqWYCvdUpP/Fn9GVtA3p42/dD/Nu8sLACni7eyUpdwr3zti5xvZhFr8ZF6t/btyJjcGANnwNPLMnZj6SPAKN82Tg06/YhOTwjQp38gXsQBEJ4b/J/lh3kdqEheoqUKUfRokmpneBl0J6J5a4TZvlAXwZXSCUAxekt583rEgiOmVoI36MInYSlL2WVT3boGKrkMDhp4q2+M17CGpRKAzlZ1c26y38XgZSTdVxpC3rVoigJWzA19/lrACXN3srWgdHMCyvhuIEfvT+dvWIgHktYNiCW0Sozoj3K9DfSyKGTCi8RgnWJRkyAeS+MRP8cjnLSKog3pi9pxhA/j7UoHLBIYCWNZJziX8Tq2v5SHJg9y8AaNBWO95OGpcXzQBXuTV2mNw6llvllGzbCYOdBy+fACH/1Qvv5lPmQ2CZTe47ICut2ta9mh8BdYHkY9wSsuoL6xz1+mfhQb8ClkQah7CnqgTDr46YLau/Foy+HGTIkOkGHKv8lc0x4lEyAlgLiIblcWX7Xxbg4f5EsfMwugzI6/TBhM9wyEBbmUB9LFVDzm7oVgO1GAzVuKKnPH4teCDi9+zEa7vRkIUIYumvvN1pMhbnEix4BajisoUBgpbf6X5Wr8720c/j8bpqZcOaTSVBY+zKHV/OtaMTA7BmYuLQRfDcrSi4WvCH2BEuQ/OohuHGGNgFQkPbgdDU1WbmsF61c82fqR36tGDEfU91GMXhZda8owMIdiSC+YZQ/4amVjaVxguxDTzHHr4xY9pib/Si5a4WhQYWxkafJD+PcrHiDEuUw2xbd14LOtVfoHFIm8or1DNmKl2uoxS6FvaZRZc0WAbTcS9J2gNhMkagp7Jrv2Naw+RvEw9MLqFiIzxzo8cYJusGJJvkpTKdK3vw6TQHjdY5QioNwB9Ezga96Zg2srBSi0B2WHpf9UtTTR8DgRcDbTEAqkdC2J77b+IoWAu4e8LskCwU20CvYVoySL0K9JH+dLAUsQlQjpVIU3hlMSqiCXxF9RuGZ+dxPBxxxjEnd3tSDI7EA+uzEAR/IctABg7c3Cqju+ejsAjwaPu+TVPGfJBuIeYlG3ZAUPGG4iLciYwrGDozs/qzri8WMWLrqZG788C83ARgQH9HYSCnhS5VYKnRB3e3Gu2u6JClz+9cpnX6HfFY2w+Hroe0XN0pejAh4TttfOinzU1UeK/0UCUirQ1PkjWl98rjyGwkb3aLAd4JT1Xi9XVcrP3dWp8dMdjuRd95ucBdmyYUM0Yj4ITO3YSnLUPSFujhz3hFXg8Gd/2AEL0T8SCPGSSUnvKwOk65ccww1gBvGHIUYJsWtzomAYXMPDOArSoJmTAz51CUavcsAJMDNB8MMkmUcC/QT0xo2qrWiphdKC0J7u1FSpcRrASf9ayTQ8DRuRsduu9ZrxRfBHmOgfGZqWaK8OkIAD3KZjhyDbobsYUWTnyfg74U8wYSGVxP14dooBgqbDq0kk+9ZsbrEECIlygfuItmKdWGhgynmgMslMJk6OwPZNcQhmqqn4bs7meoqTXqPDJNHFuYho+0DG3kbdzA+AblcgvfwXi3GcaehVLu+2jnmZavkTpPNnPmIDTUtnQ4+FNC/X4jfJk65r2Xay5KwxoTgzCt4Aso7nQhuar+bVqveErvCFfBTal1Ws22ANwM7EbQD+plugNjAaa4BAI5kAYqVdGIsU76Zj8JqYtK7bht1DGvRqeFQOqA+lR/tMi/8FRkAYC2eK1IUTS3U5rOUBRn3UwzcC9pRX7jI87zhbgil8HNTsAGeFWb/oKjsUxRx3ImrEstGzNcgiz3TNKt8OAjPtAr4USm7590qFJnfErt4pNzCHUUoTLdG4RGFoEZNZyRfGrZ9fmYAI7NVBPtT32CURbj0cyGpkOKvw/BSZ32ZJs+wCA5ZzilYa1XwOQZpvsvAZmVSrw/ULjfLkQ0LfXpAKJavUdElJ+Mol5nmNybFckjLRWp2J4ClnazhHTbES0g7bggRxnsmk5ZdFv0/ptIgKAq++PaahukWBcsNG42G+V6Yl8YLvMOopaXoGNG6Icbilmd3uOtTEtOKEx03U1KSAbDTKO8PkbUCps9821XxBnPRBZMUDvmF7hMQgJ/J4n9mKpoZJvqTqKet/03VjAWJCDpau6h3t+jb3admmmrhZ5AI4s9cESnBbWUEAuil1w8iEYYlkEJC0hGyS+zZxe8lgQ5acEnLvTBNV3D0ILVdcZXKDiccKD9ORKb46M6zJviiitzFB0OQP7EDelPFAJ5CKAovAmeGfPFAkIiGp9BkLy55lArHOrkfsrc5RcmFHGk73iSBJrwEsS6khEoti4l9eKz9kS+1tjZNDUZxbJaV5kBa9IyY3UaELr54nJ5jOfB+MfdzryJHGx+0Cx8XWoyxP9srhPQiMw+w8eou2F17cf/A4EBbk3flRnKvA4OQe9UXMrMoYlXh7efCTfZKjH3RxEnqM8iZzDsAbhcWX0ih9zCzdm6ZE+mgMfYcG1GIVedKfHgKvcqNvcIGN2TCKwIfYYsBVaMSpP+VdVKjwezuAQzA1fWVCMcHLUDuJYC2kewBzO8baIGDFit5Hw2xL3ujZdHV9K/ZsvYSWB3pjVIbn3CIZJJWEFtp79oK+8zYBeND+ymCeDIwGTHGR2HfxSPP8snPUKcIdrmQ54O2KBJbPK8G7unHXZNPgwUcLKLFubjt3hEA8R/dzbIluPNVHnnZHpOdWfl+YydHejEtnNj9SL2hCRoWm+sOoE9UkQtWUu5YrFoWjX8iEBUx+qIDr990mVtLghU3Jp2O+owItaxjGFYKQ7Z81+56VNtjYPzHX5iMvlsOPYEOEOi1AQ2WQ1isbnQ+vcW8AD3gK8iOGWJV3WcXG5xZTrXEfhS4CLQBvY1fd4aPp2SqpgeuFYkqkOyCVqUJ+ujN6esBOGwXW5NKoIyd4gvAmoyoUMA9KdJ0O34K4RrcFJ9h3FCXsh6UrWL/nbEoJoWJPYQHqBXRxrZoqMd+lYQp2PT8Aad8oy3PTrdkNF8tt0nkinSRkUUrmMDwyTO4+VuI48lWCshTSJ7jb1Sczv+FVs/ew0+EuBWADvOm5sH+xrHyqOPVxIwLM6tj+wb9AO/S6sihZ6OpqTRoRr6c79I+BIEgJpNJPB15ujruGd3k2p7JStEDHiiXJEKm59CbHex1rhtia4iIXXfpQvWDDlL9sgTeHklk3Ih1MdE1ITJ6+bjXdhKr2vxUBreISSqNjN+VoZlf1oxSmV5bX4KBmty7n4pq+eQJDGEzXGx37BsyTN5NTUBdHR2Cv+xkhCLbQ00Ou8twQLpqQso8w7ELe31HLbBiYurna5RXNGSvgxqrNpCETr4y8fstRJk/AoHPZ6Kq2sk7VkyMRXSoi5k7ktPnj9xjUx42XF4oX5Va5B6KSfc5/sG4qAzKSx23JHdl6yPHcUnaMVQoPm1c8ACMCMfC1bFcUdS2pSa2qCiivUsXzd0mOUk8gfxk9kI0/57ytMCODR89YilFBsW/OF9t+5SNeSUw+fsQptt2yC///xfaPcwsXXNmSD3VXRWkTP54UZf8w3xbira7MRNGLJFV7KOMghFF5aZmrkVs8FDoW/mlZmaQIVi358LPyUUuh21iK38QavONTgVeWe+KHos8YAqU15kUXV4czKbUtTlQaupCQLAGnKDBPyxSjJiOOWsTzH1X9TkB27SS7psFa839yU+lK1iqwAJ6zZCQuptIsRvyKTR2IjfsCwx90sT6sTa+VEubWyI0Uxi7RS2AXzjTtvW6roWkF2bj4OtbuoRa4fs1VW1JW+xs2xuK/eMkFJqgLPLj4PmdS78B/UfrCx3aYWTKvPXunQ4bWeYbAe30xMP0/39B8N5QNoLlD1QE02UOn0KOyMFfv54GTs1a0CRX6OKmlc/zDs6e1XKjxYZ0vuDZGzoeBaExT1+OJQUVyYxLJH6ZEIDbBmKO48yjI7GPuzAaDtnrzDy27/odY2XiePKxrRNf2V+XBGnzmbyGne9chPQex8WlMWToDS7Uw6py/X98/SFIvWLfIjsyuINynjiEXhoRaCUUF7PlHpabzS25VdJQEdy/7Y9Ax8Q+sVcPQp8V3/yv6XDj707DMInfyl/jXMhpCB6yE0478uthyuomz+aw7M6RdGLSLBBTznfAdKVvhVBJoiTnjhLh9vdSueqfq20/4OfGDRPrJiPgxfVJd7G1cEd44l8ATPjuYL0EELU/aKwiu+N42Y83F3BwQljSs9itJ78Wgph0/JNYY32uKWOia8w0WzvPCIN8DBbB2+9KypKfY6Ru6guSIR89fatem+H0L2aE/YmM5161+D0AlT1e3lpKZAi2SNvrtmO2I9m8ybSMYVo5Ck2cYHO0cd9yNbr+/lwLy3gzwyCBpOpINAiHNATnMiZxQFQow3disml/94DX2+Dz5kUsBhdvdTIVXHPFLZO2lCXw8eEkEaLYKn8QysGuTcqMimZtLTeTmraaZLXLF+R6FepbqHvsg5zUS/Qy6kqzdylozq8alO1YsuFQge8GI0ogZVQ8HrgLfnQfNGIyL1ZxcE6JXGMa+92Yjwrkmlc4x6A5uBf20GYb9kgzRr2YzB2+wVoogMhDOx9aodfwe/pS2VJiD+Wc/+frEggGrefCVbXsks2aufOV+UvADuM6YY5/UHFMMUKUIeOuleiPFnCks38s9I1bItmXBQtEe/PZQWyJ6oJC8/HJBxvqPM4pQUQJR/nlDWW+2t6bufGVQ+EDay8MREKFSsxcDyQDo4rNVor5n9063mwYqwRBzVFxX2TxhRVk8PoIyvsCBzPjniVkwDzTn5GtxnyOT+j+rwaXMc13jtoc7qAwjvF7Si+6AaeP27k+fMm0REnlnW90UbjrYCbOLWjl4R+xPx5teIdhW9PcH+VZsMcetQDe4T9z1y4BaYXCvFJOKbmYsx30s3fXYDxlM0JPIRu38yecAHnke/HcZAz+HSSeO5rAP+3YLfg/iNnVmJzvfL+l70unjfLUeza7I09AmuIhJKFf2KIV47xlRFqRug55vuH4BEwgkYacIo4mCrozf518cdTI43P7i9SUUUKnO3w0qr9Sl3NWmbs69OWv61zA5H5m3ovYDBBgpBlZRibvwhQAB/fUs7ifoyUvZ+WCdb1EJgGVyk+Wji2WwHKhikccShRrJ7nAUqJ/G6twA7Yblvmq2j9E7B7I5PsC+Sk2RsgPLttTrk5z+ld+yuqw20R40NhCER3WIiUTxDLNpQxZItxah0YNcNHbo6k7COL7jW5YCFBN18u+3TCYYDM5aK0EVbDNKO4YF1oqMxRdb8CwNAkOZ781ga8QUNrDRPOWZOTQOcjDc/r55A/8L8LQG7eYgFnzae+HsnIqunvLN5AbHxwOVtiDJ6alVfz9gWx5QjS5f28M83VMBxOv0vbaA5bgoPoordMfFxtjXE6QYhUdi8apzOaifOD9udlu6fv87zaMiKV+JkKg/5+Jmum/hiHaEBi6b/wVvaa9R68dmibEYfzk276FjMb+dWxShZcbJJOqHWhA9VoRCIpsl1PR9saDDOsrSn2jfTiNbuWATmDzo7ROa6l1XyGJfiZ5W14DOjHyesXO75yHDv9Freke0b5EQd4kh2Kkls/LzE0z+wvZd//ZKK9WpAmbMdrmc+xL2lbxdfGdCYHFPESpiFMvf15zu7MfWL2Pp9oOg9RLE35+1MFmuQ/AKA/9rQMS1jjOZLkdNvJLMGRcbMcq7hUxubchCctXiPgapnVQFNtnAw56JIeNb2V5EvSvECCh4gpM9vvTMsKF7tDs0HVMoDcLBLlvF4QRWPv0+LQO50zIVnKz3DvpP85VUvzrogOE4K/FTrLssiGEAVhiZuJT/d4JSHxKCN5HEc2V1aOD0w4fSVnFs/Qhc/ZeTsN1TJiPt7iRmu/ASI0gA4cDvOwdhslfeuvNmygZIIjgYG+xcYVbd/Wv/xyzfd5w94vIu699Y8hd1PnH+w0TSjjCkxx4Pc7B/5I8gn7UbGdxh2sMeiD7/OMYhxi5f/mCkiwQjMfbDnbJZN0f2ciyYPd6js8vKfO/BMo38GtTejCy3adHGgE/wWrFSCLm3/FGFFCHb+JomKFCiVd2l1OVGwRNXqnHj564u6mffWFuoWI198uAax6iI8C/ZkvI6VJjwTwwY99XXUIR558fekXzEexLCJ8p50rUHL4HRy9uxOSg1BVkZUXgTUjYX6v1TigYoqWplNLofwSD3kGHJQwBrXiVF4qKnE02Bv6FzzyoRf+4vR+TS5la7kjPh1uu7cIwPRSv6A3jTOyJjDbzci522cY7da9nTYhZMg7mrMoJ/N8Zi+JT50iCgqU0PmaY8m3zVTCf7yO3741egVUJjb+25Wkpzj9i0pRL/sKyKuWsr7HfWI9g4XWSKbOl3SBBtiE6uW6x0IS/MgpBZyQf71CNxNGep7RUuGk1kxXFuLwgiQDTCXBG/gFEQovm1STiHeVfxiMB9G7Bv7OiA7Ar3zaU1XTfurt8K1aewnru0GrVulh+xVGg2qGO6PoQeThhOBF06kN/osBflsJElu+QrPBBsQA0nsoosMn2W0OnK2mhMMixyhQ3McTweK3ICPI3q5oUarkYWtZ94CbrHpRXsrO5kzjgsGuKyLn5G3uOQvA/kUe3c77rif4YJKXQHJLKTDOTDNFRPrric4YOGUV7eiZiTtIVvs2ZMktHvHnxdM7vglxlwVP6/y4i4U7NZL+bNbC2zbJ21nbPvl6p19QFjokAaMFwCkEXI/Wr0V0tsel5W1JokkYSENvHRltyWvn1WiGHLMKEHtUxcvHHz4xu5R3Mux9HjgZDx920Xp9b2A7zdKI2TMQsAVloL10gRnLJaCMXjDeiN8RyL7gtXTFk1RCHrUdXL/Zm1t0j28gjyxgr1ii6ziKfcVi138anK6jftWdNeQf32ChNXUqX5bgR4uSb5fcz9HfJxiKZM+dbceA4czqhDVqVmcCWG1h2i83+pZABSAlQ69urafn21uE/Dby5LqMwRDeNJCMB0sVZ8/RzLwd9zKZFrv68huzobWSIbY8JThs6FWrCdWqTdj1QQu4aj/XbCpKN/531QnxC91ttbS+mQ5FFw6zOBXxJ+l8yLt/YBOM8TB1rEg7oJ8ASILX3f7PLRsIAhA6opwWaMzEFkVFtr+4DTSIIIhGnxo4YfBlQJhpr39wvE/2CZkW5beImdFP79g9nQGkJW29tfK1waWRCtQIcHGUYvmgg1Y8Q5ATYD1XtmPVkQf444E6qvEyzS4E+hRTgqDsvimCtWn5nx8hLnuAnFHFoPAcx83X6ffIPBGhIwwGwum9Pvg16fdkgy9lbAsK5ZwSF439LB/rzsn/zs86XBqK1PM2McuFlBwIsn4l7j2D3j8LLU7mcVBR89i4pKtNJwTerSjLy4EQUZ0CojmFyyw73HZR8ODZkovEaxx4WEq2jiTY7f5AtTwsU3CmGdosNU7cTb+vzc3bzPKY7HgGahQObCvhqqq0p28UfztDaroQnFA/tgis72gHxiWRZULDRf0l1hWXkH3BO8TPur0xSt64rh3Yqr9bWClqKV9qL9cll/re7qT8UdFpmywv8Ovpz/LYP3IuJ38j7kDUnyUjK1YMtci/YJPs3cgcUbmYxNOwZCHyj9mu/oA/aah/sYo+yTMoBznT73rj31x48zzuDijRxJ6/h10SFf/hKfKb0YazfgfEkYAuSC3li1VVRgoN1n4Tw1FVHClHOyULMeXiy9povjiBkIg+pQee5FsiIKhBwEWTyy4DIesNG5RM+eNgckPcJ+Bl4roZrV9iQ5cH6vvUJoSfwScM7+Vv/BDRUnwOzJzslxIwU/ucfv38GIykqBqbxCAhgJY3W1RMwUciyh70TGSjC6pLelCTJ01eRvshDppFHNhCZ6qEHkI6i/j43PG7Cfbv46Gm9s/i4R476eJwKgI26ohCapQmEVwZXfu782law1T3SaFYg64NB9f8eqVBUSrpsVMjrlG02Wjxu/OIA8iKBou1uOELAE6uWjzk3+fFIg8XtaXT1+ABjIPQbOXwPtEa7/UTVlBLbhKXlT3eaJcLqdPvDzpaK1LAvCQkdI21PiXNAq8t9DwI59tHRxigHufHkGxG69K1u/AhdFS+kdqIojMWeTMu/3KLVzSpjnTKrbOnOfAgEXMStlQZ6Vp2Xydy23n93w5ktZ32vf9+oDWjwNDQLW8Kx4M7qw0VmQdwYyEMkWj+gt0jbnh0x1FACF5zkNeTKNDB+i5Jd13AvsGENlXr3h0ppNcsYr9i4zuk2bx62J1FfOjQj33BWiZ36lH8BFDlq1OF/tX00ka+d8bH+fEMUaF8jUn205ljEVDYys1eDmqsQpKK2BcRTiXDBloG/bwfQ+gzFQaIE4+Ag/a5L5QRbfGGsQuzs0cIb956s1b6Tx9+UG8UIVjskAsn6UULT6Pf2RU8Ach2o9pmF0pbbonmfLumVbhwqJT2GAH/W5y1uoTiSA6S2ZX1jW8IsMH5cQjuQyBlb5VKNWg1sxQ9TRP9Jq4j21h0gbn6RcvG1Li/HgtQzRsJlQIwFlxPXb/9Yb53EgVy91O17REE61pJG865l1PC4spGshryTbF3Kyb1R3JuTnEguLRGPPPpF1+gbqT3e5KJH9N1FrmP8wjgRh1rMvGgchGceWEWXYdBCfj0GAPJEiz643fG9AT3TKS21YutDk6Bkj9ISGpmocJUJlDqWqPkirgz/bxp/+w6dKiqQx4FWIRBgmobkM8ldLzCkRuKbz7gtGN9z6XS5x3kM5jKbDPx0GDLB47BRqVD2ChIWcWTKs1T8IH5UWYx+OMVuudXhuEpSNjTtLKzqFjh2Idf6zcG6/r0sZXBWT7YvWCo57TQoH4z4umXZduNcQKWSO+rjcIL/OLyHzIDwZJdXjGbPcusFSyuDH2IIVjitsV/hdFj6adt1dCmUXE0DPMhwdbCL4RgpVWEUY/LrcXmMncLyC/RzdbGld8uUw/qVt55udV1U81sBxUUebpWChfKWcCFyjOJpuUvoeP86ZkpTkfansJ6FCrCIrPTqCEThmtgfveToUCnBEWcRIuXqrWYiptPC0yrVYbmJphzOQ10/Q2giyyajxFL3FssQPatVMivw91pmrZuajt7bYd/u4hC7iLe2GXXG1rBDYDG5Vzm/5YmrpQ1/4Dw+R9RPZhx2l/7Z61Xj5I7lMV3OwYoOaNdZRSpDI6jVlfO9DGZ6N6scXvdZJvDOCW4Ttz2iJR5YwtCVvjvi+fmKGrzt1nlV19GvBQLbAAKoaGzqIuJQP6c2YeA8VxLtjmlaNGtF94/5R0Jz75ZLmNPcs1kbWdHMHs6B84pALMd8oZ1IpjhSQUeNYWOSVpeEBOxLm0bDUwL0HABaymJiE11N4AiQIfhQRkCd9lNIVRKiVwyj2stNILishB4qawyKCYjgCf6eYJ5bCLHvB28h+pVAflBVGY1eSrFMjkI9KT1Mqa7pK9gh1LUZPSO6T1S57lssLlnDzWQdAADCnkc7AQcQC8+7Qe+hgnZouKaAMmpq2x/JBMYS1o42ox6hbfizFt7yB24r8nZkBtP60SmwPjg872agiTmvrbUvDH/iUJ86tdFZT82KB7aHB1P9jv8CQDlrxRffoGFH00XWcLeTaUGLyRyKssDbPH6h5t7wjcXQX/79QzKs1dFW8uHAbPsxLwbOCB9Zg43TW4BiK9jLefm8Uz+WXK0a8i2pUumtxh3HbKNWKjPG559256LwY8IVP7jspfvGYk2MCL9xSmOyyGW2urNucVdnJRbho6TvQCKCnkrnRS1yE+VoHIY+KjaihPxFE2bq2HK/qxFQ7wOyXzf7q9fdPk6umxZyuhGSdqPCqJy6lEbwXV43YXXFZdeg2EHmVqO7FWUoLgGq3tDVKd5dQgv7Rd/NiJ7dffee+skqnD2gQyE8DS4x3/qD7wxdrmhCrOKSekiE6n6WvUSsgD/xNLkl4isRIRiLal3Vjlk5oNOU7vcK0i5dw60Vn6bMvxc4y99x8wc30ym285h4ypEsBavEcOv1qjpLDTNnPE7iNQJMkhR1E08V5bDin8f2PBi5F26406F8ClgGdeGVl1b6hme8SVzxTVROjqvcjMCzFWbrwVIGJ5mMy7STwQ49DFzsxc/owpbOk4eenkEJ886rZvoA5ZK8DQvzr4B79HpSQktLq+Lfpd6r7fYLAcFe82vVk6DfeMUWoQI0FkmMnkstBgq1ubfXlPEUfFSbEwOsR+rFiAvxe3xU6sSgZzHwERDZYm/oHxdpYdnlZxaEGmu/MaXGbOc2et5FYZPkrpce00FA53Y7J1WOTb7CDx0jJNy0tiErTg5Td8jPKjWPUoaTTnZntUFMdb9lY+AtXTf+qXYUNDE2I4oo9yusXqCg29gqQFhyGrfG6mHd00KFUQ5avw46D/ODKatpw3vEfWk3N4fu0nOnMofORbuJ8XOhCd+m2GCgUhuxjRNSN5f1IJ4j4c0wa957zQf5PgwPqai6ywEK/Yoz5jd/Qx91RC3rYV1LpcV+1z5C5Dym9+c5BwQRU7wqrNghixUx8evn/7fhS3ir1CHB13GIbvZ1JXRUlW0jhT1aIKKjV4TZh2b35V6X+nS1MZiCr6sOQL4cBdribO1608tv2BRBiBv06j2V2UsYIZlhguZuZ063JyTPz10wbjYxljt9w47NHQ5EkX0nRVlRfs1wGaQmnWdB3ly9cHI4botDfaMHzEtCNaEWtqMtA6xxvqz4JM1fc23QxikH4juxAaCN2D908K7QNqtObob294BeNIQrA53N4xXkLkAe3dU1xo5tMrfhLDA8JsQguq66Fl4z+vJdeZUtBIFvo2X7tsZzfC1tVlJ8rZEUDIOT7tchH7jVWIHVhO7FSYR4a92J2DYqQWa5yPmSP6p5EDez8G/60uD/y+ZBYzH6AJrVOEWdpgTn4=
`pragma protect end_data_block
`pragma protect digest_block
a74d180b2297570d29b65ccac06e226798da191253b13a525a71e9c7f91a5b90
`pragma protect end_digest_block
`pragma protect end_protected
