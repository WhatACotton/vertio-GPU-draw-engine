`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
Jds0xET2c1r/a4sdkSiKccN6HJ8WgoQkDGmgzU9O50JPG9ioWhuR9X+nmc5kPeZ4nQbuWxFsySmfp817BfcO7zLZnhBLvax4+78E4mWykvgX7CcPQ/tCF8JwH0HgaA3yCipJkkbTUAKSZJvxseDWy5KIf0udaeHWo9174Ggyq+usDr+2x7VGXz2eWdonmFWAQDEENYSdNtDF8ohMFzHJu6IzXqbeGR9m6wxdKrwYvE9ltyJqrTW0MD59SW5AS0TqPMMmDFldiB3yi9PI0+kpsqyFMqZInc1jpVHsxKmJqckU92DU/oSmO5ZS69ydwRMO6nk2QBzFAi1J3whjfO4rNJng4F+lacxhzHgpVS9OUFjfA33fMp9fsLezNHan5IVPcadMiFE8CCsGCE6NgIL040xqlJjOmKYSs7WVrenKKEtMf/VA4kFQTdtfUHJirZlVa5TGJlZmqEbXoIyr+DyGI6kfUQ8X98wwI0BWjkfdc3Vb58MpM5d3un4TNyEtCKbZuYwoJXkIVaZLf2d9xoUZg/efbJSiGZrZ8A35a7pshbFMSlwZYTShrlxHYBl9TechReMLGVbPSPB3XCqgYbaui/BjKP42LfDipc9dQqwqckFxyrhbLP/BpCX9+071PWS3NOoCFX/B/SCl6wH8cXn5rcWbOV+j533pWQlBwVBSKaZjfbHvQr11sE/YF1vfO/T0ZYRiO+ART7A1y0vlYujq3jDttll/hk+nR1hts3tq1SXwraoEVPFpW9+6QcG5vuc5ucg3BkrNcA9KEYap12mGfRVDO9iEX6xCMmtgdJNogqFMMe7lDAreGyr8Eu8k7Qx9ArYc8LlbgXif0RAUjV3jj8/vW8OwD1T8yhvmW4ciQH8/y0+9IKgzrsD90CALLwNw2rIeHf+1Ksb7D2fgf7jnAKOWGlzTe1lqRvLindQ5IvnlBuyK9aTtpsilBDv4GyBRPFAB2W9uIcIuwAs6Ee6GSUBFHD9DoVgdGnf6wp0wdg5jsFultVNoMNo+I3bklEz9gLb9k9BI5hJSI2fANbD5MCq9LLYlUVJcHfwuZoj1pXjSeVkuDsG/vB9uQTlAL9YpKKybv4yI+VEf7uTc2oXdqt3P6VcAzX9ZVv+xYF8oua4tGt2dRg+kiYkTbwRwCgll2EktZCCDTZ5m7c2ttH07Pa1zF5SHAoHTJ0OpErL7KNBTkZK08UaFgqwqa8lYJWBGa28KGfAwuQy3ZhxF7EJwgFYZ/eVKF2lAwYFRrK+wYm1fJlfa/xYEOOALyd/0uZYkpXOsbS7S9e6lY74wSelY/QvGvvjHrOdiNEUVVe00szZcibdU3umJlEpZJc84CxwW3vkUJj3ESDFGWhcdyy1V/TScOfnDFtDHR8rCTaQb4Pdi+KFqtohlXIqCjH/LJo4zvjRZzj+Z1kC2+vBX5RfaVgLT6F4BfwavVBJUOQ3WpiwDPCkk6Nkx1PDInk13sc3TNJrhoNh+vCQTFGc+BYujNkQ+yK2+d+CJwzvsSkolL93kP/GvdO1H25YuPcJzl03RI8iTnz7+z3hin3qVtZ/Y8z6SlVGxyBGUnaTyro2WvW0sT2xYEemiU4mP+w+Iu9QPLhB1Bhg2YEt+W+xAWESnZoV4/cMjC8BurgqqhngnoxZJ3vCiiPNlc4n2gV79VM6802oiZigRiVK27+j0womCQ3v6ENeK1ucbgcIW8tc1fNXmFRW6dB+AYxdGpoy1rCYnMuekUaJNP+SDsefmPmbRvbnHAFRL+/deYMpbd8YC6dfmkatvrSx/mB9qW/VAfSl1pgE0Bsn8kH4Na+ysLfURRu5a9M1UdCaDQABRIgLFGXJ8MvIoQF3R1Am9eBJmtqJvDl8PR3jFjPt0ZFioxdpoVdskt1NX2m8I69KGl0pct4Sn4ox7VtZcW++cK5h9HIuKJWXw/t5AkzzKF0/TAHtGxsup2zMHPWyJZMPtuJFckii/MiONVitO9X5u8LtVIPsy/8oi7CVwSCzqmSh/6Iv5Nopb151qgsdb0mXyd/fvo+9+I3Cv/gkkcM/2ZCmYiES6ibcK47x9/ygWG1BEc8NdRl00b0szsek4YwtUHgLlp9WBnm3s46o4/wT6LLXAAYYNNAmL7ezzSPVHeF57DWsqxiCr1CIOHbTZIL4P/glBhIrbknjYRLaU/6kzjBsAFObTL6vEzOV+vse/ckz3lKdykFcbA7pPxUPT6BKuaGdz2lyIBH/yHpcio+0AYJwt95ov5iY6IPdT0QQ9slicah/D/AUAUde3WmQ1XGETnxEcV1tvsVWSFdKve5GZ+OLX0J6gO1/xdf2l3+J2vDax+9qVS2Op8MZCDq7xb/KHcmyEeL2mP/e7igEE12J7Gzz3iNqkEdtKw3AJyPNUN1eCMUzYJ6Tq0taqu59ihEBySsW342WZhXvdo1Q8zF30a/dsyElKmFjH21/6bDFapLs1Wt8xTovbc5PWS4MpfynOjkdApHXCPERJSBCo3nIzVXgePRhBRQ1a/57tV2+FCj7RZ2YOY2wCJdz/hLpwYkcrkgAcfbwtAeFlCKhoyl8W7VPtZaYbyaMhaTERi0lItwu+RS/BNnf2uGOrFN7It5jrGQ7MzQbHGLqUGKDmkwnos9Tum8sWRiVM7/xdnEs9eJ+3Cn6QyOa1UPRraE52DMsdWdWoMB2pZS4jeK4mT/9S2xTmuaAYBxcEpLcTgYpCaJ8FVeKhR3BkSjpvjOZT/K1YWuaGe2UQUoOtB18sAxFf4elnE+m/pA7/2c0djp7WAgvwenHcfsHVPuBKqqTrnypSScOr85OsN1O1g4Lyk1JRtoz3wHm5qmUkeppEapOD79i5G1Mi0cMY73fzHOiIX4GuXE1ugSRlOyzGLvR3M07JVGkm0WjupG1nqQ28m2AnbjPpk24uo/BpIot8aThGzchdbggAR/tvKHHwuVrfvK8bm0VI0NT2yo65gxci/D3YILzLE86f0UOXAj+fZ2p8CwKvv25avHgfjyPwvZmNVjMppzF3yPfphBN0tmnGGr0mW02Cj3TMPczDMNOLS7xo0SwR/4bU5OQqD3bTe8jp1HYWOjmGYBgtQduS1wsoHFA60/TzwaVgvbtF6/PnMz8+woa7/tpaltptg00KtI2ekrWwC1DixP8BEc/aRB/xNdDtk7eKcN1QYQm9ElLQCaWYOUzF3uvdfwCKqgdahX2npmXmrS5FyKSzzbzNd5RR0QUTEi7nw58UJ93bvc5wrQgPQkYoa8u8y90XZR6PCza+z0Z4s5FERpsZ3QjEGTHoFtIb9Zbt4CcJzMfZp9vDrsn9sd9zg/zgnUgdlc/7FAyzWPCriX5ml8S5W6O/vdk6fXdqLYnPDd0BJCHys1Vpcp6yn8+d02PeD7lx/WjP/O6i7Cdho6aK/A7NVhbW0oWIVNpe4QaxRUEjrp3rrcagYfl+XRRM6mXs9Ry+rCVjwE7/Qb5mHh0QTaNV9Oy1w6tNueCt5/2eF3OjYLgYefrVci539mnM+AAUIe30GbUUxO+2LwB91gNCX7djqE8+w8dcXuke/P/3cWJU26WgdrJ1bssMm29Ocrh6jS7dI4H+LXiiDrFu5/U1OJhQta0hZjXCADWUnqXzi7YfUxhcHIQCl9KyH/FFWdnb31Dd8uWrYux0M1z705WjA/k+aVmW2p5KccAsPKFr5aSYyXEhKOoWWu9hTq9SU3V5BZVZTDfh1DxJs34j4GVlv3MS9JaqYzV62SRnNPvup9h92U8jySiQWIT8c22l5CZSDy8MT6403WsvFJFdrswHqE9mvuxllf0rOnGapTO4/70Q62ckxzuXunMfO63Xc9LGrsMG7ZTWjgb2SyxcfJud3XrzE0dKpZ0SbSi6eTFlzLoyHY6aNK4vuGXnTOpT2AoZaBB6oDbYCvc5ICs3W9pBoNkW8oW3Yc0pPXgeL9+pD5w8WLeWmV2UffQ+gG6Co6t62jpUA6kzbdDZYlp3/VI83WYqcbuMIs0ppdG3REykB82+1rs/DMxJkXiaEEWiXJvM1qOxp5kCDBQTkWcYXKHKRzbFhFbgmu6ltJLSisHesAMo8Ux5nQdrrwkHzjD2Ge9dIF8GnEFTsR3uXYWYIQIwlEiaClNcJuQGT+7pl52MPPx/Zh0dBpCNlyucTXiZsn7ybBEqB5nsK6P4eSW1EvIM63HfEPW6aPDknJ0h5xO2t7yBzFmwJjWJaQBAk/FJr+6r54Q/FHDh/BkL8knafgVNYBw/GB028aiMFPDJh0YP8o9/vGrTgmLsUcmFeLKvN7Mq2a22rvzo6cnqzR2xo2DW+cqcxP6GXceX8A9iTmkfWNSszvfh/RyxqUwz7lJ6NyDfbUrWXM4cm0jLH9DLqPGyjSmYr0yue6R9OTRIgvx1DTDZuhIag2L85qhpswusFfHiAtgxyu0npaGd6w1X7k8lwUNHIC/aHxdm1McG3CUun/SHD72I2DHEOotzFZLlQvjy68nW9OA7nIU3ckQzE5LKSBJ5jRTA4BSxTWOyo0JxgaLT86Z89S5z0czpKWCYsRd1fYjd68emcF7lXK4V6N9kkXlHl3n0cZKrImTFbCsuS6wMoGBVZibticjvxnJxg5Su9RN/7r8JKIhcQZkgn2e/uQVYe3jAjcFGtheXltyBnHR5LlxiN+VzX5Ve9WSp8rYgARiDTrabkBb9DSg5+CQSvfVySbYIPRerzOrZXHbu/19zJ6AcL8ycl5/UPP/LDXkL1rS+WUz26VZGgx07xs47HK/6e5zbwyMd32r28n2+u+M2oPGcDlWYeB6SQHZd8CizDHvVhDhPpuyyvgLkdYYcCrDZ2dSkP7fuNi7WlwqEPqJCKVaB7zTmChVrdqPFKRvSeN5pEaks2lAiCii+f0BDRtuKFjjaZiR5sL6lxIjz0qXHXCBQCOkriURGMqmGEFnkXaImLY/HFmNQ55uikydN6FQeYvUEzHP2ccqYpXc3/u00SKIuIWu4HxXLYI/8+539vTD2KOp8eBV+MAlUlC58yrYGr+284lSNdmALFiaP7i/rpxdxuXR8J1/J3omtX8HK0dHaBvrUDL7++YtoxnjQCNkbhVzq6l0T0reuRbmezsM7uTeJpkwoOtQJloFXZOCnMh/BIJBxZXnCBFG/HW7nxjsgs7AhlBYoqyVZXd3VYMz52hJzNMLlrd4Mndw4mPNrJRqu98mz4Bgwt58AkkUv9vbcimnoSbRzID/7+FVHmbZKTNeC/yqXCmqoUpCZe5uZySjkPJP7Gl49Zh3bDjqc0SaOLIxaQvTgHkHyEL+TBKI7o8LSUqNJChLNIQ2pFjStyb6rkggLXnCNlv/nQxh0cwgwUHTQ14aVOZN47O/kOKtUnQwEOc7oBcLAyw0n+FEty+fXU0Cyp5pPhsmsAfXwX2H0umZIXaEoyiHUsNCI2y+XcwKwAlrYkqhJ5lFjttO9Xb8YF/pNvj2rqbNadm4vngkypOg4rn8pm+3ttnofHwhopwBG0PRddWf2YHF7ESiaMuq10Jte1rG0hCw2QFBxcFimHBg9oaLLcHNHL2gJCMLfwDP+PxBTUQOVvxt5bdBb3Rd05E0JKxxE0SeNBs/sK8p7Mkl6y06cS8aw4YcC/csP7oSdrvZw4Vfsn8SrMc3lsuTEU70W53HO9SX8Zerdeht0Twx9BwJOCwFDjSrbzGMw2ycMnsxvu0ZWlZKE1LV0cJRrx8uJFOJiQ416ZoXrXFTVcupqb1P5ErTkQIC6E4qsbWKRzM+LQaUjFaH1V9fujxvBcptMmfSKw6Ddgjg+ZoZFpRFgq1U0QPs11oFpBaBSxoyU8xW18zZB0bmlJSlDjfiNLAeT3rRhTs7hRGgqS1GEfcMtIyTWjiA79UGRSUaKAnuqx6rAVDTsTJ72D4viL0Arlyua7sgOXpqU6xZn9wkKJ6EBGVczqC2qJg22AVT7gaiQhfTzNaAQclAmhq1SpxnEYPDE6BQ+dlSJvVthqB2f9fGY2jwPgoeEfu3JpXr7zH7efZDBOdrWKJfr2CsP/1jpp3XqTrlpIaVpc3fCI2kTHowIE/AihyNKky7Di1A/gLRDnXq2ST27NDg3d7sy+z4LEnanGEnoAIniTJZNzVJPA//nr9mrmyB5up0DWJ8MOlRUacuGeBYU8TujHMhakn08mgoEgZuOwb2o1vJiUtRzBhv3zh5y2CkKElqqKavhIzfZClQEncisq7sGSk88p0XQWrlcA9+JFnlR2JiL/fI+2TwSVjolfXoC2W/qELgNac7LtMhBVaLroW6WN7NEF6mvhXGUfYzxt8rjUoZ4qLDmEwyM+laM8uLqYSTWJP2mhiR+dG/Jp7ROR4vlVp4BqE/WpwzK7xAVf1pljFaQQi/ZmXb5cAnidZ09GPGqjBJtFLGvPsdouHdmhe1gWde1Iu+N5ffpjfCr3WmoR8pPjKuwZdSwcyinSluT2B28ShcbarZGgY+rT2oITLbSbV1EOoz6tb/f10cML8kiAX7QrfuAZimJVtfZM1KO+/0M+UMw9TAnI35m3Z5aGj53fdCMRIW3kpKlq9pIdfTDeq1oLK61TXVcP06QTQGT8EddAj+deDLHrl1Qt9+Jn36Iqe/gB2zRBTc8pLc0f8ye+r/NkzLEPeJRD3NZDk3mekALoRR65syhn2VKK4/2/8AxhO7tdvC+sp3oNSiZEEXXKjftqDEyqy/v6lXnLLcYr6N8stonRp+NUn7YPp3GrqmjfS34IgiKQBN2KjBWwdldjlMq8qpFQzRmD6jOEtPzept4bq9Vc1Vkwh++Y/C53evWbX9TjXXSIcQp/HLigiD2DZZAzb+vu9RbbvU9YwobtYC1o4udbXJsDG1yyjSOiK0rnBoKgXUu/kVI3s5Jvg8W3QU0yk7EDo2CTkgCjejthKd8EWqxnreduXHri9LYNkDo+xxACTkLQ3UKjq1GXTMF1H2vyGI1bJlEK1liE8eZCJ3b6WtznrIttCqnGIDGw/+m3EAzsWTLu01EH1ldfDWzSKMl8gm215qkLSoa5rlmKzlTWC9cGGa+4bWVqC3+qum7wG0bpnBn/eI+fhB7+zA7WQYQC0QQ78gJZv/I+TFQjfoomRFdR59TbYt0Nxx5C0jcZBacDV/ueoMAsVZ+pNOvVZHiVD9mNcT6AaHFb5ArCNj0LweZwt05PIvGkMRdOwVdEsCBp5A0MO/dOc/tQrJVG4HY0DJHpnZy6z0ahvDGyZ4ODBC2L94m6WATHKvVFFDBYLFES7zMLQVdfmuaCeQeNlzfpi2f/VnOKDl/4ec+vomDoFUJcT/t0dzszf1s3t8X40r5lY+J1JONDxtjHEmli08mga6uHuyFb/ctQpWBO+RiIs0RCgaen9noMi7VLvpLcQ/gqBUp6tRSeIzgicLFo/lVdU8WoxupDOUM9+OQRrcEF66XpBxK1RYGvbbm2ZOFrzCRy3b2Aw37BXyWUQEVPN1qOJm5Usfr6eTVo+j5tgnislTaXiN1nrnjMoDVPKpHoY/heD/I7C/cOGpP+JHhzR5ePSGZX5LmSK2e0VkUAeZXHk1SeWY4WpuNhHSNZ6mDyAJfJcfVJY7yFxD8z3XtXSkvnxaBkiIlCQSY1+gYJ3YHNPYw8g0rd5g7zaPQfqCz9gx01KKNZd9BKtNZ+cHuXISQwGPBvdp3SzxrcUDaIimwnOcwvUyYJtoGtXwGWhgdYPmAIk6JGOz+fxzgrF05tCwlXz1crEF9RTEnEkFu53d3ukXuIjewRk2SdxFNy3hAmdW/PX0qK3GfTYNtwW+JL8kW6uv/ROWJSBo/SglKPh3KmuuZ5xG48Dm44Wetl+RPI9qgDaWER+TlRy4zX3OMYHIYlr9qcreG8iBwTzt14mQNkALLjhhMb/qDcw2AI7Ye2oMtQD+ExPvQvUuv2Ib/kFIDAuA/DRSnhxfLgLm8zkTOPWmmg68YukMlu9ehdojDy8DOpFnNcUXBdRkdoVVyN5+vOJ+WMERb3RcBMNTI9bgoNc4sWgvDJtnNumFgjBipq00ylrHxHUjaqLxWzn2mbClC48lNVhJQ52JnCVp3m6A/CKQbkFBKgRBUU9dYgLYuxAEE4KcELqTUCYP3q4VlN1iMwvNXah+u+S90byAdc3u22jb9AUj8oK6L57nzmJDs/2sAs62a8lW9Ev3vw82Dp7xkVc06VC4pReZ/BiZEPEqhRxAy+m6XTdLIPafIWIyIZDud0U/Cfgr1yiNDegc9AK6RgDJ0dM3ou+pGVF6DRbObebiwn9r7FZtbs4quXOMID0PV7w3MqEI6Dx8A6hDSRGCJ3B5YhyFhww3mXOmdBgqL/buQejlqA5nQeXyiTA/LLvwUHGMF+h/2U/EAg4n/zTcI37xcZq7TQr4xOD4sMd07kRE93JT11NSUpWR/FTQUc840i9q3F/NPyEcGOBO89N/YYKfA4eiBsfAuliXdx2UV9vsyu/mIdG4KkAnneUxbz1VyQmDnZVkuJ9RU4hQLW+JHD8iWpA/LVdxZrhiO/93BsAU+fpVcSvex/UEdxJbGMkSnnJQJsn6U6lsgYLuLDyfl6pb8L/6Y8DQX4UvVcie28fgS6CZ3cTfoKswRk59rA9P6FswLKyL+xmFzpvbB0tzBj7ZHpFXOdVsNFDJlyFM0APFFjskkxoTAmCFaDcR/WMIolL56ie0L/Eu64qcYYlSkeLzVgJSrqO14JFiDv90hIVtlPcUEzp+eJhxn/W57TgjSnhfPlEuz1wZVhiGcUhdKilMvb5vfje/Da2PB1TvIAA/1pflhKB3hia7CvIggtZhwq6cENxbiFJF9EQ7xMgc/J4HQ+xLpBY6W+V18MIN/bkZg27uVJw3gkWHrjntI/jG8QEx2Frvs8uqu20tgQS6ROnVxL55uU3DpMI6szHvWVqZsELhurPP4IODOhsEg5ruhCDI9vPYF+jeijUjd7Ema5AIf/ZaBdvEkZ78PSu1Cc2Ab9uEkgVEBdADKD/Y4KpF1qBNLG0ZbHxmww+Fap6YAaFvJrHwipMPq8MZLVvtPJjZO7nm6X940XRa2fNcfSCguG44ObAm5D/rex1XJSoyf/wlUXwFMuuMX15cZC6QGUpX+lj2oat58+kfMCpXqUZ1vvzMpWkMNClRlsCW9oLh5A13NL25j/Zuglr3l7irOCQRMUK9LKaqhliC2JFP0gg/Vow1E0BuhqSN8UOTrN/xMtO42VAjjdlxq38NA4dg55Fut4+8rf+BjbaRk0f7+8x/qla11H4MGQsAA3cZdEBkU4u3j0m6CrycuPUXSXlIcT0D6ChSolYvyp884GDsbK2kg0uhPSpzZUanJLyMif6PHYErs0GHOX5n6BJGS4b8pmVqSvCSyEQ9UCy7ekTrW8InPMNPtd4zqayz1/NjP3eYJoQT4n2YvKQX6M+fno8rpaDBsMGjFkL9UXHVREtWlhwZv/yZI2Yi1KzdPKHNK0/8znh97SP+MwEXof7rZ00F44T+2S9AQ1htIdLrQK5rv25Burf/4MC88x1aN9sVzRfsigK3doHQj/V5uIBVu8mO5UETKWsZOWiUBWWHBdOnsout8/4zj4S/62HD5fxhA4LD58+/uZ9hxp+S6IZcepthr7HRp7E5ZLRyDQkSvB1MYCmjPmlqZQg/DbbKGDV2XJeCXZHB9XikL4LDNjWW3Go4mbkjgkbtvK3tpEDljjTfNbh2NJYLefqlQ6PYUFGEH8c3Bogs5lUyiPrP8tT9vY0cdhILDJ8XgOjHn6BphhdSSgeiBISDOC1Csk+W6PT/yctaioqjsRxHbb0GycF80Dl1RC4yNkspF54NEKqE0P3abrV9wGEwsDe0qSYwMi+ZOG+g9624L15bwJ4s8zUmFWwOzW1l/E50j1NHqkUt05Ku3yMayPpNDzUC6EG8qf4dlO56NVvIKyWhVKrlcpqH9/xRUpyRrpR62DZvLtbrGEroQDscnT0UBtzHfMFKN1wJWj+cUkORSER779fv9dH1Vdb7zRZ6/FS2vOPhGG8b+SfFrLNCnuTBUOs39/LRpVt606krGcaJfaN+BKJPDgUQSBOx0NwFfcbPlt8FjgWZxjb+W/taCgkzw/ssDdHG5R/jHcEW59wqP3GZ6BcGW8CJdqtCUO335R+UpmrlbSfekrbE6LR+bQG5XHhJCQ8/21QcXR5CVQtGEIMn6I4kbDSQK+ZM5BAdk+zD3EcVfb7vcDumKKpFK4ka/MlQA0AF4ksw/byI0eKAulZ1TSiirHYTqHepMhcC9BuWfdMFrSo1hjzm3+Ovq3Y0icwJH82cZ4uqKVQ5H+Hbyfbul2hwjTPMF6UCoCDhEzsQj8anOd4+bffGQyFrv8CGddvElMuKNDKyMwv/UDFURRMDpau30s7nSY0U6G14QIRS9ZTlL6tsspQ1thBIz73WOreigXPp/yaL5ccgA+icYnJ00c8X79rIjgu0VVqqz7SQ4jT8j+OHyKdNlBil11lfG+lIxYK6X7R7pPmY+Zgssy0ggGx/B5IRjDHqoUVJwVZ/QWsm1YWod3BmBRczTKSPATTSkp+6ygU9LoWiPZ77scuFDS53FB6VF2D5HV43baqgnYn355WO2Al8hk3SUgoxjC6Z63YSimG+JYCrnf70z4t+J/73ImSAIQJKIrNdUGS7uvrGbzli1ksNyPdIm+rJfeivK637XVtdLrH1I5evx4pi23MWNRqLvw1ibEbXRvMEdvZDbYiqiv4EMPu4RlzCXbDkls6nhpQyVnF0U/3Yj8/5lbsXu2P61Kcz5Q4I6QO2g1DhEhVG6ZolZn+3WJPwlN/O68xMnA4oZEyhJdqfvEknZf83y4ZykJsaf6uqV0XzdG9b4Hb6TVtj1mp08ST+ARhZUDSGNOA+vh/J60DfrRPMsI14iNA5ITLVFCNl9tZI4T25iEJvqHujKT8mQx+muG2zeOxgVP0sCgIZ3U4ObN1TUu8IhvPH1q0lrDxMvQt3dryh64BRpOAzyo47HSmUPG/HotRugOm9MPAasZhN0PkUcQdtJF3UUG9PqJ1WztMl9Zbs9UYxAONtfcO/gZ5lIGUqJmmSZIHdyRuvjTvDY0vdVR/pK2gs5svybMU3zQXoYzcOzurRA6co+wnLKCjB906OzytxF1WZHG29U10kKTF37oXFudaPhRe+5+HVlxCzQ9fweVK7gqHHfKAuuGWQalXuar8bHffYLVAvj2fSqCnFAbRrU/ofN3exH9ezoX13IC1TXNhV4C9htPcUfFKbiysxaYWuR7iFV09LORwlbNio7MLJUkjD1oUs/0T9aEqdl1Ao4Wo9rtXNliogDqgVVAZiohDVqDfVHRQ5V6Rzpd3T6rPl12ck1Ytx+2foCBmfzvYBGlldxKMrH0g2OPxlNZNXCH7vtXFmVVYCc42lLVUqivjuQQRMgkmOZNaLp+tbfSAZvg6bR7tJlHdX0nrehaBtgQE2eh4N08jlJuk8KVoz1ZKMnJEVWbvvBxEVFmiy5h6Xi0TzfL/IDdNUVQ6kORX9kRliZSoXv9z1+smr1VAECARhmoxdt57PzccoFQ0Baob473Kr2QTOb3vPGu9xtGBKmviDiWHd1cV4Qy8GD7bZvfd2TA23+1cpUqJCAeXBTb9jidXtIl2iOsPKtRILzZyFrH1tgnE3G7V44LMoiPAv+CDMDw8zozBLgvy1W0A0Er1y5PqlWb52Ii2Z+LcSKt8LcXiumQ0ZO83Acu/uXDqHAg0M0IHT3tGkCGLbXkDaQK/8/7cZAB1IppdPmwl8A7EqtRT2FGrm101cDXBpb0YrqFbl58Jw5DTKzAHohV6up3tuhY69PlqNzmvkVkFvow5xoLfwAPVTLhHgnY4WTS1qvjB5hYVSroF19xTCdoryjQCu9dOR8yjKhciZm+LZy2sA0VRylSMZOVNZZ2zX0Bq8jHiuoQOaQUF0Zt516tLl8sWSpCFhYpd9UlPeAi3ventUfTl+q1eQlInsH2ZZ9IsWhwux7UXCihkSWz29vWxDd8GV456beI7O1WrKofNCRTZQdrnT242IaQ1mnOLexsNtzcS/yc+y7Y8c5tyaoH/sIOjBm1Ei5VZ30n3eEcO9l6QFOt8/z+cglKKVJb/f5oOg0W96G6mPch3zDcr1YfmZ7K8eOzRK/2Gk+BnnuSNQxLLSJcpVeGJh4aCcUV1LYdbnQmAk7VksAkOZdJCoH/gEngbVXJH31zUazTGkukBw+rpWL7TwXk34xyjN9UvIheb8dgW5I8gyoAX2a0F9MPOblWwulAf2WPaH4IKzENBGSfZ68ElcR8Fqio+ebVi4tMU6UGOzu8nzFKJBxTqkRCjZJzHXmNxuq06P+u62ipt7Hl5rkxSpKDqpCC8j8NAMbPPhd3WlNlhngDw4s16YibRPYLfgLSvgkQxSK4VYiK47x2ocpqYzNFhfEIe+vTuIUG13gxkSBcPlDo1TrPo2GTTaQprIsleRIvkaLDN9pN4TtatDwjp0Sn7bWQtSLtWgBiDHQ+W4tC4FF/Ls+lBKEb559quhQqxEMR2Xrpgy2zCLDNro2Wo3xtvVexyOHS1yrG8wQvzNYiHrjT+Az4i7Q9hyBj5nqongoXyuAT4C8UeO7J8mdz6BIr32ffT42NsCQeWZxslTTyoXPHVicSb9ctJcwIyO8u/+e1HS26UZoQm2LFIj1MfVY/qALAuXDYeUVsEEieqfu5yWBt9axIA/MuMl1cxHxwWxo8MNWIFvv+p0ZFX6IW4Dbz3tPL7yXAszp/ohKwiTvYx6uVlZt96dCY70DY6U/gmYEFfR8YHGqst5eJvhP61hZu/JHCLD326jygeZ0pdz/I9Ik5HBPRpIU/xai2bM1s992oZuADrEvn0dBrlkEj5sP68Uu8Unkc5yT5/qSlpdVC2Ng1hNlKEfpW3sfYqb6woo6DGVmmPhQ1yj3zMcto3Ewets0egm1Wehbawnar//8hRiLn1tdAWDNWFz3XSvyrfReMRkYGuvvrJWyn6QAUXbutpH/c16IYhqYsd+7nAhXxUd+JN2Hnr6ubTCbv+XbJED1VVHCXVaUeSndin/0MlwiTSvF/uSx/st0498Te3PErEl8KJ9iv4nylSdLhWRiMpv5WDS0Yn7ia2ui7J3Ebol4Vi0wAUlhs1wCTcyEOfxjydJf+9bZMjaSDC7GWXIXLPDJ7CNbtn5BYmN0xZ3nAzGgMT4XnYcC3uqYGNkmgFbIsU1tvmRX8VRcIHBAQoMLqUoheOllbAIXeV1CrsfasFjwZ9BLEM8VH+xfylroWkC0Ux5RITtVa2WWUkkpiXCKWIFWb/Sim53pRwJ3csHPfSNSk0J+uaneIuoa6YYscQ5L4c0n+MR29T0EDdUSop7wEvdBSMhYFxaLnH/tc0P90eIgCvlE/riKaGGQ3eEoxi91Z79/eEQqkNP6E7Dz4hfP10nMdHjkNkax1C8W/qrRuUREMzfG2aV/jjD142d1qKbjAhd/dv9JU2+dzRuWNmUYl/siQyI1r2ZY4pbtUMoBzpd7bDjk1tnwcPVDPZHJfk7PpP7EfpyJzSO+5TVqIECR20cpxEKbeP5ooQBCJyVxVa5+0YFsJxbkkDoVSRDQZqQufOrQD3JxHIsfYOHQmRmaNDQz13/spHyk2BYrpRJE2PquPoJLdSi7mrmKaVV/r5XwHziaQFjS7OHTDh3SN3xOS55uHFjSWy4mwORu1Yv4v8sc4gJxz7BDRWgyWHgHmdRNJY0ksRC2W9ceNvo7CYzL+z+nZFLXCE+JvmZ5PL1MRjJwM/itk6ygF32CkOhbZMee9SdBE8LcdFa4tLs0yKYerxoxf+xbGzwy8+CQ6eNvjmpiX5gXSrRNTvM+rSUG8/an8kR2561TWuGETAOnl10ymn/sGjPQeARLdCn0UGcOTnahCFZPdwafb/zdGxExf14iYqRvPtmOZRmImidLfTMs3RhrVIIAXK32ELlex+87k+Vd+OOsvrAF6Hio+TkxfNmbMMv0whlEsg40wxOUGJickXQ4wVj2aC1fGe7nrDXfhSuKmv5UF5zwGb8lUk/fEE4XSJa3J3ZYWpu2XDadv1nmhvvUjeqTa3DxCGcVVTH82i7H6zO3vcbs6CIAHRgSVwjXddhwbV1FBDODS/5TMeEYiDu5fYuw+ad6WsembI9d0Gjr7oC4fLn3msZ9FFgvz2VwXjXYa2gwJRiBSSKLO10dNAF2WA93Mf3NGZqjmFOpRocivYB/LPktpL3rq/zhpCeWTc9dCK4b3p06o4IdffZGzuVLNz7nSC2NET3fFqLpIMsaLgz9fxYRd7sjJ5gmOZqHDgkj43NhANd/E0OXb/ujaQQDLoQkvdrvnEDU5x6yeK5GTpB6TDjLiPEMLt17Gv20ormcs8yfVk1Bjw88uc/qEM9QK5sbmM0492eqaM7TujZjSqrUqNQGAU5V/hlgmH1r6cJ67ZloAWYNzjQp9NvplPW+0uI/ogOZf8hzfVMgp4FghD8tdTQUzclCanD2OXw2XMuwftjEjCUIRjdceE4dpsExZXFpTjo0PlKgG9Q0E76aAOqZoDMsNF2kRpvYKS/uugnI4egwyWXEzP56SCg7mIRvSjvunuExqvZ7W7vd6+VH6liwPtFAqUuYWiAPX16Px2/SS0Im/g9RukGyg4gj6jTR+E+nYivACfhs6kPg42WAbne9ILKKlF1Nh3D0EFDvHmr1elvcel0PauSq/F06QA0hXkJIS1p7l/oEqL5y1wSO1vkwaERidCucxvST/fuiKmG/WB5jcQ18zR8DAuY7C6GybdTAhrRdCsZP1eEaUNlA6cPhZhnssNtygETSnUw8iuDjtl27Ea/i1B+7ytlbXREDlTQQZ/wh701YyoxkxjhRajl1nfvDSyd7DXMnrDeYPGDRwH38KFv86y4F6I3QE7POQUrK9qyULL8nzCgdTPzaKEaYVTEu7f3Eslbi7L9jADLZNgxhex0LFJtj/4gyYuId1+/tqads5j88R4gvy1ais/QkBOf+c1LYFaLkN//+kuLlWvmrIQnezILo3CnPpynUmLsB+Ts7JGyfoOl+i0cc6uJTnI9dmDf4dVVnDLDYQ3+KpUbDPw1oC/8R535R1eJ9OFLcb7m7MBvSy+DBL1yoFnD89t7wXvKbFd5P8fcFWZo8frUzPFDE7pkUj7brRgXvzNheh4ggJuavacKeenPVxx4u/4GGmjt9YDd02Bz3H2O+eJagh8w8w/wgdXPM8HSIFIoEkM/zCDd57S8TfBIrWBJVIRCehN0amvxJpLKFlyiCX+6Wp5IyKgXtagzUaYUDJYGK8Hg+2HebJQxAvQV2HdLSN1kOxFitrYFBAk95eVxXM6DRLuXYKYmrQvhLmdQDgeflcuiTBnVZNZ+8Legt/9cbTyznllkicnA7VYzqfPiKfGLpycOykYWBQ5F45OVBxuDPFb5Q27cxhWKJFjhp6mfV9w1Ninv9LG2+7femO08ZJS05R2ULmuwbtS1eo7GcI7SDSj/GB+/wRRjfuouamnaYoGkYE/aldbeRj1W+hNH9Byp5oJsBOdsdekj1odNVPOJUhaws6vOK6z3JLybUZlFag4AYy88GEspURV0kT7f6ALhVKjWClvuAr46CSiXoW3EsctRxMPi41nPE4tmlePRccR19r/JCTmkd3ZcneRZqf2o02WCxxN8MGTJ0we8CTbIUwfrURLMeexF9QWiD19zFH413y3PlacZFfAkX63Ok/O9RA+6pO+N8kU0yMRQLlTeQEbHm/lnIdfdTXQVOVOb2DWAGBJ5PW2Zbvm3qNuYfLJQk5MKa8Ewy/+Gqz5nBZb0+u8hT4s4m2Rq7amF/NNri/mZIydctU6ciOPfIRQHMTmSoQiLIvyKEmdSjWRITk418W2cRstpTafsXsuwb0kjRNkvcVCbItqb7WFawu9Cyw9AylVYd2WF8TI1zTwykv3Ykk2opd/ojX4nwptpgvmuT2/PvBXkKbSLXb91JOafJiw/yAnp8qxjBe+fUO5k4V3utKvLSjNb+dUXW2oiWpOBjCC99advUmHneh2edBBxS1394EJ9pwBeAb7Ex4mRTZ0LDx28/xK+NIMjszrMg6lYXhk7a1neIoXgQeYI6VFawXKKlglLkmmh6qKHIEvGBK41lXg38ZiILByLx/4FmNOw65bgIzqv9+MgLooRaNIWS+lIcTfv0LwX2RnbLOui/0XzBI0SOvK15Uiv69WIEXdU4Dj81Vj/YwRt35d4ugr4bjh69zLnA0HEoQnEIoLlK8mWyAzaLd1yimY1mAUkOUb2rNduwOyLxO31PQ8e3Nr9EV0DmeXZCT0rhJsUrJbwYfooQ9DUgJct6eGBSgjyf2PSSN4kzt9TCaV3ZwDYo5sJ6avc+ObPX/h3ltbr8hy67otOT/V6Acyz8s+k7Teh7NTOBo3gS2Kzkfbzq8ituHb/rYj2cbHglKLwRS3fTvyN2FmJbZa8kf1PiHxAcw0LSGm9SQo5uLffWrYLQRQHfY+9iXg7IQL1W9EILoj2SJ404TZmpCmtwJ7Wnbj1v3ubbxYpyj46ythTg9umpwcWa5IjEr4mW9YAGno79J31vjraAm6avJvcJE2MK2YSnn4GC4JL/lOfP9UpobY1cE1zrXuZ65gE/NsbpWAH6ZEkqaHymHpXFZplDBLjKLu972kLeuzY+pxyAmD7Ani+8TU5lrluUDk9HBm0AuOJ91tbEgLHlUuw+SGdRLN2DEJzPUSfhA04jsz9YUz5VAt5Y5mfm+nTJN9CxBIIFHwDn77XTU+bVo/3g5AVC7emtfPEtdtiHpdyWuUc4m45sAx4AV7Sh6b+LIPsECyOqY8IkMsa3t99Gj3qwenHaxxn02Ga7MnCKcRgaKFsRxqagov9euLy1ne1TE7X2E7EVyEibgQFUFkO2yq6BSEurRviDJS/+R1bigPd3QQScP5ESoXyz4cW9Lq1aGHR5tb6KTrGw3Qb3ibfGvbUn+3M9Rvf7Rv7iIzm25u+zX5vo5e0U4VZBFVtoLEeLwxxpF2l/9nl3z62hVQEYYI1PX95JnFi+7SpWIXuJFJ0vUQyUxurKPyoR252cX0zy93tLqF4gyBvXbhOesxtgABSNiSheLFa2uSoBfN4qdruXCiYP44Z9xe1rZRWBirlCowsLFCKg53ybqlkN//FEDXpUtSsgb1xHVmX039fvH6C/V+cpDokLN8zYoUkqaPQaaBxIXO31aZ+7pqXbVXVtypd7LBNTjU2Dj/J+2bh/sU0BF57gLPx+hEOybptzB/aS3h+Aeu7FhKHhtzxAkwroNE14FkyvnoT/Q8jbQcqg0nAcyEo5jL6wIlnorhsb8R8evgfe3RM3NGdrIX3//0qjPBzDG90fzXE+qpuWb+i85nkT0C+Mk575z0K6K3jz/oQZaFaBJkod9u0C9t0ipWvd594monrVr04RvPjYcY97vK3g7r0s3E0Cz5YE8FaUzjipoHux5crcKLBAv0XKEwIMdHGtTe/p38O2XfB6mqn7VBp55ApGo2XjLBeGVJ7p03xv09jQEP+nqrFWwPYOPdq54SQXkS6krlvGPKsIXimSAFJqqFnlDYmZnkKfhPzpjAFQvoPJKQqVp+nQ98qGGp0jPXOYtJ1O0cCqTYIpNgJ8X1+ZDLYVgiwEFoUScvaBBDcS6tQ2LqlzbgdMRvOBTDpUZY+YmAKGwgfPf7dD0rxTzpqwle26yWkWOiHVZDW2xguqhBIxoiYgzd1B32DxIkI8N+ZX2FH2SKxDjHYYbxU2CI857jDQw/qrN2UvnyHrQ2or73pULVWCVwj5Wvoqm14rD1GtFTSpGsYIcULpURaqJhGiAE/umNqPrHjTJWkbL+vr+plbr+Ysbfm+msuz2FS+WlD7h44Zaxg0oP1HLoAq3QpFwpWXGdutWMbdLErWrxI1Rin3+W5OCi55shZhZf8GC2JCAyYDk0hIlCZrgRPrgsKiBko1AdoxFeGQf1PmFzEzwSPc/rs+kBVUlvInKnJhaFZ/sT4O86lGqRfpR8ik5AJcF/WYgZQ+OpPC9bK4toDtpKz8/p1ICAfF9+M9c7QRrZk64fchSwnEze5x1y3UhCak5X/8f7NUUBv/tqN3DyeUefGJ5IStiMAKLb8CaLUT+nf7CZ5m0aO6T/43iQy5IMY7+gsCBEP1YQKfLnUQDAC/vzTLokLCItZmzQn4u7XlCbYpGZfVHCD2gfFXYxKkLam+q4MUaEAiDHJ8DH061JH3+Wa6bpJ66StLt4Its+zLNdYY2bedo7oGWI6NPtlioVkWVHw37LiNZQd0CUOsfvGSALfIPUOkRLnjAo4/qTYOt5FE+GsFHniuASotukNOZMZSTnWo/4rOGCTHfAWgKbKQyMi/M/cbqfHYlfP1pdqzRRbXVWMjU8hPXhyOVNrkMaFlQxTlpaNHs6NNfV3Yn6Md+64bwHt7iB9ndW4Iu3M8yxl9QE8VB/HB8lcgZ+ff4TR2s2wYg3jL0Z9WLZQS6DR+6FbYe2ND19vR9yF0u86U3gn51hdi8yTrHrYfDYzZyaaJCs+prfynwLWNjJLFbhoLrTILqKzbI3FVQ03gtKP4Nu38en0XVcVG8tAQVU2s4GVfKtGBub7mWlauhamBz7dovN7dFvDg/BsjFvOtTrzB2YyohAWLb3EJQxTJ/5jPGzjrQ9/AoTFdWVV7Wcjyjpf596VEjFJMZiKHR9C9jKxDuOUeomx20L9dFu2O6qs5mAb2o93EQaMsUDkpeteGMA0IKvBAv82A/D47Lt0RxUI6MJ9+dQtgFDDsjODRq4lpnkiLIsnE1WKwHFGsSJTxtrpDKfIibT6qotrh5gxaI242YnwP0m5M44o5yi1Hcc6vgK78FF7rtgTNUvkcB4K97ZLW3hs5KngXoMoVJ3sIW8sr7gas+1eo1KtLh7d+7+NqKUyjk9u7Va5iremCLaa10JZcJUlaNTxWNaezwqqsM6+C74VOUeMKSqVT+dc1mX8WbYxieHWpZUtPUoM0Dlax9/xqcBdj2Ais+Vh9GGJ/xVLJh3sf6ODs1KBCYTzanAXIo/7/aZHeXkU3OCEgEPTFKQd3g76O7lZ8YnnnCbj10mfr3aOzXoDYKGNhygf51l1O4ov8hWBo9KLEoH56Ui2bnjxZVT/xP0UYnmRSJZW3NTfyz0W1DmjFMtZIveEhqBcNKNjGaUePuafjsIzayBvnlSi6b1F69cxTxW0MN3nfQS3m2xoH1r8XhQDPG1t+MgrvQO/wn4D1rK3rQ49Dqa9790yzi34Arlg53aiYWtsxuO/5YIfWH+xUwokXJFjve3FlsA6RftnSx7d2RifmpEmMdyF94qHlmRvF1ZUbc3VPnPPktplhmWBKgF18m9fIdxUvg1J348TAhWO/7A9wTNmrN7h/ZKjVb6sn++38JeGT5EM00Q9zsFpiN3D1UzVwpd2Lgcb2DlRIHKQaT1QD8UiLzBkMFNGMgF2wXIDqytWWTesT4x52bvVD0/G78g9e8oLnkgvFIX7F9jbpQUATgta2OdQtaa+jha1/JeaeO4t6IEtoLpPOZ00kY1PYbKXMi9L10Duxa4MJKyxmrKCnmPV6yZ0Nz0+0eLfCdadH9Em8c4wZtVjJ0hZ8d4TZ1hBdxVyycVLoHRBNdREooXppftP+Kv97zLaUvSP//sd75jKuH2Oblsyp7CG/abCknoziELYj5Sf01NCavnn2Fu3jB+Nr4w2URAR1Hklafn66JXhSmEY8qGjcTPZqdoahDbJnbMRz/riS3r8obD2RnqrF1idUMqO5ctC1E78c0UMZue4PZlozgJyJzquoWrc6RBojvDj2ENNYk3gyThWsWEq3krP4lvXijmKJMk8isnLwoUQoR3XpwiOwsa9sLZyvrOqvNrk+0lH23xZnb4DKDZgUow9XpOQN3cV9tCddIukjrUZaVqgoydQkiMA3pCa0nuRs4KA3fpYmOfEAkNvCde0R68s80124wx/xXNOWa0IEudrI/i0G020ivMRHdTd+1yfapusqBs7oUDwVS51iXYkLLlv4qvHOttu7ExFGKrlzRd2IHv4O4BnYKkKPkOcm9cvh1JNxP/g3zXt2mZhgfDodcqsvWYdK4F5mbF1EtfBDnp+J49Xu/jVreveF60o=
`pragma protect end_data_block
`pragma protect digest_block
a8178b8c04bc63be150f3195875e11c8eb557030d33e0493378177a28cde173d
`pragma protect end_digest_block
`pragma protect end_protected
