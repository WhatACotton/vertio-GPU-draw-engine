`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
bEn99KUsnFHQG+RhzfgpRwu0aucnHyeFC44YpmGU+NyEp+FICBqdW1kD8Hi/69zoc6s7q0pMJdrc2q4PXSdRZK6j5iJcVLqU+/nqFy/qtmPHOoKoSITuj93vi5GL74MtSae5L2BB1Wjv5hrHTm6iz/hyc6lS/q+WI80a27B6xwic/Mr4HEyRZZ6DiEXlaYfuE45CqZPqheBDyg6bXBGlt+kwX/1SUhSq0flsNvy1pY34w4enu/p2/WJlpYABAthy4/+YjwXDYZDBq4FXCpzwsLyx/ZqoaEBIQlwNSYvFfU4v+Wpwh5/LvNoSwwsDxwAiLUEJEtn4SS9lYSxUEQ29Yvok1UTLvXoUdI2hTZqSWv43n48vKQho6f6k70HgTkX0AjWIYPR3vxjTUVxK2UVbqvsUF1Cnn1FD2KVn0HcMoqHzvmJNHAB5AgLzdDvtqbyw0OeZzroD5w34uVhSt8KPAXDeYFmGtkbStX4k0NRVfA3F5DWWWQg8aRAPDVepM9WZw3tsJ28A/kUdgHrHK+7+ipNQYhVwk2UpUzlq+Q0PVv3tDP7W+mhZEGblmNDmyASNRum/OHahuGo7sTejlZLGkoNSsDDjVdGwA3NNbiF7H2lLuT3DXF1+25jDH83QinbP9A/jIsndmJRSUh+ER/NgvldEknrM4Y3bCcEmSZtMWv2G3uEMBnBIYMwb7181CAjeC/iVp/Ou+RlVpM9AEYmL1gpdOGxyW7UiqomxVkk2aUXkwZu/aW3T+PG1B5jY68XoSlxfVXDD8w4XvfjeHwgbRj+WCH07G7812t6nBmonXrpcUfZ2cMCF/ZNuUyxCBNlp1srNeMFPXGtWUCRe01SqT8Yg1+TT0Ref2gfYbyLEGtOKlpZS/AYmYZZZWLa/JTbdZPjdkiJkfsQ5QVy+T3J1Irr9oeO60hh8UmajItW21bvvF7sugqFFd1K2ARQYtSYQX8+11MIgN4RAhU0tG60Vb6Pu9ftu7Nf2jzgz/YFv/qe8o6HJz+fhgtbI/v7qezU58rk5ObGKwJHqeGG/cShPYCg90qiWaAtlNAWU2PNaxVBXXyU5FiatBVkOjrA1N5pjF6JwNMzLL3/IdelwG/L6wLQuVjKie/hVj419vx0Qb2/Mnwac4XphxOzPzr16knGzBr2KmD768G5Z92cBGIs7Cl/KsdwtkTnpS95b3uBW2hvOG/DYJJKYzxYt5u36KRfoSRDzqYenKYUiKpSFi1zUlhcEb5cHA/r+K617z9g+qOpKO0AdhEPSyTE0qsIoBctY1FY2kSM2VtpbgE+kqaWozkDOkbP3Uuw6JlFImOUqzNrzS6HtmVWMj+f4EfMYQswZ802XCoWYMh+V0D3/MgB5aIgs8YP9hApwRC9uGUuPEzfDMCQoYXd2Da0IDvA8ljejLlXFDK3mSo+WdVe2RORMIXeqJ/lAjEZhIUpigYZvL0NlNbAjYmY93ZD1Dj//PeV9yxEL4PmNlqkY36lrBNWpYkG0o31pb6UQjDhOJ28ZJE2vcpYjfOREHdJESo9WLtF1Z7wRxvoaLfIaDnd9w4Fx3Qo3NgQOh7CNZ+//TQTzpgRM0OBR/rb3ijEDW18x9AXbww9s2bUfU7ytaxyClLOnhVho28FnqrUoiBPFIpSE79pNOKWEipMA0QUwR0nN6SSHbi56bWrAZsNl5wCkU4ge28zSLh1fgmfRchMyayfB6n6VnsO6pfudEjw9ouaPG1Fy59lElZ7nJNb0wVguyYkg+GfADnPqspAnZ/WYne1+NIXzsj1Epm9UwVDhRr1jSZAr5G6AlGjBCyqbC576eOvYK3j4g1OCdbkUlDjpOPvRNhbbKQ1GMSjJlJK495e/kxU1i50wozBlOQwM3w0B5GgIZpEwkrlx1Zu+w/6ythqbEtcoYvd0NqEdYsdXRQmNd44E6x78Gh2NMMK1cc20/8MfjMIEaB5bgYMKg7uVrYwrkAQN2ALKfVA0i54oit/az/DVNzVihFmeMaWUW1s5fiNwdiK0TSsPekNV251Yml6GYziOzf6MW9dEgzaH+nGe1FAy7GlLtrhxi4VSyIzabMos6rZ7BAqlR4Au7I1Xqq1HGBuNwYFYskej2B333jF1rqBNsF2bKq0ZDYR6iL1pfb7+3YjZk6NM5xuiIBzfjR+ysXbjv2O5/bOoox2mow8KYgBcEJh1XROr5mhe4lDkac3N0AQwlKp+CM9zFiIH+nUF/DU67h7ggiR17Aaro4L14agx6bPAiSq99KrvGikbJoYxHoMA+I6W011NShhmcv/Ld+Sj94/+xpjcbnbByuJf03JidbMRjOM1SuoyCW4NnIdL3kwmjfY7fHZwE/LN1fuQBYRaXqa3chClKCndJGKbLWj+5mqjS6F8W1D7BO1smPR/oPDpdFAC4zJhm7h0tCF3Xwk5ScEnvykEdeiqYgz9XSSd4o4GVFgaunylG5MJ783WhABaCTJ+UzUQ8j4KZxY8JWqXaQHOGR9/kn9ClQpwJXpbblOqnKg2c1wP4b31RIWm2RVOWc4b+MjalclXrrrChC7vs23RYH5VjHAnS4rjz1l31B0yey+1qnnf9jEBLBtZ+1LimVFiFeciccJe6X0CMrID1LlimHwTt1stqLRPFrz60fWpaxos4vawm4WwI/UeRWVuJuE63atOWimjkHHsLi72FNuwlKDd255gV+eFYwyBnleB5xe6FpMpJ+XyErkuSfSfV0RP1i2eY1slw7KyMJOK07OUnPN4F9CLuVSimn6kjvC+24QyqzP/A3yujEZggycEf/XW7Q6OCdOkq6gp+3ruKS0BgCxf/IsMcRitfX6tFAxVZE4DxoUI7QvLpW3KkIoCYL2IHrI4LQCm4cX3DvZ4AFzAMHA6NJfeCkEvNlgUss/hgmH/DONI9i+B0uoOooKPNr4M9t5GZhPgzGP2tGMUQKt6+GBue+UYXwu8ESbrxiGl0rs6pCR25mYRBI9YuK+XoCjyETpgccqBReMdBH53ATT5UXq6oI2x32wtuxAU1YjcLsHultEQWRZbKdNsfBx833aW6ryZ2Z/amRQYBs1+AQcV2TOlAxyneV67q3PLUzwixfdR8NnSW+SQgZRFPEsaFgbbz5+V2giwAMJITVv95A3f4atVLbPmviuJ+/0wWlSyA7+CcKkCRlEyYp2n942+M6CqeUGbmHNfwpOmPcZeDUyGCs8Wy86xtAsX/4LXVnEBKij8DvYeMgz4xzE/YgYGi3wUjWR4zCPijxlzKl8amD255Y8ZeTJSzLHkX2juTiY46DlD9vNP6FxnpBQ28YyIxFlKlaiMzJj1aNZ2qEpeMudDtf1sRVPMUEBpMRlmFaLTcSb7NjhZ0D+kzjipob8Cn3dBEmifINCXlKKBUnyeYTtbFVK67wkYkbVpbVA3Wif6LDaai9Ry0Ld/QhkqOJ6L+NnjEMpLLUdjwvleaMlF8h+005DnHTJe1OMK+9AHmW7ZolucwtDW4BZRBTc4v7/3lHhI00kpstWXWrSjproBP1+Xe9+wcXeqBbuGUg3swFYm95TkbrTs8AN5A+U8ytvTYa2EdTME2WnVVchgq5Ldl5h/WfuoF3r2Nh1JV4YpUGqtozWLiGyjk67gB9l/GLIcs3DCQAeHkD1p6fHFh/MpRWEF5buRWpXC4FuxhZ8LJ0zrOl4nNorf5V5ElDxFfeZo/n9zDPmjK157i5OWuN4DuCtUS6jrssNHtBWF2n0/8a/BOYuzEjhYsT0lSJJKHdk+1fKyKlTATudsV8XzI4OYjxvyPU4L/rrrO+UlePmMQ0YwSM273njIGmoGB2Cxuw7Orski6u0W8TnUn3pNyxgBb/VPKcKD9DNwQFOOBaxsDA4zDhNN+Tk17dD81mSz3CboUjBgcyo6dhDmItKMG3enEf/d+EAQKMsH+O1/HwjKuMu/48TOVkV5fgb+ZpkgiQ0waKeWPAVF4p1IyREyGi1VoR1tLn9F+sVlFNfMcTWMpiSyShE79FOBjzAQCKC5USqeP2lNSj2n1qgcJY5LFQmfeLQvttPw/Y0kMMsZe9PeAT98y+aYSfq/g0TMofa0W5zWPH8hthOf+KKk7LW0Ryo7hKv4N28Qpyi63jGXgFl6jLPuI+IlO5b32mQWa6KLZST5yb5J1dGwDTzUMceyRiR+gkzo3cjhaRfiwkD9a487PMQCtFFFvOcYCDXrgEmBsSBOrpVRKHnPu9BxTz7QHWRTh2nbQo44uncgBWI0729Tk6e1VnsWBE1yP499B1cd8i/b2Q96W50iFdEl0Wckwxqqv6gfA5wIuKqcUsN9G91OxyG8tb6FHKgT0XULbWoABOr3jSW+z0Rh33VmKCTMn7wtVeQ9MI/Bd/GL6H0/zVIXYnyskbXHx7H35r+my3+ewEAni9WNK5r/EQoUIIcaJ31p02Me+K2xuaJbCTsEIxmDCg+pORmkXhf2+JYxy2FvATZgUNbDfsuxHfpYP2WkS4rEuFyP8wkUrspWnCRnjeAbuaKyL/eCI1cOOL25pLKGdYjOvnmGxZ4MVHnfz6dPylhfoODLJX/ISQu0jLo703eYVnTo67AYZL3VTmB4kSMgjmCstffyCmlUdUpr5Gd9k6U5URypXJaYTVd9sZvfj4eZ8dRtKeGv8kefcp7XnRd+z7vY7xw5/ePZPAee/RALbLJDjMQjydTJJY0EpDJbW/6T6ot+nIHkuCUNbnXZlCa3QsbsZbi3XuUhoOYs7xmpIAxSnoU12RWB53OJWaD7xNV2q4jN/BZ/Lm4CMKKZdydP1XkXXv2WR+XNsQp/bVLKRp4oHGw7I4sKEVbUhP6AS0DnT9vpjpQUb5t9NjxnCrxNOnkieRrvR6jzqT4OLWHVQPyHnRoPh8yZ0wK/3M7ziRjqrQHqBxrtPAw6IR00Wykg4ZQ5WmWEEBlNI49J4zdMFPryH261/5/TOea667O1buqxbuvijOCYF9sY6Ivj19iWTfvSh3r11i4xazTCsPn/mhVk1YY93SfYx7APvXNbPkVHxsofB5JXMEFrYpDBiLun2uP1Up8rF/QgB2AFHo7leEeOl+XlPqzEAO1jVfEdZtaMD1gaJN4Zu6Hv7mdD/3FdfWyu2a75Gpe06Jyhth5rhFVryZBtFYYU4W/XxJu18/gfJdNyZ0Tr1QliTXNohOxGwIs5ZV3GgDTc5o7x9j3PaJuvNTByzsss4vQInynqAGRuXZNXa+DcydLAM7vvAWCV4oLjLd55so2vZdicB/WU/8a6yeqBy09EK49Ft3XnOhW6A5qYUpOFBLtTKSqHXafAgBTyDZYWAlWAwViPzC28orVdankTACYqem7QivLsNtTq9CLJiSbDEYcodjYj75rvHCOySB9n8u659Iv05PVD3S3qdtjNmViq/HMPijPHN/54Bilm8IHW3rzUJcmOjfRr3NQzbYR1Pg+yOa//685lZWvQw5G+MReLkMKjD54ynP9u7jU6UY3YN68TSQw+8NzAu/jE5gQp9cQrhvrn5mHSIG+qeOiHHXDNMJxK8Ip3Wmh0Vr4iW12iFKZ/JEbNb/uXKmQ8tVmtxtM2osfLOX5qV/OwAo1wdQrNthwwReGCMXtoNL9LcsWkvw2NrFCZ60Ot3cI++H1YCHgcJY+Py/xaTilZlOqJPwZg6N5T41kDAGeWwuBAWeciMYep9BeLCTmO7i/Sn1qA5eLpVynJDkJlYwoPbuk0RGAUFulDXKKZb5d5Xc3Sbk6AWmasugfGcd9h6n6+QZwMUoWeH0tJuWHR1Z6Kiytin61w09ON6APeZC73TOd4IolRwjJEgU/j2vh7vB0Qv8pEyIc4XpkvcHCIEh3XsT1HvJwbYaXesd0svtSBuKdyd5Y2D7iPi4CmqJJjOSQewc3EfrG2XX1GEP6cDphrZU6/0kwlbDEHp58rpV3Mi21R+K6oc64xjTWi/kCXhJfg5WJso/g9K7rFvj4TU5QdHA+bIS4gR20v02wi9NzkqtZE+NiauubUuEP5wvhmvg0+/CH7AEEQ11ZG9K7VlYye5P9/Crx+7xItkvejdP8SxbcDT3UwFRuDILgCdWRzmO8mVXz+zDkN6drIGo/sUrpibdI/FtYN2MJtIdZ7W+aC/jq/xwkOYDQlOFmjizu3AmutiyDF/6Opz22UdB/okk28TqzRVWtNoRk+EDFyE/x9WMd9W7lCOFnLnPAmTkyuZIR+bShu5s9my4G6nv+FvCwfNLVI3yxb+nLdJ1ykoMdyesG1rsl7Q8uwhEAMLI4h7i3OXaNVvZLDM6lPjQ+OeFTDB/BS7Dev0vta0aF9d32HRYf5IszIBzl9nPd1x8jrsmJF9rT2QpLdwf00WMVZX25iDo8bTzp9gLyZXxEtCECjUfBWNIG/XKE1TgMSguKVaL6tJMyef8hFGJdqcMZRWMeJTQb8gfLvi7S0q3C7wXIvh8bIKuK7rN/A/mrsXgKLykepXAauiwBgbM8kQUJHa3QEJ7T8QUtdLIs83uUnTSmn34bU6qE2Q2Zv6qZK2isnr6R4cs924UaazBeQnJxNOwj5vLFYQCGRESqtg0SjPHa4qgVWp3koKEnO5XD3jIgL4Q19ZfOzofBhWNOP+CWITH1mRLTw+BHR0cZPG3SjnCCT5XoaH3bnPu8JVZBRLAc2dw0IlCCr15m+7DukWEqvoig6A6K8JfyGy0opZRV0Fj2wJ5CpMdXYCnxDNik0bB/ZpWWBVvs53c6c7VjmI5H23UW0/sN7uJ929QEOwz7ZBMZyTITT4RdblEfYONNkYxNx1yAhKYzIB8Kln1R/kcszPae5VWTE+eKtX1wa2v6bIEEN3Wql54fgepEtRs46p6YF6s2vaGzzcaOJi42Qr+JB4/pp1WdoF+t2trWoF/5iJ2dWJMEfGCLrGFjPeVpS9SEt2EWGYNtfZz8xLNHag+ONQ/M8QypgqdEaKjMrGhiCB+9wadeVltUidStsZ+sRLoEiil93sa9A3PHT9gjBmL6hTuRrlnmi6bA6C6M9weL4dJz4rNqD9COgvGuA/8x1JIX6lCUIDYIbOFTQoqrKiAy1vxW6LKwpyejzulRlx4Mb+6chptA9rSNNv3TeQXN/RVX30Bmvf+QgTcm5fLu0LmBfH3r7Y3NQW4Fn15oumeowvnAQQSCSZFrUVyiwCjg0UL/scCaTivsSEhaU88+ySBwTIjVYDzo8oD0MY59hvKwT7HFAT8XC3QzbA2Sz9wntP8Yv/qf/F/eTcWqMtUF/LlP6vTIBLHMGzBx2NCD7vGSgXcGNPV4rY5vZPoFhnFMCTq69trCaNKIGjkImz4MmlToJmXGuzy4zsiYlQTe6NOSJ9vMX0G15q9BuVGbY/DTLXWGEY6ePaHTNhDBe4DCSuRjR/E5BL/21sjE2zNxgIgbYs2ZqI9vHh3Cox8NTbhf42TiWidw9mPkn/1AlLTnfd9fkshN6uyLdFdvcYvg+zD26MSnkZS07Aiw0mtILhwkTBzPduYA+IJCkCoIMP6KStpkUxAAKbwVzFTWo0N6lT5NyH7PlA5GFW/am9zlJ5S93KC8fL14hPueZHLXqLjw9Z95mpi7iqJhyFfPBC3Wyj8hKofFGquOoIq+YLASJuqX2HkXl44KAJYv2MXNwV5XKKGPiso7wNPWoVWnayDU9nKzjxIL1IazpXoNfq9f+C6GTIgVTWbHU/wuf7tfpkSA1MlOR8KrJQZfJUGm6jI+ylkT4VWFnL9a55f66Reer/be7P3TswBcKP9H1WF63ZN/QB3KSAIqyrJQ4PJOzXd+fvo7dJWj4CqTqwDUjyCOf3z5anPSq2AE1LGhRKF+AkHoLr2KwQspcWrxHVJ5EMRR5mrhpF8gbkpSE90D3vQ7YGSSCQa45TfDMwspYxvd/qn6qE1fCZ0OPcDQBPO7ZJq2f/8nEls2pp7kleF8eetOOognw6AvVCEoe1bRK9W4w6lC04NldiyJiCU7EOV/huOB7ASiHc0dV2eTwlx8Bos4tqBumqsoAM0MSbAPXYHkQQqaUutUqB7Be9nz4j5szO3khVhhqgLymzERQkIeb8FI4v8hWoatHAvV7iHIauy8ZgZp+0qxl5Z9v6OGzvehWXuV+lqsiXsiWIYbPr4QxZxQObj8a1FHsxEyo+OJ9ds6gdYNZBHUNBtTFo60t+eJpGO2bGKjiqM2DU1DABdiVpsaOtT8vEnbGlPjToesTvkxqQYUHErdMALrm766P+EFlDIQQhtG46+65s9piNE0SaFfnnrEwNZCEWBYGDTTQw132PW10bVTDdWrExeF6zLfIyp9CM2eLikduhmVuxBWu9e11fQqAc632kktJ55HoWWewHy708wrsodbqvjoXWwa2hDXTVmBD0JyYBsgXWPrTwTWX5yJjQ44aB8nMSBLO2uqy4031Ts6oAYu/dUtR8/71qKGcLWR3dF3Do/w1rzMgMa5rMW/snX0fopdRJk9Wg1xONxgczYqDw3fwuL2ZRwP74Fwp6ZHS518yu0cU0HGhbZexAJk5hNByk5TtkmC41nQSchwE2dKMi1oatOF5GTE9OW08Fqcf70jIcKtAB0GViQBUUlFjNb22NAZObqq4kMYpMbiW7y3aDhTtWHrxK9hx+Clvw7EKOb4LRnlmSfgQX5BhTXAvyT2WMG+xzQnTwnYRMJbz1lJW5vxmEHZf0EuSC+/9+Hn1c0ry6Zdk+hRq9+4b0T9v200IyRtSA2UzbGc8xU3+5UBqcVBznJia22ejZkKAxDwSfGsptT5r2i+duQ3h94BlBvw2AI0mYNgoMC7bwpx2c4K1PkiGP6marvM+T77ZLtAbUyLpBwzXC64sqt9AexgBotsXHZglDRjxZTUbEJc6Tcq0bInKdPj3Dfclr7uPPVFeUCxKm29ZzlbcK3jwuLGYHH1HBin0iVyUuElwrzakzr/RXYC1DYAmI9JZSgPsVUtJYZnm5sYJXYGEvYIfTcAyG34WXGP0MmSrn6wcRItaIfP0aXbxXZGSwtnYDTS6Xa9I2XoBoH8thlPr6Tlk5MKraWqdtq6iUvnuGXP7Ya/TowACWbujmtBd5PcmvAwRxmNrlxkI04ThWkO3nq1duHOOVh6XJmyzMqEygW3+CZDUKNURVIFx5QImY/MSDA7TEr+A7bPR5t23okYu2bVem4xcksx4PmFWX1k21sAGGOgh4QuKgsv0HO/qDNQSoIyzu/27Vz0L69rwqvd4y0D/uYTd4ZFpuXBc62sSD1FRx9DhIqL8Cki3HIWNcBahwUEw83ZApozxLCQP3nNBrcQ573AFUn+PaWvQZ2NuknpbNlWLUw0/TK72aWc1WYSyHFCwqBo9ZR5+I5EXZ5OvFcgIpng4Nk9pOTg4A6Ax/6pp2c6ZG2I5ASG+olgkuxzh/8osX+AclEkLEYK+kubLjnJ3NQFldfbvScevIm4huhSEyTwXfVLtdQjl0cBT0g37UPOMuHAtOchQfPgnXTvrnOHeaxOeE0YTxBjT3jBIAJZX/LJZF2IRLMsPqY2D6ljoecWaLp4cfU+AXXdm/PWJ7DhM3BrlBo3ZmJ8T8tEX0aJVs6c5RuyD2uCaDGXPcIXasOtABzFx5rLM+MMHC2aMW+CoXTypnLGo8noElxhfz7ggahvUvKxmmCY1ZkZ8cVS5QptZC0ZWVPVujjidtWfy7VntUPvGxxbtQwiRJ1Y94EwWUIrQtHadFeXFjFiJDqqBx32jIARB6rUUgRkjMT5vA16PxsT/zG1Rfvb4tlHpZQY+drfz6xArm1yhlruNzWabQcUM558Uk7uHTdcK3lcShszBzz6UCWvqFnDiHaI5GsHxqdJzY2Yv2EEfWvxe3IN5qTK+4wh1GxHE/6Pj/c1aHoTpASM7bYQkVhqIlnkR12b7CIHZh+AuO5NXpAR8WqHQ8rVUuQXl52KjKJUqmHR43KG2E7uKCWvMaGja+k+oscQzv7jurNyFP2vrT7+HcK7q+nEoA2qSGlJMq8sk3WDa9G0FDd2FpuKqJuPXedJA1ancJDN5wLt4Buw3etpgRsNZ/fXdMcc8OGLxtMZ2Lg6m7f+6FJv56Q/Q/MsBr2GJR8PJigUWtPejLVEI4Erl3ajekCjjD/ieRdqJulG8mBCPDS8vUMMkPXnN7HVuNO2siowJjip+a4dtXNpB3ettSL9MeuxA7DgtMyQS0dTuv00A57adOuaIMQ6ss9tPPvUkCDMIOktpNSKtWHIbKby7iIu3O37yT64qy4s6mJUfiH5HUz3dga8EaR4ipR6lJatvXUic2WyaRqO0VbIfChecvCrCmhIJJxdNN3NbitaECrRnNauKRCzZmfUXhVDt02IK1MW36bzbyUX4YJbCCfLRBrHbbkW5SOTN7BO/iwgdwQrRxIg+Bj3zqDYGtAXXbAJ9KiW0qse+bfGNueAl0XUkijeyv/AVmyzSq+XTzzRN0DlQjPRPNIRS0b8Ok9yMKOTnULKdYz2Kjv0oCnvqDXXsEKp/e4dI69iiJOf1b+lyU9s1vYv7lelgc7eCjSRKkiJ4h09jzCuUVgKhXOeURHlF3zMOTjnOnKOTvjLVrYbYEkzNLephv8FE1KzUA1CHA24ZBcA5yx1Lr8Qy0Px77DcBhBB9qXZsu9PLgO3GMyvtdErns5hPMaVFDFr90RA4EgjDdmE8fNpVF6XZbvzZkTp+IgsEZt2J3ti3VjEh9r+XYPfpSeCjxK3kffzxZj2wzobS779Y4XlTtBc3HLgmV6GcA26h61Pzqf1ltq5hhOT4C9dXpuyvPJ92oleTusXhel8sux8ACpHjRcztRs7cawKl/NS5DckZY28FtxiyCAsXw8XVY3o8KvgoJgRNFxe+oca2ZkJyUhX+EO6oQFyt1v/4WAK5S3x34ke82E8Z3SZbJnDkooEtbEuiSYm7qiX4a9ttOMGhkWemqKzO0nTAQTSi9nhFlcVqXVZAX6B3S3wnIVlmRaiqrJI0bJGr1stMv7RvtB41JzmA9nY+TTm32THLBrUijvlXgshlmbWvXbiPnb8PzLr+bkdc80+UmjeS8VGj42frrTJBSLa0xdGtfZ+g8z27j/CWvvZQDSUyVqt6Olh/VV7qgmXrc5ym1qkzYYDOiJZAzpi8fA9XpnFQffZy2M9sitd3b6T03kuwVXi0t0qPc24bTwuPCjcUpz1bO46MXovwdASbd2UpNWAsMoODXz5OzRDCp+bkZdbl/TyIWRrGv4VJtlPstb4FFBa4L9M8PpFORQf74i+bwqJauhurABUAK8WTUWLftcAFP1XMp5rJhJCnnW9in8RfnYqAMWXvXll3wrr8i4Apys7Tc0wD9/9Md2/nGMZy4P4v0tX9R4V0a5/Do/hHcRC32v01q5Zn3qSBVesxd+iP4EtkTNCqlcKWwYlc+MdELnI+l+Fsbt4jlCuFv03m+7B8jXS1x57JdqtFl/MgWaGfP+C5mG/VXToXNqYNlR6zWOYprU0QaGRH0xvg4R3TzpPEkR8/HVMuKVt6LP8luYVjLPUyznLUYYmVlm2MY1XEkfiMbroNwikYL4I3VyZx9KxQR2iHc9WT364ziHuw06T14MvdhpY+aDgZtR0lu5yqu4imFPLXnmdyqJw38CRLLcaMdv4b7RWc+0IfdV+wICQGj3Gr/XDFIrqQPQcUD1UjuxV1DHO3DomWaHoSwy9lEE1oDN3ceeKp3tfE0AsfrqPdIVEEmxM4ArBQjIwJouKJMHwpa92cI5sriqbCazEKguLJzHsxCGYEfqcZ/AWEYARM54xNu3AlCLydHzIkz85027VNDRS8IMtej8eOObt8CRiUKmeseLmKV/hRkeqxMJVz0ht+JENn/Z3uiUpbD0CEj+YiziGTZ/Jc+SdrqcNwcmv5Vvk11UfqlpBK5zhItSxyHTPfDWwP18T/nzeJ8vfZ68CqcDHovY5W15Y9SDD+U8wynl7f4XrJghV/nVTuN60LY7xT4Rj+ORk7RHSuNQDDSrvbXYDLv3Q8RE8mbMAN5YyPfK4RW0J2zRo9yDlZBhGwQXGhA9b3sJtHEeo97kXjmIpvNY6HvLmcbG/FdB/l+A44bXLpCxCIX/dl75IwH3QMLYkUf+4Nw78IZXCvctp+F5X82K0Auf8smWTS2Ch5u9oJoyCFgF879o9JoI1sfD2I0hVVndeixYoA5YXpYqmCh6OU7Qkt1KpoX+RW3oamQeNFVc4Iq+dBJEn1goFrjH4smzYWEn2VusoDt8gC68vfC+RzNiuQ7/9OvA8J5mHvtQth9TZ+BkydDng312HIr2c8az1b0LmE2IfByJJ9+a+XeP4Z9Cf4po7VXP0Ymdfe46PfNSwfqqEkNKn10NUR+0Co5FSPZSDuP2jOeySYRlbDQUBQp792fua+8dfgmkP2X+VwdIzKfuPQM376rjlEZH/jwGhSvb5EOrFjKC8gSHshHf2akUxXrxJ+bMLZaa6m9o+FMCFoOETsIPzhd4f0vmZOaEB3lZOQfhrVIXuve2tdVe5YoNTWpXPTbiyUnx01Y5xwx6rOUgtaOzt72Qi+SYbwAxHge1dFhZDbINzISygQ6/D06zTq6kLwRx1fYHHsCc7iGa/Tx6ySwpwKFqTg/GkDwsJiLzTFHs0Av0CunHZstbuc6Z98ABKC4HcmFVqLOJMzwHxrWY7Tv55bquxdxyTuPhpP3rtxah7rqe4EOcwKxoI6St11tPxEspwSFYhLnhaUashV5wUMMVE+u/RD8fNJpnYMz9uQJGJdXDX8df9ikBPYXkvOjz8p6gl04Nm2APGDZ7VjFR3B8IuKXXtX3qMBd0JrA0v0AHRY880+U2exbmpha3Fqpj3Xi0ikrW3ZJqHqJZ16AscsVfe6jpU746hzs58j91CSovhkEhMhXrMgEr8eah79mwy6KynKqPR6saVTzODM2WTHPsJq5xTiWqUNjk99F81M9QSfYiO8KftI02AdcfS9UeY7hJ/4EB8hXs7CyxX8SzRohzg5cbLsf9zJDh9Uj7BCRDnC4D1YWId7yTuP9huWzvNVNNtzg9OLN8GLXXI7QT8Mq3mVCMvj6TlVI5+eqChJqXcM0oBIoFBAR/jyGeeM80c9zhNfl1YyInBIKZIHPi4BSCKKbnfp22a5S89Dc7+S5z8ReWujJ2rMGBygb4aWcrj7XHKV0Td8nKf+4UUYzz8eUtv0g9AN3DwTiprIy/14Dni21ZfR0WxhVtQX5dpE7P86Xfp7x1fQvqTPAaBzTvNT+9O2rxRtG9UmYRiV84C4fKoZN/EtvCB17go8SRxMEhTTl837/NrlwaCbvXCuQKTuIoud5jqYQUIyYr8FOLgQ60iVoeGYnfrVs1y+vufhqLtcGh9ZzRmGwqDLkXnpXfLMvkbaHQar5Sou9clEnJ6akushmMmIHWwI8oYFVlVyu2BNK+9odHy4mO2KC7RBMH2nwHSku/Z4I1NsILhjFJTgGWrfiHzzPWm5O6zSxAnzAwYdpgh42BlJjn8euWdmoQJvkhOw68CiAT5kGgDHdd33sQ03c9bAUPW9fOWCkd4J2NsMoqvgiyBWzX/iy5uzn1dTB8AUpAxKpYHfsrSmIg8gDH6nCf3HwmzQXkHXR3E6ejdrqe8AngGJ4XQBOwpBHt+QarDl5WWDmHTOn9UBVYLARJF0FxZxl2SPo1/xGPFWMXbOkcAG3MAkhwLG8C71L5rXFLQXxbtohNMf9hLVly1HURh16HBcUZoh13YvySbvnrtpohLaZ3YSaKEfeKtPKTv3kvqPWh4yTEV8kCJ+JNs4xkUWKProfW/EIgn5pVoYWjGCNHvXJ44qlFrhivMjjEYw7cuAAA9fTe0kAJQb9CV7TjKPBJ0O99jMjZW0lPjSys0znTNzmMmSndL4pSD52GM4U+ZAvWmq+ToWG77TxwFVB4e510usqTgebhq/Fb2oMBRr9wrySoZYIm1b2/QY2IUXkqH40L/WEAurjFdSc/0HaHK0JmYBispKRJOMLTOLKd2GRIUYNRARUwTTTCkkjzeFckiVnfAk+WVYrqjiFp9ZKZj+5CXmrpn7e5JLEuWiWSMn2LNoP9aT9dUwPrsKNs+yYANssAOUkUM91p0YngCtbAIPQd4HaRusqjw8/pxZpi9ZZnYN7nqqA8hIilrOwHfCfKJvBDw48aPBvRiPQa/ehKVMLXtdtKlOfiBRy0YXtz3u2lBgPCz1bDZCcEV84A7pW9eVb9liCY6NG71r7SpppF5lckFLsidNA04J9x0cZBjpJ3ke9GfFY2pBB3WxQMmXC+rfdOZfcPMDlMz/RwWopac9mR/rGvHZapFKTg7xyokqJTi9YYx7p457Thpo4jiMgHaQXihjugoyqn9Rk0BM+BfWyKPEtQZKt2iJ4xpEf4/NMnI+YmlhfL43JkdMHwc0GiIAgv6TujzX841cKupWCQe7RTIex2qV6hvVCC6lqdhnVaEJ/6R/nWe1MtSnLdIaiVmzOm7EMCsLqU6qDnKHkvBH+UkxbNhZfdhz1fbJGdP5Bq4oIy7qJtGMJY/PyFVbVSXHTezw5uSO2RX2OgPeq7sEq399ZQZVWI8yQOCGDsrc+zHqq+v5svbreyilEsJCTUUjEVCpE11a2ko3lPVc1b5qUqYEc/5+AnvvmwWr8GpEKZuonrxrUnLw21IVPbrtdq4ZNo6b5xHOlS/0RIF0Yu1pUyVciQ4c+nDOjzHmyPqB6p/O0X0v4HHGBg995v8c0R4MLhuyoANwFT29MFsYOs/+x1ElsUvoDS7R+PCzjeNNQJHlue9p1zqWSxAEj2Spa5xb56yV0euApOZ5/4aN+0f5hRxA9NQZT115REZMR+k9OYtUg5TbRjM8SfqmCMUsEdlItQvi1EY+YJ91J26zS7ND31JOcQwJ776W4kj0Luv7wiHTponcZE4dfhN78mucaJbCqS2wXBtf2nubIa/9zkGAMi4Y061bIhJOhrxY3ePunBfDMZRwusDW+4oN1b7oshwcarvx9OPVzYG8VS863o/cVpZO+igcxBv/I7p6amlbM9GIcVVeIyiCrTfOdakKBj6eLS36Rnh6ogQqrTc7lrLjBujpJFdkjAXX/ZJS7jMWzuyYEPN/yje7G9Phzchmh7Usekz7pAAnVjkpnWc6DwVW/OLPf+pmutlmAfB/SIvfLh8Q5lUF3GR90vnsejm4BAb/3EKy5yQGvqv5PAOb5FlnoAmP5T7CgVI6WNGJ4afxJCNn7U84aBkvELo5o/jGJtuwqrReWw/FKK2cgISkfk/vj/5PmK93Mr4FquogiJLEgjceghQxo9TxVwY4ryjmlExDTV8u2LJSqxU7JSXKse3kRRFH8o7Saxdz5A86Nk9/r1rLr1CmDDxpCK8kTW5dd+HKndBLINVFth0863cInYlDC8ptMrdHU0S0s+eEI3I5Vv+eJeI1+UY1lHZ1en6owYk8RZmG7dV8h3xLqs7a8OGb0zirG2MCbtb0JMfn0uB5TH8mNMdaxJYkjL/GWv/DoL/fetHMtacPqiLZau0ghexDYXmni9ngXRttsJu3SpRtLTiK4aEFRiRvIVp9rtxodoLsBjEtJbSjQY9PgUOOCC35bgjaVBROPfvz4TE6yfU6c4uCqIHp92kpdR0S3Qyhq0S5gjQ2pL9jTm6IgvvIKocovGToLP83jrtR8BUehpEDFIgcptLJ82x/ZwAdOCloswywkHqJtoATeS8GWHefShjBXl0kK9dghGwvWs0V26poo24kc8P7VoDYKZFV8sx0qBEZXar1SICI/vGsk4SkSMYbYfnC98WYKteYZ9okAke/MnLQ8n5mUVDWPCLODdZ40XUJYlBDzRkxnJhriBGaw5HcRcX5EMBKJRvTPJ49ZT+s5gdTbPiPvGo34k/xxWOic4k8KHpXEPiUN0WXQFoom90Ph8VV2uxepxvbxigh/Vw/DCDStAQ79mj0O/qmLj+eD8W6fvevVJmdeWms6FnPuqNUBfgZJqMpbANAALJulk6b9lr51pTKoS+K/T0dm+NkeI/tPJEGg7faxGIlItpS0VrMdhHEts7+U/BLAcH8+/78bOsCHucq/fGioRCFpnJHbrSJE/8biQyZao8waF95rW48Kbvnt3lp8oQ6ooq9ERPuxSRqwilnXUV7CFJIouyIYWZg7FSEKBbRn6Zj1URin3cE6fDgesxZXpPclRWz9jRZkAvUR9GQQjcY+IdfnhYEjmqp/KC3lsG3XVAw+gi/ucnnRPJSl7tWA5qxZ2tr5T1FJSQRIkB+KJlQktFENKHwV0DPRBQUduB7XuQ+Qt+ycUvg2gLFeTTr4ZXvMcnNM56HStiRgge5xcb6C0j8O+mnKbqkS33jwS/x7RKHXsyaW5pLZANnoT/0V5HlRJiXwlmt1noAQVmDKmQ9UGD+1anFqn60tSJX71wke1eWAOQ8bMN9Cr6+UPkrx30iryUMmbjRpCLRQFlxlMXMxV4ZWptLeXL9n+1fUwsMnlPL2Gt/E83Da8CaptcKWfsGw+x3Qb8ozLdxhBtJnd6FPEBKYCzrbY5loWD60Q+DZQhrB8GTLyuycITJDvRpzzXSmb+CYm7AhgPQEVy6jvp5lV4liT6Gfo+roTV/0Wepz0Q0KJ2h60qOhH7mQfukXVX51KNIDEdkLhzm1MgwO1fR1zlzsL864Wrrk4LEsG1VUBhq0loIDpzgrO7pjIWYUxatPgocOLTgxaPTzmz66vmO6umxdEOxzFPA+WV8yBrqt6WHc4SEIcBDA29oQp/mOnhaLcNSjWd1FyVzMWi5EKRoFQKU750LD1O5Yv/D1b29JmU8Bk86F326+wWAJ72jyRzUuLraTX3ASqlrZBHnIkSTWV5yNpmoQMZi5M0SNtzk0YNvPc6jsuqfE9knva9hUe6hJr8iBJa0K1hDYS0rW05U9wkQBePwGQWPC6/XcDZhQeWsNnPaKYXCGv13CXCLIvEBgHEP0TTUQ1X6VXOtQ9yLyn0PeyNqoTqR5R2GWzWQcuuW19K69dYdu0E+FHd0GpO4lEEEC1guUt4I+LkncJRSrvb+YqpIhQmOZPzfZ06VuyV82Bt1n4z6oICx7BA6V5cDTpQiNn6WQSJV2hYE0URaC7bJa4aqUB7wUCQmKCCAw2h2Qe6D66YkqDANwuLsTlu9pv/mz8jewxFv/x8CeWXFA5ITz42fUw+vrbhcFzCTYPeIt6gPkgNS0wVgSmrW2FLog5gBoJF0vF/f6WHYsWjfCPgI3cKuQrZb2ZWWo0gv+BMH6uppl/VoaFUJG1lqeBeIqlvq+LLjvvzHwy4hlxdWM/q8XXGfd87hbS8cwA/USBSF2euItv/2vxedY+bcDtNC9PTGsNeCsqTMNnXk4Jd3vnvxjVuyR16wZK2nCdlJxkNOwHWWCkDeovRHJcC3Fia15DQBvqQuvqdx6H1LEWQrnGh7E0P4Vn5Uod6pDCTAUQQNCfYjohrzbOxnaPPXzVCr/gHfdRypEhAU0KOAhm+7FwiNmWDelMPNsRwJBKQaYYvgXYBCACMPPmFt7CkSetRlxR3SUJ/LviNpypTDIsoAdUGOd2/9zNiF26afAhx/PCfEBXTk4ApzzNf9yL5jNw79Cyc3CT+t/nKyAQHPkVAJf/FNoHVnf6tn2IKzpgnE1WoEVoRdIxbqphPyCwz/C2QOoQP32DStyX4wEYu8hcTZrTBUQciu49RPY225ErX5UoT0gTcVo2D0Tkn78q1218WhR/yuTLsTEUVOzCicwMmZ8RLe2CRmMPeJcqm5c/OeaK02u3slyim0/Or5MePkrKxFjbF2luhSGLsTp3ams1Fm/LLWB+K8sRB3/A3KI7X46zTvdGi6xE3z9afoIFCcxnflC55NZ1UJxKEKRax2Jv7cvvcHJbudlAdnUyFFxZBa0hwFqhkkSCkg69qChGYJgEXwBysf3nAYdFn6PqJY15fUdkWgnat6dyapGJj2qN67+zTlClEkim1I5/wgg8ko1pUpmfcUz2Bz0LvvxyIfxqeXxkKR6MgCPzbDbUaxYMyBKcl3IMoFiL264kzFfyGRIJeouQJzq1afue46ReMzU+BN66tOwyUBt8e0Dg6exgJFQyNMlsKrjoAesL0I0cQnxZ7+3bAImbSGmwg/erh+N8jf6jDSl313o8fSwoYAIRYOr9dOzmj9/dD7yoIryW44qpgpl+aXfde0woyKsVj9/8zfUrhqBDVWgk8WnqL/6yEDi3SDebDTc1HjHCetda01yDUUhL8dqysJiSoUbVblTVH9BJAjv7MfWJwKhj+88QMb/p8/kl5V4c3jSAd/D0KsDjxLkmdyZbkrcMtUFqK2lVfsjTzbeAHHfH9QWcWj3g/3Fa6lzUI/TZhOQmM19PrkUwP2fW7VLcO1sx5ZQiOVHBNDvjBTCd5yvBsFQDxRoi8PhcTBtggCF/YiABBLgQAhwKHPeuWNvyUe52akFxcrTjF2JcBj4hCarsiKfCj0qe/h6zP3kfzvx2XIxUbGSdkiknJKI4X5O3rCvbyfLzNNiWeIQfre062mpg61gF7Yl0h29WuHFJ8jcyw9o2JK04uNtfgoIkC7tjUoS+EfMcSj1ldWnafC7GMH2YMPaZXs6MN+iD9hw66PW2VlGDGU+wZf7D6ujKRfHaYiEwQNrriMn+2CtfopOYysi8s40pGNoXDiOfwoj0VElrXEsk0YXO1XjSAbi5GS5GViAOCul2DQIW0wh3w7uE63OG7lyppJK/3q4j56+yjXxOxj12bY8pSsDHCtZBh5F0wWljSGh7V7ROhRIoZAnaWxlRkR/B4XOm3nPXZpFSyquFnXl/6l0TzjCySIsDGv/zd35UnzdLYyqSWc64GUxMO7auU7eihuXRa17TvPyOtxlvwEzpRpgzR8HdAjrsI7od93+WKkqLJvRMPXrGHUXCusS2WLTPVdXZuqwOAns3QbjbDAas/5P2KWn5JY96e0gx1LGP/8iKiC5NbLUM5oCucq+Fvo9oWlIgyQGA7KNhbqjY6UFN5x2uglFBSuUnV2GRsQAlwlwfyZ4wCI1mApfSr6NvRelzsujiKnVJqiCd6JjCO4NDWWcPybK50hpOJSzqOH0vnyqB0pQC1fwxc17EPxL0wEAAdaGFeiAb06ASN4kmE+z9EHr+GnYzTrrD+KXS7/eJAMeR6ai7wvC+4mNqBfX76gD39dUbVkZ4FB91D2elme2r4SZ1t1yNzVVKLwbEx0d67yjlejUZCcsYks9gU1sZqR84jwZejfNrMvwWtL5L4a6mVvVpY6mQK1GlYGPKXDJmpEKUuP9WwPYrL1kn6x9utDeaTM7ncsBv4FFK47z2K8AtwA15Qu5LkKqkYwinEPLc5p1bi1rM61N1S1+YoAWhjiRDRvfuj7qVrood3FpaPZayjcI7cQNtyn810+6kn8meVclLcvNJ68oiocsrXzDbzYQW8dQlVZuz554MnXlpx7p3QdUShpp/E2zMcx4d9CdvcUSPRmlu92H2xmtc8z1J32KFHvzgnGvz0RVX/qIvhmhF8/0Usp993WDzz2D2Ar0aVAVqx/T1B6aF13g+XjRX6lQj1BESnvu/+bt+qJpxRY2jAk7kewM6jgRW8M7C2i6dC+IVo8lpp80StkVL8lV0w/XuoaMALO9ZFYWKcabIPua+VZezwT7CsCXStbox6PQfMczhqPWTQwty4QbBngp7zXyiyLbMXiplaXv5xAKG1HPLzlGs/6mr/zxA2c9CM2ERM4QnlHHWunNKHFNvmpmWMULyueohc01iuslP0R4tEKfnjtuYNEr+uh2jk5iiHgMHNEkbXb85lvWXta1eSzyaSqPza1ts4YUGylGE0eSvuWaRHyTKNyUbhFbnd/dsrvwDW2ii6ik2QVLoxI2qNzRKfw8bJZUmzU5KdW1QG2E9OoRFqiovss+rHMXQTF2Atb39dz8MASFnDVzczSVeDp+nb1jyGIQB00uydzxD+as0EpXjjRm2ZaqGTNhb9ijuNV9VBQiWsgcu3ConlRQ9xW8of+zipI3t7E8ECohIfT/kD5UpLKcREAS25N8xZsA6CtYLvBDggOf1tFnaFqiaOswqeGB62vZsN47M15t2/4tVQbbqljcA6PV7S6oCHOV1SZAS8E+ZHksjna4hu7n706/HSVsnUx8dAJcug=
`pragma protect end_data_block
`pragma protect digest_block
a137ad876bb24d1bb488f2f0377eaa6208b2bb509a76749d5840b88636886d6e
`pragma protect end_digest_block
`pragma protect end_protected
