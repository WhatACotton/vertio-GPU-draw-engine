`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
tnd2LM02q9LQZ3nPisdh5Z80hqMi3V6kWi1qKfxaIcUojgeBRHzbxDLK6PQRBD03yqwCcMFToYD4Vetuext8mp/wE74NvQk6bBAh1Ya63BBOA9MXf+xOcfgHvSy4oJJDkqL6CNQqv2GmS8PM5Xzn7WG4IEx9O2XwjwwfvPilo95Q99N2ukRxvb3t2CHcGoAhngl6YGJGtEiuyEViFK8RZebagS62f34toPKbiyBbkkyWHNzgBYjg10TR/fNRvC8MuwdM6gyLXz+f2cZM9PZVn7NK8fiSSAZQIDEsSm0Pmmxud0XyszvY9cg1C21J4hoHOozMMO2Tx4n41Qaq7dbSFWdcvTv+23HNzqN9ToNxInNCBBvcrgKHirirxcvjAxmtQxSTi6Q/UDILtau3zhEsp9WGyG+KJeqYEGDpcmzyre8F8TxjWwmEm9YRWm6sSa/RRPVjpLBs0CXAXHDE3Cdw8hlqKgB4SmylAyT+DZohB6PArGFP9wLxvruKWUVHo5MOb72giCUTLk3nMOBW+M/R8zInXbQezVrUTU1UpM5Jr1np84gAugfjJ8ZmldTsQgDSjef7RkP4VgaQrpmkzkAD0VdZYwp6Z3cbJOANd38TUEWmy6jYJCliWZ0K/OoPMPmaMDi0U5ML+5U6m90sVtDvjqC+VXCjqBlW+tiYM7wqbbM7NaXGeqGi9dcxpN5eD606UKIe0f54kfMRUyp2wzZJQhKOfp/Y8PEa0+0Ci5Z4JjXPECgdLfaoPUbixr3C7PH3M7/NH3z/GVnE6pIY+VP3VjhnLbxtUKEqdUsrlXNllBuq0vBz7UqjYRq+2x+G27RbFM2RysHt91BYmauamAIW52RLlr4dxcxBLCHXHfihSVsL+xjLvVE/b5Zf1DmDutkNMcUKh9Ary1vFqQGN5441GyN/17uMDv2cpKJS74xfVwmuQ4GrhbmuBQpy3y4Mqey+s4Hrfht9X+il/6lZ49eqED6Tz2WxaNhES31HORNFlcVXGOREtdsIyrFqaGHng1qRfT8jz+ImfQWHPGe4dUmMugoGPutb/uBoqr2CJ0leM+dJRet9iS/WJJUXdWh8P1m+NVn4krA+7b6DB+T1jQLsNhwIRj4vueHoq+2AHFKCwKbiQTHvY/i33KH5n5bZQgkY5jepH5xOXYAgJ4wm0uQ+mviGALrTN1M1kW3kcC6SCaPsAhc+oKvT0Lm/H55ZJMFfHYYLrNN3lYDa8EG8GRzqMhpFwfj2yfgyQHg+fsZT/CMi/tN7Yw9/7Xo6v6EuCPlfO+1XFUMeW66PtIm9VROCJEMVyJftve4/CWxJ7mgRcm5nQbR1+F4VKXjUY99cmWCC2RJwTLaxeTnOl+F29yBUW7Mzo3wOut+miaoZln2s6EmL5jMdrhfIxrVgjFKS5gj3U+yPvoEORN0s5CoEbdWdtuNYSf9esmrx/5g+p7OOycz3L7lBs2ZU6SKUNPMPnuH4AooLqOOEKEKNKlU+vVGhuSvAO61fjixzB74+tfe3q34FB/3UAt+tx2IbMrK9XbWBi5STx8ohbdarJj8og6uk9TIWcEbbVNrze4N3oAMsZQyfYCZVnurex/JC4tGycs7c0cW8NqIKDBnp7cDCDEvomxo+KK9i9+0KIHZdOBQ5BbzNwBHo2fwcQZX1FyY3ZkkOafeurAPfgelbtA2iejmLfcaTh5z3w/+NKC46FyyDD7sijIRFfEiF95CABSF9aCnkxYaBmIp0wg7V97L9SxlQd4rdFP3KS+jMo57BD0X9vcs7zXVzRLjJBySsOpBx+krfPPkcadYj1kqu7x9N0RC8LYiCu8Q98alKOIKJC7QBn+LQTDvj/K0Vi79aDbg6C52pDjHcR/FfKHqMbC052fqbCbcHKNpku/3d2sChNs3Au6V7xDMOIjO+SJ4ZQZm2VMGbe3kuBtOpVqTM84H+lKIjix4XcxTtIKS84D0nJxcFpGPN2Mudym2S2c5ZLBBDJtGFyZM2cyYeZsdx2Y79AG1Ew9H6qVCzUyYRWiO5jQ/qzDp06X20FVSxYjpJSQktQy96RWdZgq7qrH+H+/GGZEddZOkfNCrGbYd/38iMGSqQQSHJz0l0pinVmh2CZNtwGycYzasGNQKS+F1JiKIFWSWD+BLFY85P4UksqFoJx6BsELL5T/qPCJtvCi1qvRtBBxbJzvmMa5n3XGUaaIDbyCIxbtuB3HWNkooRinuqDqnPmnWb/9Nq9u71pReE4cuEsyjj67aoJfwjydgBX4RDH9zA5KuCtNHvJAVCgYXm0JbBWzgd4mAjmyQ2rBQpnt/B2vPt+iky6c8d0Xh0YSy05Dshs9mC5MeFtf2wLw+/rNfL++9Jz1LDgGm8alKITRoU43Ytkl591iUnBuvjpIcVm3YPozMiHIJz7AX58bEr+5JnfagitI6DRArlEzuFFj4Rif/RyoJW7UANYwFBeRJyB2NNJv1M6AsZ3ASfAPxsbMIQwLn1+KW9tEvNpCyJEEhU0vx/qQBdOZ6bcvGqMt5kE/yjQMWndXXugwL3AVwfxNSaphactgUxyXDjBpXAViYjyZu4A/X3WZZRCengmadWc1Uxmoy/d9FvpmHzwJErzlPajO22uwCtqBHGcNiTaXCdaOJ4MayPFZNahEUsWV0YTaCPUkDl98eCtkXQBKLrpn1kBcy3VlNJnYb/W9Azs6IO18JajSvfjmhRKrvO6BbBiDEXUAg424QsU5Ed5wv2RxLDLUnP2F/jRTkAcxYBCKYy7HPv+9JjS9sYFNfrpTMaPcthEdO+bCaM4eJPul6j/enWfK1Z6lIDor4QX1uqjh/kzSnGNn/z6xT6i3QjVSfoLABIk48qH39cjkGPKuClJZR9IX6pKiBBIY3magucM4itdPleZcoRikYJVF+Fxbozpuboar/qpd36kvIrTvh9cSuY7n7DB0I7QPjLJgdeJ6FRDHS88tu/uo89V/rxaYUf4sg94Q3NqCmHHsLAyKQhXwsuF3A58J+gxBRI/0zqSTZQjqzUPHnMn9A/h8Kfddk6/lY2s+qgiLSuMCvuiQEWqADMwk9ZFVr2rhMVJ7+9XtVsXZpFLdVNyA+t/8LalW86EWB2ob+WU0rSUk7Y5VnDf8aahF1CinIQXGZDKRwQhytH+EuFvP6L44tbb+uBwwGn0ohk0QE4eMQau4vB+neAh8ryzkOYXMTMrtCvp3F55/cCFLoJX4lNNnakcQ/E8+ZmWz6nE8Y6S8q+A82Q1/hFMmUF7H9mN6wwYIxy28tbfoz3ZER6s7dDEdkNu4QGs1F4HER5izvevHoI7NaXtf6qSvbg06pzhb33NzxSKz/YYkdTmY9N+5Mz7BfTRXf5tPdkzAf5ZDHWFx5k6ys18lMYUAqVLmNb5hcPp9EnACq1kCQ2jwrZA4TeuszbPQCZBKf+HZs4Dqz7ZyoefI1aWzdUdeBITpSYfYnR16vHZmtjk1jKsHBvEgEXg1/kWJ6iREEBoQsUPfdMLYHKqUchepe/gMd4Tc+54SAR2BOx2dl1m07hB/d5Gbp9CEnN36gTNywcxS8nuxmjtJ9Px6t2MjsoCIGWVulvjTYfryhwclIuCTo0gEpNyTYs0vXAZ0o6qmIR9iP/wJPuOIN1ixZgK+jlkPmHr5v6xGcoUuz8x/Gw68/HMvwmfChcVUJy982p5eGYgc02BYdBM879Q5VrNZK64ngkC9jiR1u3JVlA4LbsDEjfVYrBXaba4VB5s8XnCw3lzaB7R7M41z4XcENwQVeSwoeqXWCkCivbybIfQCXTuU9jBFDJM343Gf2/vtKS169wpMRuRwe9slYC+ygvqltxnHlNzf4uZAB1xaJZZV1t4ZFdn3nvqRuHK6DrkUrXNb9I4iIST+0nWeD5oyK/OGoKO1bCkfGtSVRp5wnIJSz/krdX6YFK6EUaa4tkAW/iVUlRFLJJruLZMk5nZUfeU4YqbR3H67+3LPVLoAtTgRko0EZlflec/Yuw7vXuqhXdBGlLpqwqCwchWB6WtU5Eb7+IksFDXz2XZ68hoUmx+4/ZzBMbU065iiaunmHxpo1bSExM+iyo5KiSv+PCqoExYwSQGBiQL9CAs4+rMMLfjOWBSrp+slYm19UIMhKc/IKwwEvZWDN6gvOCVeeTRJH/ZKBAGkIlzjDaCNJFeX/t08mXrAU5n4vnKTDyLwWjb449NcHVttPVtLireiY51lz7vWNy8utTaVCDAyT5xQp3mfVO+J39DxcmPzfnu62FuTkY5F2vo+f4U1OaMIZT818VOLfFAYOW4blYP9CUP/ExYENhpfsdw+dVxfyaju+OatNcNIdqcIxurak+ZA0/1lvFmLdcg0//Pz35xzn1KJgvyuqv8UQx1ZIG9yLQEeSsJcuadKNIjlh426p0Gyb0lzV+hSQwXjCSQq4CLZwtfnpPR1oaYz32HWmYTpnrAYqK/GJGQf6p0LAyQCwfvYtKftfe+L2+GfGcH2J7+viAWb35p1ZDzcSxYJehP5G8Q4LU7OmrvHkF+W5XstoQ/MBDQd1vY5FyV+qBVIv57EtyJsCzc1UFhJeJ03dJJUKRensa8NRTw+aaHRfyEDi2sIs0LTmE5medlxC+2FOPYxxMBAQfsQmk3B7KKcJQqegzAuzuMUOu92KAMcUXoxK90PrmSRExZLW6UuxaObzvgVoDu27mbux40yHecDxQanvvJfwPhvEnEDnAi3ysdNm9Mot9Ob4tO1t+xlkYe3LDw/gezMddzHzgWh6cNx3IAqQHFlMpyeO5gvKbdUXk1ND6E4oi0CrwRJrEhihehbdq/hasQF+MupGXTYkZG438EO+cuDZsOAYK0Sx5H8F1dc4N4YLLJ4gTr6Mo5XXdVWAk4TRWvwP3zvH0HpszEAypDMpeVe/J+gp05Cq9i32LNctqn+ZRKGv7rryOQbSF83GUXDc6JG8YAy+Tq6zrEDVtIGEUeyoDIdejKrWiR4cGhD+LwW6jOuExoxFPa+rl6TU0SdNPsSgUeW9Jj+ovLmEvaQbFO4ZpSf30C892TcgEtsClaoXN23y8PkGuIfFuv8qJ5BpA0CjS+s+Mzpg25e7CYHKZsbtayP1cReE22xAO1dSidk9m3dkR/slFWGsEyx0T5eqhVranEqM3wiuZFS2vqMfheQsvnbM3E2QfpUz5z/t9Ei+8HGmKk+31vKufZrTuKS1jh1O1MnchPki/7k9rFlNCDljIOJfk/bnjyrS0p2eThPtZRXx1LGrSP+Lct4870/T63DYkj32spRzf5gfutmsl+Ea7xzF/ku3MkFVh5yWc0PDelUo3RB1Rz26hiUTK8mkiT1Uvm7LiIGuwjygs0pK88Sag7TJbLJBf+kizkxdn1ZWA9cu8Ij8hMpHg4QLL2OHD8DoS00LmWiWL2LNax6HZ75zg4YYRYomDfCxcc2DpGuDLCQalNoA/L7LPYtlNUYXIy4pWixw9ByTwJ/n6c+lRvDisAhKgJ2HTmTkQYSFRXEOnPdGNY3y28sqK2HO6QMlohXKrO67RaflNAnHfPXoslNJVV1gU/xDOlPWTkExcbo40DEWoVkye3JUXuIAYHdXju/Up1swJdZO8kZER1oScJBovkkdTPkyUuCzJZOAf2ih7SP8Ak2kpMRqTfB7Qg53+p3RBhk36+sLw18vNqVhLu+xnZlTMl7BRrRsbqotVK9WGN4EG8oQ/Ibd7RU14qBfA+dXOOJP4ImwZpW/ZxokG8s3voZbcRouKonhBw99gSNN/HabpPDxg9QQtCXG4xs319ZJEaIiUPbtPIX8+VWIhlGikJ5QDXYyvXV8SKxdQo/qlsKVTlfE57e4fiL0WNlMKntE3+Mz1Gz5f7g+TL/uxjM3Sfr/nQtS9uyqUKB39fxnaLIImonI8K/vS0I1ezch0ilbotFPhJ8zEGpisPPSZpWybeyIlVC3jh/mCHVRb6CqXd3QvSBUHKW6qsF+eFKUHu7BtJLvDKAlDi5jzvmFULI8h5KAv6IqHjeudiVRZhUT9pQhITxF+gZF/0IBjjaVdv76X67oNbDKOsHdKYUtMGfFRH6HFyUDMwAcvFmQbpGVR3UdQOq8qxP0GnvsNeRK+2qkaZYF1sdBlfkpcmatclIozqe5MEQoeG0ZVWNg0ESsyug5S1mJrnijrIzIWjmzIzeHuNuM3xz7e7w/c28rk4FCOsQf0BAzrLwyyVJiaeyCplxZBzPqOt/Bteza24qHsdv0A53Va48seQTVrSLO2cUulaybe+dBgQao4AA9g/4TlpajJe8dzzYMMBey3KknAZ4C1zYvxe8x1xnyf6RB9h9MUsbq/wIaUEEVTcj6feQk7o6iUdSCn99Fz9NZCMsNa53hu3urXOfLd1y46JcHjlHLvxOJ6bC/NvtwMB4TrFo6RHb3xPy7RkNDV0MvIjpEFoJUAihZEHay2IlbT/9Uswbs7ypK12HWUE8Y/pDPu80I24yzEALtU7DqVPry17DPBreVyWGQgO4GVAxcUNbZF1U03KFHS7uLzdS4VuIHy4f6OxoFNb9ThFVhV5xv+cgOB59CBXGc3y+rAVFyu6yxUCC4yCysT/F+OMGFK2+7VeXh5jouzRfhkHFqhK5p0kN9A2GV+JKBE0m54lqXyXY43T7fSBIix49bYbb/Sng0WPKcn/RSTlPC+71ikAPc3FvNHTr048c/IacnmA1+RTmUgAwWH/p3ywzct0mvC0ySlKtaCzQ4x5cJnkSw/RvNBS3EJ087msXkuRRh5jKu+lWYqnED0kNcv9y1NPBezFlhwdraidrRIHexj1oHASBQ022zdHKkgrFn8Tvc5USQQwLPflSre8duzL3cEFX+dtKCA3QwRYWoXN0HPUSoTsmxQ74cDjqUxZeANrSn5BUAJQDOx1sadpk2MSheK8Q+I0ShIPedI+UdFBZJ3zXRzxmjPXa2FiCbPsD8pcvs3iXy7GsnLwKLISqPBMkbfEPlYDrwu5z5CxxbF4VsuPPtJGx02Aomq5nsYERKCNo/57julSUo9ET1d8jOafvmPEatWFP40xwCwvr7CF7e+x4OnUVWBiS200a9SieDNQYQ+vDKl/NOe8G/3kAMWQmJlAJgJ2IEo6leIHgthXyvrfHnGLb+F6q4SOVDZbvx6abKakrZj5AZAXaZ1d3EhL9Q7X+OyWxT6LGQ5/lEEuoU7t2RY12ctexK0Uaj1M6JES+QCrdx41xOPpnX+PMru22u4b8E8CT3hczLWcNfAH8nKOOmaT6j6GQDOyCgtXbG+eVfoRhyDlEtBu+Kol4IyzuttSIsQgG1v3oR84/kt4LX4UUlvznFgWDjcHQq5HXxUn8o9V8pzQNwMCxcAq7z83SGGzzPTKC7bOYy82ywajOdt0h55uc6jm6M7h2GdhhQVRYSB6CN4OwJp7FAOwGLU8E1uqPHgkwqJCBFhvD8fboQPipod9YvukPT4xZ9oaDKQICjV/GGM4lPcFCVDjKVzRk5i4kplZDQO+W2taaf4OuhdQMJY89NocyUFGg6Dm2zT9srMHZeLACm3t2D6WsEahW1Lg7w+yjF6n9Bi735/KSJ51gDkXtW1EPxmXgs03UcQCEnWFszQZXcbBYOo7FvzJEVO+jmPUCoOeguIDbcEONmn2rE7l1AJ051SlVr3wuNyQrTNH3yuiJ+oyRgwX6DRuY8Czu5vlVBlHfP7i1VrXhMPrCK2URDYqvoFoS1CfXTw7OflJC2e8nrWYjqsGkdkcG48ayTXEdCnWdRha1Eocyg3bhDfavo3+J5517iCLfkTpnJmyBFz7SUGyxUC950sBbXgEmpSpr9tnwIKXPTZrcrUB+5EEtzIQHNcjpJFTyJfjXJ/je09bDNIudjzRuGxw1JoXhn4iSFCRVq7BmcahJfO5A4EpXk3b90r/557g9/g8aRFVLO9YBvvxu0QQtObfZJQACqqxqfLjpCXQpa7lvg/JtYoKJLkWgZebw3io3VWpOcI0QvUUzvugHuysG0It0T17pJYki0H9TLRB/ni1GFacyTCVx4Dj838eDiPzKd0c8D8flyGVXxQKcmMBIygHuKHMmf7yZdIyCpR+qxjtAkl3XuGWVHPyhYOaPlENyRpVN0geXp9ZugFlSkEu7YY1GidcT2YgEOqu6rMnxtrw2Aw/J6ojx/4F8/rNT0KiGv/nx/qhsrcw5AdKxHIrUI6u+jeHa8XOqDNaojmrhk7h1FXnow4crYWAje8ShwRpJgF/evbYJa+2St3MHG5zbRKFNi6Wp0pS/HLbx4yiCWaYr0+RZfPTUmSWI3mQuwpLHpXnISvVDyokzz/gWPksaT7MAY8Upu4GpYLe6aZVYzsOXyMeYc6C/FSei1x+rPiT4i6tw+0pl4E8AUka09A1S2M/YDRbqNncjVQ5P4Y7dUzpV6ntLcgHxMollWi6fXhC7i00sKtWIvzsV38/F9MGAf17q+uCdtD8UrztTHQUaqWTfgcEpWIqjqkCdepdd41jKs7XvQ5DlHvc1R9kS7JbKw+sT78b9q9eleo5Gtjkr5ciBpVgMUjd+7ZECsmzaI8w8TctkYrdyKgbMHSQFkbRpW2HZOIUjUxMpaP6jCL2rg/wEqyUi2AV9cFTLkt7xNxM6uR1OzVv8SV+NG0qk8xV0v5U33503y//nD9Edp4pjWTLTwpRp7MCOZN9XoN/gzvj2GbY8+kwJfI/dEd1WuW4jXopTto+NdaYgI3SrnH8krxYmSCvt045OGL2zYjwejH5XPvN4XQjkpXyatH5DDBxIIT8RtyecVRDEAZx6uI/rUTI3iagiitYDSQthBTCi23oQ84Tlz3H1i8lL+LeqW8kA7fCnIBVnqYjnVE5aGu/cCC0nnn0ADq1NsXySt/zkNYBoxQKlM28/moRqEA3evq8lFFGupzKCVzNb4f50gn5cBfUCitN67AauWaPLFzP+23BQ+heBM6GXL0Y4LkFMawTD9TlVIrPRfYCc/Nce7nHDrLnpcZSe3P+b7BENkrYDdnAajcvm0101454odZdOqQI2e0R9Z8mQDdm2Yudv2slMzFGKoVMUj6z+xREkkfSUSAphjsu2C78eF/CLF+3dG75IvMpISEjhqlLX9eIF9BSow3l3nZgAHbv/AVJh5p+8XYUoJ4/x8YrLixjdknxi+VrcgmaG+QV/oSdXy1uGG121BB1v0Lyho5UfrYSVN6AC49G/CUeclhMx7fxCT+AX48nZWbeQi9YmsRnszB82dD6+TWqIbarS36V5wACQMFCKCI6hf/NILQ/S5XtEvenabVeoWawA/apt1gGi+b+jWdWxVYuinFNSFhcoYYEUfZir532jTNNcdyavVjSITWnfusCXWrQddovxqP8Jaak5+GXd4p65tNJF4q0VbTOuEMnojLbGVxX/87tppnCZAy+eDDpq9lTewoH3hqtzbTysEXjuqCG6aU05yBsOG1PioQKLnwx2B7VcCLBfNJnPjvnEnai1NwZFx3lctUZwiFer+WoFsYk5y/DimMwjNjW9b7k1Fa25Z5yXze/IG6bK8z/Kpt8+Acne2KtEGDBlrwAwlHxFyuM2wHcDJDvr3b7GRK415IegodAOy8FYe7JNlv/AUFLvy0aSkLtLOnn9Q2kijTNCix1Gt/EfjkHpCtaU5fSjJB6RoTMRzL3kId/SIr2Vb0tj7BIcRwCkhQCxerz6eqzwMXH4JT8yBUNPv5PviCvjv/A1902nASumwMRtourxtvhsbwqll7t6t86UueVadAHnNJuSNcqZa5EKo0adcfFOTNSk1iwS7q8OkejhsUjU4sFhomwvDMn7W0cb0J2q4osHcfIJqMQY40lkm7cOjd/idoDI25tTWNAMSV9s5tPOwXUQWgt7enHuCC3ZUnNshE0xu/z3ZQJ+AWyBLw1JIt6PS6mnUR2+gC87UFehhwIcJB3M2uOHJ2Qzn1beS16C5vhi7e3vBei5r3ZbHXKIYCqESE+ml39T6rH/Wwbpg3pMuGS6hYdwqtNHDWiEG/bcTSjedwNYZ5kXJO0kLy3DRf7C2NflMUVvUBw6sLQE00Hzz8G2plL99kXO1cJDlpdNhxLSkhP7OMHaggurqhrJ5yZ0nuqDQB+ySCBqBQDLli/PKzEv29Z79GEaV6np52oqEvsNSB6QY+XDB20DmCwY8a9Mz5tOmMDxGy33Bx8at3s6ak2NO6vVukolf70lrk36Qz3ahAis4i8Lg6OcunoKdlGU46xrYSi/Q47v9AJ+MD414a7d1v0/HtAqv82QNFvlHKt9fjm1REoH+Jit9lvMofK7+T2mWiJcldef2Ko4qdklQDEQz/wM0zMkoHbepGcsFqose/OxRUHdHZ2Jv8slx9zw16/hSo+z3QEtYPdZOx1XUxX7XzfSnljfkxz/sWFS+sQxpRzq86HAE2rVcWYTFcErqHBU76yvP5zJTmL6ASCG9FTU9AU+NcslIdDrqGU8QLGFNjWlW2IHdYPscHqah/QY7/NPKAnHCMePEYLJVAv4f1H81xPnOmuA+zn6w06cyFavMoNWq7EYXN/Q3kQvjBm8QA6zmDCNO9GmMBdYk6dWNSBTg9AxxLGI6/YYnfXIX1S7HbOK1KI2BDcRhFCzg4FOY58PfqduYFlTPI2HUOYKN97XgrFfqiITZV/m3MQLxuLLGaWlRRV0gaBvSUcBiAbFTAAs7b0yJ1RYprYW/9WcDLAIRQCMUyk5/V2AR1H9rUzCf5mpZb3DB3ClqpumkSza7c+nC2oSgtFT/pY2YWSprWJvJvgswICa4jtDMPPOeVLxQrclLkbhBqTrAgm11Mc6JBgWtC0IxTkJuA0zR6W22cLpcm2fC1wKhm5dUvGOZNAFZeUg0pDbDLOX4p2bgtt6puOrOm5IYHm3YuaWQVLj5PpS92Bcxbk/b2Jd3jQC/aJ0dg1EfKEuYzknbOVgAFGLYvdNPXEGVf/X/7CpvntSrVkoZeJAJ4LLSL4KzZidh5m7EmiMjraxQfP1vbYjlo36aJxf//sJ2bxm/broyOEXCGqfnbjJauuy/skWgG/8By6YevsiFxQt7y3hLyBUDw527LTNkdcUfXmcIG2PdDm0np2wAxzoVswOqVm2AIjWZ17/xPu6PXAsHdB2MxxiC0ArLdmX6SuFg0sLEreGcMFfg3zZQ8WmUjWMldDWQFc9fNq1WlJlH+5C4aepY46fDeVTTjWZ3UDPSWAuxMYJwNbgrkWdTA3sGF5kzHLzc2TYs1NkMTkLJ6U4Xxfi6ZAb5+SVpXx//ZVf+KZb1QPmAgbN5Kh0GssSpJ10xCTEpkfOU3TpNj3VmDaXXZlg/Q2m5Hvnkvoa35ZyqvERsfNaFXMWJkFPLGWuNI7NRiav3g5gXxyPjFRTgESjIPQSp+zfqgooe+LrmLkvQp53dlADA+fue/LxEMj2JWAgef90dcOJ22QxhARzi76r8+NRNpfP5ghqXJxr389y8ubfmoszs7k9xw1JrC6mU8l0ORIF3BPRISrKHP5Zkj12pd/cmH/FyBH30hmNjn2F6AP0+4+l/mSoj4EHZmrzUg+KqbtVZ2PhcooqJW8lTEqz/SWBBp3JLDIvOTtxmLV8iAfKmQ7QOuTXyE+vkjH0j7rGYGiS44Lqn4E/nGoFitCxazfPQPOX1XJ1wzR0aMqB6VCIcetDlIbgoWu9RtMLOcfxv6lEw/Q3QHB6aglAjUuKT9EWylnquQPbFhu80MypaJ8SDyVZui4VEaIzAYyiONzckQJ73FsjGiG9ktiq8tJ6xJllMkBqjMU14GjwjcaRG31XYnH8H9PMOobo1hA/u/mzW0DbmmLs42i78yNoQYIkBqeLsbMLmWcwD9gmugNITR9GHhtA77zFXx+LVqXMxEjigenI6yzH0X62Byq8CRsq+LIs5aGHOlbzdPq6TdN6LEjjAPeeAAyerL/9TBqjYAqTr94sqI8LCg2pFdCJ1b5cQuTxMWCNxFqT+MiP4/EZlguRaqvRNtLEoq4mAibulCVmW5G5eJiET2RmyQVzlqRrgwpcauWuCG0ehLCg1ZOhu94l1FfYovj7A46sXYF9Jxbv4DIhS9PH1szProw65Qbe4FWFGVbo5pDOTf1q/0x0DIzVXhDMIV7ZUQt2Zec78XEYt2ckSSUI0RY0bEhumWQjeBFvUi0c6pna04a6TQysDUR1Xm6AYPeOWxMmzEZfcV+u3CbPF2YZ02XmSZNP9fCEetGfnkUcGzaHBTs/WX7u0ua5PgZ+IOKgLcyABXsZlC+hfNKxqIaOYYpu6xArVu2lBXiDRMDcs6hDx5zn7HgBZXaEfs+AXdPzAFlmsIUAEuIMsC+QCxkWKPnIxkWEP0Mu95koQD0N+jg+pqyP422MrQBK6W2tUvIqiSVyKwBTYM2yQpgguHXqF/nyUjAdeyMY66KdJqmlYImqz45GAwlbgDzFOOYjuLFzFZQ/bSuS3++TJaT9+d0/1zbZWfnp+U28spdtcKEW4LVvnN1G/iEsqZYQ86XPXom7wlg+OT2J2GIlaXJ8voumO0arsv7idLJyOMXK2Ab/WpJ7YKFIIputXFfMwlZw45N/90uKkNm/f8e/fF8RqA7Kl9EGQzj/Bt+vz9/nQguKZcIuPuo3kv4SWKN96sE5NFoIUoGzpc8f7W2GKpWo1HS823uRDrAPIOfJbftcQV16cO9dKFaNsirT3H/H2QDEWbJsYUrN/du5Q7I1qSvoWvRT+hlP+OghSI1BGwcFOds0iwqnojpmn3DepNA8FzlPQPtnTPKN+mV6RnZ7nmgDQBnujXfMswzR29o4+u4d7NFyfDlqKI+9mgquOrbDKyMV47+pvhTsjGLU/LFbRozvY/HiTd9zi6/MMoKv8Dhiu6KCuVOsTepENVkfVvaNLvYMGETuwDopVahqMRW8llCPZAdtg6r4ODduX/3raPPEtQEM8Z2I+aLncT6ayUi+Zmtm9wMFTpjIVQg7WaX7hLtWV4yL2Z1vqZWM1Lz0UlmmrbiWRpRMZEpTTSXYyDSfEySsufLAovbbURnZ61bfBgnzccUcb7YDnkfBlHzkObRat0gns3HgDc/yhXUqqaoChbJdtO6cZicZvoinBgIgcIx4o8UPf41pNXRSBAqHD5T9UmeekuY6wtkVOLJxKZ0OMLGFx3qjfxcWtMYcBaNQr0m2TgBJEqtQch+hiSC6uVdVhOjaq6d6aropDTM476qzOu7HgRcfeuKQ1zZMie43hNTt1DPjnozr/zYTpGUAcyTrOegMSDFwIxgS0db6hOsvn5kAKJ6uNf5W8EZS0l5oesPbB+HDmwxhaXuqbYqnWEDDTso9yrm6+K6JaR+t9bevJ5TB2XNOZzU87wWI5+qslMeMHhNXW36NSln0BoAw0F6gzx+wuI+HWmmLElVd+5/j2Nf6/ylCcmI2+WNln1HzHOEp/vpiPMFcJ+Ll3sxSvrci1cDttgFRxgR3JRSuz1EXwJUaiJ83+nCH/0VXiECBPNfmFRQB5pEEa18MWZ4OI1/tehtCZCYJQuj1ZwfyU4rytvCR8hcdmeUaWn4vWRJYMSAfLRcJKwtmwskEG0i8i5Z2n7BPg0vPdPeaQaRfXgWudSYvVuMfuZI5tR5LMG/o4edd5TRv5wEOH7k10SMK/5Yz1k9jjsZisaT901yCZQVIHB1t0w8xKftG5FVmofm0aMc0kbLy1Gtx+tsidQNsHAyrQYnrD+Zo+goEnXteK3mID+OLqGRQf3WnEbgtxjJ1Gh55KJUK+l3ib3KyoKUPiq5AhG3SqLJ75MvmuQl1vlhEyaAxuahHNo3hbSjTkn3Odb+wdl/3lgWsi50snIezCq1cgnfwpSudPmaqt4NNnRLnMhKe3aBPolb1sblkBdniNKydhP0jRsBgxznL2HvBwTCDoZ1EAGwPN4CK90w/QSNKHScHaBbfr3+Rqn5rsRznX7egneJS28t8Irc9DNcqoJIPBsiU90qYDWAAJOK/FJjl++iRZ/E7B40y0TjAyXAPIQ6F/v0P04/BEwR3taOYWgS+jf2lLi+LocrvmjgcOjYcBn9wognsaOR4M2kHMq/WlJCwnFahdAqt9DYRsTZpNkwTuMGTzDBU7AhBwkRec5DC0L2gSKLeoqD9x72ZB1rGGGGLAGOHvjx82dsRfxm3VDIzqbqwIWFdctK+UfOjOvlZe5ytaqzMwE0JsSbZ89p6tZ6O+CP4b3jz8Bk/MoSX9ofcv1Nl2kW3ibZ6eV0/roma/Gv9XoFj99b01LVgARfnuB2KAqFN42c9aZzc+6NJt0BF0=
`pragma protect end_data_block
`pragma protect digest_block
447b289696e0c41b8a1bd6e006cda251fc4fd4a425ca40cfe33927de6e3ca0bd
`pragma protect end_digest_block
`pragma protect end_protected
