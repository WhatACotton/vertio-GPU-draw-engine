`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
yB0madzgyQzQJpNC4+4DSZthntme0zj56wgssyUC8O6w3mhRvfiD4HrcSPOePr9RQHl7UOenp8M4dWR0DvkNfVNhQNVtC9hEto/14AlQRNsYIS12aaj2/fcB76aaugx3lghoDFcq7wup34fwHypFqLzspPk75dtwZC348vDMJBMZlQ++LuyiUHPrXiEEvdfXza31jA0n0zBPQnvBjbalUi67/gQ6s2dQxC2qfG8BzmPuFG29VKqFEl1VTcI6ZUzPssY5eFOrKeLiASgdVBrDaKD2OTon4HFvu6U4bsHgPg/Xel38UJ66acaVbQvSZ1iGwRR1JBIUHiLnsepzQ966/HR7+b5kwA1NfK01yf8/DCM+Uc6iabjqpgtp5vpoDnfbpsN9CagoROvxq1zuKpTZz9682Z8PNMhxQ6jNbX637KACpSGlWDoAAFXcRfdY9BulVMBQWbF2RDw9rW3AWzvCc+H+hw1fztgk0DXJGZM46qO7QjR7xPej9wt5Jq2YXbkU7hKjADcJeMPJGy+jUx+Ngz9Ogq3g1SPKPs9+jdfphaJoXYYU2ldnSJhhVa+4TNJaX4gr4SJi58yczPsBueg3gFdGfVAKJJgbwlIW+Pmv/kDGcDDINi1/Cs8IaEywur/u/p+Hro6jteMzEqgK05KjNRoY85WPA2FM5VyPk7WXiY1zz5ct5bxspj/3YV1RFFMr4F+6SM8A9VleB24ux7JD+6OuB5RjU3tt4CsMrjGj8Bk5Tgjm+tomZIvNK8VZONUCBptto7ueF+RSy+3D6EdaIPjg/v70S/aM3FhWF2OPuKawzvbbMTbLxIafV0u4fMBIfMWeag9Bmmk6N3heDzt8R37O1rBjZtHAvLRuo/leI/yNSSWT5nY9Ww93SaOrojyJ3V7+zDbg/o/H9orG4SkWxJ5EP6lkL9u3maB0jDzaDhTwkJbr4wAzlTsK7zuQ3z38OXaC5oMRS+RyUeEXNto1KtD25QPdDXmwJx7t2rh1ZzoItHFF26eRA89U3aCngnx6nisCxoDjDxWEOPehisyE/0EsmfWqYjf6PWz8RLZUXI1qeyGF7VQqOl2RSvVLCFRLEa0u+8bEUDMuzip5TPw8qCFJ5e++p13YFTOFBjNZvhntMxERzWfA7YV1Xly5qZ8Di5fFh3FqZfnH+a6Pu1Pb0gPIwWLf/shTt7iu8t6j4HJPDu6VhnLlLfQr/Syl17zzZfBDV9kZXKCAn0/Lx5q2umkHQS8V6iEJbj6cWxyDVnR//vyvDfMO+9ZZUAaQAZ5MV5VMoc3z3dsZW4rYRJzL30gJRo4j5UTtRZL+iGYc1ajRxj+N9O1FCbqjA2dapwhwNNOR7lqi5peIb20CkhDaq+tDY+jZqd4WmUvMlVrPKwXWwWAaoqNPSIbijMRo5F3OmJwEyqdZ6U1tF8C628+yPbP4o6k18KEtXoF+kWamEeLWx0zkX0X9VJzibymvUbVvvWvhTqkXZsWnsLn+VelCvue3GqKS+9LTZHhkEptqqlkFb6svPkLts1anD3t/pEpE/5hG/Nw6RdUAjzSdYYfogHuhyhilSpTlGqgB/Ew6gQhQfr6qAapADLZ4z6v3JeVM+nc5+7VJsmG67bbH+Vm5hlOYzuysUaI6o1azEq4VzGn5VX1XkTJXWi2JeB74ScEldkxf5rbVLZz16BofhmdT6r61lsGw5EK+NlWe+aRTmzhnc4fQhmL93Sgv3c/mn3f8vHA34TCKmHsJXbE31Ele12YNF8HyXvKE8JyjHSs4aX1vcv5uhoTgBJ0Jscs3fcgoCTvTFrXWzMmLZYGlcDN3uG8lGNjgWNBk3Vgnzyz695R/UhjlB4O7vNj5QGVuLNw28SIN+uUJsN7gpTdEnew+s1okL6GZ6/vW7+IN2Xe1wDWRCqpB9xurTQPkMRwPF55axUPXprf6xiWJ8xk4xzPuqy6ZZMJCXF/xdUGTAISqYmaSypBN4Z3mHJ3UcZRb0uRJHhMbory54ZGIGBjHWWWr4Cj7doMti+84XBG3NfUFtbHbVkCSwl3nyXSvMi/Z4zEQRvDMv9N4GVvNIsjFQV6YqIeQuiwTlRcuo3tGhPudmaKz6Ur3AHACX/EUeBI+TIpBclJejKqhcAtl/w1cFzSRevZW/lbRdrN7W5MgG3PlsPPNudlH1esErHW1t1qT3TCom9YleeNRKH0Tf+jVlIt4+pKT3Kyymb+HbmtvyrNspf7N23lU2889HODp+zaGdMw8HylmQBD93ZBvElpKwB6QrCHz8i89Yqs+WRzK0GA6L7ZEu9MegnldmeN4tCQxeJR8lxvSZuAX1tACaDpiereJc0ing0nBW+T1Ajp3IZBSSti5T0NI8mD8KAH7jwsYbNDWYaJSQd1YjdC36++NGRTltDfD7t9gJ+53Q/UUASN5Xf1OWb7MQqpQ2bY67pMv2mGF1RfAhdaZVPuWDh4n1UNZtY+MZjQzB6z9K+xSLAf1T1bVqxOuEbslKw9rqm7UIaOh2FQQgX92rKfkm4B2g+Qyby40xey+SmuX2Pf45RUkRIkX4aCKcZOFwG+XnDy7KnA4YNoWvCcJo2Up9cUs21AXVATgKKIdh96OFGEnhP/BxW7qpxCnn+yGkXxBHqizE96rEfnWM6hUr6QkVbgOHfBGZx/Xh6dRP7ReCtnTzdBLJaLP/DOlhPdJIpsUBifYohbb7SJ0PyTo0OmxNGpuAnHeAlDyGKM8QzftwFdlgCQbPjZLmWB2pXU+BgSxgODwfFMfZdaE5DGQQASa/1WZRqXjNBtXmniLS9d5yxoa5NYVdNWJWdUlXMpiuIAzPBhd79lRyde0VWxVhvgaxQYU9XZxiNb1P/y6770jtE7VinxqQgd5DkImOrUePB+QtYFGHowxWIH9JnHPeHZz+soYpwnFBbPBlOFMuiAV03Qm6nBPSBF+mf8PyjNIPzMnAKMZ6BUkXh1KMU6xwBHSXYSFeTY9nOk8ovYlzWEtkUHwrQHpxo+q1O2d8Zj+1M7pH9VZgYkuYigJ67gC2QMusJG+OXkAU53QUX2ao/GJVp9Y4AIlzMuSFYGfM5mCtIOl3LvZ4yupp227ThueVed4lI5x99X+9N8qGzt0WGWE+BkyWTzREVQbhd1UBRwfp5Z2G/cOMBMW/KmTPVTKxTEPQVVqh/wkIbq5gHfhYVkisR9jKApFTk7ztSQ4ypt1MtDW5F+oXqv1X8yNFl50OzT4TRuC0ecALOxUc2Md6E3h1zRUohcM5nN61hwUEVVlS/vASH4wAexmmEKdawjXHjxxcrXn7C11Px/o9vUDMNq7GM9cPCE/SSrpxUdsXf7HoxZ9fApHZa22tCt9gU7/lQYi9KURC5CxOKvmJUpqhJkFPH96+t7AMpnXCOOYHRQp+Xn2qRjQGoaZo33NB3LEmHUgDCZCb8sQdYTD/i8Cnqk3yrIQZ1uJybQtQjGfx27K8KYP9cmJGHDe6GphREcutV4NanjtaRflHtleFWkPtF/w126OUm/IrGS5i1HcGkU9cAHhjJK0z8A/B/8sAFRxXnxWt9KhQ8njMj6gMAwhclfSSiZqBgW6YboIyl8itR9yB8dajYpav03r/qOCE50yIOsNnijiWMi35/vjm7VUUA149giaWWBbUy8jJ9QW7pP/NbBirSW4TsmsAM2DnuHvFkJCshJMEssvpkh+5/gshBqMIn+5dDJjbiNu0DIYtUNa6NMVXji7MBYNqQ3ZEqrYaC1stanHLLXl1gd5N+TcgCRAhOaA7+P83frWvE62h07MgjrttsC2Yiz9uYz6drMVeND2GQdARFyrr6+vIxsFY1/uL0me6zpu/7vIRfV5STpVx8PKnCWswVXL36kysRN+S5zVDSjro9nktMBlicq+mMIKnO0S1Oe7n+MYHjD1M2Z/oFRr5c7OZBIk2C8sYVgs2OpThYjDNSisCGwEYMar/yLZJWEGO4NfJG4JRp1+sYOqGj/99MHn7RCa7TmWAx+53CRW8jTOZDSIaNn8wfpxiyf0o95YWWU9grBNICKgLDQcqAbyLWMsVgGEjHbZCZhCelrDYE3pQv3zY5V6InKi4fOStLMQLM7/kTlYstPow4LLnT2slWg4rhhZw8HsGE2QVumQfLOtoV8NM8NTUxbHfHYwWOI0UGrh6R9kbAVONg9rPYkbVqlKoqoHRBMo7ii0VFBiUc59e0tzEZaZDg1G1OnmrpFOjKXvoXpJIJIjorfa9mO9Wl0I52JHj2p2UBn5YodEjxs9InkPNsqYq+dvg13oipLKMe7tP3lSHNKs1yxBPpOV53VikQAf++rW+zwLMWW4O8f3FO78sg+09Y601XJwsgL81zP0xZNxMDWJrjyKdyL5RrAJJMt3jiUDEkg60Hde8tixLVBLbHS+d42CX/hUqQ9S2D4P5h/VWm1Gv9OZn8wM5s25nglCSg59fw0NSJYC/lzSpBq4aDbLwryazgVOmpbgeW5PQAGiSAY/J+uERM2n+FMrejh+lAPaYSf1IdRK+InXnLVhCQ1t7TJdCpf+tjkPRpjTRgqjTDbm8OMM5C/QeaKRBCcpQZX4ytuGM/0GIE7tCMdcfeB7YuZymufxsr4/mDMfphMj46oi/lsWw6iC94Kc7UCSb2Lz3rGlHxmukrPub8fWIwufpp7olKg70B85XezO3nzkLgqcEVMer8EVy9Lr38ZPV7KdsQ6ZKUB5tYCWnv2LcpZrzwZxnLWSEO+2MUCPRwyIt2Cf34Emf6zsCrYsFZ/gHkCTBYoRuQPM8ewr956F2FLkxsuRmHZgM00E3wLun7J89XAJ3H3A8KsQoUEwhQ7SXAZLBX7MTr2/FUtjYgK6s6y0oTjnuzEk9FM5guhUYXSBcUVjYFoqBKDF2lrV38zPVon8OflU7CxAOlkdL5NxmEHEzxACfXgzsnSBCZgU+mrWEinXT5Ca0ePZ0QJfqii/dVC/5SVbtcaManJiWDXDMvoaoio6KKuhOzrEiwzXGFOmFddFSXo62UR3a4KiI4q/N/ixCPFbT1ucLg9s/shuhjjt8xkamUs6jvSoGA0GHzpgoLtyC/XpN/HX2uLr+OwU7e9htu3daCxgFaAdonhUhyDLNV858uqqGWQGEHplnTLEu2JGZLmspDSI6Zf0sdJSEyRVHm+4PgjEZJBDlyUA2a/vG+iN7rYeAk6DbgVGKFOqSftKk0Blnzo0uiaCFAMpXhMBOY6yv31vSz2HwAPE2gVjaYqu3JFo+u8jk9Z8mYMxXEDRhkIQixU2DiWD0g7xadea4db4XFNsYeKdv2Ld9CHT1TU35U/nurxOyZ+v9Jxgauby5eKUJGNgTkwW00PxvhhPynyN14V+Dc/7XW7LI7wEDTJBcr9yGb3aFQH5ZYn31qGQE8uBYx+Wpni8b0ViRiQMs17MvoE9COExmLeeKFTje5Q+4md9Nkv77luULBq+zSJbuRECT+6IvMaIhAP1OKoVLULiKB/jJ9MjaxRH5DGfO43usbxENa2VKDWyIrvEr1V4XRQTVyczeUSc1tIAsZ9Jle5a0/+b5ROY7YYfW805uSfSs9is/hkaHvQC8cgxXSYGkrXdkl+EpT9xKfb7r1CEfWW/hbP6/E/lKJlJBVusom4z9dkjsCWRczxYOjeppGAYjXJayb0yN7zM6L8Ueg+hWVgbtLTODO2ce5pDilBlcrqTZv4tyXRP2gx7bZ6c7VeKrnra3BMpFosmk3XbiNYn0fmPo/Cvh4VAl2SVDSvzF5v4atZWlFYoFO+/rndUdPGJKG/m/4UedC8QmEMzyR11YRWl30eDaAue/VGyjY3CKxlBvJVREUFjIVNJ3Zy7+kz17uS4e+DHg/18JM4IZSNfzY5PdTAZ+QOb3ik4ol8s8O7Ufb1OpfhL3kakGqJW6X8WBlQiMn6qfu6L/hrJWlN9oM0aRUl10AdxC0fkh1VZPWcy/7nO39sfUH42yKV4Ysr9OA6zaIWYs5cwL+wS/zhpU2q4eynPW6JfmEoTkWYR9gXD7cDxMoPTt4C6Z7YBkCMo7kYZfAUSYGTuIDltniFenX7qlZUJhTXQ9WmQbP0CU2JykMia7nrVrXq1bT9z5DCnb/Ilb3LQjeTJow72wisF1RNIYx4XOYqL9GNLckdst6VXttXzD8lEcg8ip4oARPo0F7I16k6hqLpRByDwql0nSWFWHkij3XrybOcHylXY4d7zpUS8VszXP0Ln2u4MUlKdI9SDdL7CIe+qZIA27fVMxAv/Pe3OK7s4XlXpqEnn1XRR1+wm4Rv8s0IJdDhuma2UDMWmvyq3Ej3JVwt85JLIxetoWmWX0XFHrUdP4Fz6vBgtqPNXZviC/IeO2zbsu5ljh1AP6bMy0WXqdJC7dIziQFlE+MmwR+Tz8bWYN9v9WjoMknbf8j9OfFSx5J4rZ8tt7Yp70mZkGZK/QT49AKveoHA5JqL7PkM4rXrGlzJEDCG8vo9kNFdpLNBNmmdk+j+mRQl9cEEq2fLnoAM8DGN7VmPrfQt2GKDO9UgxZIpHp2Wcthu2LCzMzyfcIM801/z4JD7tiEcxG0a6JLOmJse77GrWr48WBwdTtO0t09nAttcK1GCAx+AUoGSRhNESFmPUWSA4hfP0Nca6tC+7yQayUUwK/vv3yvGXRwrjd9yyjYr1bOUl/8p4L/CyC3Jp84E4VREXLMhYeiZqKRwZOV2M8Aiz9EMUWlE7IOSjsP3/pC/thnFnLLacfN6gZBpUfvkBwgj6TKZD/BnGpNkgSHWgKPkNMc7GE089Ucy7eg==
`pragma protect end_data_block
`pragma protect digest_block
7ac303d332fbe18b5621af0a00c9ab258dc53496fe3c5c5362d186332c1e8e68
`pragma protect end_digest_block
`pragma protect end_protected
