`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
WARmuIx+ns1bo7giVkV4VFcp5mzpWym+XDgOVLqc2UhB6DTp8pBfoMDaKHN+RdQ6D/O/EPfWOh3+olV9AEZOwkvvhynPL6+XUFQSgLjCbTr53TOhlarnCdymOnbXR8CFtknwxqY8pMQzFeoAv2S9MRSDx0qygn+7s9V7844Ko6ZGYu4huhAovUmOP6J+YA20rqiwVS/u5GLmKrxwq2JnzGbvfDQogMcF6nFj9lIgDVgPMwfu7L9k2lIDwHbUuaLLVhr2zfhuRvZjnrGOHbCZnzOpfqvuFFwDePvujM0dzQeMTQGaYQcsGk6ZQ53egl8FcZGiqNTbQuzqNwHnMAdW0uryYKDoGL7S5It2AbdVpsPJDGJywGwghfHYZu9Lfa5sAXINOGxBSpl35aV1VVSWc2zWpfT4lYpeXf3Lt5MRxooJecwHWMoYfbJacWZuEjswpBPJtLcq4aqWRWnu6xs96+gQrOYH392eiXGAfq7uwiMbUu1n7kKbGIedgqQ2LHam+XWCZhQgWm4UJKQxiyTFP6m7XoS5goSrCQZPYGsXORFyjDrxScOKfF0xw7TD3Lsv47KANmtdAI++vDippT9k6f9sHtAiIc0lhDw20CcvkkQ8AvPDHGlOZ1jn/VG2PqsC+DBsNTQTBMgNNBZGNm+pKYn/De1ke4Br7xXe6cboasNqOFFiQkrgmgyKH9P/GnwX0CYcbHDe7GYENf7UG1Zyixuk07nGOWKU0tKfeGcIwWH6VvGAs2qE20QO8U4bv4gZq33z/IwX0xvJRfR4KMR4L8EVSRYLVNI+UZ023awVN4MJUFgVlRAq+wH3lYnXKhGRnfV81Vy7a2lgkJfglsn5LR+t900Xv4YaQ92Sbr3rizUyX4NExdnBIRIbT/TK+lpDzFs3cE60+m6SMK/Att8d1A2I/4NJ6HM0wNMRUxP6OIX+XP8Tb9DW5OBErKMDdJ5yA3yT5CmvesNjGFdpkrF0Oall1p7IVurTyNjvjmGl4LRzQWXPsL6ICzIvEoUXrDo5pYRHEf9MWZ3rYlyKd0ZBhiglFOc8X4sZRHnorKMIWive0pNFlF+iyAXLGcOEKOq1h4cWRQNF9BunsUru+nhlJMCIXBg8UtYoYk1mWOdFIVUlrfAp7krzEjZVhv1fMuYRnSrhmQbZDChIt6ZcGEkI964N5k4+pa+pWEmA018NUUzZYVdv64sjctRbzZ3wh2i/18dUEaOgDCLPMh/9WjRpgzp0j+2yfdLV2hWln5WUp35Ep7Ro/6TWTYV8KIhVhR0UGBIg6CvK8v7RvESfXE8s3LEHUbwCIZN1BsP2J75Qy+pnJTGGQTAItqT2kZioErWqaC3cqU7Lvyz5PSH1TlKtm5XkpHBrTERgGXOPcXENNLlzw5s9EaI6sRXVheS0FzKJI04fglWFQ1y4AlyUYsAGl7m/iiWDELkvmAZqQJGOVDmYSDZEf8yhlnKXhT4A/KLp5RTsg9YddkRCxkcRP35C8bHH5ml/qT8girJ0YUpo56QFbervx3eNIvh3XgILvFsLa9JcrYX/Sf2Rd2H/Ey5o9fxd1neJ3+aLNYbe1ck29/uqR9LFmirp2RQMzDUydeuLv3pWQ/KaD/aenBfb+lnQQpsrE3glSDYBD7YkWydcggdw1FayyyPHwFiFAI3cWmvgsASxB584VzFUg/3aFyrWp2i4HxDGCpU9RyHBCsBvNHtu16EJ2yYEaktEebV1DSQ802krxSviP3aPc0AXTURQjiyY8pv59tvrsp+CtYBKPhjWLscY29/3xdtpfinBiqA8iIrcLrlE/6QfgQfb+niZ5g2p5dAtpXq3ftAaJuPSkGl94VYwUU6Erxjq7mScBn59bsUfuDVYJLYIQAVo9atnWrNzTuH8t1cap9DrjfnVvJHP8ebI46+55oXV15jbTN6HB5ONAdxoThh5QDC6YUqJjBE1Ld/Q27wJbRBMCk+wL5nyE83HZG5nowE10mz+1pMr+EdZzBuSuT15F/fUWJalZVpkL9kK/JpuoiO4r1bqTo2rX4N0cEq2eqby1/SQo2RF/2fvk8UoFBgUaGzngRZQGpXYZm5zCSZQ+ps75GoOpywdrkVhC76Nmgr1UuuEBB8l6OwINjyca9QLK34upj19kDLdsDaGDIj6f2vZpMBp8c6+cVnOv+Ud21+KlWMKIyi+1P5KZPVR3CsJ3eego3T9X9b16zPqaC3c7LpOL1BtTU4gZSZCAmCjBVOpXyX62q9/J/tZNCxdZwLFsghuWD+psmqdslTwDYi5/Y2a4hq0WAfwaIrh42oFvXhe4Jz+l5vU6lT6ZLOq+Zj+YtjEiJyZr7IqjrboztUG3AwkQz2hDVnS0y4dgh8STMKr+1hDx/L5owglK6IWV3Qtb8WmsqBdiWrlpuPZwvMPiFJ/9s/+8zHxR0O2Vqo0bel6X9PtAEabifUlaUDbLy1BIU8orbVuWIXt2iF0UE3iV0wqcs0Nir/gcYLTXSdFspiIHmBIOGMnv2E/JCtX0ikY+66G4WYlZYN+yz5zXy+Fwa8d24wY0OxRLb+7KGdkLrwjVZnmYAFEGn38ZDr46Y17+ETC9imkDRIunxMduuOMOWTdt3RPoGGRXyytfceWSKn2Fu07X0+KMEI0cZ/fbiUEicGKSY5fbKmTHtFJIaNR2ugnkmXM33r1tE9M88df3AgDRXDWPWliGo3n1/qETFaHfsMlulHlzylFjYy+rvIz3dA/rbPGBUydi4KUVslMGJoq3b4KNjwr+1gkXwEulXOWtRJCvbDnlWQtkvvvAtxQl2VA+0nOA6LcXxwuXAEG4qmniPNdeK25kctFMJR9O6Et0hvakLFzuGKxIJFv0HEq2hpZbLgi1KVFbOq25mya0kcJPAm5uFXlMX4nO8vyrXgNnrsAGQLdYi5gIrwfGmGRMrmz0Av9YVY6VvFUwRnW002SYyIFiztP13sQpfndbQBnW9n5292w0HJFEbJkPDdfUYQ5Fxfxd75jLXysndQ1txneuwZOhBg36P9b8ExZtUgKIfa1ZDyBgOlocPCIrOMd238+xGkN+Tf6ABjuXKyWz7CASRJETXNwFy7e714XmC36R/eeKh1AjG8vmQxKuPq01AV4TLFD42QiSW+GlWrt+egF8yLsjhXrPZ+gIhaqvXuHh8PfOzay6X/emrs4SW+IpSHzZGx5MWhmDmepnHLSCcODtQCVLCv/qoSzMX+SSZFSWvdIqkV41pRNgbxPPyPCZjb1evYHdo5FGQ5hHPEsBgRUFDsaZxvrJQXHIUpQKd6wtE6Mq3eMjj0EUi8czTS7yFWekcoQ9mKwQxRdscfihlw4xCevACTg0ABXzK9/QgetcEZXSylfhhIaaifm37m6M1++L++T8s6haULjFBLkzTRaCghxgWjjdbzQ83Dl4PGWjdciFZCo+SU8At2Uqu7HvbsGOl8HloZd4Tqs7xF7MqCOByki/TqPQVwqznDUJ+1PsBl44U1MJmTX5XDMH1eyrsjOH7lZo/QbfHw5bzVuFdtueWbTSHgCwA8LRzUwLY6jKoPIHrTY8X3hKI2CY61MbdVG9dNT7FAn6jtrrVwDL3D4sTkpqqPoztmYjjCz8nA/SsGrkWw7JGQuXknQ9iP82hT11zZOfN9+HEwdbKhNiH7Rb3sTlzAqfJS6EEiIe8P/3fj0qTnJvWdDlVwfjNqaqfQNHz3OwxmKFp2Svb1xAgn6oTzyklXQajcjKLqVrb02rjnq1YTJpkClL3sSgira1z2q6bYVxI76hKwxaQb0Ozt+fjFzjHVzUcvZf4jbOHROw9Ncc6ZNzQX0THiBPzJYG+f0xqIFhHNYgA5tk7M6E8KpcE+3/dsCYycpIRV70pRhzosHRckhNZPiV8U+nWzXGyMjVtRMdQKkHyja8UUSRDKQrIy2zSpUiquhz9HMrgxxOgdnjHzywT4/prtn/1p7vxqc4DuJHNfVbyqA5eKeDDyDMYi/x8Ysdgq9GMM2zdLhoB4xTbZhjfDLDTdR9dRvE9gGXac8x/ty6ZFPcS3VH4w4B5N8nsuEkXJKQJQ7LB3UT7zsd40HaJNap++PfbUiROvEfVT/8TGEoY0tMq7pCilBbWzd/lQIcdlifm54xbEAiuHTfUjkawHbMpV79Du5b2Xw1CqANgdbrIlDJsRBkk2QfJ+4JT50wZUOPpr168YLJz9xlXk3iNYOGnqPqVUiq/fd+wqYSkOydCgnXjLAlkFWe2a8Raytx3Zf9Hur1Q092nboPYQw8GzGsYBqY7samrhqHJ/9s5zdN/tf/kq9TL3otTU15HEB2CMgPQZ152CO/JpgNBJs27EbTK4+POMiQw0TduVxXslIZlPSYQjg3In9qRQOYm4n5LS363pTcguG2JF6pWu4yCjYpXXzLXZOBdg2wf7CX0oha4Ds4zr4hYssPt44LS8zpST59R0eEIyD6CsmhS0uvPe2Vc2CWvDWLx4eNqIiNn8Ttb8jC0WEkx6Wol/GS7zg0ArxKOytlmN7fSA96XsWLmB5qLFl3dOSR48Kwo92NFSCR1ZmnV8PIiseJ1J9CWn1tEMboagvYcmej+JnGNDU6pgtQR9YaPL/7W2V5r99bMcJvT5MmOEMEAciG990m0Y6kTrDDfZH/N4tSKLjOUkTn2neyDWYby/+yuUgTpCjRHlja+z0wjsFnESE0uLvynH0tm1H2NYRQsEpWQB2KCH03pUleZlXGMPxjWUS8CXZ0Fp+lY4OtLf2kTt8Ttgz56WOmEWXx2aBHXJOOPjpYJhipWmm63RrQ8pE013vdRS2Ysdu6jV2niXTf93EupUQbSEMUebBHwqNMy4Y1REYx5tZkR4e4ACGjTRqkyPBLiFSe1SpME190/NRZmdA3n0pUyQZbtz+tTkqbySe/JykoRK1sosIbIzNMbjP7Qsa8zd35Q/IRg69k9VF/1ulTkKNQdzBCs6dXYXMHf5CtR1TM0m6+57YHxzmRFY8i19/3mgtUhFX3qsYBVztIMU5A0Z68mNpacxbMhmhhTqkvXzilr5fBPrDxfaLUOHuytZugNgHI+k8iYgSTwIy94YecD9VYrhFzLX62cVNaTyFpJ3b+zj1Rkv45J1aWgKY3RNTLGPRQIy3R4jT2GsQRbmUo5jrN+BQ/eTbo/c8ktQATLG3qw8zunCoFSWKlYdgyWV0Ir5okMNFasso8BWsndwlJ5zaw4maZvO1jAIRVE+h1EEwOCnyBIqFLRjGcvLwKMlXvYZdu7jG0uswvSa5bc4EAkRUkYyH8O53iTqpdryOzx8WaOk9rOvr094Z8mga0pfMu1l4bSytk3pHH4a3VxOnMlp5flyMq6Q5yl3mNb8QjW1LYOPjKFqQ1L4AaY9SHId0QSXvAmst7Gzpq17cVba7qGj98gKJGtMbFXTaJ5GFBD6MKqpIG+rePxqSgHGtzhgYR2QYX64DteyjZJCa9n8nT0twqwzqDegVI0tI4Fds+Qz5b6KIzEjktL6oP8DnUJPltl6jw6jpM6B8b9KwHMv+JhV3ScUTehDaWcMt9Xhs9zwyi6JdW0oZu0Tnf3SA3nZIFjsJ6iAIl7y3iRur/bWno4PZt+bmy55duNxDa6cFKHKZLH8IKhhpvxbAchWneDyxIM+dazol5eoWPJ/R8A2Mu0mq2gawr5Hda3Q+22NZJ9/7DRYRBBnWmpFez/ytM2kV9tg51rxsFkZwNk16RoPDNLVZtQ2Wh7LCItC2lRJrpMryiMoJa/I3ZB67iosM+1aLlnTuIxJfx7qBxhTB1hF/W42YXlqIagi0veaRLp9TzueKwvWHXIzbkCI/72igfFjRDNCQJLibxvMgMkZ8E0Wz96fP4Ofv94ohVo1iTHrGeQ1wLOqC4QB9MQEfnlhONIFs3zBUQAbA0faUp3o4N+6dLe0PIOAw56CIR0SJtsSeDU6Y3HaeM4iqRAXQ3GZBMVnxfRPpzWzpNcuCFZHG6DM/dW14qzJm8kgslyYllgL7mntHWsKea52j9yfWQ2eyt/VC+QQnhguhbWVDjZgAxDzjgG7MwyiqFMWRY/m1JTc3E9v1ZI+o+kWH27NkmFIDs4uuUXJxmfxkDbNc6wS0Wl/CUeTqKUvN+uSPgHkTVgkKutsnCM0IjFCAJyMX6ZK96u3SUB6YWaPUu2kZTx+uEgMevKIQjbLNe8oRHbap6B4eQhNAbh1s5n5TVsUPJVbJILiiqcW+lrGI1xLlbc67tQRGOq4x2EWEMTNudpEXLk3oRwYrvAnXZTtbVNyfFkRuBU19qsUVarvtSUi3DPWknummkrgllGrhIbozCjBEXEA1VYAnBMqwR7k7cGPefNy2rtCiOd7MplF2ZvYc64vHYlCt7EAsEpzdgkXUjbi/+kk0u5PQC0PVwWuc/ahufIGObMyjT1S1745rricm1djTqfpkBSupIEz+JfHnv2spqbqhfdllU/OZVtf1Eca+0BA/BDUjg5vWrg29KCiK0TH/Yw+9Nz0VokYinCN5Os3DBFEuGATXG7E0S/B5p2E5xr4nMCc4Ag9SRldKBSxwmPHvaiP/D9u5Wp6vGY+F3in6viesJS9Kz+xSQF9qvEbHr4199Uw5fq2b1n4zrdK8fk0LbzYp1Nidc2eE6wj1AnXiiUwFUTDXe400JLn+ckqKvybXa56jdx0ymbyMXev6NhDyVnJPgBKXLp1Qbn5857/rEVfpuaeDtLjhGrQSIE5YJW6qmh5cl6vf6Q9Cd6Huo2QUDOtYHtqDeknO8Y6+XhprdwwXRbSl9Hc8IA5go0SIUI1BVldsdrtDPwCETfRVK2G5WvXDMUc8O4Acn8biIjYhWXFJMvUwifxn+l34y8sCTQQVXOA14Hu3Owy3cZHHL+YiUwvYm65WiqAlQYncHiYMYQMV3izMg746C4YxyDDsemmqs81n4gEXtkwA3Mco1+xysofJYsc6lhx97RMWnedKSfpeI+iD0K/d/13Z4XzhBUpKR6oq9fFJpR51DO6je6MOr+WXDm4+CtcarizQRpcsZxjZcGOzCoNxGMbE0HUMtJPm7OnqSkfL5Bdq2zn9be/bxW9g+IsQUzye5zV7r9OvZlFUgQ1eTm5u5CFeX6c6QC+ZoJm0WBQyIqq8nmgnCEVIb6lZQp3E7y3UvzYegir1kKahuQYuMRptxNpnGVCDAilAtT3y/WaNBjsPrMwZxGYhlV/+JVq7RPajF8cFUJy7sIhbvn72Ub3/pW6cMr//b0Z5HNFBLsmhdsXWeaf7dfx30+Wwczlq64MjocgXeTQE5+FJP6ECDPLHgH7Tq2/bYlQ83GQu/gXrYKB1ipwejjwEn7W7Qn33IDrjVHKo5V0ci6YQYEeiS8negKbcxNw7hEcOLHMSvVLu4dvnBPZiSeocxKcH7ImwKJu+MQ/lJDkH010rFz7rIdY4Rjk6L2mh8+ISxyxB7d+6yTY5XB/OQfLKoFDmsCipkpleUn2j+J3YvLAQXJ/WIR0USmMemr4tjyzjk1yiyibV38eV/OKhKBg5WXPb9lJtgr6i+DWYSyjy8pKtKPgQVv3ldBay/ovoF3btj1FzPYJR4T7XKCJvNM/saQ7pUxh86l9NI2YUCEf0Hw7vOn+MwqoAT2EFhv54/qcpFErmQyvxKqP9VGD6JTk069YEq8rk/Z/kPO8XIxJ57R+oD4inFjRaJZHTD0POgqXsMPUP6rE8wOz58UdvPxvbA2IU4bK9+H4vcB4Z45ktZCg3Nq9RQ84j/73Dy6UXAN+cX18X+3m8oaYRXsW7j+GRLXBJ24inik2n2eJmc0S7SsuHjXdyY5G+m42/Ff0GiZi4ensr9vtXpbuRckSduOkd+KoqhQCFH9+i56tiqIMiYtP7xBp3N0uqaogM+LguzDF95Vl6v0jv/LjVRo4Cq6BBsNDRFb2DgS1cZdNNZ3hKskU1e2u/NnrRQGUimkXJVHsCFt/uMggMjF1l503Dcjsh8Id1GvbJ/C101mTXfmAbykwM4b5JYEIJB+fB6Xe1sWTRhtLa+InU0+ELwyGlpav5aJhRlV/gZ/+oArfc51jmmP+msNHBYtjPNIuPNAT3aVWmcL14mJ/j3MgMQoB8wRW5CxSg4O2G30zlUkRgScQlePt2ptmvsx32i1J4wLD211i2ldlOYCVXmDsjuvRnJGlX1IbhZyBjlXEKiCD/F0uw3zIcEeJH2F90OwbAAFJO9K0p0rT3G50WqhrOPCQ1cDJ2VWaKNCJ2GmwmEUJIX8gYpXEKgXRfEYL8bU6ZN1P/721yF6HTGE4O9/6eLiqyua0AVh/K28yyNcOoAGvdmBDhNtvxDDlU/hWIKFOHcFPp4EvC196+2GV/je05CzhtIvEBqCpLhe72Cv4dcnssLwSTksRcUcNHIvTFEFTpXbN1QYnPd6+2IEGWke/yNr/16dAQEzgodG5nRvHL563AFFnsUEXSCmeYO329CaZ6rjvLT0Z6guw2KaINf+ZikYGT+YQK1pNRCdld6hXNUV6FeAOzMowJMkPTDRiq91COCalwPRFWFUwJvL0oKm7wENiJsjuDViHWdwHEjUoYd4UThuVjKwVOO+8HxhhxZRN5NmHZgqOgi909EI0UCVhcN948gDP2BM8r3+gF5y9dAk5LjA3/OaO05A3+K302++vMYycBHU54ALxQPtj5whtJ0ettnR3exp2oGk5p7CgnJeenfaM/77vWB870FbfGrIQEMdLCv/1Z3tBuV/+tUSqsQt8wKod9sJAoQbwYMS1EkIA1hb3+6DUrGCBbishDIWOJX9G43ukgnfRzteBfIdbyReTeBaQWR6FPSjnCqhsrVVABow9WPEsGFvfnIhAN90msl+WWz8zDI0wn1AjUSgdA7XB+rZXI++4Cqu198FjEAHKxWCYfcKH8TTnz8JZ4gAI9iGXG3dau5KXNyOkd/RAdB3sZGeqzLQmG8pjjWF8cbQVa9YxemCRe7aNuLdnKnI5E6ULauGEiEeHVdkCjc21Z3yko2Qgn+kGdiCFE4Uo0f2vk2J2gIU8kEEmfzL27Tt8FNTvYdl398xj73dcwidIjvthY+Nh6LHO1CIWNGpexderYWpNaaQb1miKZd2vjENvX8/6aqC14bEwmip8SP3dlhbBYDo7/gILKZKL96qC4xKUQbd8mYO0/EJcHe67MYlOOzXYYQthA1DWg31ahwGmi28qwnHvYhjypaDmch29Dp2McoWeqb2vNyctTHdvCQmyTkKBwGDtC1h6rDmxdDFuMgwxswiVb26zm83eLpqWM5DmE2VD6YCdmjmiZkuSQboy52RFMZdLIW9NNHizrtvvEya7kxd9ZbjNEWglW/TBOMyKPXME5/DOsVBd99lBXEOSc+SzRoBge6zU1C4XezWKD3tooEXlcPfHerB6obowNlicsWR9fgd2bOtZVRtg0BXijCu7Vi4RK/Yd9h/XjgRsnjLGdZRGP7gkH5Yst5gSNpptxhSFRpCTgMdv5Bz9n7t+93mFrIqVkUc62gu1MreR1YHWLyiNg9zcKTXV44y9LB25ZLahEU6UTkbFe+zO0sD5TIsw9GSmeAIFb/jqrbA30O40wg7CkFAnwxOBLYubHoeKUuKxoZcV0jZBFpmW52JNpbIDs52dLBkasNcNhZAfBQ+DCDohT3vseBOwrtTbR8CxAwMfgWJiGyhR/GFmuw0pv34O0DtaxA/F2b5tJMn6lkuhm37Ppbxi4wleFQOxtSMylmLhAIUFdKdaAkVXBglRYmcYtk1z6Ge0pmE+I9ckzhA3MpjK/ze9ThF7Ppf9VZ8JBtIRDpqJrT7HJw/RFCE9DzBINUaLiLVMhufe2gDiaeGcGQsUiuF7b3yqYOZI/eJb6NYrvoYrT/kPCIf9RkEP4ne8IcdFDdsGJpVdkm04AR2VlfBxD87Br5AP68sa+hZ4Udpo16FvONsi9Q+eCafqEtcmV3bTJYBGdXS0sLtF4HXZrd8dhzaDidh5fdl8MgCYAxOTrgc6g8MYL2aeTbg607M8QfgAWXsivwKvnbsZQFC6B0R8Z+BQW6x027lMjfct6iHBCxZuS9+AUe3rDf9o4SY8/LTr2rB+Miq5yPIc9BByx02f8tAj0u51ZTe2w7QPdO4lftPFEzik1hni3mcKYBonE+TG846AKzR/LDubtK2hJH8pUyATVOR22sLk1/u7h+uyG35Si4z3+m8W1pWcPSdRJyVlSdLPjI29R+z3I6kGO7wF57ZG8ErlHBE8pzssKpK0PjeEthsWPwQeg0e80/SNkbqDVSD9URlM7S8JGUM4BYeYgnE+DvmO6U7ijK2OXUDHBTvCkS18BB/OvznJreQo53A0RLdLZqckjCDHqVIVpJULtDgxTUc81xDyUgFry6s85fZnpEmnRZUUcb9R7KqHAH/A3JwLE54mqra8d5865qJi4G6WDBFwrhA6ghYERBuSR+v7f3A2p1IxYYqBPhqSEddeyHbUJHIEMi/mGm7T8yrPkGqowiL1q1dJro6jWoVJco8X+xx3ZcyhdY8CI2oljVUSAMc9YT8HHFT7R/GrgYthjpO257R4CEYDDYbLFBHm88jbBjbz7Rv2H2O96G1+UnGRIr8eMtEQJIug/WEjez5FlnUeJqg37314+tVDfecQrYeV5AVyH8EPO1Seid6c26AWvDBsPgHw9sBsfflN+NxmKbfan9wfQk2SBVUWCZzpfNg1lAxC6M+LBbf80L3TPfD1GHLWWr6hSfKSye7o9Z1BrNksfZUZ/s78iuIpAzC/QKdLuikSgxzdLv1YYckxIwQ9aI32Rxwhsatx5fP7Z1J9Vu0IcpJnCJNFvMDTYJy3kNDCvtBQ2/pjKTH8pWlmBzzQdT+1x1C7PMeUzfkO3BUSX2Wa2XB0FtVcL/P4LOtDwnP4D7R5ivkjxqY8IAkPkKaTXRqc1NfltflNbL7mS5zUpR9UUKAAY4ZXIUToJW/4J2ykd+6SmruRLU4zGpg2sTmgVOshGykLBUcszlRA+OVLKP0ym5BBeGI14vbDtvXyj+0Iy2RomEDbzolXQ8Lz0Vr1pUqEYdbSAkO3qTQC0k5/k0vZrIrOWWA2gVtLsvbklwmZpeksSQN2hiRv2ipnm7RsDevbGchRl8MXFpsqFdbn14s4YvEQY6uhkFm0wpG+LcucElmEEPJkNJCXUSxoyq0CnTlBeyye7R6lEOaN55B759Ot9Utfe7w1XdpU6OJEfq2zUOA5FwZA6uj7fFEM7aemgFQnGQ+3BWpl3ecTE4/QXeL3KGfSmBmXOF8aemj0xfmSPFRdFM31Kj4J6tnpHg0do8xw+Lpl3k8QrWFQK6yDmvje9ffCRo+k4pxjOpMVPM/g4M47X9bd8eH0g4Qcpy1vPp4CwZh+EIihx13+j+vwdSdaEuD5wSa9Fsmb9eM5rNAADXAv4h4vciJSlvQs6b3sQ/izICi097xTkdF5vLJJKXMq0h8tQGZdP5MDIzs9CkpR6/ztyyRG/LOw9CJygNH32fRDfMwNBwiSSm6VxUraPFYTvUc9jRyXszGRAo5f0kLbYyTkVmKgMyKMiU0O5FtuiRB4DDSVEZ3SKcnAd9DHw3UBX4wEdMB5EakVT437CYiWl2lZ1b8vswlqt0z8xP2KTBjy2pK7USFq/KBSS07TEpRQkCxYbbeCBREoEzVITVTqSBkS1QuCxpQMClZ1jfs9ysJifdIxHmLT3fRBiNrXtYppDjGsF3KvLCpiw6/560CkF7io3pzHf0jwT+KRuchlWwnj0TkcgwE4vyi33qA2V1pgYB0/PKXkLbbL//w2zOKCO5wtTH7JS3d+uC1NdT+vnN9+zQd/K2o+2YUFcROZD1f+u2tIz0eItjhupSVi6NMScy5C+fJRVFxi7XmI35DaMBF2Fvqou/bJdYntLJBNASAmfN6xCDcdNKi3mn9ZaRoaOcHGlxp7/1R3slqCL4JYSjigRe8QECR2fs0QlKj3pXcAnRI8yNPwNunC25IyzGdjMqk/NkJvs0G5k4VK9Iewfk5x1PERbYhIvXcvzu53yK5uEDGjb8hQ3FkbyrPvBtLBTgQcUpH9eL1qGJtZHgOOOoVOwgnlGSJxk67wPmtV2Tk7yxY4Z1Ysj7Xm8lG7B3C14uTgLmYAxmPqmZUi+d8RkKYz9CfYi2CSDTQ63QtPbxyWDZrbbHoaLYWeWwbfyKqqqU/aSrbKq9aepaT6NX2wngVnG069/vBvJffFBTYmKFogcb/9QgHttlz80wYZgPQfdpLHNMm/1IdeA16j1JsJhuikX0NiZx85T6A5PowXq8JhbZf+OkXngYJf2WkfvcaIL9ZCx3IedD+xxVEaAbFj3lFkzg+ApuyHpptwevii/ii6eIL/wlTcI+nh61E3jHlQeZRJC10noWyYo4mk3DEiLsI+4S9Xa+/jjAgjPUuoTCc6/6Ok3ZNpDPZ+U1dHSbmeH6pXPQXkQLbcK3+rvd+f3H8LswdniwCqIWdn2PAeaqm6vEaidaFzQ57jwz+QNAtuL6QZKeVIigU/WAffS9gTxdbZY8Nsqc8NRfuKdBvXr3pn6NFxvLjGdQlQLFmHT6O4cg4+49Vamd0AVks5vheO7GLmfxTr09GXfMJKkHxAFT6Qmsh974fOmqYTwebYMTTRLm8IzM8I7xixnBQRxitltw1mVDnhtyiAdWJ/qChTFHpCiL9Z52fOl1ubkhZYIXrdcyW54f7tVyFlGRfRZa45oRyZkDe9TS3RIDdbUDGtT65/TsaCMFkY47tpx8vbidk5LwcYPUWt0kQ/IrNs1hNtNFiqquOOgNcXVTDWfygOxNf+1+hsE4GndAZBI2TyEwv5iCPsIVCCASf1QWPV+gxwkytCUfnN1CULl3l7kWgECbRpNlwieM/rlXpj2zFMTSTondFj8xE1NtCYjSunpSKCgk+EBAb3jvAj0LeSycd+MpmEFj2PkpRqFGJpmw2oQ9iRqSZx0H4PFmkla4nNKwe5XdoT7bmXFr0N0npiI7ME4Ubs8HwyEGT/n15sz9cOU1h2+i4JGfG2JxG4rc60CS+Oqriy/CrMiy6QwNTwFh0XCWtXxygKv6dmoHzlcPqO37jBKbb/Dwl13+i2KS0K+T89srAvy889jhWB8A3jV5LMWBwxQ8wM+wQejaVZ56atOixoVqoYKtnB90LDrT6Q/9Q1RDkAmhu1c7KdsP4fngwKijba5pIz59RGxNRaXkZsBerOHW/XE40suzmsd8FWcKTQ6d3s0t2ZBvRMs3vQNVT+UgNw5Ly7W07AAWfXMraOSPFETJh5LMWWMYpHqLHGSD7sH9cy+pVLUSvZ2l8FxjhOuVjhv06XqbN2f2IXgbv1iNA/1NgXv1/X/U/zh0p6Q+TSJxdmSvaI4LXSIQ7HmUQT027AkGtK7PGpaSNjmpM8JYdHSKO70iNM29AHOyCXkhoU9FzNBMEe1VkCCu8kjO4fjTTDSzeQtFzuBrk6jJCeq6lckE4To5wIEwkmi+LrXccVeMiYaBBYZnFBRiggUt/JKaj1KI/by46tU6wqHR8zEdoSgaxK2I6U24wc2IL9mBf/5MqMRCDoUEhQhTf8yf2V1M+ghyem2lm2ygS9Hd1+iWhS4yQ+oDz8oE25TmU8hfxPvfinK3Z+RoO4frFGrGWA9s7H4NuqDJCBlESJPl+XIUiQmsCn/sDvYcVRaPacHD2X3fKuiVrmx2krQt/qkiwk5KktbRBtHd+aHNDKVNdQGzOSJbJTXWk23ULitOFJI3vor0ncW0WL4/BGaqyH13BvyHMNYlbjEW6ZPb0VBJXrrP+Wlv32Dx09Ti/mqk7JfySZB0q+8BkNe20FfoEE7Ik1bhStcj2AWKs1m/fj1E+szIn+bYtOlpZxBg6lOsbHV9I0rlTwhlmGVBcOEoq5IABzQ5qgtwcpkTPguvwJf/NyVPNqpxK88TFx3CBWEdMto9HC/UDIrmNO6OJ38K5sYI2oztKxEISg8Jz0YDPSqbUt0jVVLyOjHiUB6YghgAaT1VCQ2sV4LRYcmpqUtOTy/08mPK2MPYlRAW5dAGGiJm+jAOwX5/t3LeBhTJwBPXJdrK1NK4epoO/bm2oqBd9LYEncumF/UvVmVfiubFVm4hqzDDZy+Ix/HQuwNqXe/SDoKMTGqfOzYhS2omZD2LycfYW8DBmHnczk1LiDSi2+r1q0x+oxtxKHuBsaqnyN1MIW9ME/KdjdYHmg69GETrbEt1oxYAdxpwFZ4dNLHebTxdHztfG7vbxcQPh0lK/iaWVzAIww+Q1tySmGqNKs=
`pragma protect end_data_block
`pragma protect digest_block
3488cbbde4cbe9ca4f67295ccecce811df25b63fe3088870bc4b2fa3a222fab1
`pragma protect end_digest_block
`pragma protect end_protected
