`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
3znGBgFMVBhVj1G6YRajf0xGNYgfwibE1Sep7e7S48ABE5f3Lo5zDRZz5YkyPNiDaKmYtBrXd00FMw9dT2usXrEC45n5MaGYnglRUVPqpcJRQaj6eE1e4jJwokaWNQFcvRVG4CQ8qM/14dRe2n8MgMVUerZmxU6q3hTS+mIp2Rp5Stiw/aBWCAdk3VuT0beKpjdlY0wYQ3WUnCLpBG5rWmhHbcHi4xmDE6skWl8I8XhqaOhv+O8JLZY0UrVO2YBboDixyfIlrE4/36gNrU6Gs+55HW9J6ckRBz+/carmcsio6BlFyfNbGIc8VKzKCnWWZlU03kOTiSSfB/JM+nDefZDgjRSfJierGXbvQvVtADfvCfe/dOlP/qNoldLyNJ8nIG6vWAeA53YNq1CNlI2krgfHJ3D/A2jH/hW2dKPSTCWGCic50ThKviGababy8ptJelHXgK7qg/ECcRKBDmrnnnwQTQtSJZ85DAQVizsO8Y/RARucs3r/duN1BvRHkc1D95gMvQeIauws3GjUgGMXZ/+cL8Ji9lKuZimelSyLm7BsHRkgYMOPD04bHKZFhtzjuKXNl+qeGWeWDryBsbWbTa1e3hGbvS0TbZFjdxKPiuAV6B3mk14BeQJcWomPpTOlSxuKw6ZRHRShfpv6OzVcXRe/f8+E4dTyF1ts35IJ+/PM2k9MdoYbmJRWsP6toNOEfIDA2FQLG5irYv3O0M7hEx/EnZFHJ49ptDUi37+Xh3f4yXQb/E05b+Nt6YPHqzFPkX/e2SatYl20f1nDyGtQRCKUGPqbstj8sMCXpouDbTBx8i8N8OwWn6giX1ex6v6nw2/IqDEjtn01He14FlFV1cYf8gzGdH55ltlLbGL1hmKgVB5WqP01ZRD7eUwbmzaqL/WtmkTy5VJOXH97A8kJD7DImUz3w8bnfGiKJlegRLmQ6ngFyyZT8Dza0E6bJTZmec4UUdpFRKUxEbkxdM3dXQch2QDogw3k+jbqGPd4dhY0wk7mw6UvO7W9qavb66JQ+bEGOovaJCA46xq1TbPwh0vvA2vMwz3WPqn5Y/A56y1xAJpDZzWxpJsabEmB9MJcmcQPMYJcij488lOlKpWLA36UjQEa65rob6m/uq9XS1pFkltmsAvcSBuLff+jzDP0uu/8adhVsn6aRrKE0hxVOE44P1O8oO5njOSKZ/K3Bwk9Hou0LM7MijZTZE2Umeg3u+AUersFgHv90A3/hUTosXm8eB0zXt0K4jn/UQFfwnHT7Es86+FRSVEUqdBMYkEgr3iG6OCJnYMVtPkWDnohiOsRv5zl93i0TcZ2RN2rqH3cta350CCW7u9WZD5pU07gCrfd+4/+iW5ZucPzImf2ANpPp2E9U7w0Ez0TwSoYpzCB03jX4aifXIS9t743LqtcOBTMjAuPNucKngWkhtmdM/2r229ekmXQfMA+Hrv5dmg=
`pragma protect end_data_block
`pragma protect digest_block
df4abb2454e310b08b27571cead4e3d0ee34b1404ac54e7fe75b0c6fbe39ddff
`pragma protect end_digest_block
`pragma protect end_protected
