`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
CftwfB4+O7nAfO4fwYDfQhjRPX3s+zXkQvxrDcpw18Gw06HVqc87u4wAzjAd9wwxjl4n5iYlVmcHgS5gRFfLRj3AVNRSXK80mUXKNpEoauAzJAS78dlULMbDekQfs13/XEOo2dpADDCNVQpIgI55XtiOePiIPbYyf3sWOL7bofMnYPSm/Q0NHsBxsQlOcO0CYoIM9BCjKWLhLUoCk3qC2OWrAkEvVZUUQWlxNIMxoWVe+7cWIi86i77UoZUPEHyhWJW+D+1up7/BkNLnoHTxtaBpVOteHJSrUOFG5OzkCT5Cpc00MlZElB3Zhi3wHj9ehr7yIsiQnXFrPrVhCfuSt8Ry+Vunu5T1VJZWicaHeYpVyWEkjRfhsqiQu5Le5tku0T6IPsLTi0pfGfK1cGvbITnS2HN60MAo6EeJmpqQW62TmzIMLCllHn0n7PoMcfd1jryXzcKTWxJ3+vL1TzOeQBljylFChxkhfLwN4QF1oUnGdndoS+Wx9T5dgFBgn273OGbPD0wMHF7aTJ+OzmDr4r14OU4kDc4nNyF2mmJj76ZpFaWivI/Av4+ygm0Y9XBUN5ujueGWHJ7/VecpNJJOlk2t4GNLItaEdzrrps4yAdasb/MtWEkilqfbbGoXGXr/fj3fdePWrVhB4YBqa9uYyKy83a+CD4FsHvdc9jJ9zKZlZ0oz7UQz6ul6m2uujUl3nXqfNPlCOpSWcVI7IPlT6StiTUgX9c7Yz6PYN+c/UYUNh0WSTP1tv38m18b/wNBcuzo+QsEwVqm4tiFjv/p3xC+v2ljygH4EmfGDttcPCCgIAT/PTFVr/YI4Nm954selLDCLrt+KBse51dnOLtZ4yIxQ9XUYJULlkaoEblxo8Zrc4XRE8EFUhZNvBpijI28wfQRgYSnhnvXqnAPQxLsO+JI6XJg3SM3BlRqikK6C+Npj/YENzuG2iUMgD2dBR080qTI6GQwh4iuC3opX9gqJkYzQnKnEMifeZ20YzB/hFmO9GDJMKGNpF7RkxyNEc/xYQJlg7P44jGsm6nCQnEXHio28mEK7Da+m4IlT5ZC3AQvChkPf0Ojz0+8yRcchzpQWewZe/yHdgb8J4h76yByXRn1hoACH5mteKCNRFQEkidt5sga1L8TO5Gb0inRm3T076FO32hSUmPxjPuziaDaMlzV/kZfvjFV102jssSoC8MfaAdO8YT+WHI29gi4tRgTD1HmIog4Pjf3kAyjDeuQyNo5Nn6oClAh9xQsftBf4PP20IYCtseDdLCN6YKxvVn0FH0B0M3Z6wYhxyzrK1Q8egIbHAu/0t0cc2j41JO2ZMkApacCO5YhP6kzlL0O/e3vDAm/NFn2Ty+CEUP+tgXgIopEXrEDd/fGpRcnHEM8m1QpSYrdrXNri1JfSXAyvLM50Ho7Ssf1IWR/2O87G/NQ4uwHN3axBl8B6hIQOwkeZwkQ7ipz7+4vSC2atpA/LsrreK1ef2gsV/vFG4Cu38sYmVKxfTr39UQFGIoRONHmSuzi8u91Mnx6NH92093ldx44fLqh9tEiU9QWYHLiQR6Pseaq55VLC/wFDasZmH509VrfC+AZ0jiXXpvgivu7HENp6X/wpKXkWk3KxjTJVBlqkYxRhLm/C1VWTxnUtCNkO7aNMkquS5H05OBUu3il8vv1flSrXyK2oQdL6bZNbucZW/2tn/ElSMO9OeIyA04nnsluQCIUL1i3+r0YuqK4jfnc3B7yOeXp/I9fNBNWX/qHcD5ik1Js60356RjDul6Em+c8vt8/cx4sVv0/K+QEJEZyadx7PYL21Y2mq0COoeZZr/dkDM+lAzsSxduD8n8RrARJrOvhSVGI+q8pUtsIFn/PsVY/oK9gkSmCsRyIQ4ybAwsIYctglYPWwz5QYyIT96XN/a3rXT0yb1ObYvfI34CkEQ3025iZGa40nWrblOexASc0QSzK4qj1atkkpR0NfSsEsXjrlCP20GRFkaxxEIATHMQF0QraUSq1MRNXzmzcn4SBiSL5ZnDfuq56ZZiUEeViKoeCwZYxjD3uFnM8/Dq6jzZZVuRjuFdFiD8Jhm5n77miCd2TfNYWQJHl8vHBPOJgnSZUJS5OAseuohsmWnAD1aFB5KIiWrYxEWbIQXKMm3LH3pNBNZS1zV9cnRaWtvoN04bJC8JFZpWZf0gd6aIoMC9uGtY9AbaKtaDwXoDD5lX8QJZfOpUQstoS+zCODYEi0WdGE4J1hUfpyZNGftltDJu1m3P+f7Xqw3ahFs0CCPxJxQXeIIK5J/ycaGAgWf70P7LF9HV5hlX42zY8K1RIox5u07KHGvfnjKJyS2F+0Bfk/932sgMRWPqpXldgZ3WU1CwHrY1RX1oaWPrh3KvL2CtLTNbqL7RL8aG1SP6x+VOBFLd/20oSvNQqVNyxxFr5oL0pmgS1Vk11wDdyV2lN8v5vR9UE0+roYdb6nuyu7FdfWgN3zR56+FPdNizdnjW400q+PobIeBKxVGB0hXVklSE265VG6zCMmwZFH8Glh28iO9TgGoRlHa/ikttcjPsw5HzuoMpaAkuXXSjwF9+S9NgSxBog3Kut3xePDFOk02ebpWCo1dZv8wufjyjksPbF5v1wD9B/dRdcHBXETpUKYkd+39iDg047eFmYUCltd70OMXKy8KZ3+pDnkD4SEmBvEZNJ18/0fWYwtfcL1gzsulpHAEZoN64vWxdkpZpOGVRyWHlqP9Vyo06XkMG40paLXCPpFOikh266FS8v5C5l462aP5KhzA1eap67lpWoJlL1RAuMCcQXogtFow1XgFKHedfS9LwtJDnoWtESuahKQFiwjnFvjJrfm9WcwYZvoMEe6Fk6ZkK8w1ETZKmC+rE8Rr4XG8X0DAElNaLvlxsx7t53QhqtPkBRgh79pKh/Etyw5ZbPd53psFO9xFQ7352UlVVnCfjIsarGYekt31hlzth23kJNQxcllzfnWasak75+Cs5WXB6xAqw1SWc4ba0nyuSwQd3IE4bDk6MqY2VaVB3eZ1FskbzWSbz00oy4+0+nqXwTTuJD6croa/arNeG+3ik0uD1pY5hY2VCEoJxkTMwxW65H1uwcZW5qHLZpXX6OdvHR6p9RpYAOIGw/QrsOj6A+euXKbZdejECoaa76YBPttdMMh/vM5JLRpLM7I4zk67tiIkFLjygEsR8oxTvchTjJ/BXyB7hB58qlk4UvFhZdKrihA94xXdlJcaNTkMWYD6SY/EEtCQkUw5D0XaAuHMmPswsEGXpS1Tqfsrgx5AtS26znTq4OunejXr2GjHY1ZwmI956qkkr46Yip9is+kS45oVQMNb38gsK3zuxvZlfV6mt+TbrNqNK7l47d0Q5/eZcDW2u6d1/zoNSjT4R8yGt5/cbHvNBGn/Ubqdx7d1T9/Rhr06nf5gYRKOHXmaiTP/K7/9arhvg2DFXd/hTQces8vGjb6VhuqMvpiY/+lZR/v1sXBqP60ysyAe9k8shQVNrhLjte1MP1u8xQeQo/Gh4Lw4eKB8fK0t+EbvnCI9joKAB5tRpqOPc6RuR+qnEJ+DbZNPabhpYfN64fef7pb05JHTPMGUKiiQt5Zp2oAK/cyId3+dwYaTsxDu/wSczJzkiduhgGewfB1ykwTKpusqZ51s8+HNx26pP+cl1fSSNx3tPt1ONrSz+pIJaZKXdwhjn+BVYGP3MhgP0C2tJ4lRh/otF+j3ZqB8eJdHgyhre2licUiju0sZFz44S32o8CjE1IucRICbuSa90K8fB0KflK9xPbCyEYPrU3VLxtF7C4vZVa7vEuDxZdIlQDEcTLb/LxEeow9dmYsrNWCG/df2HYFQuIk4G4ykT42HIqk6BJXXctvj7VB2Zo8T9CYULvjo5D4JwrMiFpx8tgKlXpCnSTvmEAQYsuXGGjHFv8CqJinmx7jywoPsEVQkUgGA0AKmDfkaZkqon3zkiY9xfqCFehU4VmbRHhDCN5nM18Y2MK1DOwGNW82uwC8dRqEukUZWcxr4Zt+Ikh6s6T2wpQbYYDh1WnnhzlITPKwiK82XnZ2pz6MtdhGddkJUcS1MrirhQI7GP1NtiZ6l7+43IkVPo+a13YUPfu4WT1m4ug7hmMTwKIke3OoBmOUwqs5C58wME2am11clZnRA0Zkz6lkdQ4K38qJeyqmfW4i7kXU1DMEVkF1JxUNz+LeS7jq8jegg3CX5aiFoxBo8TvyuHl6nmJ0LMWeEMBAGg+lOOX4h7DYFh58rrESQzPGY3kd/MIZhuMwMfPmJML5JKbSVn2rKs92WNzgNKXib3pkzl3HXTBRQoUbFP4HLNiQovx5O6gg5sj6OODuJw7cMaayziXvNyEZiNGjEMzpPqK3QVFWWkq3u2XioDlIIyt62x86xOnrI4IIBcbureJ8+n7eZiq9rajYrbm07wFaoipW4WNiyFbHv54BaBYqgBqU0FpY4K6Aga5BtB2+NjQ8p6ykkXSfMr/2XV5entsi1RA7pJ3/PobspfuYk47yclWxrHg6hg3chF02SXMJ5Wv7KYlqWPD4MeJ9ft/Z7U1b7xoLNz8X6Klwzu0WvecYikA0UVtzqJyEIbhk3QZ5+RoPdNskZ6wsglFDj66FIfh8DrmVBoZlFiXw+aHzkClTVqJk7Iwx00WZHW0tMejMHyg9rJJxrkzvTYPhTwZRNanYZHEPmpyDzJJdI4fz0mIGRItA9DZNGt8biHsk7vX75/YvvjUBZZpP2aDPdMBKtuQTfnfTy02jMLnUekvzKHflkZntlDXAzh2ipOkQtmL2stijfDY8unajX1a4yc5AbrgD45+CuEeaiYLzMcSzsK0H9nIRoUFij0VGfBckZYM4dFRQQ0JcSI68/WWtrOpzo6OyGbbLvNhj/S27OAWwkrbAAQnzwJiK+rw8WPPQhfjdi/uurRlwU9o80wet8SYNNzd9rm9FA/NL/5e5GccFAnqyq6X+sTLHEsHG2oA+dKcnKfSzAdcK0sVKshcLEcBM7PyV3wkmG6lHAO1iLB9eX0aqnIuSXpNYdj4nNTqM5S7j7bomLi4/Nv3MAbADbgEcu0n5bYQLwFIpvb4Aywg5yURAX1/Droetpw1Bz6ZFbjMe6iHEW+zCUoY5nImiX5AtUXpY55e0NTCZiuLvc9CCCanP5Anw7hkZeRBzEgo3sbLCUENtEX+rxt5+SE1+HlCjXcMUs8H54vRArDXK2IfaFApjfY4G9jpQZxSO60z0rl8HELb7TdwO7BTQ7yePJloUfRCnuT/Hi9ueXroEF5+g8TQSPVcnFhvuKxBTQQEXKDJ3xNUTzIWzqbbNxBTFuUHHqrA281R3Q8o+JmHowpjmS6SEccAMEtkIBiMLEMPvSpSK8b6Tt8//7DRcndKRNGj74eM3KmP3Yn9UtMvU1RPh79ru38grxApR5w7cY3btTfRSVsnO2OXuCYa2SbBeG5bwUMs6x3cuQ5vKcXaG/GiKdshd2BydVspR0NxzDloY3pnSZFp6kgOJ7A+70zM9p9WpATr0Xl2qABVuWBk3L2ATx/a9yePAIjGZZ8WtZ2fWYZ3RtR4XcfdkuO8Q2sKni0XdX5/9A50FbimAdyz/e4b5vPgZAMYeUjYaIghSbuBUFnAv+zNLn+2+7G6nuMAh1xfxWQSFyBHkZ6jXCjLRujvfoAu/pKNQIpoCgtlAV/7AJGWfoBh2N0KdfCZUFDV7Gr3K7HCkgCmatJB3sMyiLCg5XDDTn53GS4UfoAzXQyAkjJBvLi5D1oREPwGddDXJ/qod/ydx4+yasYaoyNqXakREpSkdExOKATAaaX0NE08DvGjgkbu1dyYMlffiLrftrBR7JihWzz0lIVG1/gQOZ7mB+G1tzIBqh/4GVDxylzZE1/ZH8cu6GFZ/nEEqfebMObqTAYMY3SE9ZmdXsVsUMx4mHPcDn+G/83P3d3NgL9gtqcFmemTffbHnjyqWgwN8mKLUjKtQnuLxG/TX8xLz/QqwWQ/IipA95l/kHXO9iuytCwu2uCN0B7s7kMYjmQU/TZtFe3BcvUkNbYXceYbkronKT7wTr1GHxB2xy6jt2hiqL0GGy8BDOuXDrlmSCvmVI3ysvXZLm7uIjuF4XYfxzGaM0s5VXqDwxzZk10mrul2EenpNPCOFxCZ7c0ss4u6J+7eP+cDRDA+GO+1JK9K21n/OeIDWyRY879Ry2Fs2wViQ688gKPUDKirV8AdZ1D6zpCO8rKzo3Q4bz4xASbDwuHCx8t5LSU67kr8ZZ/GyX44pe1hS3vH+wVZzoNCf3PmN2FsWOGzDBEu0gO+cGjx/BNwlswpS5rAZrLFzBMu6Ys/j2XDxrLGxaACJY7PBCsrRN4ajmfKOeAua1FyhUdt/n4/2K2AXkqoVlXO8scRQEDOkuPAgqKWBCr5wI8SS/shM5VKHlXQ1EHju6ItKKOydzeVvZvOd+c6fbmsJldM+L394GaE1kgmnqppZD6J+7Q1DWKBY6BetovQ/tJSm52t/B+6KAzrGPSmu4DsSYo+OiQ72ItOqgkRzc71RmbSKX2GzjZN2DyrQrDsO7yEWZ8KBd90JW+XhpRRcV/7JTnf+ba6YBvEWN9t54fFGGxI+rmDk5CsurLLF9X0E30NEOT9VjiW6Y1MDQWEO/vBS+rphY/RARLqf2gklI2iQZ16W03TjD1reDK2m6L0Tsd5T7gN0kUECRZ3DYWvegVo9ZvrQWbG2hCG79jioMBqu7Ast2PAF8dEu2QLaOcH4hOF7viP8zvp+W0uAfZfaZXD1a7VDL3hRVMLUljzSa6552HEQcPCWnKAF1qEb4UC6pLIaMv2ksVaSvIEl75WPwHo3HAemHJ93gguKDEZPtri+h7CZaZVjIKAvVglIwTmUiEfCFxvsgQGrd87V7l/SAfXMEg5dsFWWSPeOPy9v+v6ixMltchGUXxsYp+OBusUiRqaxVV3SScdgM2r1V0kjXXtH2GnUZ6xa0ctQfaosAKounhMFBtvVBZodMYSh+X59c+RCb5hbyAQ2wFVkgsH0ESLAZG/pw623uypa5u56hWjD6yWW4xPSpgSt3C/TgGQEErMrWLnBKDy1xXZVCijTFY5qJvi3TsVFF/d31cSORzSbdZt7bn9NjdVtocShHYLzgrVW/9RuVdtb4Zrulu6xKOJ0GgPL3xrxHZlldMCgN6l24gNDEiLDlaIFtLIGhjLjLPU7l1fUgwwJav5402/TdiwHFoliQ2M0h+aatwWDFiJBccHT4hmqVk75ris8sEK0BcYXBT/0dX5R1TMdLSOHVfu9kOF/cdbVDZZFK74HXxLhfh2cYRAwWToqeqg2ReDmx2qSomdpNiK2dgQazcRK3QM6SygWr3zU7yJZdxnJ8Vkdu+gwZ2Ch42Fz0HLNw9tOTWUNKVVN9mi6hy/o7JZ7VvaEPj3v9cOXSUR01/uTGzGKDvBJVFgm1P0E+sgNmRhArHyJrgVkOeGLogYKoHidb8MfORa21aLv+mwfugsEi0/q536IO/gHqdDY/45M6TcvqSwwjQJglzOkB5qqdS7+tJ+sY0zR6mVgSC2jJYQJCA+nv4UdrcMmg3JY/gakCcUHXOJy0zTlBR/B9udr/A3poIzQx7p7rKxkvRIAn3rhGR3JJIuFMXL7Fs/RQNqx/00jQ6qfjbJ61S4VxtLHicUgkev7kqevpaIFVmN7iJCPM0Ar/BSq9HLruXEqHLDyhyHtueA2j2UL2Va+WU1E2FRho5ZDDPitD8KCM7ip39m0Ixc9av0UJeiLnsvC4GGZbbF0cC5DBtgqxCGb5NK3XmucGMAjLPX03T4CnVfCl3PnMaMigaojNl7SYm1cWbNGiBrayN6qmHl9eOD24fgkjBotYBnf+u8vQyz1FxVMVsVffjD5x0pzWh/ckPROh9v6J0wq6loCo+4I36iCh6nq/AZ7kdcZ9MOlXGbxzBL00qMsLnNvh3jPAN2tCnBY6ZImhpdqAih/IVuflq8NjdOPsc7BzVoNOGECGhRMktcmAQZMeNAcBWVk8mRXosnDdxaKenbgE45whg5sYP33AbX4PVDSKChGHLk+lXam6cZ0qUKOxEeTlVci+UwV6CRJZOebHDAUrqh+Gs+zEmci4SM8GD1iToM8El3MP8homTK4ORwHdwDXQv3cWGQQUz7Nr59y6dS/h3xM9VHfAFrS/7dG7RoBQEwFtoDLwk8mEE6N16CqH/KhTdqkLYfyA7FdU4JZEF1Ag/nH+r3Dexpfh3oSThPzmw0sHavieIfrPe29goMhugKaQIyQRY4ouP1JNxXWn3z4NCyabaahy5Force2ARN4HJeWEDKuj6KeViTbPJgBlovuR0AmIluflqgVcKNhOw7YwLiayqDddv0URvB3nXUDkiM5P0GfCHZHWqO/klAd/O/nbQPQ4Q9A20e0s+LlNX+lmccuXaqT3he7xRvgsQQpjfHN1ogfiRMcpLX/Ew4iU9X9eELx3aZjlvdsPMrMeRKjYow8uvn0SwV8ECLdtaMMVWf+0c393pZTtnjuLgSzqz4PoHPwYtn/qgnzksQ0GqVPP9yDZOkhMSJsYv9Gn4iP2YetxPOCoQSGfqHaDsGbTfXaaK3GZPuX8pBELnOtV5ULtU3eseE9lyku8TOr5XiajABOTFNVBEBHb40qckNd0tcBUzAppHoBVmxTB1x39eK7YG/Ywo7Z1wr3AYy+oXrKifC/IgdTjtoKoMtHFtES2c68392gnKltK+xl5K8zE1NhA3e9pFHCKW65unbNiRdpMe/Yb2qMqGlLB2AmWhMXti43pCXTvFCZf1HhMy4MLPumJfloLJaG9FApijv34IVtwqZOAor5mkYfLO9qd4l3RCktoBkZgyLEIxstZBv/waI8LQwXXEFYJ2CxWW0QNkQGIeUqojF6z+C33kRw+5cFWRGU0A95us9duHKDhCAwYTWgcb5VNoVKJtAmVuP7BPlrM2AeMIl4wRzpbr9cyqn0zc/soAle/Disk/1+t1IrZamp/Y9IuGcGCCQy047E1oX8u5SnNaDuyh+XOiuqc3W2SxmUu2fHHia5ZeY9JdwVjfA3EiL2JMr1bJOLPbmhU5L7b1ndBXZW2RHbwbOP/hFRu/ZHPwWtf6WHeHFZlbgxDBI60R0XgKJNnsumuyNP6KjekcJpDiHyBlKk4uGAKFPgfhUsLezMYJyzfPyNWAim/9vBBRUu6fRxYe6FqaXpOSW4NYcMNa2H6Ojmvd+XOe7ibMmCMy1McBS8t05UN+VHn5eVnxFrDwoDCd3eAr87Ogl0rjw/ZuD6AYiUm4hxN38HNhXpBd4MzPW+rbpDs/xo9QQ0tCOo2cBSLqhyxWotgfR5ROba0FEhOMPEv5By2EU7z3/uXAnXSBEPP7IVk2ZiiYKODeRy2VQ6a0Wq5gESlo2j8R88bpPHtIKWvnYxVEYRv7CKtZRRTajDfwV+oKa7rOqCKtmf+C5/RPFkNc6DyqutSfKdDZ5Ehb2NUghVTx6TbLhvuDaW+fsBu/HB6k5sXrAWhxLoKLQjHz0Mm5jJ+STCO05+/pDmXMi7qAvSkxDrs5CofpdSaT6PVQ3YIqtHODGw37/LdrYk8XxEj4TtzghYVlLbmz3ACsZR79BeSjP9p/I1bFcznbXPd3P2oUbe9HyC1xyqS4ZvyI0phOmnjHz0ELGk65K9UqzU3+m6cBxVN0mN2Qv5AtXaqndj76puXrTBpxr7L0+Aa8gYEnOd2nYrFoLoYe2yR++XfGIGVOblhnnQQE4/zOrsd+Pm/+pypc+3sqeAGFwMxUMimJeVIPwPzYGITSi0pBmUZVLVSzB1af0m5j6ZHnh/7pVJD9ehW7yns8pCWyqRYUhYjo/lOJV84B8O9T3Vib64VpOA5NHDZfGpE3nqroM2Yr+hJ9vGp0djM6W1O+ptQ30+fwMBBP4860tZg+P1n5nbYq8Y95o4s1xxNvScJ6uB740VuWBCsZP+nhYkiR28YvFiZhnMq2sbMEDVCOSkocCvVoHzTjDYucFgdbLFVFKpK1RySlvcU7bq+FL2S4eQbSyl0ookFmI8FtB6GNwX3PuQ2opwY0biRFRyXPvdYrjEBQFxdQgWPjzmVNDEbGbYygBuPVokRyeVpUzC4rAGiaK+B0Wam8UujT/E6cPcaYOp2Mykf1P5bkGsIb/S5or6acesoq5DbxPMm11vnqDLDanbrhOmf5qSR8jpw7c/QtGeDb2bPklgPKhX+IWL0/adMV5Ncda+GeEzW5CoNbypKm9HhgG7EzF7Ui4cLUKbDQWJveooQqOQANGruButtmKviIA7U3NYAcKJbYGnOGgjvV88iJazCh7XD5hiZtVrOoscJ7anOCKODJlXkdh+35eebHJpY7gDSM3xJcLLA1kAQLWmMFcmve8SJG1ohToTqDkozhS/RkwjKJq0ZLH1E6osGFebLx11i5VNJ8jY6ZT80JgNeVfDzLdbb1Zq5z1msTiBQENruTxKaG0ANaS4Tni5uH1EFZKV+Lm+oDJKMIMWD1b2KRnv2lz/g8ZKINYRz/LNCWx9cAvBNP8F9FP7G9UqHU8pRLBAjP7uhP8hpJ6x/A7BprLjUkRFOZLSlQs4YF6I6kbfxKR9gE5TstJBIPdozn+7On0458vpu1J1GiZe3kfGh3OSV4EcHXfl4BvAq1nK864tIIhzF+BtEGBVsPgeENhwmKo5NJwefrhRCSUds9XHw0XnBkZp6DgD96IsmBjcAHM9Wd0c07gVCvDYkBSgBgjczcvLZ9yhooPDtPPOT3msRX3CKUICHO8oCF2Ezst7qzvegIjlbrsXQlX/PSXBn6wFAgahKM95KJUM8C6Mumv/qQctoHKphvvy3URVSn/3AEfjUkr58QEPChsL/GpCMkuRwYv9MCDGKvMmHYp3uS3OaHFpKNvRMA5OJTGyDLWnYGbfiFMFuhgGl2OvE0mwtW4uYRm8f1bHKCTn0dsnUbSJPNmHcM6SUJofU45eMZeH2FyduNOAhNQCAJYEvfwwVvbLCrap8Fp75U4jjHmisAHY6ZNxnjvYMLAAouI/gQuiRjW942M1V2BwZOASgg2UDbS14nIb2D9SLpnKCOqj2/z1TtCGw3PDPZIKDhr+8b1pjE36Z3TtjhNwu1KXSS8GFOW8tOKK+XdY8klOXolLEz7AQijmDUQAsN8fpRTjFl5s8Kqa2lh8MkkOAc08HoGOEXTsvhgifS/HJ0MhjpZ6BDEIrThJbehwXiIe4y+Y8e0s23wmKGRUka5JO7PipGQk2uv8Xr2Okjx2caVTdfpb++0FjHxTG9sIssVShQqGYHEWst7za/6/w5xIGvktbOlT+oB471AK/r1/pNTQgvI0pG6t1QjndXCXiKkdWl4YhaR3e74dAzJIhhcgoLW8b2z1uV9DvgZSLd4DOP/zFLTUy3efEPPLNIL/szbI+oaJuSwyIzgT8Ij1oU2SY1e9stcX4ErAJGBmVC2eLi8eakIdKeYUe1ZgqRhwpBGDB9sH0b5UV7GvbmrxwXxOMNndby71j4Q47MSw8tUkEcsi8gcxCbwSCCcF9eVMX1wupZgFG+llcVbJwfuTazLNzTWAeHAXyjhJDacisWVQ/EdZW9c2k7hok7sVt0pREdNisp0OKlPwkxquYM56cLOV0jI3msx9iQ0Vw3yIELNXEU+vi3sOSaAUJCUJf7BD6t2MMX0WY7BlbCkhnCF5Iaeh3aSGYaTdvf6+ww2h7bK1tuLR0oZMOekxdI14b+vUpbzEF+41a0FIYqWHciFkqFQsw04G2Kf2CFZ/evGH/Kox6P6fxmH0iVJ+S98XLP6HbuhOL3UjZY4D9Wf5CDmiJrN4DXU4K7+QFVe9uuhXDvLZSqJzz8o7yOQVrb3ZrbSdIQ1Xe46D6pu8r0t2B6ZEHNEg2o9rf/FF6QZDgy7uwOhYhnFjk5vId6Eu5DV2Ynm2UVpSsKiRUPzryO28gWXpVDle/iLlZGbY6oSr0dDurbpBeonFibLnqJ2odMlHUQKNOkXSP+GDs5YcaWMLYUO/hC6dKjB9zR+qm9BGrLLMabUlOa/HmAdjDWOMv3Z0cuydtPpDgxZ6OPQ7LvYglHnUeZmz+zE5u+g8avifGE+muXmYEZ8DE0/MsPi2wAmRYi+1ryJhP4z/LVMPQIkxGGCUc+2hzIXgEREpeuao4Cxk+VTaEaJ2XPpvcWlWotv7czPEizg5xLP0lbbj/4ybyGzPxSoZAdsgomuH2KBGAzHj3He9iFjRTQkP0nXCCocr7YDG6jPrz/Rl+QgLiMrAbR1iCe9JYJcIy2PsTMBKMOZ4HJKcUQty5uFrk/ftfnLlKF05ocXPMqSoM5kZy/911bllR7Bhm8c6NTP14uRO2Ma5M7OqSqL32mBaV54uHtJU2bjOKlVZzs/wv9rluT68qImrvrNdBye1N5FTTY/OezpXUT0QdJz8k383g4+ZQ6GaKDo3vzARONIkX0zcmQgmH+w0iV0D7cVzccWmjZRnjZJv4o8NqQ8dF7a+Da/OOYDR55MEySMo0l7R2RRiHhusxl22GhccGJ+lZw54D1LGnl2Rz+NVODcgrXIGAS4EabQHNpxxstAQlSyJ6VmoDqkA2r84kSYOFkqx7Epwq0y15Fchhrunr87zJqJW802dNFU/T0G2Y7byh3cBfQBzZJIy5UktefTeH67r5EHuEfYJqbYmze20qX5kwiYM7QChIbl0H80VP0CKoLESFf1ou2cCq0oJWG780LadxL/4oIaKhVtM56lpXFAKypn3PWbka8xfBWt/nmgQ/kk/aIgQsnYu8KGAiltDZkoyKWqUgH1bArexKbKAzCgFwIm7CZJT6uPAQ8YnEbWL2hmQyXZtyLTkLDkGaX0jc8smxr4OiEfanLIIQzUbxrPM5YgU4x4vyth8hczuCI5uvS4=
`pragma protect end_data_block
`pragma protect digest_block
d752080efd2bd1780ee84ed623737961d0ade565183f4e88c50e92d9a132cead
`pragma protect end_digest_block
`pragma protect end_protected
