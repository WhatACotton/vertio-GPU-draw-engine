`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
H7ohnFS4AeKgtmU4uDWKp8qPf5KROeoHb5aascG4IsXPdT34cxlVe2TSCaWXun7x1itJgHYtLw/k/JFWB8uPxnxJl3aqPJ7Wr7YZ64IiABVILJnTBsPqBHch3uYNFtWbFxbrmti6jx/mmQnjkD0EV6JFdiDXuIKWGMYiw+wMU84TOm8wwUIwzf1jTETzzxpcxBOfACCpL7a0q0LcPQzFEXClrxQUU8kvIKpEieD4G7PqLy6rspTaSame8oWQrt+yTMMeM9nR1Fc3IE/LbzfQ5CkAxNth2EyNV84bNXrU1dFbmucgitxq12SZq0LnMne5rjDwBkJ5EPoh2gO52rDUrPNtVvDTf/F8Dii7bqJ3Aly15cNboGbpXhbIRFXFQqmLWTWIJUM1SXyLPzeUGzjbY4jY1UU/C+fM/NUp7jmXIR8pi9IvBq5YDnfVlBG5g8F6qLswP3SnfqBRBym8PnzudEBJPKOHizXYvhuR1LKmxLZV+A201EWdQCxBuJd8JxTGUmhSsSFY3dRfS7NQDxlD1c8F4p453zqSAe3X98fuq6Y+LL+peO3iPApHPrLp9gywnUofdxdIAmHNtOq4RFFg9ED6EgezVQnLjfei69GnNhqdIl+/k/ip4IRa4Vtbg21XOtpZwcO4gQoAZTMdGGcgq/KfjxXGd3d/v0Ifg/BOToAYkcWnPX+xhv4RNMUXKJuasEfffh5uC0RGc8eBk75TEu5U/GUTmB7ZP6HLwx+o8P1f0XbneDAcsAlhAYaLdv6iK+Z3tRkTuDhNSMfhBMkgUPG/RsH2mzgfwB/wFhAmHeaTdxnzMrPzQxre5Eiaw+s7JJq7SO35sZrg5fQnuDq5+JUCA1tOtJHgBbZTD4BF1q5OvREmYF8Vzejom1Y5ZAFxUkaOnNcQXkThJFWvpv7jMdeUcIhdE4MerEKYr4iqP5St0gYlbduaF3nESR/S9de+uiTO0hO7n3et69w4u2RzdEyCO7Zl5JgILrLCnptMT7ojFWMXqJsKda45YErtuK63KEU+iX1Tw4pfc4p1K0vRENuSpL1Ak8czBNDgYQj9dz/0vYJCSZDtkJr4B7cUxj1Bcr879MhRCkCEVI1gz19BzjeIgKMPD2kXhATJjBJiMGOBrxEeto2TNfHeLn1zMJeo2SaGHNBMIRinqqLcxp79lUFoMUb5hucsd3bWTTOXnFknl/o+xO5kJUvQqe4t7UMkhWguvPibES67dfROXVjnyl3pzNVHlDow8ITe0bbcsfKK44kkCGnCc4031glA9jkSIWpA0RcJ2gwzD8nK473avDzwIhW4q/Z8pOFI7a+fH7E5lUgFAQI/Ws+SZJ6uefyKSmhLKqmayj15cwkHtcbUwJchGfMWnuqCxeXjZrj1YdlNwj6pn/bS9w6ed9JVzHiAJd1CP8d3Y46GM0nE65HmdNlVxX8fs9zHQt0t8z5LuRLZbIFuqDfdds10FCOvB8Lti5uNydKsjWtiwyfSMy0uI3rhkuFTRRljvOSlCxPkrCARpY3TCkolCgKzF+lZIToqwdGSGlilC5X/30kIv1hEdhmXYjlHnple7O+HiCrDE/zdeNfj7hChi5G2swT75HNMXs1X+QekuwCCv1n3LSpaLSwSVw6XlXRbhmFZdA34fDu0Erkb0HbzF0MDcT5f272PfWJGHwvb2NdHlL4cJuAc7zTXCKE4T/VW+qf80wothyrJfZGQoXki5RjH1iHnWsOxHUDfZhQ/TvOJw0OT1xUCcec2RYJImv8zw2mkEpzsvFsOterNn3GsY/XVbI+anPBMskHNccilaGVTrbYVvy6HLF5OM8RCY1vswpp9oEJDR0PspaqngagfbZmKewFcWc3fJZKOZmdfAES1PyZJt0SqREfc6aztsbqO3ZVu4vwD7hJ4jA+ru//zACikaqDDRV42hN9Slmo+wzuQ7bvpoS9InN41U2SlGWyS9/XJLiS+Xy4J6g8y4LI2UpNTtEYS/CGTGvZYSx5zEyU7LQ8BzScRTIqpC8/QRAuF3XbKfXU/E0JrT8E/ftKEvWevJtx1CcNHL+VcFuS2M0Ma/mvPRix0wUxseO8fROicvJ5Z3/fy/nEitOu934Amt+m4Nvkveix+PdBfpTJaGd1gP6qhIFMy9QIn8T7kgl3i4U3rL1SgOIvpEcX94IDGjmjsMtTvjayiIkz90MO4+k8x7KQepFoRPDw8IyqN7GDFVgLlioE8W0uy38fz9CbxlFNXLJ9qGR/Op1iLhttCsTUIw7Q08pa4kfUztOUqv+hdQXHZ4ATCc/6AUV+HR5okCOfJHeA2O3F0HIEc2HFiW4+ny7qF8HJKBycAEoclQObiTjIwhXV1MxZUHQFWcZkQ+/cgMmscwllzvGEUvang+XgEGMtEV3ExbKMQ8te3Xr9gRl8E2Ymyc9d7ACefzrZ3nnRagDe5TnfjOh4Ene0D62eUaO7qrMP8sW4OtdwzjISwEO9zCBfy0O8aa0pkyXbC4Hm1UiDuboiXX8j5nTN0YZjKnNxto7BoODAI37QqvMBjFpZBFWgXfJwDwwbJzxo5Q7iwdGSxrucKrhQRYfUtwv70KFVKAqbH9F+r1GZJj080v1EdmKMpxniO0nhhLttLyFQVfNrdhejd9/5F8ldCOtws/Howb/zwnxBZYG9Q9n/0njR1ztaVreP7t/q/3UpBCGMGra5UURUq47DzrbEgaH5jpyuUopXh0TRBaZDi5e/5XQ+q3+utBlGzCMDJt6je5O0OCedRqzV0wBECC24F0VEM/0o6eG0vAURPg4/H0sljEq8g8vMOdyrDFJyhQqOgdl37QtnHckbdfPw1aYs6Ch/2DZbj/GYYqNDw17EdIc6wJJlKCPFnFILIZIdx4P2Lz/yAPkFiwUv6Bt3nTI5bXBoOML+oFnY76hdK8lIZoYfduuw24X7HO5StUymapmT54gZ1gq7gbqF1oBLfW+/BKOfK2C3Q0ps0ua0u/dqk4+JR4xuJ81Zh6Tplp9ZI40Ni2A6wMw+DC5F08ghmhxdlBRLqcY2C8l1x37NN+ixzyY9Gct2P6pqAKeiTckwYFULn1Gp4XKdpHpDWuyX3Z4K1hrIGpw1BBbPPE2a6AzocDcwZhr6B/SKTA9j0DSosPfj2d9f7slw4/0d0xSWZmgAARGlUg+dOqf1C9bV3yI+cK6f4IOLhMuCY1x9LDli7D4JVMixgq5yQ8eF/d9vUT88q4VFWfqp3qc9tbjXXScyXPbahVHZYkYqFAXsfecOLw9NUfsTcIGahR2f7yVHpyyoF3vNLIvn4YUSRQRNeNh5b0cbc+wrfprI6yVpcRNEveBePqOUd2Rpr+IoXqjU5IvZ7BeteBD269IUdKek6IhgmrTiUsoEcKWGIwPBEpfmye2Sus0Cw32k/iZ9+stdlwGM4f4WYTctvV3CiNNJ2wWJwpODk4SWxmJZVP/kZdbladRwNPkM69xipb4/wa4bd7FBuXwvmgcHbglP6YAUi3Jb4wt/djOVyxv2ydIuU6NJ8NwKP7AyUrtAeiqVi0u5YyoYr3d8SiccoCf/L/fXQEIToV7/6GpbBxBD7m6+w+vh9NDSDwkX+2C7cKWa2ybJ3c0nWrAROhSCo0rPVBZUMeONfJ8Qoni3XrE2cVvL86dbZSwPvUY7ZpB+vN4u/rnLT0mUzy8iIsMsNNL0X8rTK65j8dEY9cTDwzNAtFtP7melHvItX2sinpRno0zG4qWewuueL+nPifk95quoBNqoJ/bEAlG/bVbuIrNClTJbhQsLglTzZ3vnORLK91+p/7UhplvR7UKIvcoNhpfvZxYEkLaif8BOhdEfs/ZzafQTFa4RRAFR6eNFbAFpEbe8Cb3H7A7q/lIxfFKZijC8hpNlc8X8Nb35uTxh3zPf6a4QxhqhW/DfiNgEK3MfGrsUKbZkzCLVPO4NvwK2YBGpWvCauspRiPO8jP9oD//OdgTObd94EWtAtCcFGgs6IrtKZRa0Ztio96Rm6njUy4Ki6Rnmc1e5uOU/PLK9BXU4vVr/d6+ciRkGg+4aY0WYqCaaoupZ5Ex1s8lbFeMaJD5gunidJTn3aW34z3kq3kMGAWhwYkIw0l5t+RkDHp2uAmH6rbOt2g6hyOeB2poVoPmf65f3FAjWnPiSiypujLZrdyv8kkvDV9hpaurvHIiEoYBkbRBmaTa+JpKR50F3S649CWNwz0HPZ0Mir84LCyOMjQXEB/CMDhTcsKrspR61kaVgiZ3WRfNoR+ALNNDEQAAgp9AzxiTiqQp64Rwygw1emNa/CEum+ZOihAIqveM4/AIJWyQw9V1j4Dzd8db8ZIbCtSJILGzucZD2rEH2wLUpmQ/M/v7HimjIth3AdoG+zTdxhFZhl2hT5CqfGbxqkafaLDrDA78+lqB6IoBiw9Mh2pYVSO6k3Ul3vZ3+YylDpYWc9G0fiJ2XXyEu0mPHXVrBBpIip/N7RdjcEoALljTH9dWXDuGD1qRYNfaTdgODLcT8KDuF7qDUqehFR+KbS0OjqEBolLNCOJvQuu371jUzBbV5snsfSbzg84qAKlFiSUUVbh+KQ2ee2UULph3JSJZNVgDldR4NlO5nPQF/ccsUFJ3kHcy+mKr9H7HUBnf6WL/kxJMysOHD9otIMBMoyNJ+S21SHDNg8yDQ/N9F3nAaBU2br4aFbrHYxjvaZzuXNzuCVH+ta2VcuqxlJRQEMwnajLS4xO9w+Xy43zQljKRBgkfefzYJlBA6JZoyXyg2VUzisXDmUQCbinjVZi4I2+hRjWyRGmw7fZPLHL0xtHUPxQywIXDvXEsbg6vTpx5yC3w4XsP3YK00Yfuc8bnB3LZDBdmRkHJZofeJSRHr1JcnKF0CTNGHD/5JFUs2zBikKkYJy4cGAcgyPHcDbXNtfsFdY31R5aff/4IvzqS4zbUDg5BGxkrp1dcI/udd9V+xBabIIZp19/glkFi0GFJkyaqb47/XgpbSGyOoAikhMUK3jCOkBbR0KWDrHbm/qrqh9vNJQ4h5d0SgPW4/LCysYDkJDxKd8w1a4lkJUxuJfvfQApmpovea0hyxhLFWJLsvsWG+tFuQM4czw1u43BWKRrzaWuY3t/VhPHudVBmab1WqRwA7w9cWacM9vFeulkvpsk1OSdzhJjQpV6xCmFLmAZYJ0jrGT7oRRW9HE49Z0JUmGjFm9Am0HUwUyHTiqSeGwtEhajd57mKOWU+dHkHW1ilem5XWszDYD8nKlQU0h0Uw4pOBGwQx3Gb7yNbPlbF6hfLvoqJIb7dfhYupE07F/thXPLfoMc/vc9FITBAKxD2UdXrOwL5of002AE+nHgZ+Kgm2o7id7YpDyy+EVLrBUS6F51y1AXeV0e/PZLBPoTtipke2fdKuyVSyrrsPmOgj+VmrBShmKqh1wHrnQgmDrkUHAfiv6mcDaFvJmeC7zKLpF3LNbN1CtL6zSzJPUz9XJGL0U2TvGaUMTDB7LuK9ohUdeknf39pjs5kfvSx7T+ITnIEcM2EX3cI3+o2yWeVsRkmvq5PyVZPjyhBeY56LDt8jan5SM81SPiJF9hIb/dkz2AFLOCBVAcrFOFqGaUHgomR1Cp9ACr1MHW2tCSXqPn+NzYtG04Ze4cNldZGdw05Dga2HZgLgrwzFlY62eqzxI1MuYeFRVGUTdwciJVc90ys5nFDAcleg67/FXYfNY/Oq7X6eQkRAa4J0vTzkFMi4u3cYAo8NDWV5hnxXrRC0nRLv/LJ1cvaDJSQIAZUgMVpSzj7RDu0mW1TyA1fLTf7Q/lDnJOgSznOnT56Q8Kadb0ex9t2Yrfdyp6hpp/wAZdYET+QUWx4OsgNDiWoFTg7rF/ohd1SPx9xVdLqx0XApUOScQ92G5Y6eB8qUQhHRMVw9Bi+3LDN/buT1V7oCpQvRgg/V6qLMZd3BQVX79LFORSUNSRnChtu8ExSt/yCCn2Go4cmvws7GzWJw59VCPgd6H14I6BKcmW7b3RTRVkRlbbHMKiQa7bxLiBO4XKCqZc6Ot9W2lcqEXxtIt/mZT0tDVjFhucRbVyp4aeOX2p/jtjfM/bPsgoOurpc+DNyiTALUIh9vivNQFhnGvKSZi4WynxUUmQBJRvRY0YwKByeBDZddSnTSTnTz4aJWam02tZjpjTCMDzINhSQIfGDmCXPEPeUoknIR9wESn32X3/EYIcpPXLS0NpS6lyZbEdFwv1r9VP2o1wDdWSX0nUmrHwHKuMhNi90RyFBBpVPWw83ba51BLGek6KHRCiDzb1ZVezsQTSnSukc4tAhp9RmIqf1toEQNhAha4SNaF21NhEdXrIumg4BCtTeKyjtQL0kB0jmb3MWgBLyi6FVFe6OrJTeRVrTOcY/oqoz6hXdTsU4wdHUMH0Yx0Y04aLeGwZcP8t2NnL3w/33hQYBc2U+awvDa429b4HVjC+iKyWs8eSeJe9Nx3N2TAj8J9OMEu61ZbX+lsMcCg1cXOdoK+PBjt7sPzwswxErUpBwRF9fzNRHnSGX66sUMEcUxPvSK6B+fqZqet8qWYfSzoHOngE81Z56Rypg9oN7zF6Fhe7zFCgU7TwrNTckTOomKeM5guBe/WlCBRokpbqTQzbl7kIBN3XIaVp0fPBLXVl28avcI1KEFf/TTTMl0M+sSudD5BWVaLwjum8vgXsF+5RU1GGvBBnUb75W9w5ZwB2sGhdSGpo6hUPT0eh86bsEJu6Tf+ocbNbsSrO/acZnMka1tZtgOTsd9+gbQ+1pKuIAtyMOIpXorV0iHblLy5I8nVId+CtNpSzxsj6OqfZd6JXakRx7tr9rq9LNzAwKJtb24xrfkWUOwkVQ3dHlLqosxq7mKnBdKiT2jLqYrqK+Ea4HCkOrTl9QHs6J9/pNtOvqW+ix6vJZzklGdCvGO+CsbL5XsVKv6GH/KXib3bd8QqCmKrbgH/L+25sbrbwaFZOFQRsYSaq9lSqo2cPUQfilp00CFAfRvt4NU6BBp1XTmwXQ2sTfS0rk7vaxpvxBLJodHacRUGJrL4R+Erpl8+2o/zSxLqO/RpL17IAHhybjeKDdCnZ6xMbXPCi0gS1uzI7T7RHsA34VasxsdBcAtytK/LBQJzBbaolVF3e6Kvc9eF7vF7HVbLi3fdI1mXiMwoeXkaWNIW4nhiFzIkA0OO+LG7MnjQI9XtCfCzymWKPxRiYIV8aqvn1OeIAQ1RL8b1ZTc6mwGEytkClY5Byl9NOTJqPfnuPB1Y+Q4JJE3ddX/LVNgnI/6cBT5MFhTgOtRzhrbiMwNeCb6OV1GeHHWgu/7+cxBW3GqTSSHqljthMCl4mJ4QCPtUZCcl8g7hfaSKbbG9Y3JTaDJ4jO5K4hzCXrgViRoQJkHIK9f4kcbP9n1epVKHX2keVso+dM93A+iyJtps4ABTwmLOnBAOlJl+HuGLSWEYr0Yj9iHrwyYeP2w+lCiRVUOUdWKI19cjCZIRjTsx9PvZpTkTS7nwm+17GrmC9x1MNmYSm6+738tmVx7W3AAvnVTW+fkPnvj5M9m1S5SQnHf7D3tJ8KUlWjiVf07i8tt4mYMM4+/PPosYhz/LCTRNtCiDxDjWu1MzumjF6cCrLSMB8QT77CKKBGlF04QPr3b6jFXd1RgqIpZL0ldlHbTUIaDOHx1MPs72Ervq2vHQoOyuoJSsiLmWxH71FlAlRJvZlGT/MtP6A3afMOdufBQDMZc3P3FicSAQ4I6KMS/2IZxkp7qfq2o4oZ+qgsAshVxciIHe/ex67Le29rsPxjsgkcDa7izPUkUFWMzEgduaBX6QfB+mCcUa7ITKfcvpg+Lw8817wX3OhymkKxRLfwDXo/2FYV/d3l5rMNAe7Njg0OZJs+j8VokXPbJeW6+DAl8izTvXWNiLoIXXRuR9YQmEgsbtZ7SEMAt4CnK7NrgrZgdyk05mYSQQjI6oNy5Z7c9g9JEpG+TNAt08HluvYUT7FNiJXnW3FDsPoxDsc7MVeSbDl8R5kWg5w5FhNc+kbi9LvqBf4HsJeUn95mnRg/iRObSxsyEcqYTcTEVcRdBtF8EW8FaF7WsBgImZKP34U+BrbBv95zmJRf2xlokGU/q1IseAiVvzLWKuLq4woNVjZdp0+hE/mz1AiqALZpmLyb6hEPHDpWRsXv55lpo+k/VUxAa9VuJqvlH6PhzTvkZhZKISjEBE/e9SpUZnmNtJPlcQJScB8trfrf8VSk03Z2yJDjVk89kdzIonp1wcY2dkTrH4lEOFjihyAPLIgaphIuRfmz2uxTC37vU9YbmQvTvnp4HFHm0eytS7zFDuLz/vUJfSoWCuuU7iqFNwR4G/tLFdft5/e8Y95Auj5dOc1ldZjuQd61I5SzUNKq2CC/jce7qlJ6nr67iWmUnsqw1X2gwtFDyZE6ZFvfuljUJVKLPgq21Evbx2AceEQ3RV393dpxyEKFexQ90ZxJpBWqbGQ/wo9JCWjY3pZRvf/5Ce35C7SsY/bTQL1FJD7d6f+ce64hwEw85CDUUIvhHtSm9EQba2o6jLOnTxG7OZw7Uo9tsEKf067FWG4qOi7bLKCK+3NvurKu9a847LO3wIWNlI45Im/8pAU+rgyhklS6HJaMYFoo0VgGYpmBSIYLP3tVxPiE7jwtoPbTzyRpXEHmtyZCRbrGRVhpdJyoY8LgmbGq5BJoAtsdBgRcVsByOOBAQlFFpbZmV4sX3ilWlIYIdIMQLsFX2T7m8691CUyzoLWF3z/Q6NVUXdzMMA1duM2ieaieboONNqxHCa1MhXipIqTkqO5qBRIDCpqiitnVuYZ9MZ5v3E1/gJPmPFJU2ASR9rAWWA2u8/JS/IbA4YoG3o9Y5GiySAy7l7HDoyWfBSAGKBP/CgtIzsEx7/YGfQopsRhG37vshZo7M650DxJBDChuZGKDZXHqvSg6QzSiq+5Bp79sS42qqYseAX6gq4EQbiTjGqvtvKwC23OaRQr9ReAbTiBlnf5YOUoqLbGMVFQIagb0wllCOiALfUBckiU80vR3zkQNwbYsalOvrQw3w6+23WLWXfU3S/kh8rj6lZpvsJ8nRoUbNNiXjY84VeGQdPKlFVxV3bFg3e6c08DNpWCmiY2+BL1UKpP9aGkEB+tbdhwEj12QdklI+FjSX5YNdCg/Yigk59MOTSSJs/q+alOBa75CFcUPkLGfxvETqDzvf90uDXXb8L2tDqaAGV+gOjlaBDGZVjDd2Zcycyw7KCxR5VtO/YlaXKErz8nFkwBS2nrM811kb5pqFE3MTuYNU+TbfcxiLmjlS8BX10003K6vAKANHPTamJ2KLLqsGTm8RQ3d+CmLZRB011hHdPG6yvbHGNPhQ9sB4wHrbaVCZJTOFWC+0ust9+8bx5nnDoUwyRYZCqxoUrPDzyVPatrk+uQHT8TZZ/H5nga8jxQLXwWRjxThE3NtDWKqVPzMmXAU9QhwDRM9/Q1FRhQTgNimk/N9p/doQSHBYoOzsaulBUpXOe6NsJwBvZ8FM1JHCe/H70PWDIs0DCzVaaFjMTuVshb/bfKVED9Fj+gH9fRaewOHI1aBPXq5PeF8+Q0ratbjzyRNc0/SqZkCe4cncTTvcg47jXnZTdSajGa17gqSZD2LZY+Xh/Go3ApA0n6BDVMcb1wQcOJJHGvJLl9lbUb+AoSLU6Papxn8rrkJrnUJHYzUMjQ85PgBtert0pkhmlZ5aWTpbTcQgPSmovdHE+bmxwX9EtAlWQM0EOZIUzgIJ/PqRugTj2pgouc5koJQprb58a13AXtRNWSWp6z9xw5kxH0PEUfKyGWT09fEKuk/EPhMgJoNaJ/lsCQmyqXHlrSRUuoEsA39brL6nyDNujd2zmmbodyHH3e5z+xQzgmS5Oavw4U0CkQIakgr2+afNjEN1balRCKiy83TOzn2yklOU3M/0PQGFvb1JJJrMIfPY8WUtsmpPPejX0bf0WDpe5X5AoaGjDZFtBddYA6F6IL9w0dxbT3ejwEVdccp9iiUfjN0QnwmkUJRysDt4OvUvhHUpkXJpVBeR5rx1cWpm1NYFPCx3JZFW/LsAtdKbuSmcNyFnlCK9pOlAm6hvDPvax6O9NYaQKBJLhxG1lPx3iWsZ1yLFjD0xkV3U1mZBaQhjxrhvtrBHpRWaPfMZqCMiYSLEqrZIywgj8GsiL18KVXbK9hN9sHuAuom480aN4TCQKZTVJdR8jeYyRQ4jLl5k3B1IWq3f9Ws+BYh4VZ5Fh9iNlJwCJ0CV/y3nsGYVpaIIK21Iya60z5PtzaOGeTQk2obsEOBdBjzb/EPpHgDn8BhQIMkB/O/pW0Zcse96lFBnzBuoXqwjJbdmeqK9vkxN0c1uh44vuBdYfFYzc4QKU9NZvOB7yIDnPBh0AtdI9qHJiLX+OrE4o9/3XGwlcG8eip+gNDicPsBjB7L0AIJsDVAhJaH+yU+s5ZSLhnRu38zsyXBjvX2cUKpdKJbXf6CXuZapAVZjK43XviU+NFNadeDjkC865z4zn7Q9rtKg1bTW0uUTnGz8QgCtgk1BuaJNjCvyUswYEui++B7j7YF2SYfBQHS1A4VfstK4dYTns3vqGUl28IqjOelKaNvsu7c75iCYP3/8Y8N1QeyKBhbWIM2J0iisKSZlcn7Wr5qvgz14QiADXgwK508fwRgzRLq/UQ8JRHKsAeYwWGN5qkkDuEELTr7Jr9r5C3QPMLOkR5XOmyye+KG4T28XzEogrVjM5e161lga7BagG5phvl4cpVxA5GJEuZcodK7aOzEye40h1/UtIj1Nja7W0a8bH343fX3BdPkO3Kktr+C1VGdQIAH+pzQNCavz+OHur3T7kkKdkBqNqx2uIi/AlRzHH6l2arVrfUU7M7vJJqwGIJd+MdtdKpTijsunzNgszKbzdGeEph1xBbHXOStb2WRe7ZySJSuaSGMZSNUm/ailrEz9AHJWNCjYbKoOGEVZT8p8bMb+C/0r59W+B95rpRr1BO2KbrhbbE+DXt1HtGu9yKoNagApz0HpA34W5MpcUJwkaHueN9L2Iw8C9Ds8DoXpFsLVrDrtuxJjO017wrw8lbZUOxo28T47/nw2lQ20c3cAXINf1RRARz1rvA4vFgLoxJ057VibIXNRU/bnWJ+BPRM/b46hQSlHUMoy8ftvBTJVivxlUa3ZjxjiUqKHeYVlDTm5Xg61RiCgWulljnQNbivyUFI0AujrmET4kf70bbflhvnBxdGCAsrQimpInvuaOOA6UIjZsFnn4bFCQDcuCcQgcyJN8ERNNWRsNo1Tzfi1TQEbd93U9NzPJIASE6IRcTm4C7lbbMVl81+ETqyjGzsIlx2Cr6Nb/Tj/7eGKNCGMwNQL4KnayYhr2+FNoOtFl6sPkauPQfA/r8T3GOrkUGmFm9fPbJmNgFRmhZECPj1CurdrXsawMl7D/L1eG73/jasdl3Rd4/I3IxEvc15b8pqehSbjgKSUMWsJQ0lcIJ0eui7gO7GLZETJ9AlUwkcC59utL1arouetPFm4IMvLN8WPXLSQPlDl8NnPbFLg71uklLsJw5Epx2QCYI7hl4O5TSyUf0ZVhPkMPHoM1lHLKQe8ZlbsOdk2r2BSvDQ4hQwugSEDdZqFUG+pZJ6aDxjutLQmBCD+d64Bzyetcx1kiHiwSIJqmgO9xZX3m0Na/HhS/w6ooSDxtSwUWXOwu1iq1S3GTDM8CTZHJzcPxaAy7RwrYLXi/WZtbGEAJ9pxA3xQr0ntekAzPbF5llHmGEmvSPa2Wel0y7ayEewqp99rM7RrDlfxaBtsdObrurzXyFHFO2dEEWHC3SC7kcjXOD3EBU9lW8BoRx3pAZ8mMYAkNEGYuNLqw8KwHw/+MOEbLxJhavZW5qqJg48pMWerKdmFC4wLmujIdhKQaYqXhoWqxA+dy9dB1C42EjEv8KzltVOU+aXdVvJUkMtePkXdYviZS2J8jo9RBDsrybEXMyDB6ME21jYBJNylZ4OQg55yY0T9YvC8O2ucECxY0uDSG1jAlmuurSDPGPNPSMosRx5sAZGxgQfNoVpnpqJsCO+9hYxpky9TG2Ew/oN0/MZ6rJCTxVoDPrwjS+c2tjqU0qKoKyZ8slwCXE3M7BkqDHyToIsgiPoAQAc24Hz1L+uAgk6h6ljewHLu7xLNBFxxHO4wUPN4o13P7+8TiZr7q4MS+2Or++8UhUS/UkmKS/WHPJ+BThou3lJCqVTkbvc7EUIEdQ6LDk1V7fsvyix+JhJgpbkRYXJEwb1+kY/HXT1GO8lgFpq9rSxuh7b5Lya7Y6UecNE9ku3cpo0cKGGv2WavKCkVrUNNNEp+IvGxE8J4igBI8H6cvaRJvUjx4lI6mf6a0tT2iym7g2Z0wy3fOEpUUB7ha9NPtGi6X1XbVXPXVBqYPVtVoRQSTHachLt767vNPFeFlVlBNUGTZYSgprEmcB1meSfTvQVQmj0HK2/narAPHVGixJQJnY7UVAAaWW7GzmN5gS3s5co+qLotHvZwlLpM0FhZHlT7ngZvtXMtazaLmL2ovShNMTOb/FScKRLHeCDSRuYqa6pAGvdey9QA/xw5w83if+AvMxWjxgEQFdu+Dd3pklp7E3xlSih82eKbeImpWjAJ1efHMbAuIfDbvAt53VfbJMIoo6HruN9R01aDZMmDGZ1xFbQU5dTtH65yLout5MDQSBEuyVBQyN6mjt9nWrk4NnX8fxdd1Lr/5vSdNvom0yI2O2zipskyq3/oBhSIWyt0tRN/M/cPsTdmK1xuGQ/qQZZKKIBXhjUH0sI9lrageqhwXD1Fe+xmPSr2v3Ilfvozik7kfOTNFghETgTYT4J/Me2VlmiWdQiU61Cg8ULkTyki1AMscRHBLGr8U64NVgngFF7Ig9qHa6r99K7RcNv+uxY4TpnmwheF1AkUxY2tCqNP7Skr8h3Z2dltwZ0UtZXI9iBHxvLT+cWZOi/WpJix/1YMSvKndKIbyYlO+wWlxqOe+c8GEcB+Inde0h6PgbMAlkC7cRCO8mC+1OGKW06K2pzUeigejRuvNY2Wjbk8Koa3M0yRHPqHHMdXYkjlqXSTtq3sh1Cn2X0LhEi1ZD1sD79oByxUMZL6Qkh9xv/SQJs7MNF8noMM5PH6AQvATrOc4IY9ke6u7Aks2e1S00Q7vVo5l2RJaA1GAxnWYUsQPzD/CxpLsNB209sS2bT3QgFYkUtyVu/N4HVl9olBMs1Q3ITiZwFvPjITAmAy3VAx6SgyXuJIAJ8BurNB88eLOEQtGW9jfE0D8Hpy1aOrf6KIyAlHl0/G7SDl2+AMwcDFXgD0TA9+Hl3mSKuV0a7yygfDIwxUHESYm+M5kBqN00zOnsbxItM+wErnujeNnaW6ZLNazABZrWRni1Crdgb3KghbjdUaAQ0GhgODGNZDPtQcNS8IPkZKSsOl8bO4+bY4rpE38crMV3NQfx8YdxUnfrMBuxUhCLsAKNspZqn6YdZRuhKILiHx0hPZbyaeyYp0jj6UDc9mE+Mu8YGwrYBD+DsF1kRQqzdeZ1YhKM4tH7Rq7sW4ZnzQ3jbHfKE3RFqiFCpYg05Iklp0VVb7CqS3t0ZsUtoDJ1t8y26f05IkzHEv4GCqDXJJRmRkDI2qOtPs1vMouWM60jy1f6oS+k3OJb8t8Y4FYz3LJr9z8ebTatBiCRn53S81cNwBkU7z8c3pkKc97MW/G+Fvoq2cYsSCmG/u4zAdugTFeqLoIMkE4u9w8cGPJeHhsr8kb/P06sCdqWR4rAj2dmmXrRy9beT8ZukkRQbiWdMWphhxILsifVmvfL70fWpO5kvd8beUDOM2txEbFkNFFXoncK2J0aHxCvukdLaR5di9iRENZPjAFy/DAM7axN6sjeieufp+7i3tZsCErtkjcINF4SIT2uHBbDojlQiUy2ky1KeyMBM05Y++qIVJbf8PaDd9cb5HJulsJdRMyfmNthcVztfSux1DP1qbTdPqk81LHfnisU+u1/+/M2f/e5u6PFzsVE1363JmMpbhPZEtaGs71PH3KSCi6y9IreH7N8ei4zzZEOTihwsjaL7/ok2YjBc2jLp7s82r6Ngx7cvzgCPWaBaZmuG86SP6KGZw7BMT9XEQR3o/muC6Zs5DPGKGY3wPnQW7Y+B78KOy4mQK3q2gRjI9izFkTm+6raHoN22ra9H57FO0RMpm4qMKgQ/HSn2+dp3RR/lDDstuyc/4FM8BvnYyUAJWf4HzBIM8xVMaw4Ll7jkfLRDRL11S6aAuY7xTrePo=
`pragma protect end_data_block
`pragma protect digest_block
e5c5498f38c49e30de37d83fbd339c3557c50a4eed041b968a28fc7c01003d23
`pragma protect end_digest_block
`pragma protect end_protected
