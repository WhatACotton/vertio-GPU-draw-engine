`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
NLZOK3LL1xl9e7jU0GaVttXW0a6TWMuzxtTHuYtJEKIidZtofD5cgaqOX2oKQYWDYhWKTfyVYSpCa352aAhJNwOO4/t409+HQpaYILE1iuP5Jc2WqJE2eou+Ys/MMksZ/goR8TLPIzsZ9COm/e4vO9oVKDN3Jm9q9p075cMH58kFkMuezBcc+oXeNFSOc1jznpI91xkH5LEG5KtZGX+DFgUlkYpmqin+h9D8nSKhrN12dk9mzmEfTwTKicrmV/KWaVrqIMZhnkdbqANvoZeFYIhRJ8SiNRrsw43KSI3nYi/AASMtG5frBOZg4oB0juB5320GrH1nLy7hii+7RZPVfQUIdKL+pBECFGnSAOzhWvaP0SvXS73H4l1JVOBZwVCFsJ+ZDQuU9RIM8sanW2zZoxiJJcIab3tNod4efeHgGL/g5YSY6mIWNPx7yr3d/JOwkFpJI5CpEKIYWMk1dpc2VvXSaJPphM2S+a7RkQ7ymAIEMzUo45Au9dPHWuplrONo+7SA2fH0u3mDs8orhaaBGUFxRK/cTILcduQOFQJEqfjpX803C8wiUvfO94VccS2TkQk13FcAVDVWV4UmFQUVlsfq6FkE1UgtncUQsGc3/DOKypFnf5NzQm40jw/885ibIUxAi/HZ+WVFFd8u7Tc8ffZtIntNyAHEYsslsWR8Wx5glb1qpcclc6PxofJIOAoNYaWcWetFJH6yIzokpyu/bEst0aIFFdnn/7ytFPHjd6cVOLp+lRjEgPP+iLVZHLuUqwxqMAOEiDQmnmv5vspU1aKqUWaMbxrqNX2QdGJpcjXUj8S59WTSQvoA/Gbfkqre8LYg2nCo2c+99y07mO7PjZnZSUzjcWYDcVoYM/5Hftmkwkz1GGh3NDMhEswJf6UN+CQBx8LCG53H83k3CCW/Q5A1tRflCoWTlolAawIna5npKG7hzuCgSVM8Oc22hHuSA2SadvoC7nHcvZmPjq4imQnYJP/ztZEaW+wxjaUHJTAE5NypJGWpxorLdTamzZmISb01LyGD5YjZVhkLCQ5mM2j8Uzm9zbEX5EGIViHh+7ntBWAph2uZSh07ii2hR+s4phXy9XwiZFdOoGc6xueGImdM1qz9J6CDtj+dd0AWDLDOd60CoXnYWzdWyiUYkCYLp3ofsEI73ePILNyZuj3bigiAMpLJLBArPCLdl5bqrb+X5KLs6B/fHsaJ3yw6w2CsWoTphRXeOWeDbgv6YVo/VGXtiBd9u0/Sb0/X1NxSa+GE8aNV5scBdtCEAQzMFh79Ym9i5lrnAGT7u5BVLLBTZaeasAsBwkwAvwN/VXhwCUzshMbyEzgjE+xgZ3AVdPFI/ECPbqWZVu+I+Fhg/uXGFM75wTBawyT/LELAv5XW7EyQb8Zz0JDT2LFqXC25+komjKGKmUJlqCQOeVjF9bmjskO9T2QlW4T2MqrZvUOj6mESSUJ4kjpDZiJEBXwq3nnO8lMX9K5w5bqMslaWOYE32cqB9uS7hAdFQCV+HUVQ0EAu5dWCT6FvRtRMTVLDP8GsAIhBKWKawMjJ8vpoQTDGRY3xkqfW11n6PWXGSshlz2OzNn9RP25VOGLDEzqD9d7oDzyyPOwSYMZAWNYqamHB+sByq5ILbK8k2QVkRFpSBaPG7+9scjm1wRlRFRX6kwAM85wOQphm7AVu/BNE/nFga3/qYJfjspB+DgBaNPrwtm4u+yB+hUoc2Vm5l/0+v3MW3S50EaPCmhZP9IMFfAnhv+Q4lbwOAxp15BO6ZUgAg2M6z8KR22jwPPTT3P88CChpV7+LQMrGeVeDOFwlaH3J0cu7ETniqiyRJ7Wfy9P7QndFDlXvaKLYvZcxX3/LHHC74H7MJagq5izh5BNDrx+9zjwt+0XM+oezEf3wd6LBKtnGpOWUC64KQm6NN3fbPAuVUrmwhI0f7H3KgxpRl2sY7N0SZeu03mmrxfH5jIhOtJM7ZGcHltXL2gXcUuMwTFdnHyt9+itENqrJWv3Qec/RKyMdtxo01gGoJ3+s6Z3cB02l/6N3eQ0l79OTznOkbwTgsAjIyg72WstjW4w7i+s1c1rPphNBrxb9rfkRYXqv2CkHoAjcH2XtB924gmue7MmtP7ExifGWOLcDnfA9MenX3eWLFTY0XUWXG21S4BVMTnJfqGq3zT2dO8zlQ4SRiGLDU7u8gD4MK4R5oeYwgMPvr+t8E722hZuLoiKhWo0CFtFj2LpnAsok0WDLz5FW91m3Op9lKj0G6sY9YlKT0mIHDz27vPsYQVgsthhvhazFD2Sxl/QRaTk4hPLp0rHhZSGMaaoesPLPQCi1S8OryC7Q5tgCIcEa945uaVr57ZL+KNtlNGTicBs+41Ne5Edy806QuMWYFq9b72BHgepPDwcNMcnUVKfxdMa4Ay6YVoqYxEclQ7WW3/buxBlhaa7T4d+zDvsDcXjMm5KP4yKTbqE34jRVYCvwcozC3UVx6icUCUb59iZsiyfVDV32T8G2LQTjDI4Z6tg/NPqXWUo4xBJCJTthVMmqNLf7rku7JbLf3Lkkl6BXVxx7kdhbkv4qiSmc+vKSm3gE/0IQ02WNJsxC1x3UbNjxZTFB+5SwwvybVgqvvyav+wDWNdsHkMubl2F+MfonYg4HPs5rqFAd1Jq8oVmgzBP4fFxLN6/yztRcCwAe0+f6x1BYrbVUgVmNvOrhb3jMD8cJQ46PItxQ5zDWDyzRRbbsKE0M4inoBuhBdcsZNXOqQe83k03PZj9Q5kZC9KfXSPxU9jqbiNrPXxR++9vXD3hFNFdUewGbE3f/ica+WkRaNi0fRJ9gW0XT9j9sMejR9z1N8H6TcZj589TENa0TuKe4Bxd896Bn1acQbttzHi5Cbh3D57zBz6lbqsz6T5+YHHWXomZSNNk8KAAAETQ7QXDgWByBFgQDnPe5hSTVxL9fbbf614T9kF4ey1EzBg/6oJGu1I1bT91DC2D1Z9AvCeTe82LqD+C8tVxup4To3P6A7nZxezZKC8s/Ip9EON+/J/gRDXgN3XJXlgx+bh/ktQp71nDr3bpBfV5rnLDFUJFwPCzQ0M10P5uKf/o+KTSsgkfhrGXougTfdtQYQRfuEMFTExKrfKy54zv9ML+oMso1i6xpz2cbDYdRm/zt4wZTNFtZq7SEJQO7z2BTkbAAPUzWnXdq6ycHiP5KzDtzV4zJRcG63qkLm9ceg/wxNvc6wZLAOUPWUJRGcyD0b7/bmok48O32CJ1mkP/c3eBUXDq0rui9ARBE6c6FzNV73MVHJKEjdy7PI/zTIMicI7Wt93bbbYRhzLzKmB0cF7t3tSAG3Dbio3oDNjSxCptyw48PlbGlK0osuUY6wfYkRNTP3u3kO+lg6lsZu6eJOUJsP2h4ihc3phwGmjrzjs+Im0r1g6TIOkvXudOlxaEzSvKPj5PulXo2qLDubUuaJe1jRs8KO+0+nsIwjeRPQ3RHH5nTE6ewKf3L6BG1ktrqfEbYgNeJ3zmDMG5qI2oV+2S03CY5iECEj31wF2BjhycVNTjJA/pVks7PSRE6KA2Wu9v0d0MQLGQYuZiSzUj1UH5eldmxkt9jh7nAg4rk6F3epheWpmT/ruRvHSxQvbuvsAnE9u1JbeJtPmwqb77I8JJdwlRyAWkuzAf9Hf3vhcZ0rg/KrJz50euZy3IKWdBApWMaFzZb4rga+fXFU+PernWtkT/2gTWKTxMFZIHU0qh14eJd4Az9T42j9XIZTqXtlMLP0yf2lxqW6crwa8/XstMdWPvIO6uh2lvRzN+Xhikt/OGwtOKEwD+SQ6V1Vu6VfTpGHx/zHbt9ZqRN28IbK8lypYOb5qox+Kp+62ROtj022zab9/KYas3yqh9h/tuAu9auSFGngdO9eGc7ACpr6pjZU5HwsOMLSJ43g5UXmsVTiv39lclSlZWSW11eUVJi7kTiA8B19zJCU8LeEU7m23NnNh0Tr4Z6v/lkeQbVkiB7oZ7l0tTZtHpYt/6s8XW1v23MswlNv0FxC86BdHmCS7KhDvsfHjrWdB2ab6S1c89zxPQh8gah2Zc+nrwSTYavr0ChNia8woBzKNznNfyZB20TQ7Lq57FRobN25Hos9MNBIzzwyv1aKf9TkUJLXQI+a8kJT9jLHwlkWFwqk1nz+P+2gyYewZOlkSM2Pac8djrJj4am/rJFC4LXr8Mu1J78VGah+TPc6vSGuoFvhcs3H/aP9HOG3HVEB0/nisQejgeSRhuyoShy0HcgexOfmUkW/ONbE8D/UEMT7E3hYReK56gColAU0cIjpDgD9NGiYQGVm0paxNqyzbpNcZG39xSJV9xjprWiSnu+eMXw/VaKy6uOdaMJ3Sn7jXtRIZaNx3A0GFq5kzj+cQFLrQHKBx8WYBNbFq5DJ6FavxMswFPn+5P6lJdlTibpx3dJoIyn/nmdbZ0GUtal5kNN6T5SiGZPBMe5buCT98PgKB4hC6pUaEZGRPsuVVPhC6X9B0JLWxU3uXCY2Zkh2SCIlA66SfszGn6eE0uAFnJ8Gd5BlmivTAA8zqo8FylLR1Cqa3ITAJOJPkNGNhxf6cX7URnw7IkDw2WjecFKfjCLi2eadMUMDiys3PwzgiHNMyoFVYc9hjioZ0TdW0oDeB6/djnEfHasTaucLGIfZgTBKaEEuiztm/23L4B+3Zhxm9W/Icadm2Yb9Xfwr0kBOOm0hoSRwJZNMZ3TfSRKXHIPqZZfugwLzmgqOP1xEoxsQqXarH47pwkQByGYPL/LUpkYIC47XWqdEQg7p3fBMZMNt/L+jQEaGDN96DDHKkykXnMoN59jTYvzotCtYn1FOhgcHvESJG1LjUyX0Quii4DeEt/NkNCuYahJb32TtPJ9/e0L21u4hnC0mIcXbqv3vjGjgGF80srwpXZYLlFV1+TX4KN5/ZMhCQoO5t/Lj+NU+oe1E6m5r6Geq5n4XVZObIH86s3a3Ke8Qa5E2Gc5Uh99apL0TvU1AD8d3A7gV22LzC3nkxqSpslj2KbJu+zw1ePKjIb9h5gz5QnSM5D7TaaQg1eVWbdbjVyZM3lrjV3jrO+4nDPHVsSHv5Gf8GXm5tBlsM7ZtBTjo7TtimWJyhRcSi7J5/fdqnPBYy38CWojtJ0o9fw94r+n3Oic8Axes8KVUNKYN8w1Vg99U6lhwIkW/L4ewEK4kkmVJDcSalXtL1TvRY3zorSVKS1F0pdWvjJ2+LA0wKMDhGJFdhrwiBESwfIXD/phrgbFKH/DjcxwyS/X58V4XDGv9sSPDaUFPj5LEIlT94cZvTiuHR7PWWVNV/mfDA/vsroOiWlnDQgMBxL2V3pwLd/56bmIbPzYp6xxv7D/X8xLbnLd6boyfwTGctDgAI83csheSnI9lFmssOoN4X11f/UWm3yJ7dYJnUPGXev6n+R05KHdXNXygvv7fwFqHG3+dFbleTquPuuhFGQvzRQBZAfXYNtXZHEFJwxgrsN0wMQt4CAIDP1oh4HzckIlFhi55mlWB1YF1X3z7sYZpQ23t/1qJJFXmi5uY4ALEJrb/na319D2Gd/ec5bIzKhGq9GArWsmTtreQRGzJGlpZ1edcLmOqqC0chy5337/ETMu2W57ZCrF698/8Kk9q35vDu26aYRZcOOhpvy9zG49sFM+xf0g9+/Vv9Z+CMDDLxVNHUJpcWR4VOK4DL9J2rrcv29z5JTaEqRHtRfPBloD+5M0qlsSs98JmniDhqmE77AOa+Y8NtmkZPNEmdcWY1XMwmF6mYrdl+ohdOKiM+IQg58H/Z/sYo9ahQeCdTfC/MDa5FfVcq3XDMi9uezXNtJePvOlscJGUbvLDVLxiLKjB7G8byEw/vR6fG12TROCUch76d+L6kAyV9v2tf2/Yzv3kdLTqlnMN1XljrGG5bGnAwRXKitfEhoFQ4aCQMYD/TWOeaHMcRqZ2kijCy71d8vc5HookOXkoTNa9X/4ejInNwtOCo72Dcq/Z7gVRwnN+wXCin3gRuQwpLnqJyOmIRR4geT0DyYneUXiG03QigZXr3HiBlI8n0iYxxGpYw5I8+4RspfyXAHbm1kUvPd23bGJvIo4c/nAM9eSTYrmQo202J2pjyP6AvVO63g+QmWr2is1svSHTQNNbZM23jwNhhiYqsBkr3YCcgBCKnArqWM/BsI3nLylMHmCMWAKTU7YHbezftfCEclwbsQDquHV7sAHTulDkNsDHnx6xArwHSHDUXyhWJfeK1pW8Ho7LcBOy5uxiWJTb+aSWQYNNrouOXZbA3IJWUFiiHJzLxDQmcTNfGryfEca1a8xUnwcn/2NGl3ejGUPrscBDh/RFaMPi8QPSCF8jREEQF7h1Io8J8yO2UZyF8ZqQPVmMl/cuXKdH9XaD9P1aW+7gvsqZUYQLrJkjDS/Vz4MmHyjuwDnul1/BHGtcStQvsOSQJmrE8o6qRxqbwFU4sT7EekjvDGiDY5oJcdRB77Fd6BkITKqtYUTUWhB1nVeQ8jrRyOub7HpilygfGTbc0sNPuMtzHEkdG5xSkM+8kYqQfBv5ajjTAZ9yBX6zu6yCp7wQQfIsmycaqcdqXnQdtfj7uZA5Y6PM0Q1EE+fuZJaYwkwxoJYokjbD3V7tA4kBq6GoI7oAZeZ8mgasIPYcX56M5rxd2UHT31dtbrmXAcaPdv/B50f3kOv1bHTmlFh9wDWcm53hQcEQSTM4hNoHXzrGtWDFcJNzOMof7peoOujZaQvYG57AdIohtigeCLjC4RCMK32EsCazKW4305Gq2fPlS/AcEaDi/ze7Ma6PSOvYhyNlNTor7AryjEk7yEh9GQyVmbrsQgAPoOVl9EKIoEsvtozSXjR95pnu6ciQ3b7E+Oc2tOXIIIOOjT60AP4QjmGcLGpFNPrefR8/U7o0yacziIhxv3Bt6OzOoMJHjEhmbYNK4HkxHVfSQowfWYitILWPwC8oCcoGRJhKs6F+MzjqQ5OiP0T5sve7Z6TUbAZgl1Ua7AUF3ECxGmPqFeXjpeYmaT4xHeeZNQMGknaQrCC3xrxF2IKVsk5yHNXxeeEO4SDU1FRLQBjbWnKgB9hBW10msBnLkDNsuA2+L2ab/2Sr8M8MP9yvmn3AyN5tGDTsTMuz7GlQvIqaVVQ6EqWNd5vhNiL+LYlSoMypDKs4o0r3hxF3iF99rHqCov+Pzd9AttGHt+eqUY9e5Z4Er0n1+oWE18gSiYeqDrK+UpDzqtZo1ayQh2sqMmi7dybOQT/oKKLhUmvmedJWFZjUH5+EBhuJUM8UkqQW762cUYOiGfNgw62j94ZAHcx9WrnM+pavrnC418x7uLyP22LeTaRn3cT/OVYT4icd3TpfA4azVL5lGkz/EFtMO8u5fx8q/8P3JmA+or7k0D8xEo/adVZTVy0wazxFVvzDCu/dRscNJC39va0hColQZ9VTqsaE34bI0YU1owu5z1QZPUP7gAHOQbTpuRbVcEuhSlAiZ12CPAWd0usoFiOvS/s0/HUGS1fImtpKg+yRO4SJzJkQW0rSLRcC7uYMUHZ6Ndl0U2OPb2yv252CPjo8cVLIcNXD/ZAswT+E++j8kOqd+IIy+tdNYbXht0kvyZZ2GQccw5TArqrV0CemJa1CGLyTHCk8hejfm8TjbDs3FWRubTlUofAsjHgZF3GEGjnTQ9lz+njSVH1xjjfUe061/eGwfl8nkJf4QL9BviLnkq3pTupl16H3qCSK3HGfBinWdLdA1yXIVARtd9KvFrRdeB1v6S+KKPdVs2/JB4DQrVgMb4xsefQ8Vh1hwA3pMeEJkPMmbuZoYtlzjb/oGbirZJjeiekK+Zhr9tNwwyCsoPMGpUmzOyTAoXyOc2BY3n5NoorqNltJN4t6fwnocesOzqTgIF5BCsuGWnUUQJHiAftG+ohDATTTx8pARll1o2DaYqoM0oP0Nr1HFf7NmjUhtJ1Fo3xeoWr6/QgLd9sYJR15pAg7Dn/+4bR2JxkgP8PWHcwjIZQcZHjwWtfKcbSujMBHG9dNN/eh/jJyuHHO46fnQHNGKZzRV6dZBvK3ZFudmxM1Pj9uGaaWp3D0I7AFHnAY27/vVmpKpJVd1XpW/y8sg/LufMrzn3M3YtwgWfTGddtam/uQHpEK6Ne5Wb3rCzanhsjVIpGtZJzmpw+al/Wixy4m7M5eBOhK5xmAK9ve+o6Z3tgRYiTNvBk89TzXhJx7s+HNJNAPF9VeNxvQtE1yUbxvx1gku9W7Zx17f9zKNfj/eX95pdEqc79Tj7ZMY7+7uc8Q1KdGnJvIWxG1Q89wAgPd2FpiUZW/Wjp32PjF/J+2YTM8Ny3SwR/Esmc6d4+2b5nuU3YjT/cL+ddNTzWPPYmk4JqGX4bYN7Rgk2teW5rpitmVa6AhyVH+4THQtbx62RW6sdU0reVHZ0UdTwEnAnKgjMNP6fH2EXDs65nzt6/a3zt2LkyGp0e8jrinJdnhmgMpp4lH2ip2pNSzfVmxcXf0rkMZzar2vkKryHcB0AFQbXnLaKRCFfghPGpxMLpLz7JQR8DzcUcAlbIwGPJuzT+VD67rDBzWKzW2g7ZNf0YQkusAkywHOgbQJ6ip/ZvJ9jKFCJanO3ainL+YFgqCmRIWi9kFswe/R9/QWFZeimtcveNu6j1T00FHfO92qLwMCPDBIYdvZIN3iAvypTntw/PhO769PfVI176H9UKKF5fa88LVDBO/RjK9Twm2DiYjBMpZyoLvhV+JyOlFcJopG7MXJaV5bku6bPcEeWjxKnsdg5Jxd4vivhSBjs/PyB8mC660AjSSxBp8zCmLkPW+A9WRrcrhbiT40J5JbCsN5uEjsGbegrhtk9iOeM+zIgX46hT6nWoTjklZKikOdWJbBlB2H9qMy43PZ2ti50uyeoXryWMIe3f9C+6SXVTd38DDnKtri3mrnJh/hLDlqcNZ1Pwqb2K4E/fbd6hhza2Wm8OuFBpxShxVyDfSZC9ewUWEGYAZg/VP3H37Bhgrg030ABs8eWA5WZ3aKa5/f15aS0DToUz+H2Mshk/Ar0PVbWjxKv6YliW43UCFe8mFjL6X2WUHXqlGf/QoBfDVodL6LCpgI80ilnCP4L9tPZk4IBLJeRQ6THR5C0l/INt5w6QiXtl+akJMe9d862UrgKUSaEydtNwT1yvym0g191gYPZ404fPjLZSR0+sU1Tlck3PSqR6QJ+D+/GtBZG4ey9FiyQhszMKbpwRu5dYC2bZPLIz1a86M24/RtxQuhavcVEfY3RMMRyyZhBp49v10IT1JkdVZe2ywxBqpH+qnYsKRaFgwpJtb76Q9oiAbDDcdyCDYSMh5VL3U1JcoLXZtA3qPh0WjVaXSIRERDSWCJdZLXvFl1OdUMPszdnhzx4YhxSBtPG1Wa/wOOomhsSRbhrWWRbyRtvt7O1rXi1/nzEi0SWLhZBCs5pfdc1UOXk+jAl5vxndT6XGJh9EAK13UpS8Zdj1IGeGHB4l0YSwvRO7fLZZyA+DxuYankBxoJloWn6+hmujRgp5OyexGYgl+8avPE3fUmlGoSodsruGPyn/HfGq5Fka2RPR2Sz4vjnKrp0LtksEfgV5zPQ1envPj/CHouSj3MPn6XpGp51R3cWcYQDTPLGH3BV6h2HNP+2D/ubZespufdGVTmhQHcGSQDiW9B7pHur5P2NVoqYI5Bi4AeKRtHKrfi1inovZNOwUsOSAWWRRdt9SAGvaSgmuP0DocWFvArn/zNts+o38G/GBK8PW5C+H3Y851m9TrPCqI7ntm847gr2+eLABHqkav1p/z7uWocQsR2ZeKqLSuq6Mczx8EzjdnG2RkLetJFnq8BqBDoDb5YoqZ6p8hGd5aGJEIZXLPxxgOnxerv/f6DWASUDHlaxzNd3VBkWTqNiW/zzHGCKY4CDFVTTPhFmZW/PCWNYGkCt37APjKnb7pfXZPey71ppPuzboU7LRB9bkjtObFcDLsdqNQBk97SYJxZ1ZjhOJoClz7k69oSlY+DWE3cm3BO82cYeneUOOBOANXnsALqiOB/H5csM+uY5/Zp29zOBXV/9N9N6cjlG5yST4Oy4n0wCz5EZhypy8/Tb4oepiHIImc3K5VhODQNvR2uxt5BQLyrsNQ1hCDgBEwUsu27Ih0dQPlAuZ5mWyZyOohx2N6Wnq4mZrD20HrE5BvApKk0jQ/PTYwMonMH8quXsr93jHXuE+c1N2OgRE7szhbjyHtoNUbFjfRt7wNINobjzb1RFg0gu0v+nghUWzgQm6bA4+yPjMqUKE8A+Ht9RwDbjWn784OzOkfzbg69O1BTiWkQJC66TFKqVaIDedAP/honG6C9ubKXJ5RHZvM+PewJa/iROnkiN2m6ZddkBp+GYFDUDhyuGVAmRnpyXz8pUL/iouwpu4pjnKHcu3pLbF2OMcNdjMZjpXoNDC+jlwiYZWMh8UjZ+ytjTu+KNalfezkdgE7hFDS2SbaX2PYMoPXmPlUjhom+GGqJc+VOSgbtS7W7wVHEOLfVBeK5Vo+6SArOCretoEr5YZHHi7ko3EiLCWkgTNze/scKaxTIn+307Zf8rTS7/KleKfyMDnquWWhJWo3ybTblnhZmDYZfDztBFwx5/K/wJJILtQjBmHP/ux/dZHpS8HizGiebgW5teorXeMKSJS/Cbfu55tZmKuAEeXggQ2Pe8sXQzoifXqf4lZCfyZ7DfoP1dLPvo+CMhZfFgDTv33HY+Wk3XJuC6dflv57b5+wExa6CYBKrAWQ0yHYxWXm9UdnfRpCpIjvEGYg0f1H8to7rORu0nz+aRZf1y4XjGuFNfzdjVAiaS7d2RTS1nghudiqX7fb29oh4hBurzxxsbCSg6T/Yd0QCUFzXunAxCpCNaAeyQU+J2Df+mQcAChf5CjWgZ6uA7R4H+FOUeq90VaqJxac8lWLaAd773p3BAi36bwsEEe563P0LAfoSl0z51cFXMVHWcOCT2Egvssf1uEo5F5kbFNtSHmXU+vgPimwp8GVPyRW6XPRU/sf61K9sZ3u+DMH00wMIo0RhDqXOc0Yln7fQi8w7AriynfQRIRs1fw3+HteRnCQnfCDI1DsHtpbjafkoF/BLUWWmCt4nv47CUF60QsjXVnsZcMj9BEseNXgxasnOX7uWgHcnFeJfLZB/y+ry9ZIOtWAT4fbsStoNKTL3oue2AqvFG+fcMBuHw3+YcbzZbhE/YLiT5mu2F4RVdT1Ezd0SADGQGjbMFuohBC277FXBQMaS3YZoO85LzHBkOYv4r/b73phYw4viPkhRwhSy2UVI9Ne+qKzDjrxDjIG7ZlvgSRTUnHjwpcHZibO1/dGJ0wRTzxMR6/ZCc/09X5knmGzkUyN85kSrq/ZfzAjozvql/wOWi56Nn5VYR4u7pmZ9t7P2WmAj4f5GQKXTVcL/qGC347pIPY4QLp1ny7SyEpuaEXP4D5GJugjHJJ5Ef044+taT++ZzZlkZCPgmZ3POOzORxk8QFs7TDyfQPyY40mbiiL0wKooShSOivRzohHgvHxFFhUnV9hfCdZaswtyZNQy992YsukUuHTDMMVB64Uu9jFtTQzHyMgQ0fHrzRdfq0VLqeiMgt9ENzGwKaVkbmmmTDSpr/WfgY0SH9nC5VEBiBARnlmGigBPJDqtIEfOaV18IvtsFNDxwNSNmCVNrRfUXXZr5PKSzfd8dLPjdL2qbNXErDYjgLJqqZPIqnx7++vWfuMm4b+CQYmU6wjCkysJsH4WjhlGB/AOPTHIHLNfDGQlwa//xQctfjvkIX540wgSdwyyZN54ZsZ2/dASfyW6O9MEXRfVuQffp/W164R6V2+i4RNaAieU6YTSaPuZVnhjLuwzN1JmltS5boQdIRxT/hR73y5YK8Arl0hljpDjTcyvS3EF5Mh5L8rGgNNUanLFKVsBAoRprLstVJ4Hp9LUjST2ZVAWIiR1T6l6BzWL1r4wlz2bJe9i5PeGneZmnrZcT8w4eXnQpNDYOXmBV9ayhqITVRCjqgNsvpLKHgmStgIGmvonNxwkQZyITyEyZK8fgq+CaCigDHd+Kvo6Wx3fI6Fmwy4ICZbyr257xemVfTIZG/pG3k3FvQNGKke9R07eKzBP/1bBpAVKYTMV7nMn4p8KH5nb2g9OYiY7PIgZ98y5WibRaaZlJciZobrcEYb/76Yw/N8HWJn2/xaTECPNKliCj50XWbtLh8AW7rmDDv2us1ndvivHCXkpt+ZU4wWfKrmzkWCZ6X4GoX702tSoI9dGzpWkNb7zjF0eFPRz+lJh2ROcAD8fzrwIeyUYy/VaGtN/bv0794Gt9FpJg0qDvjD4BV8mO7s+W71++fIRUGz4gqBqGwS+RRWy03Eaei9vZcg+M9xGAc+SxrX5lI6CWe60uJjdNDa65mcxJKju9NcOqFJ/lyv4ckOjV3wIJlnMuNpo9NSd3nqzMDIeFzfvXsH1JVFORr5ee8soQZ7ju8VYHQZFxl32/OjZFUL/lugU+T2skpiIxnq2Bch9MQ30bdPGKKWyf+yfM1mfcoCX38t680suRKs98IRayXakLK8qpwWij0iO7hkzAtZgClipGNoNBG8pGkXCNOhyWUkdG2vvEZrEbwYQPQ7E6QBywYoawGPm4ayJCBJZ+l5S6xX7YlwqUQS8hLg+sqzDjWxABShLtrojozvYTxbGttd/90pQMEEDIBkZFPgsgAiG9PLDK3gyN8gXrvbd8VbxRGvmN0YGrqZzGWcAfcgEdqH8/ydZCXHO7+GWstQPqBft75PBhE9+49p89ovgQiyacDG3ohVTVW/yF2sMtOM+zomNBlDC+HRIi4T60DYy+mH3vd1AcgcEZ2G6ZUWn8FjUEsv0IfKyZ7YYZd3TS88LVt98s/eZp1Z/7sBEgZNYloxRlhu4W8unVd9rkCfhGlDO9aliuyLrr/QsDWNCKVKJlnVcCmrWfnl1M70UfCL5csHCvTnx871xHjH5JMkxQ5N0y7LsGJj1hImXc/TfdYArUn3ZaMN/MfHrxlaLavtNx6/yL1yidSZuBbFPDFFyX/rp7RASV5eOHBjP56D/yZg9VEpanLfNgd2NBRKWfiGWimJb1+qxiSyyhi7AppCcfW5oJP8HtjunJYyeX/rCmirzy1kyBWk8s4BMeivARkmBf8xcZGTT/uRSV+vPN14mJHll/RFbi4YxGw8cCrkP1ZVTeb1wGugXrjD5jW2wM+xeE75cNTfZv6O3CfnZpKA2eNhH21l8F7eivim93t/002UJCetnrS2JaCUbFkfrXJDH4Knj5ydZ5QdJHch5eryRb3DqJANPnrqL4jqBR3aY6iRDImBQHcvJK6ZvLmuBQYVoQBw3KpLi2DAU1NkFBkhXogjkXJ7qSdr1fSYVOwY9Fozv4YXCUdQnYo1N4Bg8McMdN614qX5XOdwCFk32EFKRJkerZYH/IjPywDcZJPIzhy5D19yeEZ9cgUP+IEvMGJlxQtSWKgjKGUrZRIrl0Wf7VMY6+B7oDvGabzXAfznDZrzvXCeWbCH1yvE9eTirvN5SJ+noNcWaAWQvJbbKX5KPUgbgcyIs4IWP2WerB69YtKAaXfyFJAwfgWqCH0AEINaOqQH3MQWoTBDY/9D8Q4hEkZ74VWMtwDBDZjaRST8ZBvYSQCqtNJluXqwNTHhNTIpYm29UDDRMSTfvbXRkoksVlHQOnktFhNIzUpiJtk1eQk+RwJyXa2jEY+ucWo3ntn9hZ/nftEQSU9LbWG3Qk4bd+TJn1jGG2GVgB1X3pzxa3WkS6s02LnVuCcbpSgxb+RKl3KflCosd86z/ltZWhT68v/JCltpjKieZ4aoqjqOJR9LmgpVkfdXAO+L0eCCG8s+L9QN8CfAxsGhj3DklhG6W2EyNweRAFaurmh6Lqc+Y7MqvcIsN6KucjQdH8p0fOSuTJ1UXTd1BsR1kBcGY2+BpT7e2BnS1um8xNpyuNAo6LwVk1YLacQF9AffnTTufO+60VkuhknEfYIcvNhvGVSbkp4dSNClnnjCkpyv1ONOGJkDcHlFq8UdrSNa5ZLOsRjJU+Rp+yRKf09WNKDpB06QQpb1Zhrgl4SoutkrfJFJ8gN1UyYErDpQTIt7oZBtGCcXDCkXYltGH4NwUeOlc1av0AXjKLZXNJxT/mZSXPamP/LUKZ1FMdh3o/5tQlxBQXj5rtUqarNzu4CHE9oVI2cFtO3LTgp7Sc31lTz6mWNSRnswykjV/rXaZ0Eed7C/bPbS/rq8tHzM47CjezLvdosbFFvfYd9WiZ3bWMeyNG0T8rlqDCQ4TNv9vzhUR5i9a1h5bbKGAFLyEPyajN8fBd/nrpR0v0jida3FwlrQqhuT00hblCApOwsu5f+c+ZRyt1M1A1xDJL9aP18uTn/FQboaO8pYeEoa+P/5RKRHT59AtRSQKhL9MDSkuneoH8bU07fdUvLbGRPhw5ig9dGFiP37DohaJSZsJ6Mdlk96bYD3YWgG96XvPXKajqZIhYYtqRCEKlU0ROtdRkGepUC0Vsv7eLN/wBtP0+2/aKmfwxARsCJwt8zcaD1KfjrZkzzj9Sg/hFtd4bYroJm8GQ3xbmXeZyXuKmn44eV03s/yZHw1FpEbClHlOhRGUTxek4YZ1mKbI9IRp+zjlQHe1wzxnHjyLIsJgrxUbEC3T8UAHsheQGrphFo7NCRlAZTnRMZjvo7S91G3zk0MXTiWr3T/L4iTQh0RqjiAPuylU7tGeQn8atBT1B/a4hAccr7JS3RO0ku0/zP2lxRC81e9A6tVfGZAllGUzwkCXYnkhR7s9fWivPFzg2rR/KzRIpQ8f9ZFnVl8cMdph5DHCye124WurocQrkehJA/lCII4Non8HagjByCUg53kvR+ozZ8RnbmTp4W+WKM+g4txtf4Ha7Ajb2boMl21XBxpMKl90MTpEpHl9pb2sA8COplHz59mnGh08ykpAaA5lZyYAb/W5qUqNgS5c5Nr/AnfN5h3p5mJBBIo6wNAjdsobNRy3KhFcTBi10f8p1IIm3MNDFlPTLtxTYOQk3kfoE3ntQ8GNq1wwiF5cFkwZbIYo/sXl3yn0PnepmCurgAWhTo0AC7vQw+e3HwLlP7TqZI7TVtTdZYlQjSa5YgD4tfX3Q3r/GkPtVHNYGKDuOO/uZZjknTg6+Hav0TqDdLhGKhpovmkI9DydAGPRT9DUxG4cepHHMwtPadGor6S6mhMQ0wyDo5aH4ANufOySt+dg/IUBdFNPh5MApVX12LWtiPpnPgkaq/SiWTHKCVHHXQ8JxOGzPN9D3oturATFsOajLggXQMFRw29HPwVp2EAv3/9eTjdToaORaiisup+pR42Zr+1spZ0EIh234T6LotsLpBVhIXH40Peyf3xDU0HxdAUbs+clIMwZBscl+QV1TlTYdzw/yi07Uc6dEwDuboK6PPhb1IURd8zQx0xdk7e+jnnNk88CRIc8dyrB3PUQA6u5XfyGsh9uiQuf/IbbCRd79utwH71814HR5qELQxVae7d5zrnZlrVVcq/yBBhSws2Pdn2NlEojqvMcpTc6Ps2/iT/TJosow8UDXxwPwE/y5zs5wg54hsUXjvOjBqt+g2UJuTmGSjb1XMwJDiAol9bi3zXzSSuiQUzyC6bYZpWD70ldQH8BgeHbt9UV9xBzxoVzAFCFlG4OZ8KjCGitujy+2OsZ9s4nzpqHHSbaubtm1SaL/6kUjnWSZjja1buGsFSdInMXSUbsqFiOEMDjYjdjq6RbNyWWCvztYq31v/mu0zIW7oFFrfkdfJcmH+DMLuZPxNAMxzhevOP+AJVxo7mJY8D6GcGOz6QmgYrF4K2khkBg4MQZeV4K4D//b/7cB+GyJf0+s8c5EhhEqSGdgdlItMEIWRvipnRJGy9PVm3rS84BA3P1//Zbs/sHc6DI+rGMQrOBIV/Se/7xzwDhNZdph3XRAzHdGn10lsgl5n4Zi+vqqfyxc1S4dSGfhOiAHsXDWXryfs5kIc0TPb8fd1Y7qKtBMZ6XkrtW9mN7I805OduwMkvJKScsCeGGoORzQ0MMb6zySpQCBTucEmIWQMjKbmgaWQe4auQ+0nRwOJUU6dBaJTMdonR0RxfBRjFG3pEB1yWr4TsnXhIbxdQijwnw2q8xz4ZdlMNpK5tr+PSG7ZaWbA5/GFxrYyiz+mCPBZIJrmXaiFF5wgs3lfZMhHgmCeae18qslD6ekGAFjt2Fj+9/uZtLjYWKzlQ+js0r59YYtjheOdZ5hF2B8bKWqbEyglWjattxBDNGftqjWVTWiVWOAtmzKn6jqtKJ9/vvMGgwXAPKAFiGa/f07MVuCWJJZSzl0wBbsz0VyhG0ugDb/vfbGt0I0bPDNNm8w16K7OEk2HhmyT0eZeGxyt88le2H1F2hN+jFZQMhAOiDRC5E6zJQJvHCVzsfNqF8DZ2Pk/Ae/l5TlVZaNGqox6U7kizoOyM8XCC7AXoMGsA24nsDIiRMmhhbz39/QQpCeWRP46ziFYSlSRS98Maa1Cj0PMAf71so/6/RGLTr4ZteLss4hTmjC7YWQgGA0ePtVP9ml+A+Pp1oFu7LhqJP2nYD/X+7qJRugr6Rf8zjkvOD3EbTfOON7Jj3JdzZoW4TzUXkhJgjpPY3zaPTWAe5cAvmVgGTIMRfpepReN1J9wSgtnUF4EXT5jz05HJXgFRgRphQIvTJ2C6pkoIuT4Rz/K62RQMdGDh0SMSWCRQ9kJrUc9XqZDIMAbZwOyVpZpaMXke0jy6GF8ePcLgBDI6cy2/gW0vbHRnqpcAxvMP4o7NNgsf9T/Yw0OXdXBKgJlpMpIUZiXz7kqlwQUxeN2X9uemAYrALEPdwOEUQ/LVDmN+O4QQfjgP/85Vkv60y+GomPeQozXbnMc+q+assgiQbE3IE2+pxqfH0UtyUaINcdBwraQhRaF/3RMQAuqV934h0Es+ibV5N8zsm0s/vEdTdeCHl9rovRJXSUgotkHBQU2q8iDREqx7CQn/pvezi5/3oeo96zBmj1+tCYh+IToSGJxO54sUIghKioU9fqBASRQLh8x6HyCOAFDjkE3FIJq0TXBM4RXbdLap2mZZdK0OdUvHNWY/e10zAavmLQYIFpnG99gGDKODN4Bxwp6cjMCcPtnA1NYXdQ7wrxdibu3c/uYYafS+gRS/e3UlJkNqQM5YtBTR/7GASgHSNznNkwYY0KDLqsB4phzPSgEFNkPChZmpC9owXi4OHnWJRP7I/Kh07MBwEXK7voLj2iTCKPglEgT2BcMeXxypcTWaaGlClPMglDkPSQgdNRUrKDsCfSYBM4AbrAHlie2UNSXP4xvL30fqlieilcLMe4mhrRQlmmM8h3Ny3FhAXuO6QARr0uWfDnHG5yGo/J39d0vMC5WdxCbsJjAyPvJKm77hCNa5G+yLQoyVKyD2HjaB+x09CX1HkstAbeF4fH0TJfyUGsiZKBf0uuhw4bSYgaCiDb25gUGC6ApOR9NjpknNrCsXJcwqb8sqoqJiocDGW9yWOlwG6KgQELft2TGVdHSK0dcYfjTIbVCWJjn3RsW9+CqrX3zl/2EohZVgh9jTsNiwahhn61a5uGmsjEfwaA49aMLhq8gKDJcZYf3k5CuaiMIbTN9Dv8kwNvOemevxtTYqwzA1k7dNx3PfJimBvdoFUXk97uPpbcr0URHXE+p3GUVA6TXp7hIiT9uXDtHTRQD+1PEvXFlGWzX2ksorU4qoCIxyfI95LAc1h+zXsY0gGntzcE3qrAB4yV4N4o5rK/HS42Qgkgt759wQcePRWjqtbZ9SlYl2x5l7hI0kIvuenSBtR8pkPPksIciexTyfA/ibPu98sgr0B0Yyzpb0lJ7JpoFs7OUpxGHMu+CkRO6WXwgHSxHZE3E29An/mS7xzMvDd4C4G8TYXZeoh6igXJ6kadrlKZvhQNlwcYxo6vUqXQcMj/O3CY2HR1COHHldXu9cnqG2xQ0I2jWTWndVL9WeOB2eXPgBmQGHYqPPGgKGKJasMEpo5SZInGY9aqePiFvVWKOyPC1eWZkcCmzPW03egljNF9PU1vnYj23AUVhR8Ac8WVh4F6prm0zU2kxI391/Dwv8wJocgLtfsq/1p8bJ6wC+FO3RiOa46YGDf9qqVveWHux6vq/o/Im800RiWex3yenAfkh0pdBqvED0kEXlio2A3F/TtX1Wkb4SiqA1DwUQYXwPvnNjlAlZgM0CasYx2Cx/m6XaS6ejFCEJpPnbc9Q/JCgU7OkbXAOFtravGpey1uSwTsC1bWKVqHIGAeGAFHr8eExSfOzcDUhqVPc99wNRIGSmPPWnZS/y9SOULCHbR3poGXvr/xEpkj533pla8PXFuvi7PTV9qRbuYIjaMXGGNKG7FpxXO4NP9haDS5ieJarWszBIRalwy/HTecvKoznZCC+zDq9QvpPD8eSuXR+mj4CUfnjzTlKqPeN0jJuYivYfY6EVeu/OMUpdqYL/FbqZkS/Q+RDkotvBEwy3K7V9HNKZh2g5MFfxvddeeWu3bXjsrd6+2BCxK18IIHAZHVD/qfxjRBvO42HOHcLHvlGtV+NZn/WdEyPD21/JtBl5Ce6L3SLmZTsG7J1ggIQh4RdrTUhBY7NucNulTCG267mNjumnOGR8Vs1Yf+aUnr4U7ll1YRoX8CsYcTCulcfLcQ6/xIf23Wc5VsMOwAkf4iHjpKVQkT+4jHl3lZYzIIGNTeywr9OjzH9tgrNlqQmBk5pkhTlpsJJubFPm5eK3J0Ez9AOWPoLlxw0N4cEybOFRYRITS2pGaWomc5qG8/CBWJ6tfkpnw7e+0anU3vn40OQeYOejgiuKLB+zTqfQE+PUd1jp0h9kwHSJswwaGVdluK5VEEKx/VSLrNYoT3LNUYfH95uXiZ7baGz+GWPgyUrM5PYPehK8vvy9khyu2QXSy0Cgyq4BUh55F9UGE8QF4X5vNj9evlebwA+9ePDj8iTRg24ivI+iWREDMnuW3TA6BV7u99gffVXQy+lnHCOdcgnnMA1Yz5iycKSEBzMTOTaolWs+BvWoTRyaGmpLyiAqGGuP7AOxBjyCNcNNGZxJoIa+QWzDxNgnKuaG1PnHXOvPonE2rNLWispsHlPQjyps++1ddy5WttyKd8W0ozf9vQ2YldGvRSPHBMwB62ZdY7D80/PJY6UwLsLYTA4wBnyU1vwkQBBQoNgie6ges3liMft7vlo18iB5KPUFt9p1nwCzlp8C458XYsJoVLLw3iDMSPM5GvvDXQhPdI0rlIt5pFTIzOykJkAfHJdkVDd8SYTmkS1S1RFgP4rMuKcj1YAMkn2QqbTc564eDFCYcgeM+NYhQITpOrBxbC3augZ1x/xV5Bm1ipUwhGjuM/EXxC7H1tYkqnE8EFM+96P/axYktDIXylTRVjmDnjkmkSybAULUtcB337hRcz/xrNozjTTR/d5Z3JJWUUKBF3Cqp1nZ/3u91wMkmmE4arF0rIrPduvMDuSszR710XJM2wDb5uqJNLdr7fmW3/SwxvdPMgAjc42mrIZ51YduGYG8fMSEGvFcqus2I8RlXEDJnHvXf/fHj+0dzuyZf8oEf4P5J/bN9cVfWop1veAGVUJT2gWNtl7mlEOYS0DSMwMHSNGqZvUtTyplZHj3JnMS1JYm9n2NkNVEwsR6D8BrYED4FMDWrs+GcNUlHaZryLZtYiUY0uQMKdmIftyu0Zhl6UZfkOhI95g8tq2AMW4XeLnPdrJxtpdqpc3BevgJx4shXkwIbWAPTENUtDKyUBy93xvDtUeq1TJjwz+glmzg7Z5p1RUOpXawsaQM+8FNiSxlCt01tgWme+84M5r7RZb64RFoFnb4TqQGJCLPUcXkSc/fnkIzAUiWsPy1OPb/JVe+BGoF0FJpFhAy3kbdJ3sSwEIr/Cu8n3CjVJZkwYtg3ydGtZyyD0NPpxdbfCNsWb7A1oexICCYwCkWolv0cpppHRLqkyuNE/RbRyMp4/FT7+Icb0NitqFQ92+FLyYYkYW4D3cKDIUcNZkS+doOkJIJ13TrXxsIkKPXpfDC+3rcsrxzxSx3nkYIeq1wTExgBhUyEyrNhdIHY5N12GxeNQJeyHM7B7XN6aTXDjSI3ZsboFIkjFo+s/k0/RwJJGLNA8AdkcEPd86rfoxaoyWP5FuKwq6sfU8KZovyauBzMBius5go3CWJd3kKnvsm/3XxXz3xoinVE8Rd9iPSPl2vOySJPOe0bGT8s5GmzaU0bU2mEgm8yYwsCA+p55AVYr5J/nneDTpQ9nvGQvyXs/I2vX7Cj3CduuMYDAGz/jySk2YFQT9jQMgAAdSL9pFNo2xo8j1d7/jCpPUnuIwpYuuDqLVxY2L9LiJQZedgSUFvCGY3HItuRhJOMUwx7UfNbi5WYLuHs+M6r6vokLSalSuTkkJ843GQDbIUPhJmgnzkud7r8cO+KKbDsPEAfYWRvnH2VWfleRa5PCJW+ta+E4PQX8R9AOoVvqZGtGMTH2UgGZOHEdujdcKAwB62nfLp3ktApQ6c34WSrs6PXiP14elNefc2mVQQD98ebRZckTx3xMqs+NuWbkjMxnoZbK5YLHRRYe7jTGEfS0T3v6ci/KbGzGzS3Ns7KNi2YtP32xyT3XY5YMo8KSj3DgTCsY8gGOCjLOaS3aVNe/1sJZjONJVO/wkLACWR3jYZToeAMkCUv32tDjHdDZd1Rjjb3p2v88HM0mdVKF/HLDClk4MPB8+t/VjPX+kAmc8cP6NqvttbyB/2w43IabYW5im8PTEizA6hp6V9LakQlvxOatlDjww/WlRvvtWjrlnSYHc/o85KzetDnk81lYBpMFA/T/HqUpennl4znA7eIOA7EQHa4FMjR1oj7aW02rtnb+E4eH0TW6M8wngL9tJxLZhWTsdWUujLethJyPotMVH5Zr04e8lhLamMiFh+lRY7x3JnISAiZhvCUHCRx3yOpydpwy+eIjp3APs9qGJv2/LgZvFfMOwD+BVfE524kfRx0s4TDm7fIop69bDDbAzc+TTx+uD9hva/NRoYOrQNdCm0AaMIU7U8u+tNLdqWle0NILHyr/8Sd6IHHi4/l5eY+1CNDVDInKsXB3yqkIPaC2aDCBWUDF0faZjb5UIo3plYn36A/L2oimf0FSQo6qHNQNNy07z8/IAUfk97sUUmahZ0Qu6pR7nwBpoylfFJ3aFIvzGB0NJ/iIPK/3K5OIigLcWtwRAzY2O1hBJUP2XhPSf4XqtoMxVVmoTx5TrlkenMYqXhDxKo1PNn98sFSCMiFx5/DF4530lxUjNl4bWnwvfkJqStAk8trflKTkYCdwfJffImjVIAEQuxL0ic6Lozz/hwK1ZWPrIYXjeE0h2p/AZT6osMbPxpvtEnNBySMBi2hHN8Bxl6HUytNWkFrAB9deYJIaZMy16twL/QVeDHz9F63yzp1/fvDce6Z6TgLckM4ZsRLJfgsjNGR85vVsGHEC3sdTdA4hkDFhXziAgjxUlmV6t2UmqbEHKZfOLvyj7ff+2ej/ymNubJTjxGtQMuVfKIA6mWWVBFkTbxTL4L6zFvP/u5ES2Vm/7tyBPD1A0AF9dKjYve946b4znbo9r88VLObp7Eo+jp8UZGL0TgKZ8Dvopy3WE+KibGpeKI/Jnt801DcI9T19/ZQGHVwqzIhfFRBQl/taT26Iy87BEDqrXO1uqfsi0BKLL27YNHCLlK3z4by8p4keIF0D6TIP6RlfuGmJGbKOKFIwLbNVks5kevQDU4XFKAwx5WmxcvqyS36UOplfL+W51TQkWrb9tlwxIaCzhz6/oFFrb3E0PlogjYwPsKDEgdVo0jebbdtcoOX/OYL4jgBQ+fdypHdWOND/w6wm/+eQFgTBgaxWlJf212yV9dbT7mvHfktv+Fjauu1zAQXO2bUTaSxOgS0GA+2GtzU5znjfjuXiF++hUTqvJb0IwtzSdG/jZlUT0XQ6Fnd0xWMBKHMcJgX6rLNB/7HLlSTQeWK2njsxBDBUnhfTaOUVkIfrFsqM/3pfWPros7Ap3CM9NCvMpaiiOkZ9pLJeQkaoaE4c9DqOFc54d/s4RcGKYIx8PXIno+PEObb1PYlo7ZoHrrcE1w5iiPn+8hFpiqED7fSjk9B3ThQZj+UrQH6QR5y/FLIqFcq7m4aSUVCMBQNf29wo+sz02nEEs+qwzIGeN/7FdP234Ca94pugZJfIGZNsvM6j6ous4PU3fg5iZ2K/aN5NCCMsTmuE/xJ1Yq+F9QdNbQD8SvvvmUZJyhmfrbC5mxQDJrYnv393DF9DWBjGvakbAAt357DvA2jstp29qveltS8E+Wp8Na/t87AT4M08CPgq3RJyl8pGNFJOslK64alladXk8Shm1iP0PXOg/I9CPW0eqQvfazrhoEEj34SSvfhgVEoYVVaubI528NpXCZHMAKbVnVPxSrAkTrv9tCJvNk2QPRIsXUkiBv8tX7tQLPJFkx0pBt4CTqG4SbaBjMf5hwaB8HiHUHIWsem20mnqqHXeZdOc1G/tZBV5KQRtlIt8it14q5oFoTS62FgFWDY1xjDUovgMOhC2L2qc65nXFgf1J70/dYg2Wvv/eFgKn5p+pIhOlT2SbBIURTOsYQtodz+pnQvdTeVk7s8KYcQlcq9h2eNZdRK3VFEsTTQiMRz+qisgb+gwuJnE1Niigst/cRO/7XBZFKGBbRrYht3FEyYvtY6/dCbYxB5LM7QGWGeUdU+SL48Eft1as5Mic9H3k2lxlO9pqRcbsbkeIw8GS8VlbibuGWfvTsiCNSst1apmnNBDfJ/ps/ZMiy0whNGwTB+hwETN9ENutsHwlPDgaSBHigZw097jMRzO7hY/vQ9NHHc0GnwiFSUtPu08AlqgXHYJUFs+9Z3CzcIC8IAj4OJLrWmenwWKFh44zzwNDd2dOcVbJv60pGem5XWWyg2f4uM1m5w0ykc0GRhEH8wBHfbz0xSwFXWJxVSV2OIZkBp7Ejv3Ztac1UpE8NzYukbGnO4qDsQNAbc04MmBHmn+kIXcxnghn8A1MmUgTyvgscKTqSCJ+n91S57fnuTUlGjKyA54Mt5VYDk2tZyPL245O7kTwKtljESc1t0Pn2pGB0RuR0Bc30QFC2iAZbzj6WfePWBrEH/yOZMyblpQWKtHC158/ZxYyCLsij3WIjF9d3v5q9SEl74Ii+TZP2kqBqSLp0UaEfoCv/49FbX41pllUgAP3cbTfaScYzvc3Mzb8t9hGqeVqZsso177mHsnfQkoGn+IfseqidotDt8WeoQYv2VrXYO1MFOt72Nz3vDlgn7tnd46rCStm0VsgIPVjtuWUM8vv2DcflsvPDMkknI2uI6oSJ4/HyyDSBYXBH8qi9+628iQ+ILeeRktXfTZU2/siHgS5TiQzkOvtP87lqC4RW+NrwpjSh3kaxGA0AzNLC/BCR9K/RE04Ctp/AE0t4RNImuSbrtWdv0YAAr7EslmZUECk2X4Y8PIUh5Zqa+U8MuPz0hOgQdDKYC4vTt9seBQF2zrmjHbJELPHTGY8cMrryH3UN4CLYp/r0KNAijeiCwyClLoheYqYvFFGE7EQbb+xOaI+16uEzaPeU3vRAefyteK3yNs0z7tXkOAgLRXtag0gnGGeDYM9Bh7Qoo46xey6hFjZghUtMuvD/vvFbTDLASZvMIaFKLYaeEkZ1mh6mncxQOQQIPHxBGN8Vy3kVDWeMB1nsDl7XmzOcD+6xC7IEXAAb4qVEU32ACMlPq0Z9nCkz76Gk42toUV+02tNkDoYGWcoG5z9EuHDhpniMe13temPWqf9iqm0QXSt54TjD1pkj09k0hsuiCkiZzdR/rhx5lqH58RdgAPqZRHLyzHC6+7a1YyvyRADzEIGYeMOuylzsSkMi8itbulwZo/e2JiBIu7s/v9crr5rlnF2Mneq1x8HxCzQQGGt3GgM5NaNQ413ljsdm7jlhvFa8BlJ2ecm52a+TiTrAnSAW7/ZBQhTn11z5YFJAVk2GlZAl8VQ6HaEV8//sVG5BfI+/Mx+E96mjFXXKgTMQn2GH4YmH93LKeXl4/RcsoXM9E822wi+9dsWo+sm36wPIjzo9RF3qH1d/XpaRsSW+zqUW4RbDYjjloc0ltNHT7/TcVBFNWHuKZbLZM3Zf+fo52Kasbn0SWJvtAzzKwTNH32+h6GV5tkcMP7ryWw9XCmkjtbvhJ7kF78rZ1VnyO8mCnqE0Hvw/NFTbL+kAAnelfUXZXcsLE5HK8KdRqrX/RsqmF2M5RIeFArSplKVRlg+gPauzpmQ5cZWRR74ylS4Xc5siwP1iu4FWZchQA1hN2Ssrk85tVspBNpM7wSAB8vxddTNX0gYLuYqQ+a02cYKa5BXjDYJagNhe0FuZnrb/coQ4G2YlaMhetxODmqKT28kQqodENXoSdsYVAQroBS1/ms233fotHQAyBvqsApq3QgTPZvn+Yc8s0k5VejO2QvUcBpl3lDBOHqsGoOUGW9dlPTSjP2AOg1Bnv0k5Ur1h4PDkKR8wp1GS5sgWvT8EQt9cbrVwLH56hp1VJRatnvuuGe4RP6yB0/qTgYOiDYtPXCvf3R9No8+v/fEQv6vKOSi+vKZEVEJWZE9QIRysPdMINaoKoADpJCOSCk0Oq1Jja/QrwTLFUF6/aVFSXg9/+7m04EtqeFFaP/QumfXDJympx+YUDZFJFP8JWb4JOOKQCncy85VOr3ZLUrUM1Al/4W3hzS/A7wvvkh2FKLnsWAvXgQa+S80eJES9uvzhr5lUV9XgjYFC0j3WjSaBrZEjf3ll7mfBGbg20EAcFoHUGYNj7aCGLl2HXynWT8dP9/97Xr+o9gOWJJ63eEuQw1pyAquhy8CR3bgDVNdw0WKDlk5Kouhrh16vJswKPQNUBuUdfFLiIXjpjYVgVfdffK1IE+lbj5b3kzYUmv/oMmKmaf4GKptoNlMx1L2ddM33afmcko7yJQGeKHrc/hNW7kTo/z4XkSvZ+sbOH/A2Az7Yiopkj/iwRA3pAMWvt+cVPbFtdg3YMVrnllgjZXcShdkOfZWdLI24G5n7UQu403CqaidXR8tO8CI3g+KEqs48VE5LkMdjarf9jK2d8SwK42MDEfnQ31JWXcH+3XgGG7V8AM2m5vu+4THQ818qM0e/Hf7aoNSlrLJ012QRkUw1K4Rlzp7mgKE5Xqpj1LFi5TTOyZ65vHXI57KKLxrNKyFsLPfGT97F6EKxNVrBNieBYBbM0/trdqETCutTOuiCLUmNuuWqXUSod/6NKj+07tdPRdDktZxEq7ZJXxA/rCgRFiUQ3NYadWecZbBX5PmLnTW+mGsn4UbG5jL5VqwN1chw8qfepXflc5n8fryF9yOacLMbyQov4ItJB/7fulJIed2x8LP15XLKbA0t/dstwEBbvG+eb/uXN9TopY+Ep1ngi2rAp01IyrkgNyF4cq8QlKsZ3pFcAKT5cRAT6f2KkX1UINwcZ23qZ8hIXsrLo+/yA3tPg4gqplE4p3DF73kvw0cVkZdCS7N9Mz/NVuHGwD0hChNUFMxQNgNcxc6ArKUNWfPhk262Wj7wnFIPMKMxFhNk8rgrx8Z8OqjU8Tzbz3zpfQPNaNsJb2OBu0sUrR6UaTmOqNRPFQ9Su7pU4Nyp0+g3v4+RS6o5cipmZwsAu+HNX/ClmKs6KHSde8gzHnq2ERBC2Xsy43gtsq1UGWOvOiOhdiPXkpmOFhABexPhXIuWFbLinOn6VAIJayUpshvGtLuWekcMuRI+jIvJM4iLFzM5XexZABF8m75/68f0TCxL6o4OvBTQS3ZqUrTtKJEeGjIPoVQuAabx0cXkHOmYxCYqq0SbrWn+cvX6WWMQRqRNyRQ/PYj7a3SryHa9JNvBUgLZl2+H/+rt5r/Ia8kCWuG13sDR2vWw3mTb2xcZF91oQk9DLqX8lURXEMZ7XO3cKC3uHPLSIrWJu5HGwx6ZeXQhaKYpgVoOknYlprh02aimz5OAG8M5P4h9NfWWjKjV/6XzJ4GtHE5zY8bM4aOm6ZIRAEwAHOJ7GZM3m/2m6+LQGh7qXSAO/LtBKfS6GwCUvpgPot9iqIo76PPIlL32ApesMUI/4UvgNiTBERI+PCgBTVx5hUmC8F1z1SOk5A1fho4OkbFZ1YrBnR6OfhMXFRcIoG5P761XDyjQVG+z65imInIbhfVeJODyRpd05OhBXwFD2kJfv1oKhaR2lsPjAjOzqGsFlTnezeC2i2Wg2Xzf3SjFAA4l6Mh2ShhRZAuE70reAcROHtnuLyVriBmAPZvZzyb5tnB8UrL7ZinIjJxZu2fjsleCF9Jv99ofUK7Cy/m8/ZkoYrAqGj9OxO6oIsFbA9bvw2HZt88MWcryBHRMR3YxiYBCXUIyHKqfEkqsKv+khbXM6pb1aEMUWP/UHX/RC6VcV5h8SFB/w37GtAJ8AEwrog42ERk4FL8hJ6jPhqn3kc5T8UjPbDRxRkP+pCEoBuKroKLzbxXKkSviqBwiVoPCSoyh5dnLWj8yVj4/kxpBpRik/yJ3qNBdMF8zxe2lhVZJe5aVAQCbCHr0tmXV4y2uEmwEzfu7r37Sg0LS8N/BhQ0EB88nhg9dPlnlR61ogGyBIbrPkKZLHfUq1AToYiotCM5VTY0A5n3d/AVu/qxTUuoOiM9leaNFnHGhy26vIUgChIsaBXp2ql+XyoaOzwsyqS8rRBAjc2GRulBE+5btmz2GWhcBbwCu4uTTya4ZVNWGIEEEL0El9T6bG8mx3GOAjh4UcpLbjAjJ+bZ0y7EbhNt5xEmL1qyKZiRYhGWhg2um/KLojc3N7f3ZdQvYmJS2JTMDE47AwgFHazq0rrOuyY3r/oxCcyWcvauSDU5FOdbleFrPxBVOETyWDGPLA51Lxs3M4Yd3MJnI6f4Ju0sjdWt/tNNUd5CTyIvUOokG23CaX03veJ1IUs3EsZPi3edGNtnb9Ljx+zMUNCgoD5V9rNLDcaSw4C99UqlDavxEOyeCx8in32EZsbNaHi1Dvf8bP4M0vtTLBtpI4Qy0Nd7hP+Yfv1CEXOy+914q273BYqSBmRztE9odSphXnorI8F7USlCDG/dNqhmGX+TH6kQ5IRtsHMN6S5GuXSRnlCcsrv78XWnJFRSOngidP8sP+Sw9+4gzTjk6ClrpQgbZbuEBKMImM5TqQ1IOmQ8ZgRn6fqXJhLKaMeqNBmxoDyDIOOayO0OJVsc2YnmtAbEGgulJdy81rJebIBhy8/xOp9AClfKLOl5ccpd7CWxNZCVbtk3FA98e87JruDWD3HE021mKbxTNg7B87YviNlbGqXAnA4ujyYqn26/ferH9otdVu3ZuoyFo5qNVc52J0pEfosSZnlaVcnS9YLznYKXZf5QU7yxJSR5tVL3a8jGL/bmpmo72l2eGgCaLP71nNgGJbSEHYoPjxgX9x9s3GlV/T7OSfhhsRbyxCq0/TORqqpIwKM8ervWXwrzbVPeMvLMv2aTVlEDX7gHO05T+PTDGBKlRHr1fI3S1NG41qFKlpUL/5/4SEN27QRJe+6i12P0yNwnPFO2xsKorv4XNTBC/w/snu7ctRP7/86y+V0Ex6gDvxYShNokWRgkTisj4Yfx8Zih2jP/8L7iCgJ8S5z+0xmswx2g9QMq9fTs2CLa+wKUm41kbvZ4CegKoMTxWiEsGyQwZ5qFW2S7NRQau1GyAVlVJDkIoqMHS0Lye95+AYnGukZ8+tRoyQUpFi2TRldYMTBhoIIBEdefa0KLVKcqLznuo5pftYzPLk4sdY4hLchz+fcaMC4HNEKbASlW8VYder09sBiJPpRP0lw4UExeplTnULKkJHNAcoW64K4o/6T8zgOSGQNiVr433v+5dLQpV94/n91mnYGbi0SQeXrlFGTGWgDwGxqKh6kKHVMly3t4EN60dIaW+g94BAc5d62q3w3alTcj44HVn8Z7otuUCAfFk4fdQs1YUiH/O0oLSwxSbYHBkrt6/Jg9JDeEx8Dt27zrK8je+hqnRgnZ/CeXRhPILgT8yJH2j1u9yDvhknIX10Bk5z6FxKLzB9IP1ogqDttd3+vE8GdhTaOgndQPnWqSCiTtrsAiOy3fwKrftd8oSrXD0Cjz0CzenfZxG7CS4mqwgL8tyfzBz9WJj9Y4YKvVbJk3TwuTH9sJ4imp2mW3I5cfgVUBBT08E8jx2xMfbXJdbfIwh7ONzocC+yxlaCYDh985qTy5x1/kqDljSsqLJefKMjgme5RGQWKJ/MPM7wtvgpPudKydI/xBwyKdCETGoCgDr+JUs0mKtp1UWjnSuyJ/sNmwwCWJpVu0KrHo2edTrOtCvq4EqS0I4HYFMk8SL4gDcjHHPKQQT8kW2X9nWRf1PTefIhQmHfcAeRtZtukQaZ91MZTYWR/4EVFwtGqmZJcpvQj7LCeRwfP59EQ9IkLVPvgi9CfSwarF7BGOVC2qsoCnjhkMPfyFc3TVQV8FixAgzebeR8yQYY0iIJl/55tENZ+W3mg9vgE2oR+3ZlRWhwynWCAsPjtNAyZcoLqtekJHxCVH70lIl6wqyfZN5eTdgjScWwDNynZ5xq8f97is5y8y0KpBuK7ruHcSeWJXbCTfu9Y7KAGBWvSnAkxWFLfRgiuKla+hlwQDnrXm5G9a4lqTMivHeaCqyPwcdbGkXq8byxV477XObCVqI64m+pydLCddiU23ViZdiNqsvmJE3SPOHR68VBG7Shl0U3oeVoa3SDi7JvqNly9X0O4qS9PVu9EXUDlscrz21d7qEqQ1rexU20CJrOeWINa0W1tXetpd82oMa5dacZbbkg053ZwhwvNJRagghNRYoe0iXnCbY6VuMajZVGvegxLMElk/HwY+P9BxRjJ3/fUVv588+PYVPM1akd3yn9NiFfq9833dpLGIOiwjP/XaTSDHbxDViSelxtVQ/ZN8HjQ86YfH8nLmZT+CEDrtlAYrqKOULV/e7VIa1qcNJXsw4+TWoeJEPhm7YfLcnkdUF3+lnSE5pe+10l3RI6xxWAcSVuk1pUKRd2lUFo04NS+lQaKJ93gyVdp0pMYq7FqcbNG0sFMdrdQDD0kxn/b63OqpsPPxzl4OP58E3/cdSeNrz+wLa0VG+rKkiHTIx/pE/LA+vdFPScchtKohLhM+FBhuqw6YxFkTEnMLfAa/9cOQy+i7Ctdgvs/P4unElhFXTpAo+MWKrKxJkwSjsj9tBY5w8Omg5oMou55Y5Ohbm9hm+Qkt9cNQ5oYwsPxIQTHZiAEznP7Gkf3DcRqe9NR0xFiWjHN/eEClJ0koKi38G8UvlvwtzxB3wj8S5HyKBvBvpXvLrkuCsaF+NTjcKbTHZKoXRyxCf/CpAwqlfDwIe06AurmXqmjHTwmsCD56tats/2OkfPgSePX/1E1DBquAzwI4UZb+jQG7U9F3alP7J75sBt7VXcxUp4TJajqs9+l8hw+078YISqn4EFiWuy78L+u3z+bY+GlsTNLhPDum/Fv520l+uR3+X4dWzRXzRmb6rS9MD8KuYOsi496NLR1owTTizK5cdjkWDg0DRkBh6mvfrj49Rh1JomDcBJIpNYh9/VcxTtRP+sHSGjyxONLuJxmMr3NI5dUZ2FxZOfcsM5VOFIUnsV7uO1Dx//7aSFr3hkWxpVZ2c/0M9CKGgQgjjcHfH6ydp+ma6w+UQ1z90+yLiP3tbA5OAMu0tRGdA+WOjKV2XMAmUcsNQUQHrX+UaPofhW70SGpdka5CHVVJIiKuviWwUusB/FAEUdZOVK1oqCzQYLGdy8iJJzbOhJ9WzvWlebs2A36U2rC0zBGrtGoSKww0LiVJW9TVMjYOcg8+rRJYyU3LXR1ihTHy7I4nUzVTnHOfH6pBfgLSI2h65g9qOsTMJKbGPZTgzzQydCNjmIjkNXX9ULm8CLYWkz0aSoQwv7ihnOA+ihXfOd5e4roW6VW8plhrMIot4j1ydyn9Y8lM7UWxh8goCaYc1NEL6GMccT+1mfQ0n2RNzftNiyN1lpOz4X+9cU3n/h4gGExYxU6qOFtwq6bBZpDxSf6tAQkKiYOEt6kJj7YF6UW1NGvQZw6/V/oeY2AbZWJ8d5iAKuu4+sRp7Y/oVRYGQANpOujVlgWF/+QRP5CP7ol8CkYqP3rB0zgytrkaBw1ZnM4c3gpeF4j1kmkFXe8I+934AqP2vXAcpn9pptTVq08VuQtEhPmoMDgr1cV2h8zXzZHs9V8L0IoFROGU20deNGAJJrGTGHlTg5wEgbte8AIomhSBo20TaxOytEUWiRWHamRWlgrJ1RNLgQw1gZ0MnxM3ow3lkihCNk5nnfyUEAWTVDbj71XHOLk80zbtKz6/dThVMBHMmHRbL3yoolkrkHPRvrMLs0AioZgAWhQTrs4FL4rVYy9PRPkrbHcMtPtyyGQZrnSx/asR7g2yQrKB8AAmyYd0ocp1fhW1FYB7kPUTUFeqAThaiW2zxGMEFtCkT/LUbHOHb+6JmS2l0Qu4cIYxgHgYOy/Bk98oTKdcOrfsOI43TyOcXc1lRm0rryKhyKO98rzmQWgNX/Vd4uysemxZYOT7V+ejVk0q5ax3RCqDOAzqbcu/TT/SbMRcPcv2q1+trjWGafVqpWMO7sPx/hDuxFLhV7Nqv47jC45+h3l6UVh/i/nXuq9JwxybzUNFDWSUKe7afD+0mLtDN+keKtaCaMFr+t3NH5k70JA0joZ0aisYOLsfQ+v//2ONnScTF1qke9KBZPYe5cu50bvcJzwMKPoexyZF1a3N9hqKu7Vd/LC7MLJoTN0xQaCh9NDxg//4p1Ur/QUJw6ygq3ezrwHPEn8VK/b/Efn30T8ykT1U9i+vaKDyO5Dos6/tTnmc0+81AVpSsn5oaDQiYxL+2EBmPvaM9CfOERB8rmJ92A22TP6KnpXTnW1QiGGPjP4lCig9kYtPgC7QiiOR9HDloiOlcqlY/F2qFbcPsQciHe4QIZFLZdvhCG/r+fpxG5wOVbCBY79Dm6uXOWKhw1+1EWhrhEHbF0GMWiNd9yumRVYIt6g4APs8IHup1uXMSf5IE4VHRXwcFOpAxhZ3Ve1oZRn4iQ4nc5wLgBN7HF1vwtC7aqBIyn4TWkfMTSYHfg8CGtDbyUUkOx8/B3l3BO4ObojxjdxbWtrklmlAb2jGcbl4eXVEpJ9uglQpJng7ABOs9/vJZ4yLHYuvvZ3036Z1CYOeJ1EI8RNfZCjhnWdr3ju3C3Je9dOeS3Q+EAOLJWtg79GkxpArHFFdVN36icuVyNKuaY74fch2bUcMqaXsBt4EfZwhCiu4ipIhfW1bShB/JRXiYQ1uIr9JtyLbxoCW9U2cAqqO1ZsS1Jak61BSGcJd8qSjhBcrFZ2JRxKqQI5vIRGnl2BTbh+wVWkD1nNStVgcxJnNaNaBtoQTmOP0Vq99e+XSqjoqXIFQq2W09lZGT3by50mXj3J/Vj1NPjMPc75CEXW0I5wYVu0SbkZfbjepUCb/PyeZcLMJVne0OqHbbzLIjnenz54ot1z4DgY+pQnmB92UfCjkU8GK5Rk5NwIbbO1BcXjWc7ztcnEB6XcHhB7aXYJZRCt2CmgenFgqFXPxzQnL7+D1gDMuPSj+LJIIvXHTzCw9bTs9DUcKDRrsCjKAUP5YeWL/TvLqi6Rc/Wt3Y1ETcLIdT17kvLXB+3aDL8LCif2ZZISm0K5uMiL4PSBEazL2Rf5ZMA1wmMvmra9mT6yEjiHNtOMLf/dm8h1pdgTzqZHIRw1OckRYPPR2eidmkHyehCt47qUrlenABUdKnnrO1BYZ8PlSKZTJPFBtvqOQ3BmwygnmXcPzFg07zYos1yj3e5Kx411bgX5A1cXAy6jMVYAwE2XJZjyGSibclPSyG3in3cxNISOgSxBWa2wq4+SupV3fzF8szjPm+j81GPp85wkC0KMd/FDBzpzMtVDjgOo4JRZth7ClTm8HAjsXjW/H6cCtFVbeXrcurgGTWX0myVs5H6vuKYD8e8MgtQv+BuxgzrJvCT2Ib4T2d0f3rEoj/PmBLttzYjZW44BmAK+dMmsHe09P+51xIB5vMh1D+0GDjbo4pY5qib9jFY/ppPUC7pEnY23JvzwQLfr+AmiUzV0N3KcWymRfD4hoVJ8OwCIOnjtIxMTliUVuJgBhRJry4i66QaEOoVtBKziv64dcUEplkmoWr07iJDx4fTEStm/KvXSlPHfkuNDSaM8aS5yHgyBHa84BBgR2f7KlxlHxFqZ2hzqcPA1yHvRXT1UHNVOblgaosQOcHCSdMOm5cOegOkMN8Yrmtqeckw1D2gFOlPayEkhmisv5CZKIAnGcH14ggws6n+9xWsVvWE6fuYMMwbvkWv1d8ASCaGVnQ+PW/Nj68Q9vdfFhwKU3L20qqkkWn7Of/vsrLD6HmvVdoh64cLSMYb0tsEnu5yHpD1ENzm0DcRQ+fgjJWP+KTvo5SFDxVUvRLxKDdgT+QTWVtXZWoFBp8Uq5lQgF74EhKs/ql2y3nEeA7DcoZs5Hgo1Hgh4R3Bqy2VX1pVDUitAOb8a3Kp7OUly8WyEs5OiLc1RROJoosw5sS3IBzvvTm3YEzz4+uwC3wJtNMZ86oiNt4wPcWMrPlXtgUJTXS/63YPymHKOyisCDbpLZJQfkXPWrpM39sf8sJGdg2+VZtnFYA9yFyBo2yZzY597GzNEcVaOnOADOlF98d+DOgRyayntCCl7LXbrh+nJxep8R780eo2l4u95VOhuHJadqH7Gd42xOdTgqE3Py9GWgouK5x8mAPuqRwC4djaFF8rqcpCvTSbM1tXMRd22T9VRW0354TrQg6gxOVuoVbuSX9KUAJv8hbiENyAKCyDs7mtOpf89PHvT+LdHYDyLMHjDlRODjxE6/Tf0a31bO9PKH1gG7+HYyQarxJobw+zeFTCwidkNjzFIdtFcVaydeG/ckVlSKBsTqw2n2IkTIozbt5fVsTW+3t+fnoAv3DmvDVTkiF64SRGratnf3sNJoLpU/SuWdf5KJE5OsgUZRX7rNhvzzHBzcj/TKKsm1kId4vmd5SJbvvETc5bnyfmIeKrdda1ZinKZ7IsKe62gZDlPA1OYDboTyLfNGdQmfQ2L6Ps0tAmiX3WB8NNb0yP4EuOQzJS2hafXgLeUt+S3qJMP/EfCUCeqNDeJDX9f4ASni6zoaCyrXPAjS+YGvHKJVM8mR5cd6z8NmqVSB0I71ZAtlDPmsSzOSo0IrlI1MAMOJdZISt/l92su/9TVpXWUqxeRLmCHSvioHxvx4iecTQCCtuuEPQybpH2tEJGILTGRFzAvUwmu3BaW2N7rt2hh9sxkPd9vaE8YQ6oT4RZFMxg5/EMF2/HWI196EhT9m3szVJLj58bZAU9TssWxs6mPedJESuLsQAiLBfU3sRY8aoX87OjOCwhvpjsD2M1ausRem+7+d6Dh7lkysvbSHQYBMHlH/qYQa3Jj3KPOXC75M1cCy4MDLn5Q+yPPqq+bkQ98FmO12jSp9EMqE64MUnyhW7ncRxWA5j0bpxVQKyJO0S96ZtpFwiJONEPG4zMZuW7NVr1VseAxqvm2U3Q7xB7Pwlaifb3hMrwyRDgdOYI6ErMqoeJWO1fONDMpr4zBbF3bLKcqfq8ZGjDWmesfdtTW8dn/wpR5/RYmt4BEHAytt+B8a4XvDeUhZJMJYr5WOtW5P6TszZRyEFrvQz42OcW3TRNo4qJYY6Ij9OU+9sv91v9v3f/0miJC8g4SQyerEuMnBX6AlOOTEX6NCID8txkKmkIB7BGGNNqD30qi4Gb1of487b91B5+3MLaw7eKrNXi/WPpPpdgB9pGVSaAAnuFmugdkiGWx4ccKTwmcE06TyYRj/2uNk4dfhJMbzwPx7dWETo1EfcE6NV1flqBEeLvyZp+LErF/E2hiO5wJEiK4rbUhx6nuqA74kaeGvDhGgHqf1QGdrN415medr/vInoKNokpLrBpGpMZhEsUSaDgHn/29Z7wwk+grKLgjlGP7Tl8RRpq24dF9dXB40rEL4eO7U3RRMG5QITPJ/zDwECzPjmki52GqxKz7FKPxy0JuyQNNVxVoulWUAC2QlvjxDQ1Ht7soiFEt4CsI2PZbVfbUp9BZ2Xz3fgWt8z+9JOwbymIlRpYPSV/CEYMY7wsGVntioFpzTFBNId1mr3k4hF0Bwj+xDdiix8jU8z2tDDFF8HVN6QMs2qWnTOEWchO8+kJGkvNmYK30xsDVRAZ2m2sP1dUGk5ptLI+WQkkTJ88tVylzdwu0GfnJQThBdSPdTO1T2Ec+0flhloKMMEjtk/MYcmagV6zPPzx4rTc3M4xFsmS7Dfeiw2W1fAs5J/15nXJLwZHMj6GKEcWL0kpHHVjFxM11x2bfSnPoMGoRd405U/48HZ2MTeUTJ/1vQWxtPh748KIINExHfSqP9urlbnwbw8QLV7t01+i3V5PYwjEDysChQX5TNW+asg9EKWnv5uIcmhkTHbMAxMfBEeXIt7khcBQFr/29Wv8tvFS1XQ9mzwEQNGY4eAzAjIfqe1yTYbHCbqSQx26wuh7I82+RKm6dhOo7ZeCiRf/n2+tZeeJ95lSGdF0PiESgXm7tmo3Yq4KCHdygf+7gqDoo/tYqYYnpfuJjjXS+hxDxRct9TPnAhvEKPH5dfbGr4kMyYWBGe6mkM0Qv/xX8NLN9O26Qjdkesaza+P1TlmdW6PallTxJb5nwQQwiDPfG9+ASuy3Lk3rnixygoAOc6r8hS0ti/bzJdw7GbqR4NiJW3ki8P8b70TKGajwFQA32xid4L63ua4MnheR8cAB46LaaiydLrzYW6eGngHG5dBb+vucwQ5MGSyKVMYhbjjeWZu5/hfqezZVnK9oUHYKBrDmq3gjRs/UKSUscItGGtsbXOzbX6KMjfRSB5ZGWZWgJgCFlTgRBTaUjDVMsVM/L4Ijhh01VeXBCmn03FZVRZQ589zN5YXboW7KEasfGxGh038dPeMm2bl5zQffionZHc7UPjKZ+By1iXGDUTRZNuM5X3ByB1QDTHZcBRPSIDQN5V+E7XVsRbdRRs5OYG1MC2hR2N6/JETEswZbGUOHT3eJ9SRT2vGByetvJnAdPTcKRJQY1GCdBMl+Hj/N5At8JmJ6fA3/2KNVXiZoE1FdHYffXLVH7UCebrSazivz4cgVLLDsovkWJvnVj7uc1Mazf1Bi5ex+FDzemM9ZCfI5BJLjMA2qExrGVoorrOzJ+4dCXOWr/BuNRo/WIntCrMdtq4muhUDn0ZTX8cxOqrZ6pAhCIagEE1Fu44K46Pd9Ysxaps9FiEzmtR1aE/IjrFpg8WyYWD1cjtAGw4L7qtnZ6qLCrkXwBweMn28GqTPPfWIaLGBAMt0uqtXMADdAMUyEDNS8D0cOFexoGbgiGt07vMgIV2NzELCxhVcDB6rt6gU4P1SBFGbgKim8aS8GwY47rfOur7SheketmbJT/GG7Pdk6gtjnjKXbFC+J6AhcV3wS3hM8RnYg3TfIcjSFQg9S+Y8tww7eBfdqLTmwc9EYYZrU6vSx2yJuCZEaHKlfM6Vlq91P6vp2sz+SV1igZuwhyd7p5YGHm3DhZMkS+K7/RgJBDmnpTCo2k6YMLv/P0bjdLpGtMAzRjNN00Tle70zoqIFyghugrmQMmpgEWTzw10McKaQSP0qzXLd349NUHjn0n/t1rrX6gJotPAUyBhta82p+3rNMroklqMeR+PJrLHNg6pxhmld/faBaBKpU662N9mK9WbFfC3NY5SPxpTZCgne8nblJ/URQ7thMXsbUq1iGiXDpJGUyE/4hzp/OX4xb5HUl7i/2j4f2KOUStbJGKEEL1EORS7/vDycVwM77zNecxElRf4KOQLNaEQLvb9ZzgUlbDl11dQJhWt4rwBPFq/INgQXr/i/+SGUNX9rwmM22X+FcaWOSvKtxcH8+TyIYVDn9EtJbKfuf1uhVJKoHMWtWJrOjC/rAVI/4ka5AKBtokpWmHFdkOLicuXYQ2SR/iEscwQdWCbWA1L8KkVQPVPsamsDa3MeLI1byi7w+xTxzEwbgxE2K3yfS2d2nHNVo+AzO+G2Z1R2mp2mbhAKK8feKSMtNQTdPqLHi538FBefvlPacXMKDwfHzxNaM4fb3tgCv5vQG35QMgCx3cxra/uccPwQX8L+fnP3pNo/CcVOAQk1vyOSM0Nm85CjGkA6smNwXk4zzjxhDp8q92rXqifa/x1rh9qmAJn4n6XRS9ZSQewajqBkidZBBobWB3hJNf6jAsb1c8WCOo85pvei8mwy31jS9pmMuoJiLBL9NXsvcsAWWDsq5t/nzXQ5FJJaaGQD2BPzxjGSUr47MP2luOpce9aBvbdXycHre12CzUkl1tpZ3resj2wmazMlMdP4YF3gokx8sR+TvpAZmFBhfKaeEt+BCh/GAlwZda4jEpiZhDeuV6NqQI6c3Jf73squPopuN3bibkcOUEJMtoshdYfbfQgrSdMURpFfeSyJAK5Mvm5CrlUiQWdkSbMN2NKAgzQl/KtIIQwNhR8W6cVrjevhQSue/qBYxZu7VU4bqmNDKOTfZAp7ud2TVDUtP+ZvuHC6V7pyvFbHRr6uMkohpgxGkVa7GrxXisrJ80JNCCblZPByiFND52/67qZAeudQCgCN66AKJ0D6ToTrBByzFbGnHHIbPDxVMtkrfjX0Awxtysft5wauC7LG4zFyNe+Cuk/1CzeuoTeDf7oCjgzDuM6+vC5pGk1tJZQJd/lfTDTVTnTNOungK1gtAhtT1XSWhAgiilaLmRDiLZCdQuK6iUhmA9Qr/NkBG9U7s8pcQ7i0J/Nn4i7F2gjIlFjjuyg08TnwRign2YIqSXXqUkA57lhKlKqZebKDx3OFB1uOZ1uFwp0i6jBv01TeMvNxz6cgy/VkGLAdXEsQoEtlWZlL+aRdr6t/6+FMguA/OUn3WuqAQ09nmsar6Re73bxAAz9/+skV5LYL3iP2vn8MD2oMXEaX3SI9mSvtNxngQ6ydviqM3cSu2AOdKkZTAXTGGKuWRabgVECFWYl1pF7dqVkC0r2gqyVKqRY/3RpU3ut4hikuIVfzpQ03fwc7zTpCu7scjtfp7lEbe4ZSe7AVMZ8F0m6UcfIfcPdpfsqTWGrKMeZmKhB4ARyyYILRi8E7tsTGa52q2lHw6FXYgVp41VO6AEwTzhzXnV2UL7VvYFwLPf31uzxKUgCuwt05jzDvowf0JqWp33rbDovMlixC6aVpFil+K0ZRxT1/aB1CocLsDSI/U6b0vRALLKMVq4WmSdaov16tBP3ClcORo48KGokJi0GHiyCQwSSSQWN9gWGiLoFVr5CrFxFnZjDzAETZ8gtonH7867RlCwm2/ZL28Bqh7aHWKH16HjlqbZMVuCOFzgBwY3rVXR5nI74IzlmWNw4aRutzabr8D+NJc61Ebk7FP/N96nKXrIq7GTOqABaYMyigdq3/u1Br8/xSL/EYpLoxRaiKTRSjVq+T0mIiweRnaYAxOD/6uxGiLDZtx3j15d6W0oSOTtbcl8+UJbZgtf/EBoOKhiTugJh3QxXQWjnphiOUgOtUpU+E035RORo7KvJGz/vPhspXYjlZLBnz9HxOk/quEIJ9BjwTvUY1Tqdys9THW5XS8LwdwBeTJljsXOumpP5h/SM4ig3H4wAjZzVnvoABLYXWFCMgTx6O+6CT2IToWajW2Nu13nKQSW3ot5Kuz+7ezhTeEi7mllajyehCCYJW/lGgRmZaBH1AwMhyIazQO+St6IgONrV3bvWlCPxY9dbZVwqf7ofzeXTXqQpd2g62e3pIMrJDnJmvvlOy6IjuzLj++EFm1Ka4/RlV53BCskGSqk9wCEy3VYWs1y71rFjp5iE8MbCIKBEAEfcCAhFqRciMNhoE8kRb2rYij8zwb9kqn9kz489YdHiYlYm/e5Rw6ewnuCLpbZVlgAUmtyPKZcr3uG/9FDum3Ztqzp3VeD3kRMRBDCikt7fvAwkcNBtsUM1AaivSsZMmzovrLGy60GbRO3PUjF9hf64E6tWio/lkbVqLv3u7oxfiV3gV+tR35wJX4oYRQmYszvt+nifgHKjd0aedcfMmnfyjA+8cfs8PEm64VmEfb3AUEt0UNMZxwa2kJhQJlotxhtRFv2lUT1RRRVYTqdRI1LDXUnii0NKrqFbfs1y+AnTBtgmgNxZMhcXz3xndJtJOxRnjZtfxFKpuK4YGBCxnBJv5JtxgkILvsChd0UlPGDQwv67ZOxHRa78iG2d8BCG16+6zjL3+pd+Q8COMvNYUCZ1W1KDOBX5CXrJurh97HloUFITElgNF+bETURz/rzez2zAIf7y6sKMcHVgx4XvWhzD23WN8aWJ+MpKeBI73pNAzjSSvmf0UqgoHWdK3JcTv1QoX3z9FLEW7Os3h8ozyDp3URP9FjW6xfP4iEfbagxCierdYtgTFqtGMTfJ7fY6h+yqo8BaSpyWZ0/BjL2rpfJVHRRWRgXqUx1Nj3NkDBj00tZIJDgwMeHqpRGvy2x/Rm6dCICZvV4LAwR3GeinJtbXNHWlh25A63rWfJZdBrBZn404t0YYXShlEqueJciI+MlCS5njKD+ydX3mB+SGvnu6657ndpySjTkkcAEhcaYOSkzhLdmhr9dtDSAmximtmoJDjOO0iDgg1WQKzexhGyrlJrGKTyTFPHmC5bFnmKU1TcXUACjep11yeFMFnSn9VTR2kvF9DGCb9Ym1R+BjwVabXnBBa3Gb6StCH5eJ95BGDohsMbQtzPk3/aBKusbzOXWNgNYj8kXz1++E6sviv/utE37UiVS1kW9yaVQUr3vlfMUjE6jFX/4Nc08AMZOUFrwhf/6LeJWV0SLUSu2ansgRA5Xu8O6ijJOL0EWbskY4mf3voB3zFsDBiOGfGvweGxgEst+Xz0b2+uUTDFTvs2H39oayaHAHTOvv2Pd6Odj4nJ0Xtgqdn5y/Uv+3IHEjKRs6En/vw3pbAmzWcWAKGAdPdK3y+9WF3QIzl8nCoVtREs84pW7H0h5aI4QJzEAZ1cksRyC/LX8SrjZaSQoT2c1cyYEalbHdHjMwW/P1+Q9PnvehMxlbRhcqioobOJD6REYQoHN6T7MDMIVpAozx4hUkuFizisAokMCaUeGDCEYe/bmmf4UmJxPcKp1RdGOAsroIUwAt+WK/eVD3hD5oD+76eWHubi0jieWygW+5KtJCWcEctXAEl8GJbiJoef8EdYVQYZ5Z7Q19GfcC3H4HisdtDVKZ8CdhiQSA686jhDVc1UFvKX5rk8pdbWjEtd0Ztrn5eEEeD3LE/hnyw/PQCuKDIQ3JzC3Xo/n8BerdvlVcsVvnVnf8ev61bKCYo/jSFBrFOJhiwABQ8i+kGUi9GwTQYlgn7YKwGeLRBGFtim7OkpiXFQt/v/5KeEcbnm9OX9MjuUaihHo/omwCYdB2aHRMYhtNce38ln2IMwCWUSrj5z8eQ5WcSiq8JLOPPUT4kTvWT+rgX+/pHpqz+0LRoQzWNnFAbc1EiSQ8+kpu9r4/FaGNUDky2Ei4jYFXRiU1KdLc5MaWdWVz5g1/ru7+bW6Y0tkuOYr5trzJR9GTEx+Y467tvOBfg5CuDV/qxB1nGYztkIMEvU8HZMuQNiMJgLacruTlqwjy8Sd3jXDJdu1N1nT9GM1Eh++/lZaHIml8bzAaLE0GUyzEGDYwIc4RgniymBzDBy+jK6QiP2FvKP3E345H01+UHQE0w8N0TieogGs0ooV8qKx3cqF5ZppFmKu+iKtNyZ2pojfkQANwvGQMH72H676toIg3iPGH+R4j36mMrOxsbgCXNlaiT6HReX/w7JExQMS9aQflyp7xxAa9TDaQLSZNfcZH8dC9StXTbUr0sDra7C83Gr4zhEwqh0lRT9R1JBZQdMLnz65Ndg9bNsm3FBLaiJghqbSFdsKMRaQBNjvu50zR2ck9ANFnbXtqKv8cpthztvGWMt675iNwmNpa2aiF9CxjCEAWVA8KY4NrqAGRc7bPUVuuEgwkjXJyrYtm6Mqby2cAPrgm2XacN2L467JfbTCmBtr4bKVxMtielKmdDcYPFaT+yvpaeb9G2oAzxvrTEJQhZXZSFelKn5vIQ4/6ROwBanAlZjMG5PJtDJ55MdiHPFs9vCnHUxMYjgFDk7DSZ0CyfUEKMzS0wkylacC6M2e9ZL06VRxSDQ0FMtI8fxiL5fmbkE7Mxol/M7UT52D2HLSYTscXzWbm/IMwSJTA0BYZkCRIqtae2JyJ8fONTX2sfYqXOvzIh+7zRj7ooc300Oe0NpvPWvADG/HMbNrwljRQnQXj+R0yLXV6QpzNz7Q+0oR8GA4F3Hs5hBPtZrY7b4ys8RJBCcI2O5rUOXYhFGnVl
`pragma protect end_data_block
`pragma protect digest_block
8a3714f26c1601db3a121b73aeec03414942acc4b47f15951b9fe4de9055b416
`pragma protect end_digest_block
`pragma protect end_protected
