`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
TWVKphSDTy1DrpRUfJo0nXFD5hhy+uzjnoenNVM5WCRQwYFhGRNIq0OrdkduS+GeV7xRnWKPEao7qn6G3HQsTYr1mA1URKayA3CfHA5Tm+RTOxemwKAqrStdguAVOYuPqwOQYaIE2tmf+8T9WcEWR+2I1oU3BasMonee8ZcWn1AXcbtmT/rs56iZAre+7ZGAOiJIsPJ14wU6N+mbJev9PQQDuHwDztapysczVDCf1cXUlUxGPI16WlukBE7MNvuFIpU/Xpxaj0euGWwYK/7HuZSd+j5FkOJGqXkIadvLP08sz8mqlBM9p4sY97f//wZ49WquvQ/U5paMxVLGgpJ7ktVbLg2qiO0bDMkN26FixFUcrvrdfUuT+z9pj4YcNgrTA/NKTlXbOMvRhhCJ1XSulrXrjUqKIq7rSgDJdnvgMAPFW13+xLaPyFCpRgqUP/jX7ekkgdJ7xM1YZzkHPRATDhHat88jE0/ThCmPqWKyB83WGjlsA0vV+EPrEXyUcugZyxLTjxF308YEkjgpdeuECgEhGTdM9nozhs8YnkgmKCPWsOf8hlZ3BkB+gh5z8Y/H+f7d6qel6NjsTZ2cC4/S2sIpMeLNjNsZnRUHrra18DU6m2fokdv6rK46VR3kEjqGL3qCiKfyxs9ianah1+c5t9JC0J/d4EsS7WPK72hDcYuBG2UfA/YnjEtcHXjWPosjyqdbYjQLJ0HaG6y6WiFNtLlLxfyCMi3AR403QW1tCD6qElEeyvwAskZ/YvpO3ASdYin7Fu3yjFwbO7eQAHuxzy14NVAyIGa+7qyTGpjfoklVMMkISTNp8ygZAwg7dmivG/0M5/eaui+YWGVO6OFuRvLlCkE+sLDBSbv16N3tKzAh+OrhjKVLzn/zX/4TkKkAyXJt6JLNO3B6KFT2KTJV/1dYqFouyKvmqcq6f6WIYHtQVuvANBpvencOTiGrNBh/UJfGx0kRr+AEg/pKPcOZxhFK7/wHg5I4POERZcgaglEqc5W4DCzPTqpw07utCs4yP3DvQUHq/eAI7NbtvnJCFR5y7WFb1kSGAJmA6kR2nDKeDreV27e56uPHNfGuszofuDCUxJmW2CfG6K4mhSKFvYFgEQP210dMs8UFgE/e/5LZEXHEVkW8MI1MNM8fUsxrlB7U6gzeVDj0n6GLdz39aZgNsQS69eY0CG2Ow0y1fTsAsfPOwt15hMV0+AvT/KKsFUdd8GzS9i0OAj0pkDQ4/IKosHFC+pBKrAKLWzU2rH86PeaRPH4KXEI6LdKwd+3FaM+xxwgbtNektqUiVnBR673IrQUxKL1XWHO89X0JAuZ8JvPdibUK/9cVLy2nMjI4msrMUiLPrFMBmQq9F0BpxHItoIpYwNuLiNuoNyezo+c9nHgs/CMRaaCKXNP1yL1vbfaY5NRXy57ptT2Z3CgA0n80ssrj680AlbcOE7yMTUWG/ufm+gdHjEkTPJoLxz3kRbXqhtJXPo4XG07sE8yZ5tuTZ/qIPYr7xEci36QRSJMlU403rKgmDQQaN5N8gVjy01MiKstMlrQFJvWgQ2Jazpcor/cU+p++g/4UQBUEu3HjNezZ87xkhqNdovRMopkspv10veJ25iIvW5GjuvkvO+oAtiRl8gaZWsyu1ItahRNejGyMVhSWHL4AczErRFcM+P+aW/Lx/31rtbWhx+giNRsS8zup9+li7xr8ftPxDtZeO7q+AWj0P9AfBHhDOU/LXAJDf5aCKP+UASlSBrZtY+7QL09n1Df9Motnr68ssLCyGGQAZeroS+JEUEFVvq+W/UVIDeXKzPCsISAPxTnNzwn57LuP84akz1PSiMulpBpq9jkjV1/14gx5Uc5Hh4najOyVPg3pWHI3Wu3+7KE6LJq1rrK8gErRAFqTeGB+jDRESTmdk9kb5KzBhZLFUKjIzX1vGI7pAUhSKWtv0+68jA8N8ce7ikMT7WkeX1+6gK8hdziDBYtrYfOItyS8oqym8SDDi+HMGC4c0+JQQobWzPJNV2Dj2tZvtHSoXWI4edwH1JUxzrXW+SnON4UIG2HgLNJUozSZHiV3gfTQQ7tHEWaYcbjp8S7EbIK9eJX+zdvX1F4joOAt2M2c3X8yaQtYYBdL5j7CQHAPEg5a5lP9iH0oFMx6KOqekaZHgsvX355LqfDgg9zowYPf0UDRo3TK7ogg3cH39HEjjfTPT2dFEduluUrD+GWUAZ+Knd1mxJnZ3oZKMTj+n+nvcNtQSxCpoGIrV8kkdpUpVIh6c6tUkNV0sbmC8aImbjY3vyKRy5aT3eJSShMP0vYSiQEmgtzl3TBM7qVLdNQliQnPUrXfR5aFbo/F4hC7rKq5OQ4AjfT/AoelTuAAv/56KwtJ+PvmkogMBvPb3BUJd/nZNFSjJ+Z3CVQd9/SJsrho9xcnsFRB//5c/lnF2Kx2UmuYFIfNVUI4LDTq9tFjJ3pQisgK/k30Ro3V5e6nukU0ZyzSciFxqLT7TInFEg0FnwmnXBjxREDyjIMNi/oILQ7stUxlQHQxJXaJCmHPAHWIlmzY19HNbTMUlru1gFRi5xU4rJiRCd6KwPs8KYdnE/94Xlo6Ddx4c4NFJWe+grGPAtSS5MW2pa/cMh18G6Ed3XpQ2pq4Iv0LNHnq0C/ULWmHj3+M5SER6RHx3CjMcQP6r/y3+sqf97B219qjFDw/rpJtVrhliDDQGoHtNYcWIf4LBysJfbArGKGi80xm93o4Z2RmFo44ZFQuAFQay6ZjzssXYaj5rnzgMskHE9YBexg0Z/FKbIYfV/Y1SLC1QyPJFDP9jbC1a1TEgUyzQId63DzpuFIddfeosI1ExJsiYFmwG9o0PqpOSsmEjxhPTLR0g4Tj5nvtXJgF0GyuNAo1M7oB/DWTmwxGnf61ApOeXVwfFvBrrh3R5TkGT/GguOjHfFywIInO4mJSLiEdiLwt8lXHvEdmTUUutjcQPxmbs9ANM4nQwRS+nyug13cad10VoW14oDeLigJqJ3yp3sgb/vx8LL7nCgfHm0aI6hBk1EhiJ/VLC8kosSJJogDVU5jjRlr+8yp/DWEResSiP8kijcpZuZydJQh3IheEWdaBE9+XoCTazPvMjOP8KVX5n3ePLyr3nBt42BRfrppTNQXm5P+ovaeQsxtT2bBoQkeedtNoEe3EyYTYRSapD3OeCwzR0KMpgEfORXHghzdij1TnO6FP0/yrfjLAjqjh5hDVb8alrJxB0p0HQjqBMIfJOUDJje6tKPouXdOsHToK/FvWBBcqFyLMYbCHliS1LrwVWYIqyKmeoSM65SXJmOQdFIyBzfBaqJo2k3iHKdD0PKCa7reyp0AZEuyPD8lydGANqQPyVYpxVpBaBfAEz9nbrwOJQy1WIdxLNuaBsZ81XkpPZTQ4KPIR3Z6ztDtdmOb1+fzPTtlB6OzgUhHlfbQ8bHSaCCpnGwsPw9iUIa5zAc8Wll/XXzcLvhv0Z+dTgP7WHnqu7Evn4nxmMp7wmWc9Hv58L4WgI3gU6q/6BsgFVYH0MBlruoN+LP0ob4rznM6ZhmczFCDzs+k3EftakGVgXoKiPQUMry5UWwft3cYFP3I2MS6rI81GqJPaV4Ko4a4FNsCsVMpHVIMF08w//32pEf1AiE/MXsujERR9bef+DLjo6xR1LvsWMtcI+SqGX8dlO02NYW6wi/fKSBhiTx0+2JJs4xf2ajX5dxXz+FDUVre5M/oPmi4Bdi0jk3hklEDxzzycg2lAKjl1YSrArsj4ggdHDBzvAL6I7FZLE8WaBPb4cak7FoDKrhTnlMPCyZ2CK4I+lLkAShCGs9ms9smAiWHlH+2ZHm3CrVFGcGjV24Q96TiE4IOuwK5QEBVhp3q3QjNX2Rkbd7y4zBkpoE3yfwvWogaTd68WcKPuiPOQW90jvdaKa7YgedlxsiH9BdHJCwNvq2qSRkrTXk5gBz9Mw25QnAtE7bBgoIzGJNsDNpsLjBKJEJUooBXd0aXlBoXwCYNgpGbbiBveaPPqLNNdsr0b/Ig18Lr76HtbupSRFTibzYYLVLVSdhxYv+4rW46KNOyrov4fKx/diR0AbaW5/sd2grudzYNKZlTu4O/Q9eJ/qATZrHli9uWR6czaM7cQroPBZO3iDtFcEHndIuyqO9OY2Qxn7tEvJmVx7ODW6xGHMwQ7r6vVaBMClsSvxHxMrdOdv+VXRUQLSv1HcfId97LfzpWiqHaHhkn1q+Oi30NIuzcG+BKS3cNm5ZjpU7R5/yY4ULLEKwRjV17892Ne3KOTGpuQsVp9a+tIW2kK9EDSCJFF7Oe7FJaJ8ad/YM74A2mkmgWpro8pMWPkngfbn9De8/wWY0bCHyxFGoFUcWMExptDmSIfCg7uozWxgp6AeX5kUOGxeD+Q1EupAG0Sgk4JEmBn+7s1qXNa84RgWO5hmulyH01SUgj9HJgnSEwirqSg8zLcdk8jkAdBrnupWJ0EyNTGVk2XPcEM0N5yIVe2elaShRjkMJhRkvOGghQPsla5maBjIszUpcqV3O39HIxx9QzT4oOrj1q/E2Mf6kXktWrAKJrrNgGJjvGP+NGf80US3ulPMbO9kaNS9X8F0A3rYyVdmnhRQlpiHOwf6O1atqK6QRu7mCKhGY+jVm49wFR4oIlFWioyoSoWlELRTKGMrpQ1mCK6TChjvQU1aIz+PbQtvem4YUhS5OdsQVnCPBhjA3QwKd/jBH0KMbacxfBFSaWVwwE4righdze6CgvzpjDIaG0gwJsjkyBvnea/SSF8/UmjRhh1wVid9ol0lVHa0nlxpHXY2EplH67UzPycolxUPXjengUNX2oEwg0LKrdo0IIzRaL6NpRfF2rQVDOuG7iYRN3KnNIuht+PeJVtfPl0+yNzdNaOMJdT6XkNKMthx4qnln/rBcJ9468Ic8UEDln30NplJLXxUACkWlvZmdTzHtDqSc9EErSUYs0PCGsCMFKHnLRY6+T7Qit9opamvn6uheg60JtGIz+bYTxgs0LLNBpf3VnbFiJhtxflQEuYO/sZG/btEuL1c/rit5ZKmP82AGwJoM39RrTvlNZnuKE641XqQ7LA6JfJcu6iwHxRPVGLd1hkPeneI7j+zDgd/Dh6yrzOxGXBEErY+S4LTGwA1KXA0yY24EcYBNvjYymu0gajJvzjp/MEIGXDMhH9cZ4bE5VjsawCBbFwvvb5QIW/83Uj8jweAqMWT6/7oeBE7yKfLtgsVySbXIJkLOhdATfCRtt10J7fYQFkkTMLfRiEhy2+ihaHfLpvXY8BLPdvXwUcnNRJf3wX6KlGPefY/BZCaVUeeGxMYsPv5+oF+sQNKmaPGVKhzxOWwpZp7TVqLqi05VnvbN8dB2y7OaL5LEk9UBjCzJCdcTL6MQFx59kw0au//HkJqvwpkwExgmfOA5IZSBJKUi1GZQzTJnbBx7M+b3hJMaFyEKcR8D8V470CAtK6rfG+NGH2+EJ9Hh2NhQ2aBfsHfSbcmv1qhHMyX1LIVO58JwMnYxWxUis5YijFhpwLDf8QNTP0xRBhJvQRcuN7orNVaF1AQ8ZdfmI8sh24sGk1AXQ/+BTVxK0BjJVV+olacqw2db1S472NpykBCUGCSW8Ob0z586IyNES4/HKo77+UrIwZG4NZK9GwkjOvPoH5R0NqbMzXlDlEmDbuRBsBw/cq8EuigAezs3rf7Z04raLfyBFzmg0IAZdhM1pGXtkGb2UeiquLloAv+biQfv9xJICF446ew7zTBL50A6YdD8faiEY2JsIGCqmH+vEdFiALfwsZ+BlgkcmqUUWzLUyOuWaEoSj0d1hBrrKZGXVqqCmiX6Cbx269L14JosOk4hsOovdi4uIlSaM0BXhKrAdLtdwEIkYQEQqDgS3K8ElXSWbep//NEjlNSdSlPokF4MmKetggRFvt9GkhvBNvgjqz7fBX1ivcB1r09vL0SqHgRPqrVCmy1ghlOI2Nbjdqx7sIClNCZDNjETUNqbtc65KMxB/G77A6I2bkw6LsX6Bn3Ovyhs50dxl2HLSa3qEI2CX9xgLQP/JhkpM9N2SByTSWIwG0kS7xNrIsppLZPjaj90VBXwWj3ZNDKxMV0HOm9IZc5c1o2iiCK2zwl1KLhuaaylaicFJ0EV6/HP9PNuBOf32tlUmE3tZp+Wi3HRZt4mr32yGY0srukS6neLeB7DqeQdTsfHwscrB8ico0PObmes2vW0X5S5qOosGS3NH18p/3G7EZ73RkToFI3aprw6kTYsZACXoZe4h2CV1PSW3mvqAM961nz0QQ9+D5C4MAQXh+vw34qOkajUrbnZwSXdVPLy+tobePljc/7nkhOzrcfyRYUGNLZQb6jmu+wF8cL15lfZ5QtKmkSZKklP9HjpZX8y76PcJL4sflvGAr4TS4SfQ7zSU3Im68X4DBrEULGp0NW8KElUlKE6w5qbwYc2n473uMkvpAhPP7aIxdoecloyfWda+G4MStL/h97rRFcPFEYJcxYjqf6UFUuxupovmkFWDt9ogV/a7maFMyvIk6eCrY9pxaNREj13ZeahQ9K2syU17ynpPVfbrMvvG2fGT57XTQSSPWq5p/+HA3JieQ84OqGx+hbb9t9cw/+cR3+mKZ6bACsMr0jjj1//Z1liH0m3thuuCK5QBnUs7dfTh1jsDBJubJCHBUfNWfyHAg30csrOixt4X2BDyP+CwSX3Hhhcto9sfjiuKRIjNvP31t2bdQUVvyLlj3VwszytRhZ9CPv35Ykq4bOhT8q1L4772rvXcXsLrwk/Uc/9HU9oDn7HUMl2ySIPOnOvDLFYBS1AAr9axdG3TGCKR1Q6179sQInZGinabU/BKt5/p1Ff7DD8hnXpAs/EuwARXrQnDYaFJc5RtLIhlalFnfsGAkuHGETzoet80/pccoiKj1EHvUV3qclWpzsjGiYKrJ1Sc3hIGSEIoaz+R9C4GOSkKvd8/rs2r7b6Qzbd6i4iEZITAhJ6fkhJqznerkMuhH470LX3q8HhqRRT2xzCBlgBV9ipCeNzjhXduhMVoKk5ocZ3nLxCkZnYcZ2LN1ue+D1TYWUH5IRrrbqLyUK42OQOaiiJM2Sl89jZfU0PnE4iQwfRhZj+c6KxxUHJW3rl5NYKv6hr64vLssLrqd1X3impudGKWWC/OCgOsfH7uJy9UQIEcUsd94m1QgZy5fonoChHcj4u8F1F5+6TDv8CgQFVPlJNxfb6LvMwkuZFoDe1gKdHIT7orktNnriiEsv74YnPGS79ZZMsDsRtisBezb7PkIw1Lx6HOh9FBinRJBF5tdAuVHN4zJ7jxR5qrhHN47sHXmm8xBx9IDXSpGPZ6m57IfRvxUvowizxEIgA07v5SeyucEUM3DfXVOi92NPo4NoQxKCcUYE7vScthKDBEkD5J7GJ+FpksjfGMEvi1b0AF49fS7dFMTdRD8w048kG3eyH0PeZ8DpQREVVDqD2E2nELb0CzzrJ2XzPcCXtScqnC89U1wtkdrPeKJyg1WUc99LYtJijBZ8Qa06KeDwT3lBNGmXDt1w9A4sowq4KFO4NOvhTrQ2qSQhBJRy2x1j6Eyhsx1YIJYhuV1aTM+9xQUxngz6QQxxhXBMUOin0kRE1115jZxpsTsq+KL9ikmd/Xy1Z6z9rdpWK2Xuc3392pLLwFPjbvmdMlVfyIUIRNwYidsBigWutuLKU+oezSMOsT66hfGShsu7I3ObJXTejHRVR8BRxLLDHh3iXOZcYwpc2820it+9RIQa5PZItgVbzQkzkkYnK+cZH8FbQIQt1FyvwRxVEfAlPGvJOm7lPe0VThFng1+epOQLO28aLAg019NzNtLr+mWvzNj0NY4xGZfO6nrlTQMvaLbrHEqf6TcRsFmAK0a4dPj8ejT71Z/mLGDrV6YYzfH7qnAfbsL6uljIZNG94otAXBff27xR9JRamdbFotCFCXaX6QNiZHbTkUc8gxaz71UssqDXod+YTih1frppH9xEfiLG7MZ8/BZ+eblyKrEz3CpmSEEoQpFdLFxAT09FXsfZvebhtvnpr4p3KZzMFDC0eH1jhpWgT8UpzLfsHeHFLSBI1XXHohDrATTXelCE5zSOck36jKJVHuALL2vCjKDcP1w6pMdYyLEFbe1S9rAB2LpMol+lHTgGwpo3f9+afO1ZaWsgYHwoWYUp+VGGFtxQs0OeLd+vKsdFrzjlX5EyNPvx5Mwi1M2i1mzeXbltZqrqhD9CQATFdw9PBiYaqffahMwIvJ/srGcrUGdij8ic1RD0qheSdUwBMEnDNlFxLNflUPTTwTAe1pVU+VltSMVH42Bamt1ZvzijL0m9IGXuyLntz3/ykCtgh2iNKtJ/c97P2EnOXpGJWaQqWAOJ7Vx4PhkiUCJvTykiTxAUNSPMA2nIlHVt/22UDg8XRyQL8u/YCkNs1GuqXsAo2gBBdEm/t6n4XrJDVxBLQUX1FUWI75gvteKWDSnNT8b76EFdcfmFAgaxNuVZou0JgztDfib8ftycTmRrkJwqWEDT4JWfLa7ViowDD3XwR9yf+BEzWUyZJmMDLH9rftFPKX9V+AG/IlUBZFuKFFq8E6NUqTWXcDPVfypIIF/SKT4KWqkZVHIOMQAAWBXPElvQhW4rhFx4JkbpUr8KAArCHqZrfQS3LIr0pt4mgpPZRi4bveRaIITTuvq8OQA0LgrNKGlWdLdlZCNsF0a1JWoehU79CTPXlMPOf4w5RjrwohOVZ9NzZPaWFKCH9xfs03ivO+5V2z4c44fAbKrf1ipwROJXVx1RS9x4Lc6/iLjHDpRbKx6/lR5wwf262L3S8BfdXkffKhZMIu0CuEUhc0mn7lib8eeqVWE8MyyMuGIYZTvyTZM2te3A8LYPEwtyIIbt7ZpyepOY3E07eJMVCPbx2NE1WcXdkm1ugkknO8c/qwtYfrF97ZMGqxm/fKs5etoqcN55XWSDdbi4aNXSNN48I4e+QrMfWDM4P8D6IMvqAfxbM5AUBNyjtFbKlAx3Q/nlqkANUlCxAeg4eBJdBYFOZLh85al3xaVek1fD47/4D8kbMB0XByYQKljYmGHr0d2cOsZEvBgBUmI3D5JN3r48gCa3vjN8F16nvNIQ2UsItSMVTQBSgchNdodMiSERmTA6cHxnrOnhBgkDhZ+7ipO71cTKaZbTfoeCmDVX3Ux65mhqoBI57k3pqNlOgXOEHqvcV2D0by2yaXfjXDOqdmEIfy76i09H74od7kyP9DHQTsSXw3hBBre9npXuXnRWEacREO3VcomPwIK0UlR2IBchweP0Z89RacGUSz5vyvzlqTbzVY/sM/he3zv6WIOvaxlDQuuhi9SWGR6yj5N5JafvFdZ1twzDdNN+c98w/39QwNmIiMqu838UravygTtTXjbyYmSkNF4TumgeH2GONoiPXtfLPOILUDjyDNyjPS5Qg07h2zDEIgxp70FzuXFUQGQsTF6R1VzexZWwN2qag0LF8uil4XlxEz1eeS0guaIMxLdciZaf23C79TQnP4m1Ovsc0gLTrEp5sg960KHtBTFJpGnVM7gKv3tt6+qBLyvczevFJJbt9UwET7q5vFe/P6lcsIQ54Nltn2qa1dZ8zD76GI8i3VDcKD6ASdc6yjGU9KYsB4hy+xzm/H/Oy/WWU+qEGo9HAyUv62bcpOZ5DwPSUXb7HHVTbZRvef5+ZCRIktEkQiDeCeHbdi+sEO/G6ng508Vao/YkrJmvRGS53/PTngmv8XUfvbTv0IUGRhvD6CTqs4c388kpEgdNDLEppmjUj2WPVJi3CGo6Y/10y66jIsnfgov7c2k7OYP/EQ/QLGk8LJNdIrCKJMbGN4LDSblTWdSl4ufw37qhPiSbZaPbx98zhWH6O/CY8p3hpY4T7bE1sOf7tQ0XVMmhm0rBoQ06gYk6NlfJOAxFRcerVOALLTVPzLpDQ9aieA84DYn79gaL6MEWn0zGc/zEbqMukHj4m1uDzkTB1py2mDZt+jrBf33MB2gGvuQH7inftfSSCn76RadwqcIgCge70uNfDZOkwEQaeUEqr+0PtQ19l9Wp9T2Fz9aUvKdtQjvOY49oylmhOjr1KxhA62bnEyYVlWe7nixD/n3KwIzKDz0hJ/ERVA69GwJVWP1sp4jkUKh3CvR5P6asvHcSGwrcAuAxAaLT6k9oWkEg40hBZI47FpLvWJgG3hLXIix7rvOq2VfVYUV/no9JQWuAX4xy01FhJ1fG93hYCS9txKFgU4V0cYZsZEqrCbrOEIh5U7kwqOn0dagQz7U+GXZwVkd/pJ6Iz5h9KOdBtG/HzEUrC2PN4n245APLqdC03CExtHhariOG/Af79ISrlBsh9CvT1OWeC9gnfVgMZROHiw6YiowOnQKIjr86vpQzNXpNwr300veV0CBtw/jxjtlO2PFX6rq2JonzjPfmqhwyIuD3Xa8aaNxTtXCGoXLqyK1zq2LvVYQTa2Kj7c5n3qEM7HPufFwo4HHcn3IHeyHIWOp2GIlwKDAGR0nOBtDBW7Y8LKCaZOb1beG6Xw5R5AGFFTP1Xs98rOIl+PaWcNMb/a7yL3aX3jR1uK7/cFoFCKQhtqYRp2E8R1SMQePb9hAwG7nniyrRgugqcMewcwLIPmnzuOe/jaD9R4omq+q5eM4lLlsqBMMV9JSrtDa2OqRCXp1ztWTGgTV4u26X00KB0hAhwtFOfkGnYWb9mLr82XKuq5xdbRmVuKLbbzf5hUwZlR3IRFFmi8KD3vExsDHdUOZOLQhTgrirM10XG7s01k/sibLiwCcJgdzzcN1T5JgnHdO5wMhr23D5csmcsGxOKodckI+/8cqICxD+KEE7JCpjRmrHlV3sLaimqjZlnjNma+reVsfKGx0nIiNwvXzXZlThpw3eGF+9EEumwsLhhmujEqesP3bpfVwibsbDn7SuduyXWfCQuBRPpHJxK6ORW1o09O9rNawgKjjYSsgrL+UydByqc/2m3Wm69CvtfaBVRSxW9ILB25vuNVh6ZgQ6T9mR5cHWW40vR/R88Y6QHd6cu06nGw6HUS8pkVBTy1ZKsD3GqM+hjIwmf2j1DqdtcLzfxU35qHg9Z2dyiHOa/0/QliNM4CQSLzDT3hbyheVeuoknJs5547ZgPnPXvbgGN5YVVLEqaXo1uF4j5d1zKZljRqQSJFn09ZrM2ViLBpRzieh8imgeqIQ5ptcZZ9MKoOdsDoM6YNye88umh4RkbilyPRMQ1qiRVeooJA0nYniXyPorGWhHTaE+0KXWYvdL5AVhA5gsllJxxxCwvAt8WwMn1ZQHqzRYcoop43kR6VzqnXf278kDcKtfovMhAy7R+GHqEakjV0c7kqZShSKaop+NVdv/OfhPRZzfjdWBZYrR9WJM+pfEWOb+wdScauFAAgnpuy92jIv/M9e6PhCLM9hHPEAYRtWXGK6pjh1YDuJ3+2kWwMelAdyAtpbM3KowIlqbY2IYtXS4BuN70xxIcTAgY8ZkBaL37xNLSuJVD78/02PXehjMantfByMNOvtfQu/07XM+/qwd22CprLz4WrWENrzARYzhz6tMprCXCfFu1UtBKNz1hvIqAm6OkuRbomIcSQWy2CdNJRdd9NtJFC/LV+U7v03zo40g2uvvVfxZAe1fMedWBrEmUsjdv1cWBz2l0Lus3yn+1SPvKZ/JISNCzsZMCFIH6XW6yUnbxaZXY/BJCKeqm+PCrLTJpK7NUhbUAUo91FB79nRcCTC4cOkQqKft66ftl7Rqd4bzCSxZfPsl+JVTmpMi9KEsHU56dmnpy1bUu/BTVR9/SikSzvmCVaZzQTNkBMYL/weoNUjDdc1KXg+yPgo5y56XI4TErZ/9w5sUbpN1uFuT+xovBx68CxCUTscbOi6Un1Wf+7OxzWg+kRBZXsJFQgOno67Xtk96Z1RHITeqgBExOtI+iQ4px9FDUsB+Vos6pPWBu8TEd5F68gSyK4V3H1ZOZcnQYeFYOrnJbjyKY3En5ynbjq6+kjrc3eG0d6qUBvbSzkTvo7v0OA+luyd+SpOjH06XeDmjhfX7tJgYUY7mc6WftzSa3kqswMeVaGXq6R+uLIeMI21PCJ4t9oaloVo+dRW2pMK2ibgqpETIYs6xiDzhZIqB3HRsQxkWbh5BjdP+1zC5VKOI8Ntc5ijZTmgeZX2m2jSu9H7Nz7XIwmQ153+61OD+b04Uvwalkfx9vO/F2fxpXN4ewaq4jqfEIXhpqvdNhcIhYXSCXTgP74psxOABhpCc5xRJ7iEjJAH4shuNWEIbFx3YCI5Rgf7ow5N5czjNUGrLIEoLRKBMJ85lH5QfMhLyAp6sfTa7OX/vt1Hk3WZRkzEu85AO9ZRXnVWSU5rvwX+sWTcueoaLhWoF62YdiPm6oc8/WnRE1/KLunSECkZ6/xbFHh1vZp8Mn0/Mt6Mk/KAwbVpmbYxITdiKxgabXWYGRPP5VbEGX0ccZyKBnYpfMj0SZNj5ofbkj/6W5FeNVpXdK27FKerl1h+quV/oR1emeFZjbeaNfMJCumGruDqpdIZy6PcigBA0j0o6gb4v2SsgQ6xh4fk9gZ6tiJXlX35JY/z0Lpj2xbAHd1jBXK/eRPeY8ouRU6erS35AdWmPtQB7OnVr4IggS4jlpjiMrfqqigJQldXzNcUu61dj7bZct4IQchNGqEnuH0HkPjJ0O7wcNOMWBvcNdLJirD9BKTT53Al5tJ6TLJG3rIq4EOx+OPnc3xD346tCtqmtZko+h57w8aCf3JCdwo59A1vWJOcWhMQ4DVRUaUnMB0wqhGPUoIJpRrw56PETU+ShNdYIjb9edPUjMMK7BPIEFbcdmLLcXmvBw/6uaz4miO+VwzoF2NVxMCx/24OE5a0JTObfear1/E34NsA8ImjDrmT01JXMWfF/Z/8taDACYVnc7n7KV95tcm8mqXeAhfaPoc6QWy/8LNKOVCW2/W/HqHkOTLNyfJrEAFdd73XrK0AKAGPFattGTNGoJUCPGM/Smvi6bMP8rTujDDcBrAMvxavZiIVPP51Sqf/b0TyATlLKATZZzvTiLTzaCqZvit8N2va/2KOuwz4phkAMy2nArBPLTteesI1d6boChCwA3WB2H/WBkmFCXiVDf5Nl1Sqp5qq9wEDVAvu9/Ju7jQJ2yRvJAJ5tfNMTokFif22zPCMdxkIo12RhaEGcMdgZAlRpZXblrIoNSHexU84d9uc/t1oYnT/pH4xGXiEutLhySu1+CngqTmJkWfbN3LIX01+i6QaKyZcOtTRKs33FT/phWZKWOFf/YniJzy21s1TpLddvup8ZQWV3Nz5qUfu2iFCg0yW2t2M/U9MpCaDm/mnSv4NC4JEFj26KIo5lbkXR/5V4/Smq36tIH6sRWeUcgKp9ziywtcssIx2txJ4g42wqYoQ9zXzy2uLKDMiDXkoSR7HFqWlF+tHMRzATxu9/CZ5V6JetK0/wbL0S/eZ7L3x2dhPPtywCYT5qkjYfWZ/2g39WNyTeNbLzMl5Birt1dXi6zzFYSdoWqX+rSXJJla5H083zB32XToDJs1Z6S7ojyE50BPOR0FF26kq/q3YwO2YxB8DoeLjwOCzuPE1Wu1Ju5aU1LjTcG/Ag0ir77SDn/Silt6om0/zZmV2qmj/La7h7CBn6Tf4i3vda2/6Ios3UnsiTZp6UNqP/uttCvb7AIu5LJGgFWx1Y7iGjl/pi38KcMKXs6ATBC4d8bUCIFR5wKBThpPfhScQRaaqpbdwOweU5Cc0sP14Oih0/oGmBmzOcQbQFAGyUuQKMt8zlCLAlIIXmoLHvckEmYH1fgagxFtbBcJRaNkNgdS//CXNYMgGCFC5DrdsViJ0yU+YV/Bkc2BRmdP7IHbckos0CvH92F42Y8SxumERc2Iko9ySUfZ9+iYslAKDAI/4zTTL7hZJJydoJEK+S48rwwoj0eiOCnhrmgMvMazcWzM888ThNF3RHYWeFcw+iZg+DYp5ymCXiP6z9uesvKrBeTH2RiW9vN23rmheA7wvG219H+I0qv66ujjCXZkdTzd7Bp5wo7y0noFDv7PjJnJ4Q7ejuJb1P3/tPm+eiFjnZOW7xo5MALg6ebKtk1yM++9iPtKaqrTi7HnUzxwq6gcd3ne2KFhBrliRMR9hdoFu5qH7xnWmcz1+H62EsscI3NNz/vRKPdRgBoUKx3xc1rPk9hAjisWXlHlsYCGzv/LxA9uyhZUnCzIVdkDrCN7KPrZKx69D7P195bdsN7uMBi29MKr1No7NlCmFUnODannWV5bHlrt/KxK0JTPqhqarvJRUa1lSg/gaS8VNMbe+/kfoeEPC01M/HMUq/mRiw8WVXmzj8e6eQ6fOVz+oEf/bl+6FOnRcfivdlVnsfPuIvbcmNmlkdCQL0xDbEP9rNYLcyOX6iepy1QefgeL1ruZsnC2u27Y1hodZU1y67Roy6lUFPpf6XU3zTuJSSvRLahBWAHgl39y+MXEsAwpuMjyLIW5CokYKOxAoeeCknugqtjTCXbo9xHLGYIApdA3A96JKfQmQSlS48yVdj+fwLzwV609e4tnJ5NwP1BoVLTmIxGTGltyvH8j3Bj3jZaEJpwxTkGwimk2UVQNrk9Nt64kcxD6nmFNaa0ktlKl+cZ7BXyongAZl2/I4p8i+y1I20RPrWG++CNOfNx6eMhnIJMzOENlKSdC5DMtekb8uFJdxRk3IDzg5QKjQKHArRQbVQ7SzcjXLkcSt8LyDZobWmHFcw7wYddXPIFI2z47KnFuAdfk72g4Khsu5dhlmUnbRZ0MLimlMVU7WxDYARvQCp5/BySLkw9UCVg9wRcgw1L7eXoguCCHzxxmy4fq8XP7hA1UTC1l4CPYjtX+hKQV9htB/7Cx+dZv1M0lEpXUt1q69NCc+AHYRJLB1dg8hZUbSDMYTWtz0uJEpxKNWpNjL8Md11GI2DMNtNM1RJyR2syVmROjjTy4qEmUS0nKHvJzMVhaUASYpHENtfIGKzR9jr+qko5g0IH5fyg8G2Mb0bMwHS2H3r/Wp7Id+aUQb6ndR8TApHd+QZrbHQQ9N1nwjAw7TdNwfDetc1och9sH4yujxM/1XirUD86ALgKfGCb1Ws/wPxLVnCvIXbz9ode7C0c+5iREKkgWuFazslJ0or/wVVJJeyKDnDskoif8jKNVbR3zBx0o/XF4Pf4LBdUTex84SKLy9xC1qnnVXqHepVbDGPgLSt4rqGXebu2Ph/+IZ7xIwwKcORj0FWVdVzoZeiXPKKLmXPA0gvL2X8AhRhyPWfHciSDQKudujQdE+CaphqtUq2CCgjjoEtPi0RZ4HZ7eM10n61EuCvgwswooKB03oNPBPCyyjrZ8d80eRrYMguq1Fccijwgmp8obJo661Iqm9eHwmlDlh4FdPVq9aaUDReiDfAicTa+doTNFx2J7akX6Y/izI55++5GLzjQrlS0u6Zqe3HnHm1+QdM++Zuu789tFVc98Eg2EkTBLABPu13e2ad7tWKMWIOpEvINMnJocNr1Ub1WCANWPa1WInlzyjY+gFRfYDLbmmj1ui7pmGnUYW9O1bekpQoCrTMsWvZ0/hWyF2+E5XD43xnn2cIxEn2C/NLJmYZRqLkC3Fo1eVs29VLkGuLlafhowk0FbdrWOqxugEp0+mxI4DGuOGb6e4yAa6ACP3QvpDUR1BVBkC3VaXk4/2vFyfbM/8ne0wW5IskSJ2BiSyHCvsXsSaNxLzNJUkuyZODAP5vxmzeef5eI8PlsVEOXJnfoHO/Z4NtY7Ex1zUNEHoxGbIHE+fCoiDfmi6Y5p5mUCBK0KsP4rITBnt/mORHwlXI/I211sa5j6uktDDKtXj+iZNcjX2vhGmczQxx0WWtOeeor91qvCZywDwbrRw5jE2Lhgr/18X4KXMml8VoSO3tMbC2d+H0RLtghXKX+f2YFcVh9bTYf8fZXm/79sWaMy6FKnsy3wajyV/XdejCawdGc+7aWS5ezCJjr/sOzE9+PYUUBYQAkuAPMX0J5Wt5BrB76MLzhDZl65rDWraEZK2wp+YLGL52GFd7IabTM1feZUYDqdoBuNIW5m/QsLwMLBgObMVX2W3w0pe5Jqc3o6NVSXm49a6TpE70qZT/aEzyWF7OPTv9zuY5DJPXb6MzkmrbxPw+ZRAzrF357iW6Na9eOs2SDn+n8xiYW6EpzsWpWD5xbAQea2nNTd9uE7a/ovGPHIFmXvpR+WXXrEFuJ2re2ooyIaYQCddREXJTm8DSIQxRvvX/8yj2JAHn2yE72+4J5FU0Ws6XUNIVgBego3JETCx4Fslye9tB1JyHYo7ERmehFz/5zow725s2mI3UOxDryvqapgVZcU0A1Ny3nVk4dYLvFFhiR5z8ZhgL6G0Ci1B4k6gKeAa+lyFh4viWLfFO57SwQK/3ZEYcrvI7qYi6xowmbxyAYkgFg31jYmCzjdXYbvLRZxCe2HKt6Aza2aCX+hN9Ui+yd6jD79ChxNzz8ROm82BpyTR8pq1KRjgSd7RCD6CnJLmb48bH4vORJTWLrLjRQZ+1rUC1YJgeLCcjqKRFyfGa7anQF1LYI3HBW1YB4HomFF/5I50REmjqysrLu8y3AiV7ZJv/Cps3vfzpfL4QU8voVpzYtPyynkU/OrrX/wLyUWvuWw1iDhITv14Gdq1hEjjYg9u1k26BxsG1RjeUXJgoNHR2uvNEVw8WUEPxrFejx4guxYHxOdDg+qnVfwxNfVqH9dlgYNgeksmHGvGGIV3cW8N2ByhNBe9dvns1e9jgr1OfqXwfeDnRvyJ9TK2s0nLacMjTK3ecnWk/Lz2OXT6vOOCHXYRW8u3V9KyPOn2O+CSRlPfnLKSSuQVv2aOWAuhTooZHfRjHDJd0HNtMeNB09u26PQ7I3OI+gAogwokSDgdZsoGYFaefh5UWW2J3zUH5YyFlkBmRmL/Y8Sua2baQS0RQvVf7W8m8eph/kAsfuUvu4NAiK0sb/iip91d0gKhmpSJZFjTmhQg1MVGzrBc7Rsi3GePQtn+g59yDfQCfSVMATWivwTWjNR9oK3bVKvfHD4fbwOgRY8GP9y9tMxZzY0DTCCTIBiA/Z3O6UXP1fT9LTlaoJMnUU2DNtSs7SjM0WU5QPWKWZgQoe4P/U1nDEwlKhbQsMi0/8qgiKGKctdzyJ2DntOYiRd76/59Lv5D/QRIDqpZZN1vZlZIXU5rHsSO6HuMlX9akcU95ikUPBkKPooIZMCQpzvHfUREl006a19ggQyP0YJ+IIdmNKDeQMWABB+TiUIxKl8khvpYBUZCBU7Lv06xbIvFzIxCiYr81cdsini7vswAdfTrre6LKVF16qc7uV7pIRUNeSIbFNcP5WYPTj93m+m8AnfdyHGKbWkcB5+cMdNjMgqlwwv+WdQWpOePHTX/u7oLT7M9wNeEHpJ+myxJX8pOMYmJhhx56GIViEeMtLDLSEpG2+ay6gPpn0XUV1Th7FTXGo1oCc4zDixqyWeidOOe2kkaONnE6R6b8DB3RweXhummTz724jnyQHEEm9OhzVFvEiY2oxe5DAny0XxsrBBmtvdhpN4gRqEGYy4mb0lM1DjmKdf2XV04VsEVUybmCZ2bmYz8h7V5jWso0B+l4CRMhwRbz/x9UnrNhDO4Zc4X7SiQoiK+AcOXQZotPGQ9rgex6V/nSb6WVflUww+yL1UOkFJGxvyacQdvfk5ycCHJp7rpwG7U145bb9vEJC5A/i8cHaGqyETBPpIW3Pu3/1foFZyswWeJY8yWLGrSxnvHjY36mwVYFV15tOVgdoJdCGCEeV9zxndqft78rdJH0XHxYOezVZPcVf4DAkghkZTZYUzK8DdPwLy+y2SDpK9daUhGVidtI7MwrL+Gmwa39242xK3Sz4MPhAkBkpC6Sd1NV65wziScW+ZTsHXLzheFiHva4UOilZYLQ7uxWaqBMcip1A8eUiFL+zx3AVdcAmPc0526BRm3dL9Ydkwx9B8CHrHaRqMQ/gxfrCEOlOAKdJxK26c75vrB39WVTkRMCyw7lW5f8Kamu5m/Bf7Hl8o9xfmWMhoFgMUuru5wpEStHJ1ogtIvI0lgnx0IBnK6S3gWjxYOYEWSICdYYHkKKxxDrpwMv5JBbdfy0sgmX6Bzgni/7pZothz1ppy9J7GZw9C+hYB99TqZKrEurji0D4xyoRTVnTDKfBzFptl9Lm2mgT/m1gWg9e2IAhF8hc62q0QAB9ZPquw7Hgov3oohpKldNk8DQw/p0tlKOfdCIMeUuGQUeoiOA2+Iv6DJCDND0iTuMB4YeDNdPq6HXSQfy5bosBoaRXkCFGLX5w/mMHk3qNssOsMLda9+YLSWYkFGSY+NJyZlwDspq++MeK168LsxeyFNpgGZb34b5jSRdYbbJpc22wjduulHQSq1TSEN4K080ZSVh+H6cugSrr2UETFPAQ5En8pBG7bTrpuo9dO/v9t6YSDAlz//g/xNcL+jYcEaMMgpYTI185r7hyA6qQsbr7GGoePtqLOQFtEtd0j2eX1IhFdMJCX3fxuxIhqj/mdPRc+kx7jWcoCOdNnoe6tU4AibH3tPtkpH9qw17Sy7tZRtj1oqeJ0QAmMyDgK4h/M30nPi6M9gxFJzXsSY5ZxqJjPrEsRgwkz+nLXLerJ/laoxBKvF2SF3s9K8k+r6U2T86GNxVXpZCmHl/9Lm+GG/xIeP9cBQhHIZzDRd96SS1fRh1b22xrVecm7eKwdx6t7Z/xtCRBTZA7DwQBhfTC19hojHyfYV3Fwg/ljGRotQQGJ5Fi/pICLxtQ5K+ld3IBhYrArdECD56N30x23Chp93VqbAK98DEZD2Mj4hKBj53+7grLUDXIt5kGCipujyjNrc4DTEoAab7bcDiGhA+y1DvV3ABjqFo36gXhJWCcsobc8tAb+4jjtTnLeYL+RPO1PtzSHEiB3EuAeCWZ39EdBZXI6MXxJ3yOEYlFyNk5MtT7hnjAcqJJJO9S4fHJxKJsg6e2uPc4v20IS5NhDnYNsqpXvwky11XskZvHCrv+3kwUmnwMzVNcMzpRCi6EAZUUVUdF4U84TR7UsiRBo0i7wf6/9Vkn1hmKbGM9UtJzUXyJSAAnuypY/V/g7ygtLFFx9chn4PeNQ8dVY9nCB+QVfNUJtuAS0UnLg5IoYCIizdAs16FfNiney7O+5yqFZgeMvGOg2Ub8S+6vjD4ptagEl7iM8J+1xAYxXjSkW1qHuzvM1bETw/sMFgc/5kdFtocwSkBxCikYxwRyMiShpeyHqeTXOIZ44Z/5s7sQlhGrVvWwR06jNgkSwE0pq/miDTMneTJwwd//Eg6tVzxUtMoez3U6rAm3ouUmJOoCTPyPT8P/MBt5RfK3tgbRrH5RaGPjvp3TCuurwxlT28BmZoI3MbOIufJ3ymNWuNqn7C9DCBCVFCCLCc/z6JGgublGe9sR5tP9tEhawYaqAqS7k+iC8aIi0Itnwstd7ixqR7btHOg32Gy6gmInFvmwsmVtR+71AI2ClisiQHnZwp03LJ2rToC/k8Mhr8tClPgoGeDdqY0L+24OgryQIzuo/OIPrChmZsiivPzwzbEZhjkJK8Ed1tBxx+r+/khqHpHEchPA9nZCcwKp4JG0E0F14WGNqZbxFcicCfrMYGrYo5qIfJCdCU0vutjyLqwqEX6SIlm0Ta0mgbCcJKBDalizqLHa26E/ALKi6KExs+FaO2iiktd/CoaTZg1yiU47+bZkc5TSaHWQJCP0+ZCgQ1GCpa5KFv+w4hpa9dwC9++YVgA//vFRZtl8oKWyFZu+yxwiK2w+EWGqIF6urO2LpxzbLE9zlrp7Mro+lg/hzBYOdQNk7+CiqisY9nRowkNlE6vQBhoEuRn1mqoD4vwCjfftkYS/Zp0UKo2tTcfSx0WHlpZx9sHZYgFXS4jf0CaRKqXSPwBoYvygouKzOzVxx9JI1z7geunlNkilT3JuyDZONpbuMGyxnmw/J5JfCKvQYzaBblQHoNTVnQDMuRWdziDT1yczKeoUTtmgTObur2fvP5iMm9NlcsDhstYLysrgmnMyEzjzPX0DC8LYae1ds6CinbGTeMiF5vNxxQuSbJ26VMJJud+CQjLbNcZuZ+wn44L932QdYy8dKQgi8cK6UoXAiFMQpWV3laE0zYumiBdBu20GEDEh8wioR2qI9U3eVUriKjHVnwUurO0MVKdy+B3Z0cQUmZ2kbLUJAKGKpEdz/P08l4udEa9bdAlZ3yzkmkIvlHnadHibe4lHs2g+m7DMHviOs3tGYCygRTEk07VgKkYgwcS2rbYJbglwPIpdxH1AMTtwEkuxkr8UI4HsWWBUx9iq58tIbQZKT2f/QCdRU9FMlz/vk2J95Hk/D8e87tdGXAKtlANLME+EalLM3k5zgmWkQ0R14mSti7iyI72u4KwRRIBFpNm0QJv0MgKkxsXRJSTCuRDEA/duKYclbCm5iyM8+j3uAlwPt3eWxk+rWGbinj7+/Ekis4NYmR5ocbH1uONG/UDxKFzm0XQyGn+k5B71s3o3ZvynR8+gOF58663TSDvs7n51Dps9PIGsmFBFrWhZdp8+Ro3fu7NwiZi3tldRMKsQKcNwyGRxjvb8hiB1fUvZR1F7f3E8t2b7xFQnti8moS/WzdWVFo54BRm6NC2IswSTMXejV4paL8tN2O5WmxmJe/qlTAi/8w1ofpfpoiQjkRsq8Axe/NsqIscyKAfxLKxm5IrJPX3o1s1lQPhSFOSjvgRv5ujf5Zuf9Y6cHtFriOwg5FrvLYQDtIL8Mk2PXG6E8c6lzJNXEY+5UeE7y59a6PEM3BZbJjkfoOvSASs3Nc/1kBmbxPcvtQQ7WdlGcGkljS/VC3RRj9kvCEoAKtTbnwSjhAvFQJW5ZEXzVdJ5Q9kZOynWRcqdY0ezrQ86yrz8H9iwGCsRdMFeT8OhSTGDZJ7i29cLGJWiCyBuXdXTR7Sa97KnUnwIFSZLuGH1Rqt9nrpsqe2qeyM6RWZd0q5mVhWuM/Z+OtKLg+5JRzADZ6eeWGD2/rUtVPXZK0qVkET+vDYYFYIUWzYe+rkAkt0AzrsjG8sO87HEiXyXch3l2F5j82a322aSj85B8r9IPOhW1BNbFpyJ/luiY00ePhdIcDIlsYlAMlWdP45S1Jh3Ub7eZpC7SRgCoVaeS6YMjnvj/XiYTH9naYxEw75tblf2rT/AFuheC6bUcEa9QiPN3pA7ImT6c4Rqypoo84uaofIX9KBF+FRHSoChljE5LjX84Qotx5Q4yDqDiERHhiFYGRtZIPWdIJaSFEHjYJuKVrA/ysXo2J98jh8CnS/JvGAhaSPHRU/OIUvvSyBI6fvhTQMggcplARz3Bga1zGPgYttr3Gr/Elm74jgcoE6Annz3+YcsySWDAE/hegxz4AN1fF/EF78YWJUhoVPBEE0g0xzkuXsgDpBy5JH4qliZLH4tgIUq2DDgJh1b1r4Ln9PEvUXYvNmZ+1UupySXbASHWhSrOlSZyQc+Rjc9HOfgcPsDMbCt69Ch3OSVQVJxx9gEXKnCFfRpQ9f8B5UtCaVYe8q2Hl7IGAFVzPZcOc/IyoDnfYSwBieMQTGi2ZymLGPYqwxI+f6FJFEwTufsT2rSTVFQBHUb+CE1s8OgXZ5xNrd0jJyMSkN6KwoGGxhZNHjqKUUgIv+1y+duXQlPrbKhcCFMKfraONNACt/9mAFBFByD7GAvkiE9MQ+iPHO2K6B4DlA0o9Ss6VnJj6AICXaw2fzMnHCjptzamXw7CqlEs6EN6fdlgV9Ku0QxZNlW4cze+OxrH7jTCPHoMLg5Hray+yAWs04EQsD2b5HwMoY7+TvUkZe2zteEB9dMN0wl+GMjHUUU46F/0JC6YiDdid1msC/A4+683KJi+U/UmxefDJsu6BqiKZSKgjL/WAmpRqmk2pXY2NnJwQmX6J7qkrfHPVvrlXI/ZV+DPPH4DKMseyjumfwqG7rxtKwM2lfh/I5Uu17YDthLbzE++UY1RTphwbvrq5kSgXcc/C4NUBCNu0/BIB8iKcYmb82epCqlZ+ZLrELlK5FUox8n4RuCyMk9dEfgaYgDssMWKvWCgLAbpEUAW/DO4XfsJkGN8R8nba5bGVMhvhAb9ROoRCQe2t+cCWUcBHVURrGUetFGVlIDavcYSDPTeEkcNRVCelNAf/2gZ8VzY3U5zRAolczGAdZ2YnaBEZ4v8l5TXWRQ28uR6aa/7dazeMtl1vS4QfhwQrir8zjE/uUENqyZm7AwNFXgBUF6ggbh5uWghsKl2Gkqx+EvO4UIjNRiLvZdzkQGiAzxeKUrbVGzr6C9egoIo4zWKioR5bqLH+EpuU+Yc3EpDxcOSpOPoXkSkqvg8lmgMjJb2G6zhichEDMjQvrHCPMn22XqCl61zS4j1qfC13/gLcKlieMFBgZQ9OQf7I0/hCW4VvK2q70ONE92eqU+g7rPlU51BVBLkclM4CwqSA1YdOjbNLR4YtWOHglE4bV9ZDTdl6SLqUAM3UYOABB1RCQImZEas33tm4JNPVFynKKNC8jQDyFEKsCRP0BvqvTCEtGmSotaRJTTYWODtFlPGCjEL7Zrdpv9sO5Luzjtlmz0m0h6O7OYKlWeZkeNTttBck4os+mkgyU+DH1zSUH1TH7woe9RyYSM1almw54nNuEoMvgohMheSfHS7twJ77KjO154jczmktjARjZGES3y5be7gfK4mZvHEyFtCM6ABNKEM2WjOEmzfTnPhP0yLWqjGU7HdZt2IKkFWsU4R2C92cdiiJcgZikm616k6DJGwnSCvWM/IBN+wBO1Ea1eBNAmqyxDfPvPY6lWYXtbbCjiRFUATcpFs+09p5Dy+MB95XqOm5UCAV13hTf6FrSbtunTgujw2PcsbJC+Qs/CkhiwRhRKOq1b8O8OXOUq3PV//GKXlIcit4aGbGEDxovSdjgc4iYQRNRLxYrvYQtTmBRNnxSNwMtC9cBiWgPYggdTbfX3JBbVCWJ45YekZnZPhd/aQAIDLE0e1S33hNQATgG8SJjtd3BqlruFmJJrh6QyF8/EwKYwM7rWyrzNJkSQj2dQlzMR+fdkV/KvcmiL7fs7Tb/NQXmBy8h47poobi7Gs9ORcpanoHtNRSp0GUCU0zvhs/IIx1C8q0yYoFIVl0Ga/ttr0ey64py/s8zFAu67j3bD/RBjx1dyMH3s3LlIVDQwL0bx9XTLE3m38MhxVJSKB9ZLQB2po4Wq/4rP0EZKUi3J2THgpTXzJaJgygu7erA0hT1N2U+u4T4oEphD1vgC2BRE4OGpdgUWCqV93Q+J5tg1f6CVaH1h3D+72PvCyBUugpvjwGhqkkjhMGCxF+yhGx+LkJhuJFLX45xiPOcKMMhUCOSUee+OKCoprIYSV6oRKe8HtaEm/6o0ZWi3fehi9QSWlCZcCdT/DGGj3oxoNZXAqsEFKW7aItAgMAlFVu59fCyOmSC23HQM+CbsfMW7if44m+ksrNnkpDqVGGyBsRjbhMqFAaSo7WWW2FIwVvpeh7dPB+JQc61GsGrPg8ax9LwlWjExm/tZU9LbXa2JhxHQjA2/O9bFQjufCZFQC0lZHz/FRBWgWF1iFkmRZC/3xNIL+etcvM/A2uPM1gRe7qao0/Cw31Wrxb2T9JFiYLUhjXtM6emIz0Gwgc9AYvPkvEh1JnRzIlZxyJI2vouftgX0chzaQXjotQQ071CPiXbbTpAu/bqmUHVBsI85mWD0fkFXb7m+cDe4Tg5IMY7kjGDqBoageZXozXAIXahh2QqoYJnouBP0ev1L5Mmty4zPb/w1oFrPllC64X3ouC0F5JpHegLICQsDXtUOEsmUxHxpPQKLCRiFvtUStzCHdVG9ZzK/2rEd5YSvqqd7fdjmRM4q/hCWRfV2noTk42VjTsS4t5IUou0V9Oml+tI5OwogtqB+78pvRuI1EGNULek3+/8SK4z+0JHaNmiLMQTt2vAeWUodrpkvZMRip2SMAVmh2xFPAjowzo3Una/95xcJG6vYARKGYN/BlvXUlxWIs03AWBOYDXKz5e+GTnK0R7OLizttoTA4F4U/te/Arz5p9QPJ84/sU10g8A/r5vTquWV7l9MXOwCAK7f+SQ4lhK2Qjqj9X0xgzil+hdzQrK3tshLbbGpQmH3jEodryORMSYRMHodcZfBLGtvHxttSYtbceEBhkcmkdZKZ0cFvOWfJrQEP0tOzb3n32u3OynnAOGPBXGmgwvoL8dXYwrrFQukku5lKtl84HXAJn14WDjUdSPqiSru90ZviPbbPqno63Dt/IOQD/GX3U2+7zbBzgZIGK4n8LnqmPj6fw8GVqKaZz6EKD/mnMPzK0UHhOeQ+OjOgZAvFSacNx33y9UcC/fjq0bil3nDyz0o2RuxFaYoZRmsx+ExgqOkVH+3Js782QZZfL2kj++ou/ErbEIcCMeMqTfYYy2XlAo15VSaIsFbbrrIiDs0ibAz0hL4h1WqaUSaATpbyhhLurwPyBcCtmuEWMMrX4p75h0UDRu9GkfZJb72Rtr7NgVR9EFiaVB6K1xrStTv8q1lHyenurgFPndZGXfydIP2CoBY3lfUfk3q0aJAhwiJtq3Pld75g0TQKTFJYn830bFaifkx7tAsL4g2lCim8zFl1UyTvFBBC7ugwW4hOd2TZB6YHuz12wiAaYFg/pGjTVBSSiI+hQPIFeTvHE5+FM4Q8lQwxic7e05tovLia8HxqBM+sSfoj9IewtD94dc6ffaQwvzWk3dgwyb2XUMai4sS/tumZ5JlvblKqaCw+CdUgMQgMgnOYZZMiBRnX7REHO6YXD21MrxUaqyV+RmOf4TPuRYVQZprwNDQoacIvA7AQoNAGNU0WeUoXGhCRPG0uW+u5Ub2vlLY3036cnhJHvL3L0vEwWav0xxczUJ271/TSkorSbpKfCAtvQckZjM0JHAAWgj8Sm8+GL+8mUoFFoBOfB1jie8cTNt/9KF6Eq6QnFbrXS22MvBTagpCts9gqbqumuysoGxrc8HfVOhOQeF6g+92EamSNZIvwKBVCG7s2dbmaOaeHl95kX/EmVYHLYOqMCSk+ItmoVma3BoK5Vpl8yE/KYQ+leRL0nSl11RTJai6TzjDEwW2A94ZJHvCpasEBNVjWx8dJVaNYfws3OgCAAfw1TrFTPxBr7wv6nIkDvnses0MfIB4acmZvHsoHe5JdzuFKSR6ylNr9wmdwst2dZAHv4U7nJ0L03m/XSfizrUY77BrLZfOVdOJVxEYP9lOLpwT/1/hoIY65OrHb2MNcSjC7KX2xrPUAGo5L4T5OoHbLpUpS3mZkrG+DClNJ/0p/9o3536vsFTeysVszP2dM4dXjdMP1ppYbNY2F0Hs8eYNSoAA8yI7m7h9uT/6mjk/wL7fTDx1RSlL1kZjYVOuUCmQSLTKdvE+DThfyWv57QT/9u1EkQJauh5x8Md1w4+4YqtK/1t5MxWUEKeENN62gNNct4d7R2s+1ZUFp/3ZcmcM2uiga1lVTaXxLpN+Fw4GWKtUEMFrunV2yfhFE6WPnqAovk6WU+ETkZUSB2qJWMvHpBNfC7QnhXuLC1KIX8LfnDdRZMvFo0XVTqMeBQV2utLXv8OxYU2sd+o0rPVxWr3Htzp20QyjUiSIqfZ5rfWihDo4n+R12dtRqhYl6Od+aqz0eXgnNpWWjKH7cdPFFF087zR7WLF/RTYu7x1Rro7anyVOlfVWX29DDvV6mv/MUN9wXuF5x8s7OkytGWg2hYrzh3DqTRu9BnzupjyFGLS1FifLHG2kRtniJ9lS8rirsX1iLWtVcrtU1iGgJaMKErGM1GJcwXM7WZfzVB3CHPnWhT9dTotKQcTcwllcFPqj4pTrU9x1D+Up+np/l21bxNtr1y+j4vz3qck1YeZutkyNWPzAcchWK9hTSD9NuOsWZgtZzlMFsAI4qNhzrdlaXVLV36ur0Kz9GvkuSTps4CMn5X+cJwUyzwEQmtV0Ua22mZUnIdXblV4ojUyzXfPtJ20zlz+ti6FcSwd9EpD0cjPS5yyEhgJegNb5E61O2A761v/Xi3Jg9J4dcYVOCEtmgUWdEls0rg9K8W+xkhgZdX3GEzp/X64510QcyIiBqrezPSa7i0iPY5xshPtWc0nEq5DA25A7kqmRFiJbKf50MUzfLLJmw6TTjMiDdNdHo9TS3DwM3126yaY3gDOflBCC/wrzdf+uQmVPJDR5p+842jt+/ems0xWQEmtdCm8VAh0RI1EH7/zaGGopXGFO8DGD9j1ZtXKy4WrPYLkXXVZcOazuBxsEn5hvyGX72dzKt9PviCPX55lt8ylvAJSrLplzLnPGq2T8SHo9glGYDz7naSqnEO6hQZ22GaxC90YeL0T2S8M9nvakaoNivleuqjg5lNxxvdbi/dvgzZQiX7Nghewga4yz056oXipaC08k+Ppv5j7ijl83xT8JiAofA2zTimmXSdXgla3Scy1LGA9S07peK97PzHl/Ggja6M008AzJu+omZyLvuF8znzutEReCQZX1XjPYvCagH1fZyuWlX1/I7EdwPhERnlnqRjDXTBYM7XBqCbi9TTLa3fZEwVWDPufMKXvJfd9mnSw7wftIA4xINIhSQ+0VTCVkoHO9f2rtJeRNJvYYiP49KQ40Fv+dpjXaDP4ZLDCcyF2enY6c/HWJM1aZ/dr+Zt/1qKaxLhFZPuRI4BbD7eSyUKSM4/f2V6+D0nhzaRD84RhJlPCeRbOgU2OwMkXUiKotoRdtUD4Oo7oFN5kaCgy245CAEOqRMSiLLwapkagV25O2KhAbNySxtZt1s4i6/JOXF5ozF8tJGI1XA09JOtR8/v8SVC1bhco+LWFr3i07SqEx9F9EIcn0h3DmOloEL2z6tjTB2+QlQvsUC6tdkmdwjioyy8yB3+0mn4/gfDjdu1eOJdfzCz2Y7C9Zcg/RLGd5Gvg6yhGBSQyScSNG/DaW7izU+o9E3U6tQX6nK3ZsQRvwYSMVhjzBTFi0bZmY12vtSr53ZJs//Q3UECOyK5+UWj8yqQ+NJUbvU3cMknsHY22bgDkjM2XxdfKlvaGT+Ijmo/xArAMYlix0lyAWKOigdhJXtovdHAHsqxTLethuTSqFteUjD0uMUSNElW28pzCj1i3R1q97tXf9Kp8Q0lHP7s4nKE/M4/Un/EZOEAn5OrTuSMNtrAu6WK+stLudHWyWtVpJod4lfOiOnI/w75CtOoawiCQEA6CWXSaSh3naGFyQ8EMr8nS3GclTkal5kxAZ03jEGfgzxpcw7SHgtTUIbwpmZm8AGmRHWK0r+EZhzQvydciSEeB5Bb0H6qWogEbuGbGUEVBXmqSP0NdvoXsx96gQaRqflh3kDmfczKIiaIovxuPNY+36BzkKD4j4eQ9//6rqBd93vS1XAy4V4fCcskgJIHyJwlrv0jEZAyhZGt4Hvu5XgNmp25FX3D+/UEefeBVU/r4DP6O1FIaXQkJli2ZlQ0JzIUvmeFcXZqiMcK0KSNrWnVJFBsldDrLnVWfl/eXdssHafC8K+WzIQTmXHHsfelLujyQ4+0Zm+dAu5BlprG0qmnXeHrq+d6MuJSh50p2jUAomjimC3QfcK8d2uUjAcTBGWh1Se6SRkqXx4f5slwWEl32/zEAMTgBqku8oHG3ah0ld64F1hUJXg6fTMD5nBSiD2aN4FwbWq8rrlXnG63U5IFBAhxhdlzv4rOztcyhJ3tdMzJZgAsMXys84ku89/bxFcySuFHnGENNJ5kYlCJdy1CrATY7AsE9WeQ67hlyWKVQtFZLI6IXgYKAjiSOSv2RudNfZIU+VogH4027X4ifXVy7tDpi+g+yDJILrC7Nfvz6jJJ0qefnjinrtxmgPa+tDUKj4rZ8nTiQCp/J2UxlU5q6V1vKKq8FMcM6G81fbGd3KZ+mvkUtjEWZL58Pw9NfV+hH3hzZ4HJ9eVoY8+XjAd0YtfDJEzrBNGjWNXKmxwTKRBn2xRLsYMrjEK2C9WVRFqJmEqLeGEvsg7xlR+yPZ2U7LbdqqY9V1kENu+32qxw0Q5ynRtvth63G33N6hBRqEAqm7qZnoWkA7kMKGnqZe6tpI0ZiSeC5AWMJfqtZ/yt3xzb7hRuN3Ce61TSMajiCj0SqJNd6aTgvXDkvF67/rZHhj9a254h8dPRJ06rKzLdyF5DJ1j2I+NSEpdqDIJIT0t+r2rGWvt47JqZwNmCaXNfTNZLkrWbvGg14J3Ue7rQYb/aa+NmrnPx6BDPTN6D4+z7rUtEFJmqKX9SxZJ1WfcdwdCM6nZP9UfwHMqdsnFL8Yu+Rp5P00ixrC6ZzJnwb8Ky83eB8xn00dfkkxaLuYZnz1ei2GS2Y1SMF7qRA29VTyYxvxB4UpWTMM7gwu3Y7Q8/l19HNOSt/FHukIiQdVV7gyQ8KBsAsnHG8g9aJ8/Y6P+5A1LJew9Qe6IrwEM0MjHWmwUrAfqaU4iHEICxkKKLXwpPx1iYwrPOKZRcuq2pFvNHx3/iycR4x6LtkYp153eyLn6RB+DPwe9951DQ6tDFZpmr4yp4aFU9e0Mina7QUkAzKgsLF5Ofg2QjsJ9OWWEwTDkReZ07v6J4f/j0DZulJESvk2ZBE3wF7pKePsIVJIPjiYe19HqmdvzlE4HBdC/MVYDKcmSzoCGWP6HiXQ3lQ484b1dCyCH9u4MrJhMfpJ4jPleLNYjp6ElViqM+aNdGvv+ZJesepWYfJ3O9pP4kmt9ts0BZAthJtnxBdxr/QkIvL3hfCQnN3cBa1KarfC4poTrYrXzyk0s2eXuPm/oPoKRZoLuHC+fA42vV6oMOyvsFZQKmd7KGd2rghD59jQNASyQPOd8wu52eFlA/LnBM4dkiteATXNzle9TF/wWiqmNJwaMSzHYqqJH6vAETuPxZRieBew8SKMqIrPgresKBgGGVfLebmarOtfiCorH1WUbhMH+0BS4lJlN4lTUjooLY59n398vRh6BjFi8S5Km1Gkp9rpUlNGUMIKiToanl59z9+KkZx2d5FONRNOIBLYqb165wJ4abtNN3VgL+WGflGKffAAhc4ozR+bEejlRgSmGsPY2ACgHpYgLZSIXYUKSxqiFTtN6w1gjJZMGgNWjal7KYIn74RFs7CYpNkI432jC5rzRIXvt+hSp/FY9wv175Tn/WkCHm1FnGLc7LXrNgGPRTHqgeDD6+z15sSDUCBBsOyqwn60EsA5I2r4SSA1o6f1U/UKyP73p8tl/vk9ldc/wiOYzzAJyBQh/NAPfOYSGlLNhlMqhrkDvEcIavMKKyJX/zzwqFeot6WmjnzNtaNF+ZV2b6R1Vup8Jh+lPyxI96Yj6fVXisCd2+CjVzWPyPCLeKdK4BQh/8G1KNnoyBff5GfHSku26QkWVPxKu5+MWVILuJh1k4n9ElEEX1GT3Tcwso7cmB5io1zCl4Z/Z/tvQaGWOxWqacaf9DbkWoJvlrq9n11dGgycrt6imzjbf2I77XDnesUefzEw0S8ePqV5pi4JA9KB1/H6C+oKvzYSHNvhBpx28fQexN3lFvClqhMlHcyJONhm1GKeIdi3SU1+Fl4AO7A23ALsTX2AbvIBN29eKSeN4rBU85pUNFoOBihPc6mS2p7Tqkpy7knJjqNS8CMp9+bJ/AWTfHjBDCGGSRoOwhG0AAuS9uXOBIEphGkbjSbX7eLkCiQJ4Ln5K7aps8FxflncIvR+Vu0U8FwZav73dncqYGs+WSGCtSqzhuWGmy1ZjEW/TxgBXs0jGL6EYjO4RNTRWadoKKHbIA4QDTToQHd5JEd4+YEn7RIhmJZpidrv385xZmZitn6RRokZcy+1sYr5p0FxQa3+soz7Oux/iB5RVnI+cy+7lVAbGcKOuMYXV95YvjRzSG2xsMqAKVf2Qh1i5vmehYAgik6OLc9rqbq5Uy4jd50aMGirzaej3oiQxUyOhhX/icvTl4Dy5tN92fVwB7obclbGmfjWZOYqhG76eJG0qXSB32VYUZoqPhcuvDdvDDskM361HHZIBZ4sll6v7WWDfLS1P53HXWSml483fYRp3xRp2hakJUPl8u+dVYQxYBLkIrAuz9qWyTtreEJkGps2NwY1nk3/b3lQLyAxs5Cok5CN7iFktWOdag3v9cL6zhCfXdg8lyRzlt5GNp9/1Ohk/vxsnkH7G+1EgZMl1r2HROB3kE8NDlW8YYw7GS7cFxx4VqjhWQoXivxmYjMglRmPnZfR/RIT9oXrtby9F/0lM4W3TlRFU9QieEJT/ZvbYC6Cu5MIxE3Z6IcKyFq6OEXi6cV13M/qRlH8D4CsvP2u0HyWCliuhRFPTxnLtV4IN5fM8EsamsgKA2CEmjMREG+MLb86JoqnBn8OpIeToVT5kbReEmqy3fvp4ss07FqSpHPn8itFzBZcIhu6IXFch4oBccnsEag2PEM3l3FCH1N9P+Wvs/8ldUITZaaFvtSpliz2GL83c/Em+TsfYl7uLuCIMW0RHxWV0Kxi/9EXpN+ema0o+z2VByPa3u4xiY0fddFfzhs43dSBOjz7grULj2lRhELzaDinz9XnjD/I6VbEZGQltxpkHJcp2fvzfGIgFTksll1V3XEXDyfxhfaNMckrlh3hPgezax6SJ4oPPjUrWfcB2+SEEVpNZG/Tz3qffuWt9XkbHTbiTs8RWeHaPkW9CSc7PMn5UnNhTb2Fk4PIZ5GwOmDdtvWLEfdTqbzTYSMdd0UVKrC0FfEch6h3IKJ971eEbvXUI/5ivdd/Ezpkkl53AaWcwcT5YYNTwAFbGBLlLrou+tO9Vdnbj7E1GqgNqqu0gQ62itkGG6Av3WWTBQBeFuytKRNWJGYbre6uX7JqerVqEjC/ouiR5CiJbMM0TEhFZHiPt9rd94iiYHSzOeO8HoM+B9cN+4rVfJxJWiQ8XIgXyFceDnNSnLQBq5mgNsT5Zrp3nCcy2KYeUr8bZj/7ukXOEaAH6eTlIlSqoRl1EQPZseYsfW1L+7iAtkUKIKe8nJB4Rw2NqnSjsvsIR2WYkHfrpuBidyAFknv9W85Kczpd8QdhwcE/MSv4+68Q5KH+HTgsKV64aTsFpwEuvt1pTG7L/VFqEcShnQtvwp5QPLFMAwuolGt13QZY2VI3tcQEo/uoZFIgPuh8mkKXaCoh7Cd926+SQnMqAlstksDT762jWZpZsy8r4RIXatGbyNpzUnl2M93Ce0U+i+RjGMFThETlDC6AxDLFOs4rDZZ/b37HZmwtLsBb8ZcmV7ytRt2pibkYMOeX5pKmL1EX51PNK07RPPSL1fKbhtzU7FptxmK3JW84R0F37+xxUmG3ZFM/yArZdgCDq3hY49mprBcLBw+WuVNbJ2EumXGYhJqDOkRDV1tVoVCO/S4oWhD5EcMxYDgvey6Vb5elwIrqq8NgNlIpplovnHSgQf8j+WUqqVqK7o9C6BtaJjYSw5v4q3PbhBDbCLm3bKZVNNnfNVj0Igm9fTRn3tTYO0VhtjQoLp1pFOTcnpmK50ACL2sB8WIy6veeh8di+O0bjtFqkzWdW8dm/KhpHslMAZaiNAlJy7cGrFpPnrHBEnbFihepeNv9AjRhOUA7y5CeZUuLBJcIwAolsSuLciCn93VkbTCsAOvZ5zDB7H59IPhGG9oM4tXyg+8f98VwDPGeFdDxKMYDykUjWizKITHhl1a2LsDp/taGrYGQCIxvPyTSV+XpZkDVY/kyUIsH+0S9KJqbIx8HqEoVADnMdhiL3EE4K8RlKol1USi10rwrY5NX0ku/psZ7M5HTjgY8fHn3N8c05yFDRIjxJQMMisPRGygP4DH3rAiBMcybJ5pRKGBiwtnVWjXTG2oqMkwzc2c7Ytph0wQd1+WM2cIQS3QAF8M9LO3y4ZZUYLs8YsHNL0RInvDRxrwNPL+EGHm60Duk0StyVsetU8p1p1nR+BumVICxvfdxPsSZsrA4rMUqcOCy+zOBe9DJxQRqNbECkhaCH3HAijDKQfNaXg3tkVbRkFZm3mb+XUmEJLDdb+4CclcTlvHrk9EfpUBoKVw/d4f9xZhuj/IwV59jvpvA08nOgaaediTFN07juTqjcDU61GOWr2CnvVT1kmUzaWxLrHhzyWwZ0rfdk77qkok9CNDfVN8w1D9ExbuXXinNR80dfK6knjAyVdSyb4betQAfxQbFBMsSLRfFxTnGD5aEOqQVGSUs4ODZHgIGmlWoUV6x/HuJP8PVUgCbg4/gVm5L5aMRaWRp3zWw36Ox2AHw/tvhJLiy/R1/b/ElIHmbhSQwEQTvqXj6K9lAHuRBcdKQa+6CqRQGrx86MeLJMxeW2lLotdxrTfA7ZXD2M/Xm7KZo7NlCv0jne+QKjpmNeHWPelBKJzsFPmBn9WfENsc7lDX43QRd4rp9bt1KYX55ARaOXetwpM3OAIIRb/BtgrKYNce3GD8K3DFjbshCgj0Zhw1oob6cZD8fqrGIDOl1iJcD8fc/MxSxe3NgNR7rzzR2hVYGfW93t5vyZrfQRjN5uyhehmTtd0H/hqm9T6EaOF6cy6nlzX2Um8qQGH8Wo6z940xSlCTidfHvuSPmS9SdWyoHH+fqSTCrudaBKGC9sWG5NzAP3bDeDTfH3CeokkjZJ719mDB3/Iv7vcZz4TyT2roCZlqjPZYOeRySpFkaRvv42o1M4sxSY36iyvDVM9x/Ky0VabLYDeCoDfjEGpINMiDuHzR4IgGL+ywl4OzyAf8R8ZSGnE5p54dTa4cqB6B/xyUZXg9kd/ila+3wBbJMyqbqwl78K5kl0ryjd1aIavunu72MEl965oZI2c6FH/4J0PWAcGg/UqG7Cu1tt/qNrb8M68+Cx0yrPAVaK5k/eW/GC5cDIFEfAYFleqXZ9m7s8e/IS1rKQt0W096xDseYi5FmZD4miILaoQ58QzLnf+Y01NPSbJOPDIGXxr3iW2jUKLLa5oW2Rb1AGNM4QoqUl7jMeUcUbjuiiRCyRpfZGriOyIbRUNYSCvZj8NJ9uYBrmA0H8HbdSBJ6/rjiHnzkIKyd/R4rTANHeNry6Nd2f9Ve7G78NIsf7GImHDmkjrBoKfz73uSslGSYyyljBp/wZZVUSvBsdXQk04qUPN/cX9P3UDzoAZvpWwdOi38+f3QqNG9AI27NSpHh8miQp1ydCBQNzXPDguq6LJDF0H9OZBoWLMeGGGM8x6IFGbZ1sUXzImatu7QkMHVG79NXdvoKQos2CSswuhaPzTyZGHkl50l9ZIy1I7GOzNtg4wpQe+A88OsHZpQm+QEvP/WVGwEqarIzFaP4UsLL0JIH7AOtWCyAyakm4JXp0hMYy9Kwt7b/I9N9xEODPRXdhVZe//F7ZYXIGzl8PhVWGPY9kNrJfYaNYugT6r6rt5hxcJLkCYduVHwhMkCU2nNSRtHI/0MPnyAHFgz7vQJyXbBs+Y2BhR3GKiQx6FZNzwJmwelfBgeW4yGdBdddtmIxrwbvUnu88VcS1KIqHm0aWZTRMDjqjbptP8CG6CIr9rxURV8DKLYgkbXQdzYVapTtnWeg4nwVTWVhupnjMu6xUUSuAKQQavoc14wdZLlgspjW9sWBcK5wO6sD4ZrDmO9iQ3IfePMJsVTxLDCSihYQVD5h9uLIaAezU+748AEJQwlzDrwG92fIWXqUvH9ofnJAxgQpCx2De0t+j9TmZA6ZqFJB43Y1+8SeHQ1kMy245GbQRY3+Jf7ZipQTeI/bh132djcmlAR4F7Tv1p6F/Xdx3aeshEwGbRtxndczGuFGSDjZMFyY7rLC3mKXYRNAEgYWGNDdncsXGnCxh3W+VfAHti/ysH/RBO2e7+GuUJmZhUwG+FuqlJdrQ33+3HSY0zouV0sLJF0aLPeQ8j0U3yseViG0pQnZkDHKjZSjvV211pwXLNbO//AU+0GlNGSCrEZ2KFITq0S4K0bJeDNZmud1dy2QkyhUgcy3f1wE9w4m7Vw8fTxvoLbYCLQ4OvuGzgyRGMzG5G0h3SDtENmN9blXslonC6kKSiC/vcpuHZ8Cuiqq5hmsRxu9jdLTgYkmsOOaM9wtDT11MMYBTvD1AXJt12gwLYeHBi7WQMY3hBDaGMUMc4d3v/ufy1UWc1dJhvDypF/Eia2exwPzZhiWpUjg7ZeiTeFT6LhKb7EvAJgNgF8I8XzyMyREBD2/r4vGqZMFidhudtZHig6tI/izka9xaTgn7XqIWL2LidozjcNxtSPtB2g9dftwg1Ej5Qi6drEAEUiuPffsttXgH6rBxg5IJL2b7EuS0jx4xG/eR8ZzF1YxCipKYED1bsm1QogdSEkuhDxGlUmNT9Ib+w+3H8gy0RFRdbgBJz6ojqQucEfiVc2JYOF6Wuo2kYAbLBoNGv1UxFz1CzKGVBdzQCLzC1V9fit8spiIWqfd/8gZAQZf2rWR/CkHk1TM0H0es/XPARP87StNii9sX3fZ7mPX3WiWW87zGWitvlt5m5pLnKp9Fz/48aqPDy7og7+jJuDWVkQfG5XMZ1+YLhLFC3TlQBygzI/VaDe28eNLq0TszUmbdSyVIb3B12QWe5DypiF2ud916S//qw6/S7KUc8zlRRZCwA1pgZd4U5fagEHNhXq3agHP33NtpPrhJ3rmGbiJZBNQlRihrTuFe2zF9I1e3SXNOcPkCODf2uznmQckxTrEREJA/wn6Rd9JOhJmyOMQ/pXpf+iG7pNpf4q5IodlLU0/o3gUUMAOQVgci2Nez9j0bt4v/jUu8pG8pnnK8k3PyCEtUhVI2du7Kr7N6npEXB1Gud0Adeslf1oq9ABkkycNHDoROqQ5ood8YRNoE7acbu7CdRuSGq3ODEKsTusVkwCXGyBFpdN1uo3yB5M6RBw8zoGFmkrQIZK/2BI7wv0S2oOVCel67isYr9ibl5t8eXJLIXnCtIomO7tV6gt9TiCL+NyFXwqdLePByG+++mQaMAEM7Q7tjvKjNgksfHqJ7dhFxuwWOvIQNY2/aqHB6L531DFV/p0BgzVuNyeNfyuxRxMndIPZldXSRdZ+PTcbHc75BKr1fyg0CUZlcNc0JkH/RWjdkGqzIyYb3GUWu07WEQfnm4cuPhxICc9Y5+X1Zjnolk3/WyE4DoeaOifONP0KlWmnaBOBjULc9rHETstPCdyDoafcwKRZZo1QZCAWGG2L29I0ZA7EcAK4F5ZTFpByTHw3uMhSWjhdJ6h/uELn//kEP4Wd5tfMaAVYhLpROuuWe2y8DYis1iw6pJ+7QU2aBnS1DghS4kcTxpN0AO6GaB+JXLcANFgS1HyokfqH3+c0odbESMIJzYxKK/Ix03z0JPeHHJuc5+tuBe43QQvVMkEc6o28CvxDgHxc9g+GndCGtE5AYnD7cpIZ4N5j8Sei81vZR9MPnC91LYyjFHRu9vLfIn6tq2fhEnl53xTN8+MYbWsjE1hw+GO/2qoBsinn5KQhSC7kjBqYYQovI3vUmaYV+d9IMA7o0RySQhyTi43/8HoBvQwdq9+Yx+oXr0wwQmgfO8bwlt8xajcmzW7YXizr1in9vz8tfz+z32K5z5bINFimDHqvzTKRG8P6qVPXGQDbTeLaw4nVBNtXqOfNDR2aXQuNLOTkUhhf5cekmjeV7VySH2IzZaNcPGHcLNv27A8qVCwyooU2eSTIbjw6jJy9vLOgdnpmsnSdEOZjegqMyT1Dh4pxGsZh4AG6jsqfEJMDldhkfIwBZWdkNheD+It4WpYWFsfjnlNQYK8YGuolVEw9iaslPjGtX0OQGeVchXHn7HnRijfSfoEPxpYoRJr0U+K8gi3xOOFmq7kQno5xBjGuWD3sP2S9stFkDsaH58KgaHJxxjaSQTRmUPE5L4fJxV/UbKHupSjz+P83odLneqPl1AptP5psRxHrNi3WZWv1mWlnFqFzzZW3thTAzlk1dXgZ2jFr2L2nInMKF4rMOpVWatZuVIaUKtqX6JQedWfG6sPXK93Ak/2k9ZdtgoDLmFmSe8CfQAssmHQLG6MW3vCTH22j45gqUYNe2gqlfFGq9KtgFF/pja48tg+tJ439xK8b4iZFWtTNJs8CoUEbIJPSAf1Zqt5HKLnQBj0h6+2tD/CwjuO4COf/rZSeRAzh7W+xhPJZwurMy3peYAjCUE0oAa7DZulTPPI55szzdKi0LokIBvkuCvpBsrtbNUX1QTE0PEgdiA/iawPFn8dzDTqp6gBG40x+DVpbu6VeTU0Itkfidso3MT8KjK0+k+NqiSAi2tKHnKb+ucXvL+SpbhKGq3bR/CHq7bZFMPvxxoAZJgdv4WB2yHx2gceu5iz1KfdZTii+glJO/Ej8ntQX+zQ4zFWb7Xh0VMgABfTltQiSo6nNk+abZhLUIOkYA21qcwc0P/BAiE7QcpyuVj7Abt8kpD0FihcTsBus54p/1YcuzwyAWD9G1XetofFdhBH0UPdtHFkQx9H3LdgS/8Xe3eKI/uAYb3/D18rWozj95Ya14nVzMq8SF0WDdINOTxbLV+NgdCVVkdiczeMWtsyHJKYiG8+FC6pwFBUzzqGUKM+uLVTIr3tqmtGXxWKT0dxIYWOXV2mK1NU1OW54jNhdz7TJij7v7oXJpahU0L9YSs6FGEYOU/4kLZKs6rv2zYEkMv+spQ9BvaIuHSCabrdF12kUMHb8stqi8zhHftWSw2p6aqfLM0dgfSGZg7tBq6PmqEJUVeMvqHYDw2kIHpt7n3QRx3klSgx5oRyHoJmJXf0VEXAqahoX33QeJyY4Xmtd4y8G0LyTxa1BbJZGAHjg5+IHZLfNQdcU7TnUNicMhG1MUhDMJjiXNDMxcAWSoeX/jN7R8RefNbOTUAD1N8Humgl87e/EJ6PjRqvO6ra2CcZN+2IwgGh30r8+MDdaw3eeiirnNsKSyQKDoarDnRG14DXtWvXIxc7mkzsbQBawca3pTHV+TTjQJjJkG9i9A25+IVW1E/Iwv9xpgYArydLI59dfoCCs4VhWpQ//xzs4q3FhqPXGiMcqliw5TlMEPF+v1xbq6WWT/9FpZQcbs3b/sKCPB4oE64kXWVq4AoQHMHzR2O1XBi90U0R6e4mBIPUOWzmYAHJXuRyNSHXMs0rpdGS3kmI5bYdyRaMXUkIm82kLK5nroDS+9KBle2MmlmUVJ4tBM/0M67TWC6EE2v5WmsystIG1qusPHqCCcdGgrxkJuwgEDhOgTc9UDegALPYuHkxWwpmAvI4YNoyGsTKoOaGTFoJ/XmZ2IlBxS23jlpdTUGHbjuB3MRNgU1unLGegnKdSFbN9wC9RK7pjbd+hst9gkS2XvF1Zr+kExhb5sz61+ldbvm/1IJptZs2xkWmo/Z1ArG/t/k0j8rni/nL+u/XIvTEnarGQMjMSzfg85vqIkFupRTPTeUvbA0K8bAAEzR35FIwjzCwp79LiuIrTIrSF/ZJ9OQF8kCbbQOLVn9VCbO/rH7LG62FgsmLVbcouwrv/yolAu690LjhQ316/KZ2kbFPjWJjZYmSeoTUbzYiDZbcFlob04npKwmmAJYLYIQ3ecj0/kgVIo046UiZhS+dtu6N2Va9WZ5k7l8HX+boxwQSsCaCzHXG4/qSK1lByRJgNiRU39MXkksWkF1S0A8arRryd1SNFWM7JdWLpWUajlxzzEZRkbryGXB6RvDZMv4m9W9NtKyVkKVLXqSPcrNR8NRlyRQL/Gburj1n8Uu/vlCpf0c4+egoWCFcqan6QE0o+pziVrYlkStLn/KZSeRhbAwopFAt+LDOdR4UzXyKLK2RAYhMC/SPc8NefXIEiEWyimM/M7UNyW5qtZ7HB5Vf5xzdlIMEypnJ44MD+9OQCCDAlcSebhZuYhsmMzW/jboU3WCcNPNmK/WJJARZnByzAIsbyqGij4RpIKw5pIHMK/E/aK+SfhXhukYdzL04dmVtVJKVyK671Y1YQS0yzMQwgQPejrfFslMTLvuwLQVjcIHKsChf5FI/bvKf29kMPQmfcj6e79rmUlS0P8Hggr8IACa3s1ckegByZYjeC18Jn9SGrZ4d57qnfW2thr0OEP6kpWnatWQUK6+Sx8VCExbbi77hL2LbJO4nMl1jK+EkSjm7IViilHOloV7nMrf8HN0KBGAkh6oimXIDxAg2PLl4/9nCOZ+dTqoXwuT/MsEgOjs0IJwM7ToGRo8A9B9RXABc9mDmYjbMJpC/A6wfFxxOEZs8XqxLgPQDu8rYGtvacReFBJYXjVuigYSC6ORP07XDuaYTfUIXESkNLZnmPhNBut0lCHrxELeiNp14XyhfptbjW/nokbd9nBRpR1MLrKXVUnoXM8WKHRaoOjiBlRe+G8fGNovX/KYdJwYhCgeFdcckiMC46I+pUysDVcU6lMwodY6rRQTtcu7aAiNWTdBBDlIrSQ9aETU5gfNIjT4wPqcqFuMQNybWa6Obu2zliHk71gjVrTolubziyhwH/b5u5h1WSvEv7TDkRUnpk1DUqLwNO1eB5wBjTJsFi/r3CbELxtbbgHD3AIGWFYv5tjO1skWiJM4pxIV1fJRW03yXSpbFQbsjBy2A/NQMdboOoqF+lxVPxWnNN/P+59zLyjmYsWxu+0ie3C5ctEX+LzSmfy0JAaYxZuVkrMo4b07ZC8MoGhjmhRG6cVec02rNyGD95FQ2Pej8XRYe93zLcRDIU1v7dmN1NO1MDIEmFsZ3AMEKJqgqY5ffJZHD7WeWAyHnHf/HpRMGKWc5/UJ+lQ+JLwbz/xIeJSnkP4aJaeuDc4iU4Q+EcNUwLwEsTTJhZ6dgC2I4Es7CAmOQEqOHzNikIalO6V/XZq+r8MSTT6yFE35ky0LcZg/s+uA12PtuyiLD/8EVMyGZ5w8i/TTw/u7r2gViQTIH03Prcq4ig5XwHNjGQJNNqWS9zTylNSsRu5saacZ+d/GGVkFSWYLtbKSWH42QdR9ZvagpiJmRBLVj4hMGlPTNHz4h9DrZmLLxLYkmVhmPe9vCAwWgdznZBIaUwjNT5kVo3i8dUhBq6sFCmEEOvQwMvZw27TirGOlXz49FC6PJO6fTe5dlEKf6r57cSH4LWBvg2H2FcnvOwzGxgZwcJLvU7zDYEh/hK1HohKcPtQ16d0B5apAYQy/+aCXmHEtPG+d6JzWZ3WUUdV8/0RiEpnMMZfUhPrXHBOqJhpEkANeyZ7fkXDuDMGanPR2eIjU94tNY5F9xsQUx2lJrcG1FWMjwxssyR5o9L3NZ1AAQqUvmG9VQ+aaEWTjFfK3NtUKyPXJ9enl+T/+43b0KV/hPLdA3Y8XLGtiFD8K0d8jXmihZEAhY3mnYDhQqDAIWtxUV+OvRFaPcVzyPy47zW99dC+1hPrv3ZuMfeKlRh8SQgzVWVYoHz48g3xlPNTZsdz2SsKbwzFcDvR6sTa0Y/IU9cRXL8rGi5gabpjFtk1VDty/S0IcW1ItqkDwYXhIp3UWdm4UIllgsd4c7oweIE90vVxTB7Qg975Yng/OXlYa3h1oVP1985pzQSkIApIl4aerNOxBXDpG4Wjgqd+t0xPZP7Z4SD3mdWNeqnXzL6AJINj6Z9pSDS4P5uNPPkV13dCaDH8GVZ1SEItKh7p3ZC6U6wb/QN4Y/1vLaU7PufpYo+kHNlJdfv2zWZ+51/4dFCADDm+obzqk9LCaz91i/cbe6Q2ZO+4kjPp+6tgCLPiFJt2eZO692ousGbbFKz0rPjEowlrqTEMrqlcwULSvNqMGtlbztvQXounhhFJP/I1k1V18iscMpiJWnOVOPKbIOkSTjrCF5WYft1q8C+rlCqwJ6Wv2w/yuoDywfCbHRQU1RHjhT6oYVg+WEoB3KG/J+E3TnxFurbLFofEbpVoH1glkUSTJUUUda+PRO/VUc3pqOiQzyCaXnmuq6BG4NmcWVFKOS4GeeKfVUBOwfBKmrUotcqqt2WvpvMsXAF7dRu+DjG4V4xJ/D20X2ueU6fe2h7bdv4YJBsNKIaxKCv2m4JE3tNeMuVug7d3U2z4/rjkICK5YZnlVrHGtPGlPE36+NlWK8H6HAcyKqgijRvpfiFYIA00bMwGO4MD6ayPQTQukyBNZZYiQIcvIiToWH+nBr7sHxkcuJdBvVVoSxWS7AJN1v647Naj7bs/nie3TGYxc+TL3ej/fFJVXFq6FvrfxWbtbvUujzpKpijBvE55CPxrBDrhQqOyLiXAxMlZAHysjtzFk00ImGISJ8YjYDXIx9/5QIX7HfLKRy+erSoEnSa/i5BRRHEQE0/w52k91qD0oYHHnu8SJ/JCBw0f1qE4lOu8BDeC2W6NLCJihuLkSy0uZzjlhbTo016zGYjcX0SlnXkvHcHNRMm9s8/ccYtpRKrDF14q0SXhLojoxYrXTSUbDkeO2B6m4qF3ZlS0d4
`pragma protect end_data_block
`pragma protect digest_block
8d224c9d3aeedc5febe3417edadc1055eec82bc15d407107a168dbb9a1cd929a
`pragma protect end_digest_block
`pragma protect end_protected
