`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
0Ees1DDRM+AGdpvWhw1CW6XQxRZvwzoieSZn5KAw1gNkQ7sH4a/mUNpwyF2LXnCaLtMJ5CXbz2lXXcGLRA/yn48aa+Hm81fdGPnKAkiL2NoI2Wx4jr90+zWfYsTgKMMdXAKcPPnWRGnLoygSg09FR+pZiIrKHhp0Zf1XorsgKqOWWo7IcEmmzXXs0LODvNGIEytM80PZa1kIKFswa9i1wHKWlYn9tGKKcL6YGniKBMtFbTQglRYQW+GN3hCVoQpCxhWkB48GZ0W/YvEUpLrkLCKmE1O9fa+DMGSf+7tmrLAoQGQrI4RqRCr+40TUwvp50eLSJrGida/z3JBESpZ38fGsWamKVxSKx56ElKaKvkpFqq8f5LPli8GdkOYULX7Y9xXlTfIM6wZPpHCOYy97OkLB/ZXXtyCesKmrhjfVxf5B9A/Mz/q13DKueFGe51r2Z3gOuqiEa+OvWMgNEAetyt6Q5LAVn5NoelD3dS1KWRLTi2gBg9rlLt/YwyuI2SJbrUTWZguCtFJM//c7q0xkjMR3chuQm8vN+0zGYBgk+KneDVQudFKxSnVTrdm8kOfENY4GKxlSOmlyhJpKSldhjhZiQmY9TzFd8bLVaYT6JLoO1hFsgOBWaea70nbiO5s1xI2hhez/D5ClLgxpNszI8wg0oOQC56qTQ/ul3LLp/Qr5TP671kVW3VO9771qHqayi/X71s4vfoD67Wmt3+6XZk5hEou7YOXu2dCNejq5q3Atxr6om4YwDUfKPe5QxvMlsjuwHSPODayZPb+ofzubd6UQRsPDkxJ0cv6/fEUUT2JWQw74KHHfC0/LOsmtAU3n25yaQ06Djhd4yEsNnOHifWZaGmWhjEgkQHm7a+EFJMMCpdDpIw3OYUiQ44iwxkDfF7KMiqn207H9NQG3hTQ4/QyEv0J4jVtpXuRggneA+CkccHhh06wQ+OjG+AsaOuXSvP/fhEs2p/F7BkSn6BoebaTY8hTd/Ayzk+SIOOjL8I7EH0qrl7Yvb5aoKf0TxsfbeMOdmpjmOIqkF3klQDM1dV6qnAkf7w6HMmBA9QaKgyRYbwMBMmGFrQN5xRaJxNHhdLitOu8/foR1mW4/lldRYdOrnZqbDI3V1tDWNybGylWyQbWOQKLb36SXWXQuOyGBWOZwIHR1tA5JEPITRA1hAbyeJ18MvFg5C0UKKrRzgGO+z5W4G1xN3op17a0HFR6cfLEwRIBsWwvEG/qmORce3A8N/QXrLO9+6hI9LV9NEw6LpFrlPBxCAviCTPU4TWBnFQkb9r7AfvCl9nRr52jaqFKwsPCFpYi81YkBfXpdObsn9QVMB+zWM3q+zdCgAy51zwgwm192jLRBpvLZIBkQr53IguVJyYyK50pt5+f5VZz0G+4saVUxjRToR1e0vfzTtA6lRjuBkDFLUu0z02jCPXfE0gqq9iSVxFOBJm1FgYOntgMIaA/TrrL0Rhw+gPeB8FqPz3S5eLdujzEYWcbVHNMUkE8QzQNB1LMMfe+K1UVI+osy9rlusNfFdx43Py4hCg0l7l7+r4zxmZpLsAzH2V6L/6fI+CLTHjzNROOOMRjpIEMeN3wG+9XNEA+mqBMgq6LIyiNKTBlXP73fWh1Cn5Sqx9VVOVlA/6FXybOkrV4vfc9oZj5faajhSz8whoSEGgBr/xgJI4m41bdBEFQid9M5M2Geu0lU/9Wq7bvdExcmKiJj3D7dDp3TZCvEEIKmslIQsRK8RIsOw2h1Cv7p9zdKdxdC/zngYnKcLtS8/9ojIp0xXGvhrx8jjDjT/fs+61SAuZDTOxS3hUV+wO9R6EhYp89ySEgapbRGtK5jgyI/aVMo+bEXemuCYqdfWqaIGvn2y2uVBFPVO9+dWymU38wQbAiWYFjwk+8BZTAgYKDTL97xl4/twv+bEf9iYNNM9jld0gvHgVDZ7OQhr9/8EqPVhQHXjFQcJN9npbo2KV57UZuIairB49Ku3txriWZF9Bai1Ogb4XLA3NN+IUGUMs7GBj/ZTRJnoN6D+zuKWvtMxa/8UJBgixAGweUXoKxQHI9cKmrKOWuKvSTCkVXnu7cUeZcc38xa5AoBMUc2ZZkebxnF2mda8iGJViUMRCJGR5sGua/U/cOjmqE4d0SK+w7APrXBdcLGHrJvejQIWrBShZgL1wZMnqrybIMnxwShzliD57+Eg+xoVlLQ52kQValw8CEEZ+RTvLY3I9PA3ut3fUZvNbl+Nqf2f2exECTyf6zCSTNLmW/q7JOhrU20Kg7d4xVJD2K4z1bSdcQc2q5h2xowZT4i9X/EJZFYdSJqRknLy9+3bS8rJT0Wq+ofwbJkqPC7vXVImVbZnae78sDedD3/YiurA19Ique8XEeMqABEutKYfftCA3Z7L5gYZQe0VZUS2yXX0VqLJYEQSYogIIU5v8Oj7WUG0zFlCdZ2RRpMKv5Uk49ztAYDs8a+qzNQvwTnPR9MrJEM3SK4aDitJp30RmWyqHq+VuKRDZFe9xAA1P7xGoJ/nx9saXJLX5nVlyqZAybXYRLm6JicZUDdjuLFM7iMs0CJz+fJRUQ/a2voRdqSOOSVMZTxJUexgyHCkoblGbVqexT/1BZnvEGiQIkp/MogdZlkE6OdnppyDQRmsSywOT0Lp6Ax8xk5oWAcjEsRhEwdJEcZn6oySJAz+OkBkkSVXFwel1WXhoQOuLRm+5vnfcplVNWDpokHAOGJbEsn2ZZCWj9tMwZCzmyQfW2eDW7twYqlabkugYJxB5jgA4laL9tLXUhVKOiKd+8QnkQPaklnwc4uWQs/chEx3jlWCvUirhWa6CGP6K2DhsloIVHt9vA1+RAvDKM3mM+kllxjz/yqxgfuGsjQVPmFstZnGtUiPIRkVTYRQ5Jphvsses5T+pKnQ8eYobUMNQfn6SCbLXqjbm85MnM95diIUKjaxBFvvFJcOwhv+rzatHV6LF3Cfg6lReVs0G6GcADJ0tWbAiHHoscP7TGxCSNhpgDVqyxzB/tBaVrydiH/Ed2q05NuP9eRJLKPglfK9uOUPdP/hznKabd2xdxqrON6SRuBc1jh6opzi1al21nwDQG7T9neb6/zJlyAZvlXIaUPEMYT3/vKvoce47YON1I5tJrG8/Mq2tKJZVBbvwlI++sFzc1SDzETGgY5+TmCGBkNxJ+AyJpi4GdbnPhPgFwfqcnaMKTa++9t2qDUlHYwa64RIFbVAyrPZ25L5OxEDyXVGGAZpAAkBDSf6s4B8JS2j4+tQkMxBRnowhGQI1hkfm0wibb16SS+JVBI/ux3YlEqkz0H9ZL0YnQyPH1j2EYlBX67dvW5Nf1wDgetSY+DhvrYGF7WRLwHAnQOvWckkYXutxLqg8HXeVbRkSpGxAsw3VGf024SELvNSTqSEZo+jrMsAYsZzJ/mPWUDbJIIEdJ6jXzgcVkRhdHOuTr6vCpAJDZ7gBciDgMzgHS4RY1xqEuu09IgClFi/thmOs4a4cKsRLfOv62F2veKs2JQjFV3YcNG9Wdc+7S0/umhfQq0CBrHsSqgzpgNeh4FlWrGAne+Lx4cGPTZudijnLPq5Zff36xp1TdKg3fDR82ExnY8z//jTtykDRswCBoQ1iq63Y8iAykFXVRQ0RdNKYq4upRKLmStjGdqC8Gv+6ZZxZEzOHBKVOddcuHHcL47+G70915+bYtHJsbneNRD9oneetm5xMS5q+dRPIWfhliG0kOI7u76OIoikf2/xBdDBAP4fLhEP520XfWMWaz6WkXjKGfYjmLGsQu0dGM8eiFrRFLQva8+YiGeYJpvS7cKJFTZY/hvEcBJFGgb7XXv21GzWN5PFiG4J8vss3GmlhwXdeht8pVumQZ9bDR9TrLQorqmDwByn+CpHU9K1Pf7+MC08ZDY9g2TZ2H181LaHXLmHeGOk8XYiRVZFRZLXJJTZ5soUIT3WeKIjSryFsgnFkyphambZqU00aLeqA7ARWJyV8lfeQMULN+3AfvP3cSvOtRRc2CCQy6D16ZWaKTdGmUTuHo8s1C8nxDwTSbCYWcui+tP2HzvU277gzBrcy7sdPpVltvG6uE00fgJEd1eZ2IPAk8WfmNgi1SJOolJvWI7UFuDczecsf6EpCjQVlQNe/MSZEkejiZHoPVlFhe55ciqXNy02vjzqMHESlPuZeo2qUOqyGMMxclDNksV2jM/NibVPFgdErBwbxGE1QKVno1l0tKmybHd5nJZe1bgQ7ztP9Ahp6JPDnF0L0NH6BaQWsCxJP5e5RerJB4p3QpilgkywMAoy/neCTfJQ6yt1o/oUDyCdRb3xObShAlLgzBPAikxGSOUJSPFFjQNNRQCLurMkAd1BtctgWiLSNZYX8QfbatpkgdKGU8SvcSgEeOmD9iHVBXdQED/pzm05OghBnqWfk2idpPI03FEA9oviUnkXutvIb5lVKaC1YMppbNsRXxPJsf8HHEE3GW/XE7Nof4uLbMRddLmggZrR2WYNk6EIHpxCpG00JSyLPMJIEyRmcIuka8gxkz8lj5Zz6NiKzHu2/WKpJPfMa2MsvGUN8RutOS1Kl3CbuBaMrXM4qcEKhCANK3kkahiLJgyUi0fud+HBVphLido6K/CZQqqL962tLuJkgMYvJFRGqhsVm8u/MQTr9q0nsSbCSnUlhXW/SE0fEil0YnNctSEvd8cFSZ9Kk8nHPHgYp+TsbvsRavOg/cIok46N+nvYSAWmvtKtMcd3Rmc30Fhb7IE1j2KbXiC6P5vgNWnntsceXN36gCAlz03Oa29j30FK3hoyCEUr62Me4R+0wigUEDevWjeU6XTG/lropDkxE2Skk9AHkEtAyDe0You9ayW3TrKZ6LgqkrMwj3xCFVxkEbL4clEpITlu6k5Sjm5ejteLGNMkgLa3iE1B4QP/RsphBvqbIm6/eqyuq3A12faCUfGYSCU37ce80ZaG7hQoR1TR5hdpi5ndiwbhpl0B7gBzm19jtgkf6HKMxAfxo4O5P/q80cbEvcgBE8t3ivGVD+4P9oF/OZ0UPc4KSe37jqx88f6gV04AGZe2dTg9iANLv2srK0CWxPsSysDR62XUjKv9LEZaUdF7W/42IJkfF/sat6D6GHQ0MSkbdVhFENWpL4JwXLjRgSGLViPef7Bsb6PSxl6Sa3+KwYMC8ycFCiSvBHAsz6NS5kduTs4sPQF2yGYryQw/alIghTn5ARfxOj0BBsK1UxTzLnEJqwTiCiaVNiLPAQ+5lladV7zkzB/Vajlxu805C04pT1Nim28VGb9cXwkWc0aWRVAK5smitZhZRq3rIQwb90AKBrCEk3KxsvDpZcbOZ9ECN3SktZJ9zelrcl+wt6G53Ut9oxsA6XFmKwG1p3wOh3aEnPTlsdL19WttojlQ3hV2dYaGM71HEolebtgORREjgUvW1ruh0OWB+S3OLGQv8c10jCuPNvQ5ulQn1UEs7IxVtMVF3cxqCpJsLXKBLJ1MGCDx5KPnyte/PceWjAEzBc/WePgeIujU3/P2woX6Kg/49Q0UkktmCrGJZqvai2tqx2LENDxH1hkjg+T6+WmjP4lgUQcThjYh0DGPYeP/jbo6ZFTrNyg6Aaz3T/BS+didMDmE6F21ZwKyyrCH1w12uQsGvdxoKJB1fdrHDmPgMpXxknGCjOsfyRkCY0+dHV15DXcSsqQaSfqh7VHNZqHGvkKk2EIgH+ORVMgPScbhzaxwn/wP0FdkkmwoHUDjc/xQa6wV7hVWMkzE9QBPrKrKRTTrkR4fu5OSid1EecpJ2+r4O8C6hlaPTDgXuvAlnS1IDdct+k3+vQawc9BgGt7VB6pDn9/i8g9X6FCY1o195qLQ+1aZ+s8GZVU4KkwWYWt1Hpgir5uKQddHSnrPcWkBuVnqZfeh+yL9ZzG2LVHIJgPtTl11IlZG/CZgRu1Nc/HJ5hM7eBSruSKbum+H814Fi0rQvELhSOK1olgo7uF2TFfRgJ/dnY2Hyu0Q2ErmkU6JpEUVB/y+ZfGZhpdwJJfFbCD4fvST/pIuIQ0mp2c/RoKsm5aiGzVFPcF5oJkUSSPyzJcdjUSAB7RwuqDcjVWf4uH5QOLbxid45pR3xt1DD1ZB3N6QMEuozOiWT2mz2nDJzij4eQbeePx3OYDVDlzYZi86QGECPdDYKupYW6ouxJYMSy2U6kUEYzj/jEHL2ipuQRoISeQY4PjIUWauzGN3Nw0IIaRZtF/k0Q72p03+VL7dO/tUS/sBaJ6+w/D0+yqQpD84yhuz8SOZGX3WnmlO2M2P+QDSXqVXztpTh48/Tahoed41oyGgf5aRuEDVvzP85uazIvFNCDohtqvZF/I8zQWmDu7c1GedWTUXvTOlJ2hhR6h3dfUJO3caT9PrP0u4r0B83aYbbwUPGDwZB5WjRhP+AiMIdmzSC5yw5m30L8UmmvTzgJeL4fF+ox/PHY0pD+iqTZo0aho2KABQ7knXpgs0hBjeVs/CUwCEmSutzaQ+ByBkzNFDnLesFEBpDsGkYbwTOPKAtRxPxv+tL34nro/8/9vh1ybN8Ls6PVO4sy9OZt9pnyx9PzIZ6C1BsG5I4wC63UglI/K0YDAU8yusdVY2zF5pKhePmm1wVIIIcs3vVs538EMBj9O2pQBH5F/D9a5f08OqRSW3WVtKyJlxtJfelbSi4oNipaheAVezaL1NJq9bWy/Y8E/Hl+2Cd23v2PtoTpoi8uSa8OIgluK/TWa9p1DXk+g2r3yMGPmfXN9ohXRuDIUSImdKxC2rHBzG7ZkMlA5No7gPRW49MW9XVCrJrPswmOj9QsAfXKi3mRL3QyYU303CZ4MpEyHxjt7urVhtavbL5LpRmy7ZZ/RLVo456MoC3igmS+S+I/fd1pzFv/ekJS6ZvX5qmJt3tPpA7qPT81HPPU8NA1nWEIPwlvUYaWmR/rcUs0+FlLJXuUwnrhEOkeyAAbvkcN/dod85dV6ECY2V/dYL/uXNvcpEgjmOcNpzmfFWyGe3n/FGtOvuLsUJ0PpUrXo+k/QKzqVnobRevVAI+NClrbudR2MEi6PkTNIy4chiel0H7nxdQ/ND1XvBXCpKV2sENjHKPGcCQkVI2WgQJhelrTlqwJnhj9TPxTNJKHURTcS1ihGLZ3J8Qqc+h0X2MrzMros/B6jUcI1VMX2HL9b7YnYweknkm5WWlYFCeDAbbtjZdGatDGQwCf/tZmFk8fZ6Um5BbrcTMaxYqTymeqDEQD6/jOERxlwE+4H2zluaqhUo2J0EJ3Cb0hBhCpwH5D9YCv4sCgDck95VxWKRBsGo0y+AtcewzTRS0UVyFFqCJjKKxaD7fuvC0ZHfw5nuSE7LP5wyyBnU+3tJO9b/2waNemNf3ZFFpxCElvOK3VwTaCIUqvlm1mz3Z/owJS3RiDCVP91s8DqOg4pJFkXbtrM7kp862sXkp2rAE0Dd/jkQXOEUylicW+RcPY/9hkW2Rqcy7x8lngMFT4cy0pFYnvKgQfnPEOIl9CcQ9Pqpskjt/knPMATSLUxYSUAUEO35PK4MxQQj+KPtJwqMMn/4t3bTNPiigjOz7avFB8kce3jEgJFznFxX429WY9vTQeWhTemIxbqfGvO5QTjpzz3cOZSlv3MMe5/tmUyYU0x37MeJezNArUOUDD/DhATbt/3hUYGaC8rtLnShLcyxNatIAqBQxBVJByOqIhfdhtX3mdyuJlM+xUKRc597Xw3RAmH+x2MBkOi2MUhHeL7dkv+baShuYsSGZK8TbATcI0e0v0mJin871KbnjdbLYHpdNcr2wrZjfzYByjTSAORL2RBx9sk5JQva1vRkqihQK7LrHDppQ85UJ5KjGyoFiyp4Ms+ywVesd5gqNK+MQxIVoR6Ryy7/8VCpk42H8heirJ8ahUUajGxY9ECAxLlg2nyTSw6PFb7PB1T7fOKjcmdnRq0og4g9DxEasDblbC3iO/ikFJCYtuCs0edSDbcaWf6iqiSVwfI4KWVzWgVV93+lDtBBOJ08low54SzMsDtePDrPBRu8W0Ug4C7FZDqN6Ijh3YArrCG1VGhbyASg0AAEhe0cMFKMkDRWk4PLDHy2rxKSFVGczxE5tP9p4lOSkcn6gn6ktINEO02PM8uO78adkFXd9oNGcaPnCSJrv1YpkIqb75Tg3Br6dP/hM2aUL6DBgWcNLsiGmvvpZPrEFqTo+8N9aPyOUlFQ/vLZfCuK8Powao3RqGuUybYjVj5j+vZ8YOyw0foueyexAEhw/ufEvAEN2xYaQaQFObe1WXaThfHKVsgxw+ZVy+VvCOyOeYyelFdSUoAp9PZ/ZZs/1azMDlpPBlGj1Q91vbTuZFxc0+uD3Np3jdm0E+GVfhep/HxGW1cYt19U/M1S8Q5RVh3dwBX02SKccyFvfGp/zjcT4PWcbtD7Szitzv9zr5WeukIlyxbTwhBIqwuRJu1RGVthnQSeCkQDeK0LZl2Y/1v90lVmIwiMw9eXob+yQpCIl+7ymZ80lv8N9UYxC8kYyoWfbRczduocFI/GzllkaYZQV5HSvkBIcRbCgeLsfweqp6qTFhN3rRAosFegTRZtGv3tbgcXkMC7hJuS1AEA6d8QowcKivOFjE8cJtLlBs8EcOXPZYRYwoU1A39y2KqzADmkqJ21NuWknH1eNtIzXya33lZ/+95g+Rg6Xv5AtRwCkwoHjkSYiF8+MzX+lKDmXbyGYrhu0f6CeGVmcIB+7i0VM8mFC92u5zsE2286yj826WxN1sixqHrD+SlqMqzwnyqb2B2AeZ+4wXa0rhM3gK2KgktfSqgFp2n9Dd7ONlpH9QWjxyQE6yMwk0pF2+x89inj69JjXelQCSTXIY3bj9MTxyKg6QSdknn/VXoDYXEaIOCoTBK8TQR96xM9ud4g3ZUG4QVVhDLV7hMo863iGHddJqjIxE2yva7P0gTx8h/7phJo5wp9rfHeyEzpYUocPomRQt8BmMt3Zp4nPDuhFoKIck+F9UK1KZTV5/1usX/068hXJ86I4oeJAftpD5cyXWTfK2vJSUz11k7RKW4K0D5IcOiGh/2iHo9LxALgW7rd/SE5EEL6Mxno57K7W83/0mm5sZ6NvUqSeyi8LdsXffV8EMwKcAevYgZaazCGjnjclHrtdD8xPC/kinjuc5SV9DLXJs2N88WA3jtu0vRNYsn5JzNlroaiw0Ba5EFqnCgwlySA+sootzp1OWDlyK8mjUXorRGWQmN4o+HHTz77pU3MkgSQJXdaGlpM5uxGcM8B6UukQTeYVPjp4MpO2vGlz4CNBSBjRSdO9IUOY0ghtHEypMK5c67jRj21kVYHF3NwyWynWXPfIRYBc5HYx5+VYQSzKhaqTvkdv0OMWzKO8xniCcussGJZV3LP+GRJ6JZTSRf7SB7xPcvnmLZUAYmnJ5eT6SQ0tL8fHGGOu23FrvDfZQ2NRGICglcIuWShWvFU4kLm4P9Cn4nMa0KVsEySXEbgj1LDMCFMZj+rU/nAk6XTM8/5w66aF0XJu5TY6HYcH340rpozB40zwjMHsrnkPTuoRxNKe/8bjuYElJDDh4nZnNz+4x7rVaLZ7mpZmEcRxooz1Yydoh3xsOvvtrMeyU422xkoQU0wX9kp3AVOXqKbNHCZhVWG6TteTREgNK6I53j2nzGeLLUZGbwncEu3L4xIterFX8E47I0H/whkqRTun30C6EsLmqMgD7rQ+6T7U/3Kp8n1nLlZY1UyypXwdkdBiZxWQ/IRI1kH0kR3t73TmDgbajp5dOnLJhgXudycdmwYer5rQKI8TDLQuhLaN4KClqLszXIWuYVzWCffxlTxRHjtMWV1IQiKrvKhfIFxhs+E/5zYYgH6wWpVajWee5eGlBW+krh806QxPkgZtVIaN06aZPVPw2e6JyOnhfesazVVbDB05DWyqK/8y5CisQB5EerDGFNYfJE7Pi416gGm8eaBzCK1wUp7VibnI4/lZKPZ8K+hGjzwybllkoShJdsCqMFU2rlJaLPya9BHMpXwOc=
`pragma protect end_data_block
`pragma protect digest_block
49246ab52649e37ddae2a35c1bbac486290a02e4522cfd9b2b0c9e5fddb108ae
`pragma protect end_digest_block
`pragma protect end_protected
