`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
5RL/Gtf72Sb350TXWhXoXwkRCRmvKwXGeYQ2ZGkJ1mv5XZAhE2nILHO3BZCy0cXLX48qOvt+L98J7U7JQpBawmxkmg52ceRZLEZpc0847OvZ6OsyXKM0kZ4IcdANcdE9UZlZe2wpUMdlnY4RDvaj0P6sTgmP0tkipP1BapkJBB6vyCIWz/7K2AjnfalUmS9Zpq+k2dpIKC7Togo4r5wJIfhaY3vIbHuYXQRJk72S3KOhfvQqbLFQskGAdqKf6dyQqiatnAB9NJflFa+wQRNwKtF/iamGzBG1UezTCrFTznUjK5Gx6Z4HOm7yJrj7tOOmIiUpN+rqHtuRc6+MQIp1d313YgSLOP+o6+nwSSiTQ9IyQTUmvDQjHNGY2ZVj+PrWxrN12ETDiB1Z4RvezUOlLE3IfX1HyBu10fsmXhWKzAaS7AGSXZYMHkwCTTgJRssq7Z+NXW4JuCP9+15AW6SYKQKLpUzH01LnpKpk3U8oE7k4DBygI0hO55391M0lxFGhAsCRNsEAyvxSLwiI4oxL3taN/wo3MDB3abqd3a+azpIiyc+MPfpkkBNoMt/4dXYzBcHY74cK3lZb5NfRpWHdIPGzqex7xVD/0iVT8wRag/2/MuDIKqOxYeOayzQ1ANI+GuaVirDNAcU2oh9IwnvT5iXEzMps5Xzokm8BnW/jmKNma+nDGbEQMmtMK1y3YFIDSZ2xVWCu4cd8TAQMd4c3eVtoRqd87ReNjBPdOq8Fpww6hB/MH/GzRutMKuY3pHrovRmQLVxAuW5eTra8S5yavFzXq/80gKoQdcCCikE1dyzBG16i0eyuV3O9zt0pLH4kOJe/WbYctR0TIk+Uw9N8Trlpp1cCyP/pFPgN7ccaZPY8RUMO+zLs/dGrnQQUJSNTiu0H7WYW7/NIX0WQFpzS+ekzGwsc4QyyxTNfflidJh70dNACUb6Y5PDtaWxPONickd0Hev+5GnjTiBwH1RJgrWv5Y7cLoQBzMHt5od5lVhRuK62GVbXSCUmc1jchJD/q6YjHXPmIdz7sW4GAG90HBnHr0BAL+u4Y8rWj0ZfBweOrBOGkF8kpaCDoaKWZgonYz1ATsSQejGlEjjUkczipmBK9IwpxtMrTqOYsfMYbap7WWzCZ44TpU+utanIsGafhW09uK0KbG/NZyXiXNtGDQ04AHTQNs88Q7zkYOaQj6SroJ/CBw/5b6r595VBIniH8Gjzq3eKc7OdBI9zMgdzrQ0KCKPhHTznacGAktD74JrmeOLCoNWygtZ2wPUbGRsuFp9h4pNR6IGsjJ22NBzUF/exusUPtzqeB91ZvrzzW3IFEtC3q5HLL4aSH4fvIAO1KzVWUK5Nm9gH57TD9hOUwZtMGEzUOO5/ZSrrs0/ku0zIbyXvUJJ5sgmNBaTTetSG++459sGp4IV4pi2LXxsgecvsEKrj5AJyYRM1heqprUNxZv/UCltC9MFbWn8Gr4sZVzAOYsudO/BnRTXMVpFaxptadDVSazJtLtz/IRbeCbYeJnSNSjtTezNprG0DWwQFVNN54NziYmQSBP9Y3WGp35zHt0sFaTsCA8fNYVfOjaokMHUlAaRhAUNsbh3Jnk0L2LlSc6YPmwQYzg8jJjqsWqBegCTuE0DqmYBbeGyH+2v0IJ6nAbNd1iSAOJsZyairRWOWnWcHeG7k+VKmWnlIE/nTy6MuF6G4c0ufdltXOGNxhCDFom8yFHE1lOCRBWgoo+KSPQxNjTKjRF5YjdRmSSa4Q52Oo/LFFLVwttIhcwEOK1x/zKlraEXSqAzbU7/7EtLuBrh4waIDyan7lTVeeIiEDM3fLJuc4gzY8bL5vPM3uytOo0DG0fA9YFID5Wc6SNC7o1dUdiZSydWyPSqPqRPDN+nIfGM+EEy8IOccGr95KsuZCeg7X31aZ6p8ifzdyWQhdTpxP4XgB7GZnLNAaG6xx9XsxcGAl1+J4oGhBuPTrlWQGbvLGcA97udgEDllipjxurpFFdfqukbWeFVKlFX5UzOPHHXgajxpEJmtn31XcidZAxj9WcwPPb8HcB7OhfAYIl4tjUpJK4SXxyvFmO8XCNjgy5UhV9HC4Joimz/UNheQIY32NRrnz/3GUcRJtLeTGXfcNN+ZkncOpUUVkhQRB/hllpm4qzBpeZm1xzly520ubvkmAZ3WAanu83rEi3tiVOOkXA9SmSip/oEtC1BN3iEZrxv4GudL3Ef9P4XStUYIl3sFUz2LDheV8QnlXtxEL3e4y8x2sYbr0LI/7uYizAgPCn3C7ohdgiM+x6+z6nkRCeUrdtnG7XqjAxK+Q/tDDDFUQMXevLvfpAegJp6BoPyrrEaGToCQpAlGmi20wWxNghRZHVZ05mvbuBFm1MglNJZflJ55AmTVJERqVqF5Vv/kvCw2q3a2Yvj4Dn6d2d2yWJBCY6ZcEMT+2N3B85roehsVGSbj64knbX+r7T18Sg5obY2QPKnZReHEp9KB/Gz+lVVOb8w6ohFGZXiNk3bWY+rc9bxchMf56m8YeRU+61st+m2ICczPeOVs4V+jAmOsr8faR+XbnxuPb47GnzfzN/J5vmNOlUgWUr6jvp7PwvTJcMyD+GjIMOEG+NyU2OIf15hHPoH3d0XEVFwTluQ8nxwnJsFAY3Ey6sp9+pWfpZ3fd0r+TUIJq72I69ySvzGnFcr3Z7UMyayhOPuLNMS0LcU8Y5Vqgo2iFFba3Xp9KBmnGlSq7xtA5gtK+qpf4k8/HRSxB6RqUbn/nBkQrDP9vidkmFZo0amgf9OKk4f6CiFTEpWOrUBS5n/GVl4N32hcfmU6XEr7wY64tlqnyD4bY+mUkLlgjW9MOh9azsQi3VbCa6ZwvOwk0pqkLl+ySzrDpbHet2KCjx3ssQsig3/ClJ0nLo8ftJKiZJcr/fuYT8T+fv1fnRDzzZAyD4KDf+821RmdLg1WTPVGg9aQPSZsTs1Quy4Ub6/FccCQu2coSRdTI23Ps8k81wkg2t3WcoIrmkddleN2rRDc7izaUdzmMM4NxoDKp0cR3eEr6aH8BEQsXke0ALKbNIKW84zuEoeHrw2vh4oXDggZJT6XeCK5UkEIKoUIkZl3KjaTRjO+FKqv0sfUYMd5j3j6IkkTekZ4NULvl8u3Gzs1iGS7ZbtnRPevCfDm+U3+bHhluzuW83F5ghCepGwNx53K3Q0xByojTrRV8rTPIZ9sXfhOjqXELxICd9YQuUF5Sm2dG9kt8uIOhyGkIerXwEnRrmUhlN6//OKWxdGk7gUW5Aw5uCgjdbR4bCHcOYgwKTh2doqfc+IjB/psuYpk5QzD6NRUkY+Lnc1/we/66QCfIounqSp/IPXO7j0JU5kqPaH2o8QwWeKDUNq3GDVrzUUc6W//TGt2NujOkvWviCQ4Lfq9+aSdyNRQevB2Cpk0BHY16hCh6RrR2SE+hcCW9v5wikZXJO4bKoWSobYhrCizfRtVIMtDdSWHFKtKn+SPMdv3LdmxjxTmhcSHj9ajvNEu8GGEkTk8pIiLTU9rlvz8X0YvqGESy9j5m5t2KUnj3a4/CVVKZk1ihImjLplUYG+4etrlQeSLwrCoen/h4QfcJPoraZW8Y9bq6SMqbIWC328/hUUUayNetIOMl7TP7vJYD1Iom7qY4ciS8EZ4+zn71OyBS0WArDE8g+VYJdca+sUO3+xCCSy9tbIsZ3E6R0qv+QS+LkfpHnT77TyQoLQK0/u1BeZ2uu1jVPm8ZS1F5buABz/oPGb1uV7PkYuTlHoipDjLlGV2gYThWhS1bgET3YBF0eUO1/xvf3Qe2hdPFoMQ0no8SdT0EZUP23VPE8j+hC+Tk7par8RrFTkifJzrlyG2rCAHJIvC66P6s1YJYl2gjT8pnA6YLQzrpwrvbzSroxWpUwH5brpv0IjzPag7/hFxRuWKJULha/S0xtc2/438XbCd1ZbIUHbIGtE8FxTT6puFOuutlVwfI4eBd9bAUDVHLUwoBQYNfkpvkFfOA+JstRZQkNdNwj8S7BmthI9hxVEdjz6NAwgbQBXB8Gj8rlKNv/1m+42Qs0Yt9iIQlK0Xi7XeVVU4dnn/27XfJpUJsa0pY5WKmAMz9BtbEfzu2dbU/VOj7OMzjoegSsKamaxbsBNFsK/ZD1IImfjAAm3+zjGtqSvoewKVOck/w79NaehokJFT2EfR1irME+YekmmZvkFF/ZQ9ATuf4o0LzwOvZXoPEW1wQyslgapjxvNfuhulx4XHHAfqtzggB6wh94omxJBe1uGgAeE6Q+DcmXPK6fpZ2GXyJJ5ts7MWnXn8Rhgj3MPx1SqZAeJ+/VtRf/7EXV2HKu5CARBzdwCpSQVussniBbOHqfgD1LxUtxBsMNaFUlv1VhFSELEG/ngNpcSTm5sHZ5Eq/mSl93cNeNNV0zjGytkQ9hyVU3jdRjMP5g/Ti7kDNz7puJuh/YImCZCvwTm7bB2GOjfUJLyeUCXxrJvcORNcKpy09f9PGRhnvThM3TeeQppEXLxG4ZHFGo5Wf/1Aa4Ntx1OcYbJy25og/D4IHZEFyi06WWqeBfWSYcZoMESYSoXHD7xVKNi/5ECq2SVNKW1bE0dxuwottjX3uJVdocInH0yiSeGt2B1yUK6iEQRj4OOHNhUbKIuJDrlJtbNt03vW3cY9N8qKL7JI5Q82oVqXbgwGFU74xqjJ7T9Qu05AINnk7oavurz3cBycXPXxtMjl4gs+UDeUtqB9LPf7z+9+D2LXq2W/lg1QVu0ywyjxzEIjJt0wrak7spCgNgBYG17em00UK0+FtpNXg2H1YJ/iCLFJPYjADEmPmQeAelILCi+1O1wjzOyiJKhv2XxJzAvIfJi/RwY3WBJHWSNpPqzdz9aivJ8w/erpDeeWdKfMucWoV9/fvQLeZd+LnSSHdpvavDYKtnPEAQdoVvut3HEovoVFLx5Wn+5Y4fw3HKQGjYfWnjmvFcxC2IYEdIUoBGNrZvWqpZnG7GR3nDkJwFTKbNsdfzzh5k+iptshdx9tydQ7kZqQ6o2m4GC8unusX/18ijxuEr5bVDY05typ4rRRS6OlbJUyTEGeOb0ScYKfh01yRo6x6OGlIUL7+TOnX5MLld5FZAQl9s9HaGyV3HgCr5fNnwaSjb5cd4yFHHlHOCfrxUIaI6cXaYeacWPylFuF5/9xnZZ8PYWaZvGbxziaRxBXYMD5M2VZoOekIZAeIIcKmwghgkaQVxvvmSztdMzWtZfRWrQdAHAiKABNPbQlX6SahV5xJp93xhY6mIlIrBGCMCUlknvzL/taLzC9uHNOCw3ttLThQB6HYfarFtBuH64JK3ylLEd2/ofvM9zc18Kb9ANWDDvPvqyttc7EBVgW4oajJ86RycUNKgmpO5m8AtkZJsCEOs8amq2EuopjkCRdwrfHCQZ6GAY5EZu7w5w4AUQZNP+dhRlE+wD5eJvc+juOR9uY89QVhurEOllXpJwgVlh9xFKfZFfhhTnPqQC7KpR0uGRPtXnu1gBQyNtd2h46MszzdqeY4JbtBOlIwtvYL6ZOQUNACQvllK8phYAlJ2irhBzQvW3p2m3nTeTeDo3+YwIPNwfqGZ9qptyZ1DL6PRBft6bT28kaYnf99sYE25SaUHzQTE/a4cxkC2+7RIGtiUGcHP0/LaQ9o4KZCmhSPKY78JPLCx0poo54otA2XMnUr199oE8NgWI/BcgG0dyU+pihVfq93VQUxTkPpumzm5mfUarVpJHQ1J22mcopfAdgWKvrB4YbA4q893HdeXvQD452Q3PFXWzJhTVOQI8DRniDXYMoLR5Itn92JDRONiRKNeSRnQXd6JX6Ju2bTVYGqcELiNR6yVXwp5i9VEfYbIholv4HUlQ+53JVuxpT8aEXo9HUTUd1KRTH0CHMaKyJQaRw9RXRTssxO4bD/v7Ntp1JVj0vDRtOziDmF1Ln40E9byxTGidXEsfj7SLx9yHp0NtEIlMzscVQskXuXMXqpPSQnCGnILJYhTy0vx3/OmK/3XgjPNOfo+tCYKRYKnjlSJOPzZQr4w51tRuKJ9EDw14q9AC3kAhnNu25fkkAHdpdSe5TQMc+We0TKQnIw6NN5wx7t81hIh+fduDEGv0JuI6i8E2h2HZzxtJBf/kxuOuwSzAswENY9sNVJnQN3NUY+NcgeXUk8NhaKlboJd7CnYWpzwSwDu6PjQS2C0DHKl2dPxIIQlurBrCOfJOsgVLkYlhivRSkE/J4N/E1/BEsE6GapRp7HlXIZLnqXWwZfPpv5Rs1e1z5XfpIWOUhKyiUukPEsFO5wzaUavsy9fDcNZlyFb26MYpEXm/gWO71t2cdSe7tELsXHdc7Ir4d6/O95KerAp4bGbNKOY51QG9CaG+0xHlbbI7CMb6kd3+OBX1ex2JZVux4AaGrRSNSX6oRWELwQAu9auMm6vKXRr/gAAtCWyorjfa7uza6J4JrGLMC3xrcx4iVfYAHnY8HDH229ElY1htH+U3Ge6auhyRqxBWxCSHT0VRNL9F5mdAC0PjSLHdPNf9EGr6Jez1R6ORSjUAu6j588kK6VPTl4uhNA35tFOdrIpnUHp3Sieej1HXtnNgDS5qcgWV9FhVgaT7W17jFjmIV5/3DrZIlKn4nRG4lX2D4wekD9wE0RvE1bUvUySB79qx/jfn4tAB2kAPFgyr3JP+6j52TqFo8mxNgJ+k6MD76B28OLMR6PcJllVSSqQxgkyYC9kFG0uOUXVBQuwD1FyQJxGyRFaHTFQ2EW/qmvLGaJ3cnsfg==
`pragma protect end_data_block
`pragma protect digest_block
65259bc3c84f79edb5e70e13d2568bbedd6512958e864cc69a7121a4f9f30665
`pragma protect end_digest_block
`pragma protect end_protected
