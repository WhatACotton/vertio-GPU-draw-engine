`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
EXrp4ZvZ6V4w5r/ZC1x8Rm8KsGhVI/XevocUzRmqTOUAYk2fwwuw0B3xpKBrdcieTxPxf5Bk4ZciSH1PVMcHA+/eS8ftNnGgKoSAKWOXmBOUiaybrXYzIUnmedlCul8sc4YbZNJrRVjvfkyK934mRHReiR8eldXBvVflr7/v4HPcN4ccmV9d9J1PjP475SAWE9xgT80Y40nuUJcAcoLUxu9dzzQtC057ktO4XOzzVq8vR0QifJrCvIENc8NqYvBBCxAISRK/SuRI+2sCCXp+2Ij8n5VWEdcq4yX3wfQrxNOCZdAQXKP8UZuqPL1alw00EJsmgWsCmklLtD6tkejcqzZVUo4+jRJ0c+zKkMHgsoOjxm6Uzz2qBqzoZQN+5hofrnyi4qUvY/jpSi7SgTbp7c18gK3tHWBDJcafPO7GzVEF9/UQO+f/2Po25d+BW27e3aKWd883k0GxkgmYQCKpvpwPf6FClvEM0UJUNrEoLxae4lOcnMW3onpRcxRVMByyDgDtBx0XDGnY83xaOICVxCG18hI9ZMgrZPSwQWuGsbBBABIfTKvwkCTDz8bJSORtxxlr0Bry+lijH0mAGAHDitfh2aHxfiFVJnpy0OmXUPe46UE+Ro9MVCSYKRx3mYWeQmQW6BBAfaAIu00ErYUxtXpnCWqCfTLmuUUrVLt+8+wRHIOZIt3NNosWm7PSDmIyHAFjrlyZmL1XbQa1bxFbEFeTmTDebiwhwdUvhXxxcFd//kCb81Lq6ht16aFmlt6YJyE2KcWsT0JQn57uPdQk4Wu0Ka6IH3fK2xuKd1AkXbNwi5B/E0pY0+1p48skv25p98sQsx4YU0g1n7YrUjvv7X7aEKzMVFM4Q5cWXUN8z1eEUbxSycojgqMQ7823ZTLYe3mCrL01nJRzdLTicSUItbcqXWvHRevfMq1W6dktHS9Pgf9I66VgNk8+bRkUK4yUfRapPHdYqmmDDWlapVmQGN9gKfI3fxFvKAslH0LWXOMgWjCj+KLyjoTnsijEniY/12ZigrjKDik9SXsGaBbDxJuTCMjThkoB4Cd5yf2NlTrNL6kcJ14BfwEAEHxFzl5zGuUpSD5ICLMbYaS9PZFdhU8XJGU2G0VIYGVpOOsVWUv0hdCZGp+8q858ucr0TjGoeRXQ1E9RvH9HRtjvw9WjXu0wQrvW4T7grNuLTUH4Ro7DqhMcjf6zxFzfgNGia7R5xavnivcn8K8PimfZ0EPTxJc48sK6DfLqSJnzm0cLjyTWOSJmc5HIqOoi3HWg0lhcfocZdIU3UBmOJ1geeB5R5IPY6yRryVGVE1w5NBcKORFvI2S6gHBnlc53YJLeT3/LsNF/ddJFqu4BOnx+L0MczhhIYbVPE3eT0NMojNfLCos6baPvrcG2MmLnsP+Z6E2brNdIBBIO7fNC4Fr/REbJ7vErffKaAgMxlJzA+bMWcYaowk4NGdW0Xo9EKO6R8au8K4iSXwb6h9dAiiyHTZMzCRS8/gMS+MVHCAwLeKjmjl3roEDD//SIQhjC2a+bpvEGwvjFRQP9YXU+0cOKqwlW3dngKIQK76fSLcmtSzurtrmm8udMfIdROUNG2U5A6qYeWcSKB7nzHghPCMYZGCCElVbl538sekHhKV8cUSVsuqf/UFpDBKv5KQ2TuZaghC/8IH/kZeRidzPRsdkLh2moKpIxZOHSJ6rSsr+eoL6yUrQhYZdoFCnhC3L1QmpR/0sqg0+uLtZlc+cm8YOf7CcYRKP2pJnFg491M8FIZwWw3YW22CCyrNqx8dqW0vZKfn3QIee3t9rhXV3Egv3mLxqbtJS5c+aaoEYays/L3qaSbLUPQ1eKtvTBZ7x0pXhVXPYf+OAzazWLTpF9M1iu8dngQWRHuTzqK2g8QpsV+XpjP+5kHukGXQDXxh5A3gxp7MieHZEjpzkeLjgvCEqE06ZEMFSLW+mqRBg5Z3MW2utJQFIIsTx/APPOccZxJBHDLEiDj+4NtqSxq/kbSmMbLdiRQPK1lGpSgxCLO4aqAK1ApSW9glRnWplt6imKn/uTQaHrERFsmwCyFethAEGSe5v5KqCSrGX78OToulUoZ/LlLBkvpKxEkp4Bj2onDz3HRj4NQp+XHFouKsHjzGbxZ8OWbtsjUbPnYjyqTRcTNN2dAvmLP8fV2t4wSZNx0RNsWEHpXWDB3BF74SEFZtRs5jyBtLxUuuTrK6l3jl/AbZQCdv2KRsZpxgVvoTsrS9wYABaGIvh1TWnSFb6InoOA3qmJSm2c+FbBxBW2ZvXvVs4ZrNvDWL1trSCv6S2hAu7pPmmrCOyS3WMFAnll8rnqyimSivc6CCCJGA3BlXi+iHxLJlfx9A2XYwOL5MFTRYTqETIb2lhcX2zHH0gIECeSkXPQKA8X159e38j7GnmFRBqtUEuV/WWX0180csQ9uwWf3zEeII5KBskW0ZlO4wOjfKKnpVZ7BZeSlyeqzDo/7+J6fltVrit9FJCBUlbs3ibtr4O2LSLEkDHuQEeAIHbGm6rEBtGkF1DG31gviUvCmYC3zAj+58ZJiQ7abXwJhlSvnyqvGQHEje8Zg7+4BRXn8Yn5rBI27RyAPLhVMTmffD/PjeGZ/QJXvJBfFZbxZM9aOcvxXhwZxxk2DllLjYNAdKVwbc0Lmq/FBP9r2qV7RovlqDrf+0B4f+gk0kUUrQPLwJh1gT1SV+raPTz14cyc/rXUgRB1G12T2huLhtpSLdyOXnp2+DY6zP3Mv6dDktes2omg3VPVYiaUP7lpH9tSRLStsiRhcSXacB1eDkfOTJCmNDDqd+hDC/SuczuQYiF54DVn5O3SLpCdSlvUXVZZitazWXAlMzxYu7QX6cpDSsseFT1rOUvDOOEa3zDMjA8/LE1p09QA1EWFh4fgYyiyELO8NkM9fj6cpgnO70Bvxx3YOgZOvu8NWbOG6OyQm0png23uNUFQ67reAU1vW0cl9YFsTXflbhY3Jeb5U3lPNiXIkjRoda5GmIuW+KyJpTXbLmMwu/WWuQ/UBQy/gxHCA7U+jtEqG2j375bCAhW31c5i078pM9yb4mMRDmmWiu0mrf1CY+o5XNiUiQMHgBisRKLaOWCAH0UyOliXwCoKcfhjgHFhcshfqK3GKJE4rk48IzWHeEhxcQ94ZGkJelXbMKzF8Ar0YI56o0zkzoTj2qhcRQH7gqzi2JK+WqOrmFclHsavBmcOTnTctkkLyxSGaMCcQKtxnOSdw0kQB9Vj98iF85TVSdxL2YG5Y/7faq86kvk18Ap6OmNYYVQuQn246luN23QGg/H29aHjBPjGb8S2mMZhVnssEstdEGq4J+aMubQeGexRcebVVCZOnwsN1dewuUA6bHahbhff0vGncXcKw3uDj2yETdIsrgzPEdJkNAoV28l9/JszS6JuNtoDkchWS30cRjGlFjN6tlzOLH33NTu8RA76EJQj5z9fBNXRvzUACd+ZtW8W1b38rUSog8zc29G29z9LIYTlvOz9q2DTNeTcujmodHlYoDbl8iO1PGHYvXed8QCor8MjoHbxHsB/xCSswscG1BlNqf0aJUwthPN7p9qF+gOyEduMGQ37lFfU7hvUqaVmtqBq7nn2Ajez5uLnne5Q+QH2GkBhXYX7RfKGUNwdeMXaSPv6eGQeITCfAQHd3skr2DjKXxuB4QYvZa0YOdmBWJp1gjzTOuimlu4toB3J3v3CgYMiAeIZRxsEtMKqLKtkHmOfq37JkD9B9Yrxo05mpISHSDaTrEIfbyFFuoHiGq46PI+NrKcUoh6KLvwvgG0oStwtkYFUQokSLEFL4JwLAeXMk0NmiafTP755e1k9xLtYD20PETvoVe9hc7ouw1+UPT6dBJJ9zkbsmBdZY4/V7ZExUFgAxzyfT3ZvICG1jaZxP3IOVNvtu5R7KbhJ1pzbn9arF18EW2Tf0bxhnJS79e5VbLeWCZYyR+ZKBSKCfcO9y40vHIsp7NL8X30DRk3yrrY+Z65iVkpM4y1pw5+FtGbh4YdH7TY7X2sCbVBv5oDX4xnmW149Z3tCsta7r1wsLnXEoXtZPYkcwmdiIxESbVWR4c/WiN1gSiRcISc2Qx54aLDkoVxhxlKdt2WRJZEbQJXd8dNsOQqnotOBDT61/AOMdtP4hxK9EN5VXwgFeKpaZ9wpp09s42Ve6kxs1Y6/tstMsn0mEkDMNQT8kR6/llMuiRbMi98BoJCCUPCsPK+8fMa0YJ0+0mkOke/32QhINly5FnpQn+Aeg8kQnmgU9svQeO7ARo6HZX3DSGvbYganHwFR9+WTZ5glK9dLQq7TykwwglxtjfudpktNl0bKsvh02nu2WAJ89neySN3fqmSH4mkm1oIdFEJfhd01eKhPn1GYUtVgDLikoWm6sIzfVt89k9j4ZfExlqDTqEqY1clvpjvX5ojewofMRsL5tsRXbYn3RiFhHCdcjgJESWviSS1oLWj1VerPWEWZX6cUZnTwI/wnHJwTMPHE+oIARGGFJG3XoFlM0q8WGSBPDozpsG0TEL80TZ/9bAldkRQPscIT0mZHJHkAb+1yE+rkliwwWTTMAEHv+zN+OAY3X4q/+Yeo0MBREPWUM7xjweMzPkJhXrQFCj02GpW7n+cD1Wni4DELsj+zgc+cBtWhMk/5WqFrYStoShDjD56oFqdw0ZiU3qb5oRWCSy8bWAWRdr59HsqkoU4XtOTgtakNEVjOE1/ySrCeE6WmTgmqyHVMkW8sznRuN2jQ9EveY6gDxJzJa4O45IVF130JD79DriXB359ho5W7KNxPyCUFbFFt2UdcINa566oxF8ImhRGi5R1h01C/Ja3lpRbG0BINessDvv3thEStNrNc2N4vKVR24JA1ufPd3ApAqC721y14u39CDtyYZd0940Cb8c9MOHqLlTY2VY96PbeMCHxnWO0ovAPYSLSouXDkMRm+luZBqR/kcBYHUEX29exMNfpyvELKkaTCgqPQY25sozNFVDNl7Hzb+fF3LDmxa7RTH9wChPY0GjU6C96HDfbuLxo0xNYMcQyFgkeTxqodATdUd5B49EWP8LO8maw7rBs3RDJqkcCNLqFDyvct27s6hQWKPIhQmqpoSa0Tasg3L4k/0S2RMy2M+kWH7WbMQ5KBe6wcmAofdZk+LvZnLiUz8geyr/8eaNYHg9KauvScthMQtlukve7ZNsjgE+cypuF3OmW1UeZxOpGHK5PM478UZTXtVANVzE7R93NJsVz98P42Qu7S4FCOmZheqM+WF1K7WYg/h7K2QnN9Kvhc3U4LiLRz0AXdvVQAxyoqjYIf/NZakTlg/DxluGolLwk1FY267/Qbzf0JovH81ddHQvDMFwQfN2IxXzDB9OusMSfCffMtPkhuLnQ9WReHRWdssxzixjavv4ygmq0ay4ngDMtSkHVD03kipT50Zs57+Sfxh3xCp6ezqihKjelLmwj+QrXY7+dxmgXTMOj6sc02Q3pPSbB2la8nt7Fu1z/ErqDulXR330hKzavKCDch7GoX7LcSzk2IHsAvjKjEf+w6DuiHglV/4u6VhjMC+0pQFY9zpdLDZF0FLOLUjri3lYDx9G4Z2WbY7ucWVQxWGMGjkqF284qSkVjBMfKbUUfCFyjuouMVnzGtZvzEziHx7r3pW665o2A6TXiPTvvRduqQKlkPTN3rv5ZejbG4nMTZjIB1KqOcEBSjD6ZPS9ade14uuhOqYvZ7VOek0LNLmopEZ5nzB6U/SYF0cSMbmgnXd1bZrQ5DpWXQwJlYs5CZv1G4YiWUclNQG7By99fUvOsr5mHdedkoH/UqPpIbc3aHxetkm9+7WGz+oy/NLZ7mA7Wn3qjAzf0LmkqxvvKoGFNy9b65WRailkzmjJjyUZv8GjfznaQvNNgLllo331ovsArE6hbCsbNRsIuqSUszLo3v4EEQn4NrZg4rhKKh7jApBETjL9/cPHLH0l505oXaE2L6ANo02ZV9jgwGCN48giXFjBpsYORQ+PQ9IQOF1UdHKZh+MPK1xtqhW/8teetsnZCb46g/iUyv+eyfpXPbw/57Ha0BBZlLAgbF5Ayuio5H7Eu09cJZ7+ny9gHyAfYbx8h4ByKL6s5ywtMRJfAPVtYwBbVSnBDFdF2nOKvItFIKJDvkweFaPQZWPOwzKrS8RxH9kui0FWRn5TIzlsLymnL/0uY/TlXZa1ZJi9rgtsJOSby/UntmwXN+O/maTm2UGLMzTzSkrbCbSUUsi64HM06JH7bnA5T/nMUITxPcR4QlwYHAxStKeMBOQf2B3ugPQm/9XzM+bd8HjTutcWHLzXUtegcnTNMU33CyFdGXZWMjakz2TSxTPKvwrY4g5CMz3Uhh3fFnDPPhVjQ4z0U9UA2O7Tt9yG3fGOjqcgtY6iB6mqSsMgBbqA+xG6Psu9/650TkoYbOfCKh2YZ5v2W3fx+ou+xnhhi3AYorGBAbrx+ofeZ7D8TkJAvc6P3u2DK/+2j5XIe5roQx35MZlUwdYWy32KpEZG7mxbjDmot4OAci33PwNYvhDckT2p0ilLMDL9L5hlo4QlLAbRDFh3ZY1ZymWAYAnPm9oDKq/2+8rmAn7VJXl0rshEdiQLkxrZLtwWQ9kFOXWeGjRWJikOl+jkVhTZk4/CLiHqQ0TazYydX2PtyeJksOiaqZkR+4ZPI/QHl81j3SuozW4LmtUpjrKsqNyU2FKuias+FdYfnO9m58xwK57KwQva+fEhH2LZtEoGYICjKjewa+lEjUSe2b+ZAuEWa+IAtUF0l0poBtJ60WEJUxO7dq8wZuf7JniE2gThvKBNvUW2NkR7gl1yAdNZNzgk1Mj+xqbX4k5a8nbgKp9fxHC4xS2MSMTWjHAQs2bG31XDorhRtD8PVjKcEwlDJNzG1xRitFDwvW+CXWvcDIYnkP8kIksaS/a5iWblOVxl6q8HvfkyH7B24qzAdiuP342di8lCmVgFzVrPlk2xZoT5MZputbAoimMPTQ0gPOdRo3mTW0sawOeSCkXTii6jyOPT+5FoZetcwvsIgQHCgsg1BDpeepSHOjLe7nqPQ0gBohSSUSThpp/P9jiljaohx+ziE60W/24A8de419gPmrkfqTDHu7ABJxvPJtfqCynQlpLaTPcD7JD3VT20VvFHrzsQiDBZDZ1HO9y4uSXqm2PQ/4YEYALKOt6pD2FF+WfyUBxfURr4TcUeMuRW2PT7fDxNMSrLzQnycfTsOMiUXQdYvQD1+qg7S26RJdXNLN3rcWRmTuEfknFPOLvpwkT9LBOSUArqU8NWxz53ESBAA1C7cCTuAR2k2QH+IX1jD7VMRT12mncfqtpDlV9qtEhlvp7COn4HbxfEb2gSHXUWdfIjLAu5O6Qchyt2IeA/Y7ja0eGmz7ZxXtqsixoqL0CPlM68fyl4Q8rq9rC+L/iy3Df3LPR+poGfjdxIZiFqYuTQIVzDEn80BJRzM068ws5bM7vfrw5ozfhmHhcjl2+RtFVqPIiEzt79CUJsoxHUbNQjRRfz1dufLfviHb0sjdpL8VgquRcotFP1gyahLkebjEmO/yuJ64dIHk9SW9E10PGAU9UOzfveKta1MH+9TPW6JtuPeHzhE4aUbUB0XYLV4o/Luz39bJk5cQZsuB+4OI33rN+J5NZPw1z0Qh1zXkMvS5nNlpsP+Q4ipRzKeoK4oyQTdUkIVMuzXxBHdKGVw87shN53viXFR/NGxsbNQYLDPOVr6qjn98ACQrV/YwdXpk9nAtuGj5pTaEsfNjHdKNP0c7JhPr0bJexZ0h4pPD+I6Q9OuHjWhH0J3aK0dKHp9KctjAM26szC50t9iN2SlklgPYFn2yAI4Bizm+LKDZGbcnJxrzBHW8yA6ueXDBykGBTTOOv0poJRqpwvLgPIN/YHtPramyg13stTG+1j268MT7ALt3vD3f9CKjI+viBLSqifai6Py0pVi4ki/Aj6J5o076vxEiXSx72x/lKinZs2+bSsZmMzbQt+n/4hJa/2aLwip5l7tplvtclfz5tZzb2DyZZ9H1Oh8yDKMuvswQlqcswWEgza/U1WBDcx8LREZ5M5ylQw6Fw7WTxr4cOyhuxgH8LYpR6vnln/NakkZCRHh9iyQFlrNzj00jw9jSW9sbP1KqhHk4VQdu/QA7VEUEHQoxT2GlK8NQbl869ZRRilvlrA6T0YYIX3F/KmjM0VmrPbrMk6kRg9nAZbwySgyeS0/18FC2BlOrxQbEMZjaXW/2jBOn8RxeHusQXb6MgnLy3W963334Moe7aPyNunSpTGSbU2jlcpbzwt1YVCV8uoo9BhLdLEbrzOw8L5hN+X87I9cenTrA7PPuqYWdhgY8Y4bzV6tu4741UhFcb+p70WLTQLSxJYnPEoNMeHQl5C+gv5DdpEIW/Mpp/0PjExpT6uGqecWhV7X11bhN2GSFiP/BCUxvVfbfhNBTGjUrDnFsKwTYIJBKya2x7H+/RnebsPuJ8G01/IyXdghZTH7bEwprq+htM50fE7iOTSyGddxLmz8kfGzdhgiNZysvRR9+dpMRoAO8Um/Rox3n0+1HNLwlvBc0o/0tFUWejQgJEuRIPDtcK402Me22Qz+ug5RDCJ4qWC78B0Oxp9b3tGlq6x3cDPrUgM+rCPpaT+5qs/cy95x3llFUEDSELJxB9ZniWhCT0Yxkmha9SQEYHO4XVGmelJEKN1uA2OZ29ChdaXh8mxrNPYWpbSxbu52wXK6SNtNSvCZCFl/1DwKAZ0zF4M+1zasqej2ToQS2MIhXmMWSZDXbv+VE4+dOoK7vQdBaxu/0wnYc2GU0vuuBSDTAX4fYKbszSrpHEsI21b9TeVLpKo6Sdp+3mDYLgEdwFtyBjcWmhsQxdo4SThCrIPa97eJdWQ0UvxMtlSH8KAORjvbg1n65kcUBtzXLsmhBaWxF4+RrphmB8rErNpHYuEXmTmS2LP1F4aWEAM5hGB6ssqkeDk8pwmeluti+QS2JooJdwJHYGd5ALQDMsN92WsJGsHAKG7+DN7VMgrJuQdR+ESF13/0t1CP2N/YaU9GeUwYVlMcHMd7q1D/+D56qOgQf3b9mW7oJ7PAedeUksoSrRI/MGHP4NZjuJAEdkzIgv5qIW/FcFmbuxnz6zhcN5/0m7aXrKk5WSQXM8Qt7GuWJpRjigWrN7bPFayj542y6yoIDqKZLedx/NlIqmH9zz+t9MKO6t4t7CAOM2EKUnhjY0HfDvMErMnz/07NGM3R+Y7ljoIyWeA7mvN7WSj3TDojf12mYDfHIkv7R+4B3QOCkvYTPsf3O3BNbiE1Qoayl4iCfZRATikWA+8Foyib0u7ELeqw0WTrAYE+9UkYEO4CM6IOmn3eNXGOO6vS3FKsBAOiTvpfaw/0FuBP4Xe1poHrnv2AtXsgEi2mJvxODvXqkP6JnVn66C0iWDOfG6EHyw4zwUxwotjNNowrnoZTkYbGZgbWC73bSe5drzPv4TdSYdI5sMQLmMZL5Vt1hXRrGV9aV9/t+9LpKwonBqnTf/i84em/HR+lyHb8xlYg9eYG+8/YIi2wYMaxQV8oEVJjO/BnDA0WlprkTMKngIaQeV6M3p3cmZHuQAZ0yEVNWuvJKwyec+wuldwuenZVoUeV5Bio8VZ0PFV5qowggg1XjEpT3OYO3dQ76LpNHvNtxneZZjKlTzibVMoVYKi/7YGBX/qOWMhbtlsVmruTCGjDdeBCgEkNDRXW9EYIDMgamJJZiCr+LxzZ9dNB67lzcUjS2zm8U52lMbcD3v3b53DfNAaH39HhasHpAVzDoY2naf5RbjUORGJBuXiezXpx34CivfXkLwkG+fuTwTVoF31dSMnKIiXdGerC3nzTACe37prs7nf/Vrtm+dHL/J9sSqnAsgm5wTNLs1npFLSCv8uN8NluEXv1PojwNE3RZb9+u2PdBCIbt3/JQmL841CGNYPbwwhJLry0F4K1+LVGw+rnGPokJpZ+UhaM1+fl0bOnZPtmtj0X1Yt7BovA=
`pragma protect end_data_block
`pragma protect digest_block
72a53ed1561bc01b567514319e7f8cbe0c92bfa1b20891750ce1fbf9169c9823
`pragma protect end_digest_block
`pragma protect end_protected
