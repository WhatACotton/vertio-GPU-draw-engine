`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
UzG7ncwP645sOBH6fKHYknG5etm9BogVXbWCzp+K3DVXK8V+0PSXTocA+LFST+9+h/lSf2Zr/hkmk1Mq74L5CyW0X+7KEqyVwrMDAgyzJuQ9mMtNDV59qPELIRH6UdkB4BrLKOJoqlsGlDLHDEoJVuaJL2trkQIN1+UIGp0a2x1AyOBF6N4dnMJGfCIrwryz6GgeRK5JEI+SyAiDsjr0x/icQzH8soxWrAI01TMyfVxRRraRWTc3njxsHrIKyjPgjBK8y1vP/Qj3BocQZU5GXfxWTS7w1E4f9wlkAaR2MllpK7HJvkwnFAXNRCXC96wuk8PI9yuzxe4Fvnm3Lo9XJAcmubPb2bDJJRX0GEYEkL5cZNxD9LmXwErXbKzw5u4NLkzeiTfHbqBfo5Rt+yFZG/44Iro3ULZLMm1A9UvN4kJ7D6k/DwvdZXEkUVz4r39c2YcBQ6o5pUq83/t0I+dZg00ENmNxgpb8mUQe8m8QC0OOyaefei4sUmWen3LWLJpNrCoNT2x192M5mO1dLT/w46Ciq51onQ+0ZorbtxXVWu/LYCOFiVLtUn9YIVqAONiB+x1kp1he6Bl9XkhkA75BXfvtLc7jbskPQq7SJnQR46pAKfonHnTYqjKgfk3EXMG1fygkIY4eUX8lI1/KD5A0Z1zRRGI4u5KE3ck2rSpSrcyh9AACfGHwBzqlMgW6ZDWzGGo6mAurxxYWwT3KQPKpubSL3dgWhBqBuZSGXSAFRUWOj+ww6zHhjC3YNQAi4s1t+kEB/N64uBGpLu+7TN7vqZ6/Cp3XvOi6dRceg5sGn/6NK56DH5utB5NXCfwbVgJm1FWWVzjoLVXL2siwj6dc3N7CpMrEvyt4Q7uLOKBLQqncv4MfjRMNc3Azolwt2erjUSJbyXdwZHpO4LVCtnF//BwPknfGyc4sBRJW6O/pWbDlgWCnhZPUrHGM8eSHk0nqS16BVVMXQSJRVE7jIAeM82A9HZlmEbBQzRntAh98kYwPC2qfc9CakjjUl9O8JOix0vSfX/Gz/LbaMFvsWTXcYs3HieTwxkF0Pycwd7XScOSz5HgGf3U6vdS5UHBdBUd8WzQX2Qhj1NJNuw4LJxPrEtswsVVEm7QU1gEJPb0FW8XeLrZrlTfcxrpf3EDHUeK1Y4fDx/HBD8eIgbzPuMkvtZUckMcjwsi2KZ2VWfZL//XCbQLrCtR9yRIDzEJ4BXa7rjSHbSLHP0wqBWJllFhWx2Z4F61YIi3iigLMYVv3LoBvLwGYkgHXj9V/Dq342X83PtHTjhxsU4Lx3FCo6ZHmO+LquyRCBmEgawwuTGDhCgsgRX1V/WaRfyiicuz4vDJkgd6qI+u9emW4DMDuk3cMHNqvZ7/iwEUqXvP/pY26AL6DCUgNwxrfrsDRJhd3uGEaWtOhln/h7DBceCWTVCEia4dIAoaBlLck51Jl2Lu+B8gttRYzYN4OPbz5NM8yRIZaBM8A8Ig7iOiH55AN0A9wY1Ah5b+WRKCHSxFRC0cN6vS09v0O/EENn1+Yy+QgY5A2MEePx3p70ySS0vGHzbJ7PR9tRFxA3yp9rdOztyXVf/ASAMa63O52HcYzoQlWa6JfsopjarCl8Gt4FgR9uaezuLqRpO/l405/TOIR5sOiWCbDLe5XOSZ4xBcPXq1XPNrMNu8Z6Gm9nH0c1LX6eh6PWYWKOttTns5S352FjgPW38JQ8WMNP7m8ELhe+vAg+qlchVTwdgiHvSeFddTqD3jxH8jLfWzU8ynMdyzvwBmcLoJ9E8R49kuFsA7Fot3daN6UVmfHpS8iIHnqEGqvV4qZUXiTE/5DFYsDJfe+NNIA7dN8wVLxwbLssUI33jWaLpS3J3qdBQ48Wr2iBDB17N3oONEUUmNdKXYmqwHvzBlZbNHlBt0EDGy+ahWaDL1fq7EhX1vqrcPXr/nkwYgagLiuzUfvklc1HsWCJqcLCKFM75MlGrymNswjqFm5vMN+iB/NGmtr7IgO6THDrd0zE1u1mo6u/qClbffE7A457GNESFX4BlJlB4f2h/5O2CAwDR0mrCsBF3lZLip6ZuzA4ns/4VXErJZiH6DOHG4ZVZq/ofQNn8igdQMYwJFWZhSOSnOdPJddHDzEqd2QAL+9CzGWMxepXgnqdRPIZFl3eQtr9ofTLu5o0WWDsUhblCnRDwwkDb/prwuIEzHf6eQt29fTaekznU49Ld0cCbvAkeH/c3qRUs6PezfPbh2E7rfPrOcYoeHYMPnF57qYNpBXu7UYfTKnIkqQmkXM1ppigbbJ0/7qCvdsdsWd2EJIGV7Bcn9xLgKGFku1OQmCTiL5AadR3Jd7bpOFTLs7S6/mZzkvK9HMrVKGDAxSr8kxRVaAFFM1aI12VP/Za6fZ4SyTsZX1xQRCKHozYtUADpCPyUrpYNUumimrkvFThfeQ/Tu3Oxa0MkW+PpcXsvRbz+9krhvqYT7hRbt6i/IPlKXI5VYRATbYTL9OzvBZwBP8Z4qaWd2aGt9mO2b0F2mqG3QajprnoYkADQWq8UGepFtGSTl9jgCWZZJm222e1L8K4aGhs35zdWK1bPCcX8EPWnY1P8pMx8KuK53yVJ4ujp/m6bRVNxEI0mOH7f9QuT+qQMH8bo8KGNt5w8OVy9oOrKDz3hNQEpmRPc7Dvmh9VW31zYceml3bZaqWTZgw67qc7EPec+gfA0rwblOc29nwo8/FjzOPXWcJeVZ+XGthrRF1eei3UJ8S8D3HCt87H8P8Zg1tJ+UMyc8b3pYl3iPoMKSfz3sjJq3GYO8BK5sN3F5Eo6IvREBfZoWfr9ceNaqnmmocly6YKH7pzKVEY1xYpc4nVOf13UiMgmLI7JpSQYIjGoszOi6uESx7AkTRf7HV3C8ZV9iTkS2fdtj0qosncRoW+LqxNtRICqLJOhwzNsgKUjV5qZC1EM9+bgI0mVWfz2JhHHgDns8NxpbUpz0dzhhQ2dGYzs4flEcPS7jCo2IM8q7GWiCE6zNJkpbOQ5IuAYz0hb3UFqV7mV/TVKhrZ7L4/IAbsI7hUAGxa+aHEzC/v0062PFADl7cqDyCs9eBbv5EmeW+x3CcOqeYDwKMYFweA8m40MprdiEtZPhMHT1ZsYY2O5Q47+8k1o0OeAE+U52oDxZcQAbXyg4EszGncmb4TGXS+/MEIG/unnpzUqJ/6HhyMl551Sl++vqmpeXckFYmF2cYBZHR6xZn+04Gze1Z8T29JJZLkyBIJBMxfZPGWPHSDTGkM/InpffHoxK1F7PoBA4ZVCnZ3AT2+ZClk1d4N/FEhnCPhtY8H0IqTcdGJ/8vxHfxpSLCLbCPahXlKnTh871K0G9WjOANA5NVH6CxdUetD5K3O6bYWWyGtycEDDM1k/p9O9ik2ps3NNuj7nZYn9qsxTKbVeB9CSVmXQ0qG+wcqd8jCjs6UKQbtl3HqNPHyKkTDYGbz78ZOAFie6DTx6H/LbFjK/3WTOxPQvbdfgIjD2bBUeWjHXSU0cldohexTKemsyetmQ+K/CDUj+WKLZgCtEvhrfQz3bEjq2nrh+80NKsD6+oyT6tRpmVYC/UFTYvbrqBm/lSZ/bynNn66K/L50ogqZYZ3EgpjgfxxCt7FWL/3Jf2lXOAxThIynQjLlweps4yDTeRUMG5jNwiPcha41BYeTZ4F95rV+Vj/+QcfdZrd7AUDewLKEKKltwzD6d5QZCW21r5H9hO/A8JxYtAFHvwEPg2ddrPrcP7rHK8VKYyhiC3i+fNfmZpMC50NhD1eS/E4s96lGAhxwp5KS2hHVl8KH92vEGfTw33/gDg0LQ4WB/Jl0T+ZOdVhK0gCEzx8MvRXSoWtiu/b0mdyTJmgeQQ3HfPztSuxL/YK7Qk5Eiau/BDeGZNHKrJGQ+rdx4wNmNf/d2Vl1QJkt4nic9L0mllSaIbesINQnJNsrxWQUruYkrvz8fFr8gsRtTEquOueZDHJ/FuOmRnhE3S6HTNKMR81kmuSGqThk/u99bU+VKtSgptHbVFrZXWkyariH8ux1tkEnfI9Z4KJLt8cwAbeWBoGfR4sHH6A9W2+IQL93k3dZLn6Pn+fj2czsRVz1aEoEKt63vX+XqL5MppkkjggknHkEzwAxx+ffn0gk8U7nATW8Kg2cOzf6sQTBcVfcvuhe92qLLhLzyc9i7hez/gQnrizPQOiR4e7pRb0naMfckgpdS4aK3EGUJRPrwI4G2Gau8CIh2KilHBNHnAzAA93uRjyKqRVYDiggVxQmS4EPv+0pGlBnhdE1/XgEFrnsIkUIsla1oh6nSSNdjTHd0qtsuyJ7KAgVpzWyy7Nmt2uyIF/2CmPBWY5m3+mKKUvOHQY625dbSjKcL7CaA+yshLhXkaJPxlJDFgneXZ1nhmOANhPZGrtUVWZUrG4WPXzmJdO0bDJsZnFC2kpd3wImFHhvkcN1CM7w5Wo1bOVZESCeCNhySLoBFUszEJ2ZhaL0JTN3J01kJYGp0BkqQ7cMI5hGGJyX6Rl2lzY1oA3R6Q/5hnlMBrauXPtuovcRkH8x1lrJmWLUBnwNpzMR/GmqCjPJhNKfDzcuEY3sW3NtWXjsvWNnviRZU2MxyKRtVVj4zcdYI2LhJbWrx9CKP3u413gKph4shIhSgtjHUI75xsTPhmBJ0mcsQW4bkOGuDDOYn+9pyCV7w0/VdCOzm/0OLHjawt1gABXTej16EcYk2KJqS73hciJv60qjsrcntxbspJ92WmWcvGxZfbrExSNRSLOjUo0MuQBp0k+wP0NPrwjcqqb8xd5q40byqnpvKUkx1Z61hjkJ8Y0ZUZ6azsdolGUrA3+gIsK+ew63Mat7RUWsCDpvYkZoUL83zl6wjuJSKHt31uvP9QTM6T5D64kBnuC2t78P19Dw/pje9R+Yl5sr5IX+638yhBqjtgD+krX2qWz7qCGoFRhPhkoGtcCDVQYRdKORtBWV517qZ51S9bUDTHvNZN8PwIatUIPFB+1sAUWWg+vNrQ5GxwO9G3AOwvAeS2Hq4Zdvf6KgqCN/oZPQbgJGDqANC1J2SfGpB2sEzPs6/JnmVt8MJr9n7AUtbDE/cIylzAti2QtibAaPq3lI8T+3a1KcrWsJfHonJpw4vlCj/SmOaP5Brq0LBBHMsPvWy7E+gVWfV3YOD8L9dvAGg4Z/4D+SiyMmjAz/vHxCKHYWEIhqmVRdwAGnFInz3Fb7oIb433XmOOrCO+5DXMBoI8NL3lj2qghc3+nxgYTR8n4r3sV4aTnrwFMJkU8bHC88CQT8Iv+UQT35ir7TXayHt1Do452Shj2ZAlxDJgNQcJO2fmreCTj0awgVbWWk2EFhNtUbeX1smexFoDDQwKH4PplE3CltVgLkJ0+S88XyQ4PQWmBS8WL5aFCs+YQMIR2xm3veOrk8gSVKThZ030W5EK4zAWpLTcNylrgto1hvG/GhLtIxVxmxurxgmpJBiaIV6uLd7tm6m/OcQ/s+ivgUBuf5gZoGO2nbW5HiHbIIYIrkd+F6fgRbOMib+e+50LtZ/kNDUrWvWWRU3idGVR+bOTngZlXTWshzfFCgUdvE+YN+/ius5aojAZmAYPXU7K5405gyBZT+10umJ6FhbJ+jd+aFd1h1TNS4ZZdSC9D6y0E/4BrYyL7J5H1eKdXDxca/55R7UYto3SKk0Zn3R/j98bUYd+UEel9h7aAKOG+7ZE95o3bJEkwjyAjMQumas+U8tUaBFvNmXxAOQJajbGLSiJ/Kwf+pTYiSRdNTgyxIJLDEpayd1BiwDgqAlpE9X6F95vJb4uDq0zvwRg88ac3O23B1dux5joZciAsfEo98YkXyDxqqbY8XIpcWvNerrG3NlZzyHH35gA9huRo0aDruvc2c8t8kpamWiPjUPv6gDXmndipNid/Mh6eSDJsrsz8Hi2nyDVqWWmZTZq3Dh/RMI2nB/ykFDxrbZxd1IknJMJ7hHvJGKUaz9GdFeyGLcP7UmXFxpy29ZjL7sYsq7Fs/l0WbzxtqliInMbs1V2r6/pRSwIt/+WXwObYNvDPk1JrM8FQ90t5IHumyu0VRskjtq/+aiJVhLXixBarUAtj77jras/v3dBtu9HgNi8ouCjvLKDwq4Y9DnRXk30dbMRBzeJMq2nfWVRM8PvohGBPHLLqoIPNboz8fhush82DSNLP7VBFY5cHeWQfraKhNpDREQKEuZ0hXrTnPCtFF6kPDKxiMCtNmfPzK4YYQp7xkholMcPMeTbpHfrAeOWJgr0Pc9Ah5cO7xS4ccPISw8fkVXVDZ7SR0/HSnDtDVyTkZ/+MjdGVpbP81pJRdUjeFAj/l8wSxoJXsgy3b4RlACWvUWLotSXSCp+tet78qorZ6YipyG9rDuwS+MvOtTQ1689ItlUbbDPDL7eXyhOhCFcOG2jG2ZrnKx9bUM0q4H4pVWPlEOKuCvZxxVBUtv5QiS3F/Mybx39GmmN3JMG1n23WGPmLicdLhHcJwUFnjnlwO+9GtQNAFPKlH72P8Fo/VqyqlF9ZoZhfWPmFLMBjKLWC5m2DaNXNvx79gRsT/k7a+QswMBV9R+FasMKa1M60+arTzyGsU+2E54N+YHAj1r+mujaY23FwyUv9hTE6RtNuTpxu9WLMRi7qCHKsLUWT6ehWyEFbiUvca+51iYgoJbEtrYuheb0Mbf5vFv1Yk8lVMmjc6/D0hppNe7ln4HuERxpOM0n9aBPVAlxkkTz4ioxmljHIxJUYdHC/UJTpLdsBMzWvlALZg4+Kkx/ypKlFlglKnQI0VJKHlVjcaBXNDe15wvNyqdSTEG169rUgEPLmQbTzbJdPQfvIXdZF7Do6d6Mg14UoCp8NIF0rN3KkE0jsmJrQLlQ/b+yItTSYkaB79+9K793vbYReujNi5FeAhH61w3GxVjLfJpFDwI8nLMWRNt5c9KcUo90i60sWuin8VhVnjobUgIW0xwjorDhhut8hCMuSScpq6nNUbPWfNsLAUxlogEKtGEhdtOGpc6t8gMZkJ5xHJgfjAmRr1HIVcQAKfVwEs8gqYMbU1NalOSmfP0EUDn+rqXyOyYoEI0pJg3ulAQtVuez2unI8w7VZ2luRt6/qd0zBVJ0j/YD0JHbOFe/2yipb2DXHkH03F+j6XIcoKRm0iNfgC42F7JjkGOdKx25Q51IneELOqowoAi0JrZhXYV19G/2fXDDI4zC4W2C5GUOFa3nNfkZPyvggZhKtPDd5ezG/kaxh1FHegS9Dcne8j4DkcDnMxH4Zi1JRla7TJQM+peORq28KRyvZ73ECXg381BPUed+2V/HSGW8EyOUerJjbLMOEp6iMeAwA2I5SEX44WTq0CODNMsqMhWI8k9vs6rxWpj4WniShX1wLUnICnLlhBCOnKi29bUgO6BPikFbIeTr/l4lIrf+rXlTc1yUKDA+7b3J3znmBy+tqY+9/B+DKiBeYG4nO/de6CrR9bYi0ib02lzzgx2EqsSFA5b5189JcXQ9jK0nEaYOXUhKS0c9GuiKvLz3pvOQ+tO+6nGEdw4kV3+ZpHhy9SqQdV4tJbYI5DaWfKy01L56bYHkgUrras0P2ZnO+GCgEiOFc8dx6Bcf31U7NpXNjzu6h7PtIdbIiGJ7b1E19fn1k6kQh0N1YMhZCwlvjxRhG16ItEJWwBrgwbpj15hBWWRvD6wzvm91pIwl8iWoUAL7dJa4Y5R1bxQOKOWIYE+DWk6M5sOoyzNza//K0fE0AM2dDqQ99YxuPHT0yei9PjtKi//LbyaZWakm9nmy0wvJPTh9lqFxN80YGL49d+bQNS+k1BJ42uG6Cci619VDBROszDATKG8lhmFV6XVMC6BVbvN+6eHLN2wF4y8seB79D9t7mLKYMXYLBpE18VbSeL4bqTHQKDbooyiPs14uE5aK+lz0QTzyL2l98dIq6k1jdBWgyEhsHK9ZUYfTweohsUKWXChpfhLA0wkBn8UzdMnKVytbQ5hVDkjfmwLrrCdgp4rzlLHBYCzk7D5k/EnhZ90hRifVBAnMYWyu39kGF3gtM0nOgVgGxj4nMfe6Gox5WI6vOC1Z7a10vy+pZpS1+Bv9EkTFDwYD38J4btBnQNi8VG5bnNHxcS/k2P3vOBE45UWBq3peE16Vrqwg5NykWjz7tHzWbIbNq4FnERGD909qXOBGYTBtvM5FqFj0zjm7aDarx68OK7imYHHubABIoEGHxJj0wSpFi1EWOoawOuOCJIoMaUIUUbnM2cRrBlo2lVCiuTr8iSltPZIgv6YyA9vfS99F8bNaWA5a3OkAU51UXGQ1zoS0c+MlxgxEKbKXgtALjU8fQjvIo8l+Z4m50Sak1KSNNo2w8s7QsUe91oQTR58z9/EfyloiMmdNr6LgibceYLhS2OsmweZaoqCz56XOyEjhFyC2Q/2v5etJkdh2acJAYHxKu2/Xpe/acnHUhUgBh3aSpoi5AuammJB6R3S9QUUy/DVWz2pmGoGr7U7w0kjeZxbtHd25WLaFnE2Vy3rQMBiYIwnlEgcAeMrbAJ2sPtOjrrE2ceTRluhLkDaOf/tQwWb2UXHQIXDwNc1dTB4qeWaa4L7i/FALVWK+5LDLY+/uXvG4J0iUXPYmqLLYP82hV+TXwXq3CcTWHpgnv+A/c01eYFQwGYLX10iZiXYxONr01PULKoOTeX+3RYi4mgGAYTXAO8qXBHq39dSjFuCTun6EyNJpW/if17m90yEbsqgAZDRE8iepwXh0TsBSb6S85WssHUmawKK2W/as1vmzD5x4dU3oS8VIPjX/QBGCj1nfZOHX+Q6sUSg6NS5gvUhF61xZgZFgXU9IvPKiChoxbNEQ+HE+CdGzKlvhl68O10Ayd47DVbdAVxIG/qV0ZBpKTDA9Up7iA/kSggWyisxrfrztaGyQBW6EHsqSwu4zOXB7S0d65YxrpKwp4yT/AupmUJcgPigdLe9E6itNssLaDCqopH8jU8u2yGefKlO0XZKAv47+w9peCESu8LMgd0RxpxcbVI9O0ZG+62Y4nGK2AGORdSkk2CeMWlGQ88TOPurXgxHDPOcMPeJGlDn4T9x8gJs7FqpjGP47TVjE5VSVVZG46raw6acm9KzPb9Xsv/61QIS+73D3y0T8Tc1MK/Q0xr7qImhS9vDR30UMo5E1EQ+s0cg6M+sBUjTKJXuPMpr5Iea/p0wtqeA/cym8wOLH1JyPAw5W0dvaaxce/8amXNuV9KJ8Kzp4Jw9yjc/z2gHkWvoEnV/ZpHVfyG//fIt1HnyRdFDcavGC5Z7AAo3K8nwaxLe66HtnmmZuvZo0C47exQsDsOgCN22TMeuDs/nfkmzgVvehErf2pMt5MMw2KJEGobPxKGPtbHgLTueJ2jJT/BHhX8WKBUjJksASyl5sC/MFsnhyEWU4yluu5+79U3wG1yCG6Bm5QvOSPV2wYXiUieLHk8j12ySHyNzUS9LZqSPQ2aalvOi2HLqBfuWj8A7bmNyZby7HknO4aRQnYsVBZ3J0tx41Jabbduk4p7XmDtpKqcaGK882HNlktj8SeXz9gKTt62jgQftdTigz08uan3UQpT3lfPyD4yVQoZlcLBe2iCdqeCRUyEY0hoM5qZGwUUrXMECCwn4Qn7fCBClu801yfHvkPz8OWOE6FUu7C0i02FhnLToY3dukbapU6qGYm1BguzUeo13RHLeEj2X2AfNzV8/tPFa8Ry9e14cl8N/xSBPk6dUr6qDc15SnuzgrcVIWv0wjuJ93XbwlJW29yza2udNmwu4fkx3upOIcZi0anLlUWkm4Ys/UfOEXd6fFV8eQCiz4ymiEBkoQUo/R3CQBippO7oXqHCLdQALuprl6JLiSxDkywtli7k7+jtnUCL0+yqz5vgyCFIhuULHIMF/RXpr4lTsUIuGYQALSYAwOH/wJaADIl1jOjydKRLlumVEfLF3lZ+S9b9GpoBiSAX4iIK0UkcqVOJO5eCItUENsUKnUCfIjDavxflHMeCi61PJifkeaiX0suI3aD6blTawySnF/+2I/3igiMYFZGx6Gejb+vrqH1iWHafbUNZPAsCL+COyuMlJpCMVBDmANuhaJ7ewbZ88GxMnMh3Njx9M1Ku/GJ2TvimAcM/Uw/R4WcsKhKSMzLD8uzpCoNGD+ig8Y7NMjkf5Kjx1lZm1cASIrH8wXShreGQCXytkyGt3wNK9bF5xqMxcIoz0AhVXmqYoq+WRkUTwf2cLXzc4OFeUyQPfPKtVx/dvDpZoUoT1sqGYuh9o76zWL4quUCKYggo6g13/GmOLSCTJiJHPjFH4aFIfiBSHcEBx0PObaEh8gw8BlIilN0b/Nsyy4QhihddwnE+1F/ueW3wCIK6wEWIKq6lHJfh942oVNUkLhNk0ihc5w274qMqsznZvqnKDdFuipf1SnzSDluNm3hQvSQSvMhh1iSfQMGVQiqU8EffTSSfIEIM8/kC89Rj3VhL+IYC+BHNQVRD8Xe/qh1cv9dsOQQhqjdGIRQMUThOZpjW7s85HJwr1iXvmHfMjhGf8wfxe3At5u3qhz/my8TD3ci40wqzRQfnAx8Z6C1a/7+en9NApylpPyr0v0ayzTiqEILGMzEriJFU1Zw28SNoZkTiTchmTqxB2l0jA0a+Y3IF0kkTN8KKgiUDBE7xiiRcoG7GuSstwCF6BZaWapU5BcxalmP8Rgtu4fIoYHtJFar74yG75m7eNjq5OgjXXwF1nM9ldsHrO99MOh8+WUUnHPfW9cy0YRw4KUAft2mN+ZOpeb2DRyJGOxSYreSZfxnNz+geEN66YqAdcId6k854+LjYn6KWmLsVuW1/ITBPJvtoy55987tOr9r+woGfdLtonPSbmno3oOjadGicq62XJx47xZVo7STrh3Y/YMJwdpVrGUeD3iByiixnISvkacVdjpD48BDdkR/MJMhvE/ywCwFei+eWgX49zwVSdu0RwwDfkCFUbNyG3Ntp/SMXaqqOGwfhZ/L07sc1rMk2MR04vYroGNG4E5idpPJi4N8MQrmgK5JHf6N1NNMfu8bKyhrepxNIcJFBhOv2E4EYzFCqOF3rPRVkWDPZfCKLGrBURtmcY21KTh6J203i+2mESu4xpVJ4aWpQ5OImKTimVDDKOHonaAGvhAYGpfK4unUlkZ4G+erqIe3MNc6NH1CzpchYVENdmnTg/jGLbDxM08+l4wSYer47nglydnHc5otE3QaKFk5PffEML9SttVGZ0tNa4zkReeTVmi0Ua4WHtfr24plJ128atKYpg3Y/ByIhIDcMeYTjnLSGjQWqIZHASPUZ5uBLhm9MkEAiF2jIwMImEA5kWJ6Uub6O5kspKbxIW/PqmMZgbihaOh9hHfbsVrqyse7gS1LMFb+ZiuLqIviUW5O+ol67IfuhYSalM+RQn8C5dKQtldNPpYLTPDOmQMa1pVjkstpp0U3MhNR1nKN0UUpPd60xrN/Emy1Dv0QqJx3WZ4s6VBzDIU6o9rX43PmAz/BE7HpJ9oSpv4taM0i0gIeDEqAWmyJKzKrcw6RLA1TtYNUMvBK2+N/lHihrk8meTRC1lM0sVne3Jy8/KZbzOHhRhGxXl23qnguSU3oRuJ/TlzifWoy8GLWE+CsJEkZ89r+8ISumHqNFqrYfkOPB6L7Qn3jlZquBg1Z87rqqUPiTig+FBA4ZBzV/x/l5zse2Sxp9BTjx39NaONri0fIwdBu4YGaJq+XdzvdSKfqIdVCh7Z97E4K0BIBdseCq50w7OAP5eBZ8PPp7GpKj7/wdjEGKBUPRTct+wkYZgc3ePqy8USRDLNDEadkikidzoVAYu1sAZO5ta1pMGWRU5oPZETKgw+VyGLnBXfhQU+tjO5/2r0TXm0waYKnDJwlJjXhfUHLLZrbgnU4/KgD4Evw++WcuYvstTP1CNL8bb5IIH2texuiI0tDhubgrUv0h8xqH5Bhm24O2Zub+0Q+qY3dvgivoi97V0wYJLufg3R0QnSjfnTgZ3O5lvd8HEpEP0BQqJCes1P6fu+qmMYgEHV6AkjWqiZzBtc7yVHZr8ZKBmRE8p0f6di0BMbZlpiEU63Yi98EUOUtqvywzD6ZCLFXvXvaI0nCX90b+PxJg9BVNf9BLDBcocyMVUuDf72dRist7UlOENnvACsbQFfWp/yO+RT1/KhOc/iXHXR316xqAOkiEdc+wLWVOUEN0EgG0BtP+ga2N1pMO01dH+9RZetcavXqWpCfHSRLYjsA91tOnFECHe1YFvcWvB2HIlPxO4P2FmwFohJu9ekehQVDxmtlDQIWFahxFTEmNZG81A9TvjD3GNrQ9oNnfyrL0VSyTvF8IzoTwqKlLDI6m6kokHmEfXMbrS4kkfPkvuZpVHJWk9zxTZmXo79T1pjodb25Fc3wl7HroerJ/OFPMFYRimN4j2Bo57haLEC+R6LcmWdVqYj3t6haU0nx1pOEeFo+Q//o24vO09aQWusl787xBtINIKSdJywUjfC3k4lTrZQXl0UfNCRPWZifIJucUNB+ZcztAa8zfoIYZx812TxI89RnvAImNVD8rRHfnI4aWnFH0QWuJ+x8MxF+V1l0pdMA2ptUnQwE/IEFlF8xAKNhAuM4T1RTu4hyMmOdTW7DeSoFkdicbOzQtJrN75zk3LjhZkG1j1SLqHb+cpBeHIrirBUIMFHL7pTyG9bND0G0AjkwTN9Ojres96BBR8uTTzmiFD5DBoENmUkta8d5dKYeeJB9lcBfB/yY7978Kjv00PdJYrZAYREVFAl3UBv3mdOElGbeYix4EHttQheY0djsjIzFdW1ACR+3xvCB871nMqHfYzhFTZ8g9Qc+5xS1XOlqPst8DLuc9eVMXQ/iExRi4OMvIqU29Ei5LDJg2H0i/sG+Sw8tIBLuRS2xec0ohT5HqEquFPJgT2AsQfZ6+OvFIrRrNsrRPZrCjAkcSst14Rn1UOnEubwpYO+QpsicCns2gcfQpcbU8+SVHL9IV5+BF4crSkz1LymyCR3LCwIOc6VkeOGpCNi8R/xgDaD7aCU1e1TsPi0mGIM22zuxroXHCn4wL62KghH/90fFLMIJ5t+s7/o/uY7ABEIhQ8MwA5bH8e5F0I1WvnuGGMgJjtEU0OcHCidUCRaa6Cx+KlReXtRvmYAodRHpLPoi278huaGAz2YdJZkDbSXAPeQhBEN3c2qziHYq3WA/2l/9d6dVbP/jJA8RxBUlyxeb0kt0Jr5LwEEGhmGmOwVjuciWNOrMymiStIfk6Gwg48fSFwgefJV70zgcSE/X3dhzeicQdojj0Zc07mwjzRR6sHD1KBoEDnwHNLJ8QMy7ojEloAn9b3kjQWDCRQXZSJvJwrumLA+7QCThE7rLFtpKmwbwq6pk1OJN4wD40LNSBYVjjwFKRSsgfVsOSskr/haP4/k+KbzJKOwecLUdWwLF+sX9UzeT6Cpa8eEExqKOTkFYdMW1nugtB6hA8sd6FjWj9j9zeSep3hkoKK7GeaclC1Nafsw6xH0cAqHtr9xiCqjACifKmK0dbT7heroRoRaAXuSiSN1vIGREl4XAnot2RRblBvXa+icOQkDXexHnFK43UHy36HrMSj0jdIVSKZCo5Et/m6xbG6WDHzy5svMSdJo7d7EvJO4cKhZpOYNaTEm9Idk4xaazY4H7oD3lcyYRSfuU62SXvaRxvOo+TpbU2z1Of6n27gyczIQrM6lxFbEtKbeFF4s/fSs2vG7CR5i5BzhhTBmx0yufuxA1Ve/4QzZXsZNPPjVEneefrOxa4l09O/PhFNDOhVc8sXkJDNrf07V9I5WtWSB019rfB9tr7XmItv/OXtT6O/O1eSJiicz5DHvMcj8nYt3Ob4dazrL4zo/Peh9mehbDVtRdu0oI3ueByxcQ3ruta6DTHyqmOp4GtbDg0PswfH9qgRXIHTqt/rJi0O8TYzkqdVoRmlBEm/VvMYWGqvO0DmQscjcFKUdHhtpvgw/D7gLi9gmRHassPcjGO1zTXcEmflA7hutV7wcpnhFtnSwNDTXsLjET0Mk1SjM8uzA5pzBqJGw0BsSC/0aKKzmNu+8MkpJG/d+9iE3EjzjCb7eix3mKn7sRM0d2wGGNfDJqUFV64zHCWWuz8POxpI5rif+tm3pgihoNRr0krkwA4pQS3yfp17Dh6AMCNAoitHQNl9MjqZltrjPcWJvcXrm52OfXzAb4HM73g3hmyltt4/Hh4IOfufdZ8bOHzmaY3d8dMHPl/2OlAP3nFbZApS8iazFfOO2SxzLssLW4qRghAz8m2zaQGaq6M9Bxpajy43CSyPMXXy9/ZaY7ltrzP6+BODVjebPALKOaZl4Wf6M+sSXydwnguxao7yOruTe2yTT8A8z88B9dEL1r3Xhb8gz8Acdze89rS/HHatnnqRGHB5dnYsvJkw4fY8+1zPPSzUirBopZd0guIrYcLXTme/AIaSOLp43j94QYrz3xtINNkK+DsrK4J1tw7wTJG8kio0KDHB1LN9saxR1Lxohrs2mX0ohzaAzc3RKhtC9xG6JKzK8ewJ1wrVOfoq/kKt3F51WGw751lRGDmf1MqQZJ6MBPPFf5lppKcln0duhq17Zxkzc805FSLVrnCd7s4+ax5GbT4LWhm0KWtu0qnNK49sow9dic2NsW+fp5GFza7rDoVG8V7vzksBlz640WiejAUAs52aAemI4G7WoHoRHRtC7yguPoR56uHxsr2q1qJbOEOsNUT9W8MyqTvRo80kwAWgivWxnpKm/5bkYFOKLiVFzmS2xYpkbGVaVTjEHr6wlt/yVFMJ2YG7+9ZHmg4Mf6Kwe8q8QlXc0prHHXZFwfEZLJuIyGiPymPrUa3nBp7fe3FiJ6F+P+3HNLcev211h8pq1d79j6Nb5/4MHXOjCRchCWeBFmQgAqKsR7k1zzRbO74vZ9ZW1bDQoC6KooEiLTkN9ffnNUTBjSgHzSF2T939VZutQaUyMav7KLT6prkt68qvi0EFIuP93iWPRs04/XP9PtAXlvbAFbeA9wf913rtuw2eaC2PxVe5J1tERUqEjOvNhHgUIkTBqA5werJL/1T56ED0YsVM54veS0fe1Ruv7QmyYdSPXzZbySISSCGq9gFO1x3G1Ud0berH308Jyj6CgX8roqB43PEermr7EivpSXPIlpSYtPigSqg7517XHxedLV/87A08FRtk/BCRILkark5R1ztTS6KST5MjaN5iqFlefPGEjtazDjpkbD49vn1pTnJeecfwI1GgQEhF2nN/vnw52gqmasbYE9HVSZRhkQ2lYwBbHRcsytvU/N/mF9j3maKYh41/+3iiKIu0WlJLVuE4x5Rne+VJAHytc+aoNug3NQqu8iyqPnJwa2YZQE3s7zbwyS7WrwGyBNPO38XBXeAJlroC7zdd7AXJJIBkxs2B0BLuoteOpxlHumDq9Jq1hGHudnE3SOw2FQ/V9kk5zD/TZh79Do6G57pdPhKY7RGyJ6DuqM4V0ibv3D9fcr3wmHjtOM8R6kuvBQp/NroSSFGxbaA8ypTILmEabrYacOZrx157CqyVhMoEu7kzX43n5BDwi4RhiIuTetmI02WVHhg2PDXWtKgGd6joDbjHu4j2QJqmHn3Eiq1xyvgd9Xp2mURt0LYzwK9ikBym78rmvX5d6PlcXQMQj0kQvD2k9yDUuWftOQX2T6vAolnvlAWpIJycOJWOZF1IM43z1eXcdfX+QNn2RSW1c3kVLrA+KHFLnLCV0aGLP/RIu+Ei7B1zMX2gIjfKmgEP5lwyDjMmi8hi/IUqEJJDY7Sn0oXe4nakISHWs=
`pragma protect end_data_block
`pragma protect digest_block
6d70d323d72376b62ccf966d055ca2c86067f22dad8287f41c6805e81ba1297c
`pragma protect end_digest_block
`pragma protect end_protected
