`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
8or+SvCcUHGeC9iYX2ateWQswmL1cvQzGIsR5faV3vejfN2rr35jy95qxF9TJ9CT/r3iOvOnjL0382d1pmnVXFicSNo7mqpzzoeJP2MJXNq0hUT9pHkCkKRLqLaMbSRIHnuriZjq/GC4ekRmWjVxtW7shEdhVFys0/vSet4FTpua7c7IgxHA8miAdmWM9Wwhy0WLDTyVykG/FD4qnavpRrrq8W5GMYK7XH6scaVoBy6REPxJ/ZgENoL/EjYQhgusnPpb9/PS5t7iDk82HYmmN6oqcJRsp+lyhio2YYGpZoTl1kwcgqoAvR8mYV9l5xgAjqcgkXdvovcKED988nyJIW/ikeZrPi9vHO+nmp8xBjbid22wxh1Yn7nXPbEv+zzpQRsZ3wMC1RPgJQryX9hRXHx6DSzTQ9GgHuXY7z3bnO5NauXRsOC3XYV2G93T1dR145pCWMU0lbOFBfJYQWon2MqQaHyo9jcZb+EJGXt5x99aDlI4gpuftjn+pw2KLn0M/7FVdVrZaxWAU79rIOMfmvrDkBCj/Jn/IfHW2wWzVV8a7wWhYLhaFVNJe/Qb/k5CseQGKeGACy8mxptwMceSxw/4mBkD50LnGYagy92DDB0V1r6wjKfQ1nVsUZOf29qIYjNdQPzoVvLqzXJeZAS0YIpWy1LmGljkz2E1TUvR7EnYfCDreQ/RwFUUTtz+XFMQxNGxK0aXO94/7y+/uQiI7L4REHqHUyK+hVduH6iXiqiSKXLpvYAWOKXUcOboCBxiuAWbnzGzlU716HNEGC5jo5ErY702AaZN9SMvqE6/NT7bxwCVDSHHOiKlwIYp0muZPwNlJbeJzOnKaMbTYgGGZiIP5NngNW8Ic2kzwAnZXMmPEtP1UfNmsf+9hDkva2hTKBip93YfrEw6qpoTFjhvfkYy2U5osWI3eGkWxwNLTUujWkDwe1cGHMKecXpg1I2Q9lbIonlN1Ru2YRwSY/JN1qvIy9NNF0ysZx/d0w3ol/ivZw8B/vhlJgA/BBpzjrIOZuv4jLGjWgsdujLEn4S3w9ebZjlQS8DO9fxaIGIjo9Inx/OARIwvLdRa2TTb/AE3p4rfI16R+EzplWnnieaD9xg8HxQsz/KY5uJ9+zM0aub11lCtIzdY8cOQNd1zbWgei6kfKs2iEcGqkFiK6/QSbSWeeR+dnSUdbUVRP7nza1fZo7ownjMnXJqYl7kUdzBBUmxB1NWRyzRJNcGG7jdVpa//iD/3aH0dVTSY+Qa9/InQ3pfvtgcb2O5ff7CQJtml7RBlJBGT0JQz8uBWqtgOEOv5fur7s52oJ2l+r6jgtT8TvJdPLrPkffDUn2iOKoYTIa87a/7L9XKv45iMa3c15gMgVzN9AbhiBoZQ5DMtgzYz+1rhihRxeA9Zr4YbQ54o227YbtR1JmDFP90Hs5DHyXohsKTJHbwF+7uOxtNxrgx+NPE3O7lqzIfX7/8YiP02fgIAmxphh7cdQYJOOsQ+gLphXJGLRt0an953TV9vn2sjg2eeCuHfRKmnYN+kgJuS3hPX5KMNQ3wX69hh5hj01HmUBSezODvcsyzeNMXCp7fjzJyxMwRO3zB/gsKuz+2V3WZSArsaEWKh8qLSEHcjCnuhXJfRfj/Dc8lB3OOCUGdels45L2P52UH8DmF7NcHG145BZYiptCsrsebJxLnetEJwf0VhMh9XpwikusXu1w6w/25W8Jkbe3VRiqgmCAdXgJJCv2iW5/sLo8D7r26L8sVAnn9wZ7vFSeCxLckwDDLxBDyO1/4lbp90/MxxAUToQr/FoFNetGEp9n1ou2XoEv7TR66Urd278P+egosUVxyib9QBUMNwsARqDY+VkCAqQxc0MKzW9zRvYWma0Xgrlp0IGHFV/P1O95fOKWkAjo7RM3FoUPL4d24Jaj8JJtnJ3L0bXQhVLPgikDXUv2SX89NNW+tr+xp55QUrDhRJ4LerZuNON67ELgReJm8XM+NyQLaW2SYN47neCD0J4ANLjJW8Ms+OfcF8YrSp3z5vGt+qBIXpQYsM2BOCuEZULnOafh5vejFr3S8zyrJV2e68z1ZH0j/jD3SsUwspARW6E5q9gmx7UF2Cdye3SFE66HSWe2BwSir8loZDGH8wh1PnoHRqqDdtKA6VSNz29iMN8HMYPUTOCxGXGsVmHeQWuFq8X3UPA0pfvP6/JjgkwCoIDitjEDM19WAaPthsC3tjI1sLc/jlMgjgXVHg8QzCqk/TZZTV3yzs8glBUpnM9bpQlC+1Ir1WQQxUnsvtwFaVarDszya87JcfgnWOs/jndDJxg7RoFel0tgooNHQU81rKhLrPljcPQQjqYMEd6QZRqXrOimD9VnrrWab3V4apf5JseL2X8bw9Bh4HA9kQGfYfLYA+Og5xcJXZLDuPLGoku8FEASj/WtJSV24HlBf5i5V6qsxpXrwjBHJb7VHEUV+BmQwGaOM6MRqE+cKjFfHiIrEXuuOmA+z+0O8HVlttb5ArLDvi4tsTwBOMr/wY2ZNqYklzlX84KtUK0bbqdtEzRQVmbYgZJrGQC68fWxy1PZmdHINcWQ+K5ru3QO5N4EbvsbCDqcK5xAOEFDTMBP6ZznDD2AJHU9cYBoaV+ciJr4XKnjF3NnPgYZS6Y1lbuSs5QsJxAjPwsQJM7Y4PNHetrbh8QpLAc2rofnMAdNcu76/k78lghsJ1BrRxfjxb0jU2JYxXk0UwznqIDDaPK9IGFv8z/TD0ovytfnP7eeNgFtEYS4+xLNJlRH8s3uXsrHlRQgALwspoEFHlVPgUmUmlkKzDZVepXQ+cSpg8iMOjRTYDo8Omg/4D2+zX7QE/c/JJRfp6TDtyn0JaiEoSJOIJdru7ytFbOT65hjOZoh51ctE2phMALmX73LL5G6ErS+cojaTOxnRE6QR8mcqMvPPM7I+b5EyRWlLAz9bbbxwMWOmtEiQkJPy4WCbMszCpAQicmlKeq5KqjnchGfhlmcE08sLpQ3Sbo3UFkqFREQuYwQNI/cq/sKaRTWq5gaF6lEMn4sGOPFYkABGP2H9wV3HzLaMcJp9sCMTIJ60/yXEGCD17QEhat2bEV4EnM5SmaTQuBMocUeHPxl9sbWi3EFuuNymMEx4Si00EOlpm1xYCwj6rPYOyWz68jqq1SulD6uhRQ76+NI23LSf+/3NLvj6C3O0Gse9lKRVwZovBFTun0ffcjJeLr7M5v9r3qIdj6iccBeMnjpc9ay03hbUkHE5cgKLfpcIre5hJiygzwopgI3g24GVM1mfioT6BWMu6x3s2sidwVqrDtZfhxQ9h4hhZ4EpNwD4q6KBSUxUOwDH54g00h2X91eRtfqRJnW9KvAGGS6qRlCLa26FzFzTuJJSX/QiNQIKDlDAHmnx45PkQpkdO93EepiEtlV4rusp/rqK8Cb9WK2jhwu2jWdxjKXd/J/3+e7FMiIhjJJPOV1dwmpIFiYOnWtULgS25iQLyN7UlaBq55EEv+l9c/wd8E990xHrgky75oTzJqd4X+R6NqvYMHgs/L62r7e7Bh8weUOfbL4l2O6fR8DFwl9BONxPJooafsK5SSLubH4V19LSYLRwy8WJ8su8kEwwI3h0AOX0m06eRU+itFTqo87iPY744DeuwH2P2sxq+/ALKuYl/H3rkuAFZjDXUA5OjtbjWYx4dBUgkwCjAMrv7GcVopBazEi4oLHn0dqga4DQz4QJ1oxu4cTmnScffwjdWaUW1XMOseNwcTtpYTXklHpivqjxOhk3ILKxxFopXDye0iQbEVRe0mFvSXpqIrD9CDYyGAFWVcnY47FlGCAybvWUS1ygb+/AEAWYptHXvUvTDwD+10BtH4zN6JCPbDAHUzme7P/JY60ZXf8AWa9vtKO6Cb9J3zWLYBG4+aWg8Qc952ahyFjGZOqWhh0d18f9k7B3RF23YjAozeysD1SXFQx0MQ5QQH1G/UvR9XFkwln0vjMk6Olrccj0IcBr40hJ0cCiS+c9acN2tQBu7JysF/WfVrdv3HVbz4WJKJ83IRREXekojwXp0682KZwh54gg1yvcrSYZbblr0peAXHU9U0tO3uR1sSN6fKEaEjIZhihI6tHH0lnqRhOqRDo56PxNmiJz6GPywmoTvsA6uy7fvWkO1/+w3bWXojMvsNywSvN+3IytolQWsCRleEsHaV5V9ecsepwiQUhvCq2ixNzK0Ve9rsxTeWnWzBeAEdI6YsGl3diwcCkf2J+sCwfz0r41kZn+C9LwJY0WlhjPL61yLoXS/gNz9zyTkWSubHeAiqSvd1LX6uzvHSbeer5GKPNKowpxm5sZQSXt8RFqsoA/C7ACwD+OTALxIIPk7Yau06jPyuLZFazGzBvIzzdU5FNTARAX4qwSKFLjOl99ju3h2B18icHynYOHVjAN9P2rc3rtIXGTZ3fVq8Ud2y2YUmElRT0GcSzZmM72YQUzv3NzjejSOK8orYXfGfuTJsO6TcabBGyhs+KRISE/pkFcUx5tB1durONmwcmzU44KR1JWtGCXt8GSGmlTSk5M8fkoY7934+iS1YttRbkzhOEqx7byU5UlZdH1J/tbRV8ejtaYAQ4bRTAaRwKwS+q73LfDM4ByIdoP5E4n39Fiq+nIKZ3712quEAiuQ3AwfJZmDqeFFe4w+2VhpWlQGbOgZ0wX8/j9lloOLD48m4Rf7hPu7AJArZ85IeatmkDOmPTYZWvYEKyW6AemhaqsVwfKSvgp1q3YRyLnF3fqAN+Hbn/etUhnBZ/6SKnPeuJ6/Ve0+4UiX2p6f1kuF3t75d8OQhszKg5r34P9Tn6d3/ZvO/bF9koGOBtWxAOdUz7MPv+cX+Th+vmV6q2zNeXSWngCVQvedJHk69qrPjPB/FYn2OsSAtomFRskRwROCYeR1eNT5xcp59PEsudRg7zCpqjxb59Mepz/vQTGE9uH9p3ZIHqDIsPQmD22iC5pn/Sax7q9kX3OS8atxxliqbEFjCdMk7ksd/g0+5k4xZ3cIAGhNYsycqFGSrVMqELxtW0JZSffZ640EmBP5B57MG9PI1Ai6P2rfxROR3ZPn5YPjFsSqM4ceyYb8ah4uD9Fi2MHKkn64iB5gT3LcEMa2jSHG+kK47DwlK6ZDa1UClIbTEDlIaz8FHWgAeg0sJRZbZVfZRJVYtn/BBn8/fXbYCXLEzQpcp17kssNT9GH9ToBLGkq56HFoHQoNW3gFYXxnimM+5APHUYMQd0xYpO6oMyZgHjSv2Af8ejf1kkNsoTwn5bVFWqP62eOmXpPwfAcLR32R/dxT7cAjpPdLY/K/xW5P/oHUJk7y40ZfnXELFpg4y3Q6xko3IjE27y7mcFwk8/qtArrhk5MOKHg1MB+bgdd/rPQyeOughNbEArPur0WxpKifc5uruOP8/9DVKSFkv4P4ya748in3H8h7nKyzGw0BfrqYFhHk5HlO6Qpmace5PEcOcra9w0E7oWcLyEfvHHtl+kbnvf/tIftah81SW6iWp02bzrjFnULAW4nn3TPD1y9t8cWB9QW77tYjWzNaocC7w2gZFT3GDKIVtHlYulnJvzdWtSpE4ZRjjaF6XX4XPwgpyg1pNBqPBhd3UiMNOVYbICioKLHdR4oZpbXZKfxeG3eMSQTKj8eR9O5Zp1PR7YmKwJSQKnTkhjV4W96b4bCchmA0D6nWth31ACb3/Cv4Tp7zqdz7lDyUDnAnF6xY20UsQ8ZsNTZy8Yi51w2yG736S7EwZNiIo8qtOgB4kvVWOroXBB13me6kwdoXblpmKGpRaRQr+GXK19oZ7osaPW0395LuRggsJNXpVcIoxEKGLw+K5DPWyTBclZRY/Aua1+Q11Ubh1U88WZFbr2VrBnKT425yUoLXii84r/+9TGnyKTrPQuNVgpMq5+ZAQQSwlNGq1xZwfKpeVjlHQSnhA3HBBMx8YKRfW7HgpJ36TNsJpH3FfagCKB+0eWgn2xKaQdkRV0Mq+pHBaccUgjfL4GKgjFzgeleAHaxOZdSaGULDZj7Zer5lrHsdX8wnhOYu44F7At3XSXYp1sYDJGD/bxONyPPRnjuYAEtRW4uXb1IPP29LfY8/s/We3+0NlZf21lPIU/sQoNX5UfrEHS3o0x0VwymBKUkrCzA7nVWVjvysc1f5BQxvSTUen4239Lq9aqw2ym1kozO7HqKNK9lV01KIkf2zce8msE45zSF7G5c8OlcNmo4tb7Og8AgY/fsjb9RCCRmKxhLrzvFJ9+Y34c05rG0FxbUs4yFuKY5WAsC/BTwxW3q5s2cta6OpMYdMpwthcYTq72u/xvV5XTjPYPugEfQ76FTzqigQeKS0PRGGOetYd44ocyl5aHkezQnHO3m/2gFnrAHgHoMWLLl0agSytLOIzx4slbKLMP8OA1cQRgFS/4bz05QM3CZmMquj4Una0XzkJZ8Qwo1riCW+03gjMqlS2SntFJKlWjb5rmp3SrfmUiNP9XQb18j1h1VsrHS4mqJL8NrXvhwpnFyarae/vA8G6itif6ZFUuxDRVlK/QypH2utBQ4JvKGHLwfX4WQnSiWQE9Xo7DyIBvxHjtGe2UMjKxdTNxmaHd2WggEujfHPnkb3Bh+sW7xWogLr2XMZwj7lhGCB2OEcWl+oPfLX3aIU0lFXO/R/H47hJdRl1xUCU2FEG+xk5F5/IqXx+SS6XjGlWM04rEY06S33f3AdQ8xGrp63oaXlgsY/6TguTnRjYZenIHmcYsBYDsdvtK+NnY6HQzPahWiAHa9IXEtlwNBSzRTd34XtI+llakPbSCX2xBNyK9OLNIiDxy5Ac0UDbQWJHrWQwhmY2UrL5rkAC0o1zHd19ysWN16nh6T9F978FOcFatQ6wTMb7A5CBT3GfUWT835uogZcS4hPHJPw+V6L7HSrJT6OanE/4LUImbIsyl7UItski/z3CmTAaX2IF9GTJyqwbW3BzyF3kygVNvkLwBeJqe4Ey67Sl0ZQ+S2Ur3nTHUtkjEt5Ze1MyCpZLgjtRlilKmS0ukZRyunltm3/rFKMDhsVZS7w1QprXjO5AnHk7exW0wZL3uKsMH8SBuYVGsAmmOsRo0zRF/Fh6GJ+TIwwzlMJkIi4W1b71pkqm8IsGuFFle/4+wM4zGFdgdS+/npSJfEzdrBFAqPjMThuaVS+S+46+eBdFaWr3wfZFwWjJbln/3+D7CinO6p4yZ8+Rte7r2s/AcF6FlJs4edz88a2Py2WA9UNTfjlMJd+7yDWU7HClOClZIS+jnswnUKUenznVJaOb+zxRwCxOeOf0tumUMZXFUrrjS99YTlQBRGNMhGO4xuYuAQEjkPtOrlt8xJ/MqPi7QXkgTGRk5tuio3qyO7cz1lBQnIWjIXSsCK7oJlfNv5oEJRFLVOvkfp5KtpFrZCRLh5p9ux/uyggGkYQ/NIdamMba2DDA/B+qS8RVpvE31HAW/uFJzFKunjoyqRPaRpQ/+2nb8UdmG0KR/9wGCslsF09LYSuUeuoJJcpYi/GNNpiNx0BOb/YWQxSw+6z6DYdMUUDkn5wtAOrxM2xwKPIbkrteDvMNqsJL/7OUoOkF5kjo9T6H2ZLhQieO/MYgbirLMX8BmTidXmaYBSOGromJtCVUh3T4fe1eOilp1x62I1zkg1R6grFOKnZaM/EEAxqwAoocPAkzpiT/FfMLEmZlrdnj2G0n2qB2PN19E3g563VCZNaYaOslFyQVHaORmQw1U7C5MldfBCH/QvGX6wJgaAGivWbyt1jJwnmoYyPoGb77ZrjnCLq97M9xMhz3OElu6Y5F1WJQJ0GayRt/XZ24tMkeSolgYTbXtpgqf22dYfU6gr95U1jcOSgVlPZR3GvK34f8QMIH803iMAL20Sa0b+u1sCurEz1AIn3qngYof9V5wwU67NusnZCyaWaVvOfzxTmRFsoVkfu9IoU3qYhCMZn6JdKu1yIAQsOudv/BqvVK/cAeigDUCFOQkCHd+/McGS1SDBWo/M3kLabF/8+QcdJAUsMThC+dmIQOzeKD1wELfBYKvAUOsJPjFLUibbgZHjmeYRmMO4Y8vGBxPycuA/5mqJQi7LFzRZi2kF2id1Tpmabcc2Yq4YtLrxZ3zGD7q3WSWk1xuYWM2JpppOWJxjGDXZ8ZLVBCv3dIrypmEahSqqlTd7+JsOAyRnuvgjw3h1SLypvpTpiVOE30bhbAnIBXjhyklqpk0WaLuN26mp35tQG1qfD36aIV6uxF+NcQSJ2BhJ+2B4Hw/ytrVNjt2xjBcrk2N8bczfRtl6Y26orRDdBe0Z0m9FKs4vQ0SLDhtGbb/Akp2vUZiPr9orLM61TbIM4wUC3Jufy4besndlO8KVyCTUD6t4J8FN3zCRv6fPDLQ3vL3HrCU9EhvqTYuKN4Sc+c7znL4fTlx23QX4KTdNsrPrz/n6HoS/x8OyJQH8XwqOz8yN+CCBM/CcABRUWlEvhDUke6ztcmykmib4kIbCEkR5/Aax5gmvJ8CWdohtITD6A7tAz8UXY7CXwl1bViUJvKa4J80d60koEvKuVYmDaTy8gRIUPVso/9FbAmQNjwh2rrzLOKA7dD/MXSldKKadj1ojq0rcQ02Bj9QSTbks3ftRrxPdi7YvcFOklQlqteiw2ntSpkxO1anMhGE7IZz+xWve1bZnUED3pmrfoByxiF3N6RgKMfxzK4+mcMMtIMOrJeZ9zjHbRk3fux8XnCMlRQgf+fzE6OqgkwX9k4tevZVtaM0ZkFgY1QWC2iJCNqVCj/Wzx2IgbL8YVOYnF5KspgXZ6PAPYGz69EllxPRzwRUPUfi+jdVBatsOlB/2RwylEW7nzHTVsQchy+zurNd3WsFWBOGs0lkd7Q9NFUNHQpOJOabweG67KEhvZJ1bIjfXQTXi0zwBBpeB106jbkl0eUeSXG95TW+3AJxtmUSJUDx65CmWd6Nm+AG94AxF3Tef5q7Dc6vsuvKM0mOKRr+G8CRX71w/JLPQXSwjD3VuUHdKQ9lSppN756OjBmlo6J1OHs6jH/QW8b2IG3noyqJtVzn1dSd9k1i7YQBL7yZkXIahlflxmm1j3Il/GLp2y4W3oGc85XBVIozJ1LJQlJd8JSlENaAjiXwa4LAScSjByRmuW/4OmfU/XnLKAyl0GyhelHs02BbVYadmURLuumxPdmx+6ptu21cR94kHM7Tf+80D7p9f0VpQbAXTNN6LqLtuqWZPbSR8ZPGAitLLHsZw5a2uvnV5IYc0kheb4mgg955kALVdNsilrG7+OLoTkTnfWcb70nJVY0lRfDtdkl7/GQcA1A+IGWGJc74+TWwAOqaUCilcKYBRSPe37k24NFqkvd9oJ9/LnE0B7QvUgPOE7vwa4gSsl1HcCDX6DLRuyPE5ECVCXnrmQFqwBCrW0EO7Z7Cli14ibWNSCtMmpJl25sSWpF/10GMJLGEhPU8iOMWMHpQ71wpu/chYN/DtOvtvygTOpjQgpQQqGP5fEVGG6vziQvmOmc5BZkVV5YCDnpp44WMhRhr+LuCf029F6PbTRJqCryzyfGq7tAwskiZ/nFLNoreJgMeRZ1DBPi12xVxzHgGhQ+9U4msEPDmFVmoEwscFdIrED1URzJK+eDMNSQZdbZzptTfSOnp78P8/NHYKRK3dznj0DMLhGy9g7Jr4dGXzxSvciN020rRihWm+URbvhhGXxn3zmSqI7UfappEBjC+3BQWz3Wa+EaHVYrUCEnJwU2/OtahLUBUdcrE+yo252JyyHC/N5Ao54aOyFKtKr2d+Q/Kg0aK9pAIlBLocnoIWn8cJbpmTwlok7wLfcVgA7V9vIbC/rawXWMtAOWsZXhcnwtKGutahYE4O7/b/Du070RqEccsGBoNI4s4v3+FC+j8dCUMZTLANvqE4GKGc9L6tjRwLzQQA7nNJ6ObSsQZwxKUvZHKuD3hOWE3yEQQtnPH6Qu0UqTnltomcouIMzm5bA7MVbQfxgDym+JubnQxKXvlA8x3O2ePhEiXuQrxtz+P9FhCJ8XqE8n5i/BygxG5DaSuSWFhKDTfq6uUEBtQFw5PfQGlEsUroBb8dNYwm/ru7Do8Hy8WubDnfJJIDYMHKxx0evvQ1EKDrdnYBcsoiGgCBtk2J/Bz7oP7P2zQdE7q4B6ztBDH9DddBjj6u6HitkA2e4xw9rENztJtmFhDzEcbUmmx8ISOxSmN9FNXR8Y/F/As8HhcATqz3OEircZfdBtY8uNJcnNGUXkdiA1uRz+5CKmXsjfM+wVm85HkMltTwU0XPgNEJhd0C0h8DJtnSO+jodIcmAiJbDIm1yiWTbZdNWci0FxJEOebbH3QQeLKHjmokn/C6wwGrE7queUSFC+pNqM6Er5NPLoJ4wnSNZCxS4LujR/EuV94ihKjuYsZEYDX4oLzZAZh4xGuSBNZH6rgdcRmzLid0GsHn2gtNcdAU2rgBDaEtzJq8b0PHtnnE/vMRiHhOKJ7c8yHm48RUmAr+iQwtVifcrbgatH9osSIwjxiFmcdWdIXMFtAhj1VCjNUjXtXlrqqZA/0Szz89TzPdgHEXveKBcAAtwFSK49tz92sFihZ8wbSWHhF1+yxLzQKBN926H/lmM/TknhExzV83wRQfygM+PogpJOoCXvHTWURYMj1u/0rPT/ispWoLyHm93+3U4pLTD8eK/YQ90g09Ekt8iV0jxbNPAKU0bVRWHs/xw6aZPa0P1pn4BSHQQEMrMyWhPUon+5Ob7VUvnp9lwMJAx9f7Iqqkew8yWbFdqqGJMTopsANXA67zWxTihormnoqWrwQGhnOUSjwk6JEBPxVN5U5d0in2mPprDdbD+e3n7YRmYjVeugwyNB1Lg/tcFRhebyt3W1qPvfgdQC7LTU6GUHZ3+6JuAf6lh+7TVnO0mMLfVfyiPoznh9RO5gW3G+kZHxFsJPFUJQ1yUx89SNAc7cAmHEwjk62da0uAJlB4/o5oHmDBlFGzSaOQkvYEdzJ3dwB6QaB1rdnJmmgQN3l/toGgV4eqmuyqgg7kbHkqm7ahkN3WUwpp+Gs9uQrJFqEPTMuf90tTKkGYfhNsFgyMoZutKrm52pJAURVJZxhKadbZZf2/KF4Xr1gL1tw6qzpSZLChzPX2Mc2RpeeTYEvOVDPymqsfXWnwYBZToIjzbzN2/UeyWxF+3r9lkUTDZaM7bDEjzqKcajO6e5gh59Ndj7cbDMTeAkqifbhKzVaFO2XLYXHHuGBzb8YTpEW0huC4SbbeROWm6Wek24fkpL+Ps+VKiwGjt3QWiTZsXg10tBt9giiQ6L+Ga8bEC+OgM+R4O2R0otV0aVMSXXubCrNU0mn8R+iPiRx9+CWcz2f+ir7IVg+tU6f268ZM5BaJ/nzM8a3H+iawtIy8AcUKiuPadn5+OP6yvPuBxgPGs4JQ16gc7R++tDtiBxPOEt0pjROVhAyluTi7s3jnkjq2E72gyFfkpGqDbicoIS+fnCezf6eAkvUK6Q6n+tRa+tqd6mWCpo8R94cPV1PwjD5azh2KZxcIZHdmCrOY7Lr80IsfmLgWpJtC4dn16SGMnr9lr54gPTPo38y6Lw2YquiIyqz1JH6Yrume3Xg/6Z92Czf2IqWIjoa3g7+jnJIR8B0p5f8PYgUIaMRf5lc2XGAFjSRRuG2B/LCb7c7LrvoYw8PBOnB+5jpJZ3bw2zCW96KxjIgbbeyKBSJhVe3FGxLLUw1Bs1jyrALAyCUqDW2esHchNj9kOdZvSOL9OAmu40GQdpaD1OxbK1PZ1wxtEnVXCu/AV3NoJjYyAPhSGcbEk2wCxm8GkVjjiBXJeQFU3v2n3X5YsqMalZqeLp3T3p7kRRVo4+6oJyCe39RjdfZs/36B5sFk8yXs=
`pragma protect end_data_block
`pragma protect digest_block
6c6836e77929971ab8719c66986159368f5cb0635753bd7aa272b332c9184ba7
`pragma protect end_digest_block
`pragma protect end_protected
