`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
NGMXSVzXpaMoxql1KZTLnjWg5Bur3eeqfFu25fgktvdsCUK/I1da1wffwkhdQmzgssD7ADIzYGw3NM/ILXWPNEEZzcIR3OprcYreNwhNUloqoyf0SlcTU/fxupV4UuKKfYjV2RbYGg01q/ugLQ05Gi8KEU1LAuBHZONsZHzEtlD8nxpOIm9YIivzRDQWKtOPG5vAu/MgtYkhocc+L8kIfInfnaND7QdKSh0gTMxYlflN3TfWCA6osH4vFzXasi9XeaNXB2aIijHS6j6jFqp+SO2BvxsKOAbDf7r/ZoCBB4FtVduBQhfQzlyjkHFwMFajiEI4B2HRkvkq/8HfwIVxFdwsQr94MWWOk2JpWjgM0y/tEvtzVa6EUocAoMsLZsCF3outuKU729IL8WWqRXPucJO99fIGckzZq6M5b16QVYSTMGqXyQOVwS1GjGvh/w2cz7Gk3BRvhMx6uTfZls5erROhvrfoel0ZKtHJIzcpT4Fgiv10zbN8MTiSS5b7kGsDscsxqkZ5XDs+gJ1OD8siesOFQ1jYQAMPNjHJdMbu/Tyx/546tbxO1X/uw4kjPYZpfI6dcUqUrMh7QP2Jgnn6ibooRE/roULNpPaiTDAq6ti9ZyTf7tsAfMqKwI2b5UNXVEDb9MNHoCQsmSo7AF1tjkoYPad4cTVVuJiNS+1OSvfZFB+6HTYcfLgyEc89ZRvE1dAeJKn+Wr765Incnt2Av9YP8T8JkiMNY1FyD4OkJxwGb09E2ETqkYBwrgR2redZfEJUBgIiAJ7KM5PpidzAWltiVtLf071ovODwNlvmodPWQR6Vgbc58iU5CqmUKjyJBxi9e03dPcKD4pdgp0PsqwWc409JGrSZUOBpsupQNg3cKWO4Ra41Sk8zIJeIC0oad0ya+jBwC6mAKBuA3oWEVXZhInKVlodZ8oHKfW5yENOJct5JuvNDk7B18UVq7v8sP4chY7mERf3Qr1licAt6tA/lhP/+nGD2tHpX3/K5wFdIBtSM6axD8uIuRWZDLnJw/G+y4x0+wpOyVauVdJpbATbEKh1zJp77goICKnjDiD+psb/o0dNeNFzTMs+Oc0kZkraTxaNmTin9VHdxVKfs+fmxwlW/rS9aUrNf2XGeBMQTgWr20tc9yU4igVWw3WuPqhLY9wKB/i2q+pXb13FW7ArcHYPf4ljONeq3XJzJnZusuGSJhTEajEj52gYzTfEJYCQsxt+L6veW64iCd0tUH+F5KK8wq7KUg4WL1SsptfHI0J8scCdn5mj38rTnOhN9QhU7XVerI5tzUMF0Zyvvk3u6YEmSKDLm0+hyd/iLpL8JZAGas5Dp6OMxEs3BmnuKpURMFX54MqXEnE+ShSe4CRkB8Btev9a2A0xGnxoP84wSAdj2j3btgM2BBy2TA4T61lAzIWjV/n3vp5DG+bY5iPuia2NvYJUON4BvTJ5Y2JWxoziw8hjawuuKssCtCCv4O2ZhNvEPHvxheRiDwpBznAmkWpWAH+AvQaDhC9HbAAVXGyvbGbzFyq5lK7It910pJu6ADdyKPeYVwkSXDy7CedHAEAQswmeI4sA74VwfFaizorAA82WWU4Xl8aQ3kGexLvIf28YE1CEwgINpefc0+fF8ubCL26/0EHHLtGKRrXOFnvaL8Wd9YhzDHL0T5o1bllxzXmIR/mMacy3T2dRFcvPSkaaijoxIBCyNx0YR0lfXdL0vYwHXkNG/XV9mzUwl9rOluyPnTk56fINGPWV4vDO2cssplxy+VH2mdzhU6+wzGUKx7z+39k04Vuvy6mjRoK2wyQyedscAPOE74k/LO0l6O6pwJoSp5TolbmXbKA+dPD8h+W7PLD6NnpNmfKg7g5KfkaEQawWpE9lbm6nirDMf0FiEVZShD8FSjpxyVHU2JW7sOkqoRnl6M5ug4Vdcu9chMl3BX9SwssioAOuiAjBmAQzk26no8oWiT+BXzxPZxn++DEfzkKp+0ioC0r9O8ID4uvg0RPxrcXMKFg2PLF3uZn682hH5nPJMUv6apAwjTFDgrEptzDnUoW2CI/JmlMx4cgzYWw8NFslHExUhIM+9942FK0KFU+INzQsEnDji9WEUsNfMH5tKV7InQnl/ryDomq9eKQbtRmja5nb2FP67tqctHoxD4gkdBCxh6JOYmdSPaJbdC2cc+I1XuzN5WFtr8TwDa+ybQOZkw8xo3A4lYCuOpsFWpZhAwqZEd/2330Po75Y/yd8ebpY6EzqNkMPeRUBj8cYovE+6JSzgaKaF20vDUCwycubh456Kkdn9NI9fQpcdCeeBpKrodgBf8P0bSR+Kf6QVQW4Z7ktP1eZ2S/fjEgLt6xgTrjRHsaLCqY8dTGJdA4x/TlrWJzXvhxA5+XGjlM8HXlO9FmKdLa+Ylm598Rx5AOQRIQXbEP/TU3hErIymzcTbShrQPQhr/9E+n2uAQ2bi9JkyYhLM9mFzmKjMNBmylBLAkhiyj67JYsF6MA6erT/3ItkHHgGxnsOniH3m/HxeIpabG2Y1uyadRbjZIk4v1UYRtPX1kN45YQ999kTweEle8q+B33uCAC3nZ+4CqUGY1F9BfIi2wQQZ8DeAOIv89bvK+VQuMsdxf8UmMIWbo9jjWSZzIe9SdzQS7IC6EZKNdK3YKg16BEpeI7BpwGEgBvZg5aeSR3U3gp1veNsOiXoy3anGgbCogNjYzgTEHZO2yZ7IXjfgwemlzuITCUq2afarBufIcAscnG8QPYLYfcxgxFVnc3dJLjDa9c3oDyz7B/CDE/ee4Sc2WxjjCbGmRG3CRwyY4i8Dhs62biQdyTe/SMCA2JGS7DIIB/mlHpOUDoir69LR1rnnegprq27h0I5rc3ewXkgt7+JIS65ofsjvD45M6zmWArf6Asgy3H1qw25VsxAxKeFX6DhJpi95QppFCPzFnYKMcRETw8lcjT+cjzlZ+Mi5yJDSbXyWxlCX8RAu6XdSKPS3sXyVA50yagL5YRqXZyOkyhwqXYmJNjHaiAsttKlyG7//9mIqvU1kB5ZRwQ7i722s1x1EezgBc80wlIkCvol0xl6drUctQWn0a4+i7vnv26JzVWFu7cV6Nszq3zddkA2GAE0NiVNBrbPZCvQGDnkJ/uFMcrCRE9wr+HA7d+wk1tEb8TfaClxoMoOILfkqt4XSVMXxmaAHnBSE/xeTXd+uCkSBDejqCUXoNqfMacpfRQZ/c0yDJ6K46Aiy1Z69VjTHfzjJIfPt8YDUa5ZxHvtAF6nzZfVVH1wySJFJvJ7ChMHw/RQe+C3iQgcegVycm/3K8xWkVk0iro7aiFSudgqNj51YRGksJg3yQ/Xqye9BuAr2mRvSNk2ic9RZ7YVnzEvNvRj0Tfzh3EUnN4Gu4wK3kWS0k21fJQdZadoSi4HD1T/N9Vl+7C9uyB44h+c/BF4rjtEkOZGd/8Ck6prYbHr/Gc85xA6tFHSikO8PCuiYZXfvQyku6N9rHcvCyRgyxEmuLE0nsN1UZHCagE90IU6qxSQc2Qo1GXs48cUQpee8p2kWC1pjZAnQKD4Yaio7+mA7O6FPgFGUDmFWWfPVt2hX5fNTeHNrXjIhm9ADmdlDUsUfd/ANU55mIgBvqjetUeirdMfONFrOABXynV/ujUIf0IPnAtGNllX3rMzN5sSWIc0q/j6Ji8t8kXYlmTnQ3HSKsz1gQvI36eMGLOE6IvyoBNxGBz2UyyGOzehshANg35cyVwstX8KgxJNaKclKnRMG1UFhATDXk/yPwdl+ALj7NB6QEOQq5VbtmXfmke965a6XeR/1mtIz1pfOtRD2XLqE9CJF8i/bdqACk80fz9aedOB8jN7J6FayH7dHoP280ZlvHpZos6+RQuW99NitBPzvtqTqQlNRAP39d2XseNnNZX2mIRHZlNG6Q7mUSkYzcvgaQ8wYG7MktUmDbQV2SgsPcxUr6iBR8n/2ZqzO7kZg/rcb4xBzlKe7Xpd7O7Guyc3Xk2hb3K04JMLroe16eCxH4esASz8Gxjwf2UV7vocwNZ9y6VWhRPyCL6ZRcPM6pzKHf17HOqWIobmxXLO8219ZC0lemBLRTtDvxTYyRqsJ2Tyksupjg27WdAuv56odC5Z9h6xyazGF6QmH2t0I2r8tkg9rsptoM/guhIlyksnMnp93cCj9O7OIr9V/7knwmNV1Cw0cFZMVFtVl+r+yz9/Gz50pVY17SpOSnWuLJuIjs+tUZ/nYpSVLtM8mCN77ABds371dQJtuRFjgTcZYegRDWXGSIiIR5bxLTz1pioL8CRPNaqE5vC9dKoy1QlzsyGpz45ZVki/BBcCy6Y880i5N7SfzLv1aM38xrhY6cE9qywo0mPvFuiNEYnzskGHJGqKCcWVy3/Waq8mvTMN6knh3UfScVQ7BAMeJTxKBDX0+RXA7u3kNJFbxC0cHdzq9CQlxc1ddK1MWkhgaWirfUBdsN4Q0L+7b5mOikjW04jjea/Zl8pWxvJCcpOpfNFlOmHmyNOAYCZKgh0LufI2lJ04d9+tcWb+SyL/Gnu6doncJSNmXv/hqbcXk3OnGr5ALfrLzqkcKvnsAP90pCEybqbSaQyzFnm1Y/Uj6hukOWZqmQ3XZvyJTa2QV+e8ZHIuqD5FhsRkt9Aqxd8DtITiA537zTSk0OyyBgjI/y3kQQFG/KwImAwMwzYp8YmxrBHnTAt4cDBuqLRRj1F3LOUY82WVg5k5ZVMz2NgkegcOGd0TiwkDYdpxNDI0A+QT1oTDEcX0ecLwIHlP8N5i4Y+NxPHIctSNmm/t1IDX78yj3Kmmhmy2LBLsnBg/CmtnQ4adaP51enOeAiYcsoYgJ7SBd60diL3BIUHug5KqpYHmC6qfOb6WRo7rDPwLEgnz3W5ht+B57OqhJpIoxeA/B9kOhCpC5WaopySMFcnnG5yeyCuvpBSbFx+jCSFDioy8AonR+aHf5PlTM48uOKp3e3GD1v45MbYt/AIoLBo2vypUwRDnUP582Y4LUXFRHWY/51s4VRCa1szWK8jXdtgZFKGIByrN2hAYmJqhljgO96NO6nNZK5Qe5DNgXdBpxi4KuT7GgaqRkrCcquskbpIQ8Kli1A4ecoyTF26kqDRHlqPh74t5JuBSZWYsg1Pn7qhM9EgL3V0UM92VxlSrci191a4SRFGihK4I+rckk/nFqCpDgkX+eEukVjKcrB2by134N24ogYqs6Pv2kc56CAs3m/XTXdD6kiC32RahzDyPf/G6nyDyDKvMl6joi+Y/Cy6GC3L4eueb3VH+jQZzNj4sNQoELEdl+szpjHJqyfA/9q3KN4anvvjXTZL1aVfieA92PFMGDKXEpEH/nCzwFuwgNt6DCy+25gYoo21D5ta77vLdClAIx5GBeLTaYVZlapeaULjacAq/KUXAh7sGVJbQsWY01suHzXiSQ1o8SZxacR4nvoI5ngpkKCrnhf3fVaSUYm3CBZQ+f/XXkDdMtrPLLeOeScrPD7USt8balswo/iAK5MIkyq6q8BMR4+l9bBO3Xxp2M5HSa0yvIA9SUn/zlyfE5PWvXjQP/zh0AV0oe349lfkaHIOIIPPFSh1Y8dN+NKo5j5gvnwdF4kp6jUOlike7asZSy6OWboKKVlweM8UC3La86FiVyNBZVo8nG2k/g18M6ZH14DB6UCRsFeqgT1e0u9wVfkr0KUHVcSJJIH1dHNk9q16pfHD3LIaTXgyweIve35/Q5XDM8CD70Ou+boN9g5D1Lj93HUcbYxzhI0EwJb0t9fJ0nAwC64Wcst18l1otPg0yI5oWeAV1jOcoVUC2EeP7NDAKoZDHmU2DNcLcKKHtpSo3Px67gdNGmqvsl00OfY28kRF2kbXFxIf9lrs45eu04B79ZyvnX5xnm7kd0hN4zQdxVaNJvzabWyuaRBCNxcbOaYpUzsNgCW2dC7+MKJUeVrrvYOP3WcPPjNeBEz+glwyTsn4LwY2TlAv/LZ2s9wLb57TVDIL7qnac3bLNeHiGsfyuwOkVYtas5jZgY8LXOqLm+vUpBXKwBUllWycb0q2mtKx98aMLHaQoZqR8CrNQSYsMTyyIif60uGJYqsuaH2ATvPEGyvgiCUNRDLD2PJ5VWmZChZj2p5CXAbTPF1irDNtAQhlUaL3mFtpN7u8LgrQOroXxOVFLqLjNritvi3RfABhCeaniYLJp8EXfYbY2Jb4p6Q/TE1yoS+iO97vtTp0rczul8s6a/I7oOWg79j6qk9q8zIjD2PCXV0nFlW1pbWWWD1RHP5N+C86TIkZutThLTF2x/RmAXlyjRE/+jf0Kj/MCrKUwquShYi8+trPEiUa0LBS1kD0yPi5dalo+SC7ZMJeSDp9HS/2vOhnVqf0jPrGSTf2mkFFA8gzpBdIZ7ahMQAubKQMV7ec8Ov5YTEMG7Ww0RtQDvHcTU2RlrU16zvFNzrj4iMsFK/5ikOMbce3ipHTosSziPpirR4FQXrBOHoynxOIccUtQb3/EoNIeIoXSFX+N7KvDGpyyUwytnmYVwzoFCGCfoHpRzKw5bwcAg5IxsrV+yMx1FIANIH6A2b7N6rt78PMnvR7mMP5HMwQUAEDgvQQnids8bU6cm5/6ZbpvqqMZhU2yvTEK6CZYsbZznxdwxJikBEYx6h2ypkGqw/6tTELRGrocRogf0rA815QeM4vQ1ErlN3FKQZYOHemn50PXoflDkHMQXjz8Uz4iWYjDaB8lYOu0z7Jy21+/JTp+jEosnShULdjsivgu8uTo0GVOD+KsJn+LOEBKmacig2XUy9Olcf3mi9TPfoyVTLFsFn7MvuN9LxEvUPKQWXsBNxsw7mvTvk7YimPgVeJiXlwIjS2BwN9d5WCAp40zwlPWy1kZiqn+FuSkt/z/FjGhjtvcMTTcmD1DYCOtJj0Bs+AJ8yJMvxx2A8b8n/5LE7igAVEwc6Q6moO3VCySd0A4lgH8s6u0otM+uoTg3eWiBoNezzfPmIoHvUmOOshyzAgrb3nSnM+6Txofi1arrc2UzXxTf1L8m1cdzKNvEaC15BtNvqaH3EdY1zOt+Rrlu9WyvKdX7N6mf+pxsV4pgAV1oa1IE9OTOqYl9EGWG/x44rA5e3C0RNRHirpWOjn23+N1T3fy60I5s9YSxSaa9uKJtkNh2ppxFPZojgy1lGhdX0ikySqVqPYpgD0F5xbcbqPappvduiDJ4jQ8mAqE2pTUgkvSASQ3DkRkBSiFnf9XBvhJcPNxSS/B58ghGFDPTcTea0FZ/Q4KNBMgL5TcGfglkaMz0uR9VAJQ65mjhfukMFoRdppvlta8I2jNXcU86NpLZPkyYG2P/SvFCecQn3owF1EOliV49KRM7FcOSeMAO7aFuurtjYf9HqxEoszyPDrgo4Nupo+6mGb+nSyltyFkLIu2HITnluxeLhcFL/fffOcLr1ZC/9i2VMRJdOfZaN/E0AwLXwjfhDpwy46oZfXVQa6fSOdAvw0y/IjklNqDWyn+9fKQ3mMbHawzL70HJrdm0PxeuX8Lg9yFsMLAV+icuJFr+d98MrqRS65UMWrATk1npbx/1WtI2B20+VLgyAAXmyI7WYEhYblS8F7OwgMe/YHoMCsCPJXQqpMZzuHHTY6M+jv3dUwZMyU5dWtQ2XCcO9Dd+onZumOmi7zzLlF1xJWChrQNy+b7no38ogvo1fhOVipIE7uHBlaODHAqAEJQzVZCxC+RMGE2M2vHRPndhTr5n7ww2G2wnT1i0ty4u0q/rcmrZyB1fkAk3mttATjQN4c9zu6bYimEM/4dIt1OQDsXZOV9ipzMs0+CWBDPc4YNmq1+4r7RbiFl4jt+w2SdYLkXYIVSS1aAdN7hl5c3ZGQStY+eEa6xu5Hr36EFXt0Y/rkI+O9vXV3Lk6WnR5jpVbTkOrXkiTku0M5Za/l9rrOo+JxK9g+MfncFmFAeEEUQ3R2WJUeHI+rOYbHBMdCrr8iSs6seih4rMKOd17RngGtAREEghKhEhwgCx4K1CvQ11STvgPcus0Ugf0mHChX/8Kd+TIQpTxJDM3iKf4hjT6pamkAuqEIJyvi7vUjvD1+ZjcbddnrDho8sg6SMZtxKUuTb6iTUuG4AZEgVVPpJ0t3k4BCjScjawWjoZK/P8SnFfQi0ceRm5GDMIFvBmncbCSHHnhwUEN+o2R/qrlMIniv3lXRv0jayrWziemZWDebzQJzTT/ZpHbe7DhU5j8n186ZL+p0ehuBQXTpcWXnqLIfUsVbsv0WYIzuTF2Tlr+IrIKL6RYAoePBXwd3Mts14XDML/HckwMlI2qvNwOsUU9YKD89GFMtgNr8gqGidHIdsgYwYrfCvCiIQ1C0jcf5iR89WxcjqSrqpPSreoLf9uOzwOzUHoJcr9vHQfwGEvwshZ7rM2WESYn/DXY4P+tzGFV9uPDIWE/eK0F/TW0tY/B4oeMCD03NIQ3DFIKhfkpX2K8KCO+I/lX1LoppTNzQmMkmnH9VZDd3JZuyPnOUr8QcugjXY7TX7uFlNudHBXUJjczbqVaVGVjzKAy6GqchpNz4l/pJT99COb/ZnbuMIq75l5woUlp799YIopjMA7H/Jfd3ZPd9420vE0LUheLv8g+uxS9sb28UPYDVJTIuQXA7Y4Bav8n4XHYLo9q2xhvye/JYFHLqTZFJ+9eyFiU9q+GD5MYNvhtnBaslmXTZwPfdFXRR3rcC0vcjj9f40/t8QxF1lTCfXNPBzETeC5+XLSPBWiStXcL3kvlgArXbF/M54E+me8MLhf94Z74LzR5cFpUQ6+/XECTlOBGXAi3ZsFvIvz+aBo04OR/FJTzDkGT3IX8LOdB47GlsVN4dXJ9owuKg/IGw5vJoERdLnmmllq5Pp+5EZNAeU5w4DS3Hl+WFVfZDVEiqUnb71By1KCG4WRu5Gk60EmNNcgOWfHcO/nguzkqxa8LtpGk1PTEHGNnrYfU3+iwY1q/iqmboyGHj1w3+LAWXDt+3bvIE2TU5POIIR83k6KrKBNtKlmzA4w7f2eWM8aknc37SqgaDjZwXpuSGdUh/qpr3Sqx8m8spctqUbFPA9AANUmFya8dvTwXgqp920jOMq0fkhlIFzn30OU9bUDi279vUiZ1snn708xjMO97/luuA3qjysNjKIdUwLzfxfHHrIpTz2hfi2n1n0vFnyX6UXBCNhBE9WykL9vZU3xj6mmLYHNtX7wTWW6FIgS6v2oViMFFhkHkYtk6i/Kh+fI5cEs2CyYnoiDlw/Ibjs4S3k7sHvIgePdvv5Sbu7VL4hqwa7zosY8trfA+bs+3m9N0CNRXDbqnx8nudjYjNnnLeT0ipgJlOTinST0t7ftcUc+n9SIRkbSzjDO24NrJ/nrE8ojBqCNog/TPOUy2lsePdJVikval/K9mr6d3bbYLGWMdQCt0CPw5VSeGya4apKznkMauEVftHA8xTdql7nlK1jukeWm3YQrS2aYNyYj3wecfUhEMY+6yYppWD/jwjNvcIEUaUF5wgqwnSzYBeXN3dykhBJIJ75eM25sTOvirA1RZ0HFkM28WzkkC071Kb5gyCye+rIhAcw+a4BugtDEtx01AuSNe2sUzaEjGF9wNC+URzJt93bFq8cEJHJmo6iat/0ns9VJJwkR3YPB1yHugR0gXhRdzJh1v7aFkk7+v3JPwIvxwR28KCOLXJnZ9WaoNZYCtTbuwdL/iGVVB3/CVnhFO/3UOXDRbAUKRyJKpvfr3EO7bBm7HQx2h8SstRC+/ARmKfjtwtPuTTOPJ6w1NjF9cjb89LjuUyENI1KPn4D39x1POdyacYEbA+9vQcAL8w4W/83sqBfQKMCS98Wxz39O7V440CAKuHMxtgkjoeaGQ67lsIeVMz567eN0HMEZw4T0hB5R3XLx8NCEczMURm8hfLlQG1tHXLf8E6zkufUee2V7LySS59OHtnmn2aV/nwCEpzcGat5Y38CfR2utuRZadSPfN3CRMg3b9Mt8Nygg8/Vj3S2Zoi9zLZMOY5Osj+CFiyvh13DM4mLU/eJgxYF0Hafj5fijN95nuKNnPV+qSvxAqXgVfirAgT+CLkf6PG+74BH/JpiYGu4Z7pv5/9agwOqKWefzbX1AKXYeHvHd+jUflNhivDLOUBD8rRQRnA5yXsqO4XpbtE/a6p3bA++gXh+ZF9r03Q9zMnDp0QcNiLQj6aSJC4bVOZqWo4TWq9pLK72LNv9YUY8XGlw5AyHUVMFOK376W0NW5HCz1JuhjxQtWDesjGosElmVgeYMbvA9b8WNMZYX+mGuRFuL5WXKVlOIZ6mXGVVNl17fQ8QwmLB4lbeLRtK/I7ABD5UQTdlEySXKtKy05eU2l5fM4Ogq+VpPOYK2dqVJy21vnoDO0/kHzEYU3xVmxgO2pVEZW/Et39NJZGXSNXt7dG3Ep0UVM/WUdeXuG8XkVJhZCV+QCznJ3fjSFhTICW19u9Wa24t3WziFjS3LgUZwzHcWm9EfbdZSBUtqMnsSLGP6S3ris7BL0MRvyVwkCMtiW+jvpt3hHhVcX5LWxHeqph/DKeqrFMso6MYDsu+igKhXRTbaGsaZSiCg2Wq0YTUCNhkx433nMpNj1aJScbwaNoYd2yF/NZyGXK/r4XOK9o04YFRljd44wj2fHMUdFkcAMb8+DoVyCkQY2J1wFJMsZ8jpyG0KH0/vcL9oHzciMIxRoR60JHW6FfYQjrYfNnyjafk68RKiok6OLHbkmErXDZmLTyiK4+cA4ZcWEMVBZ3fVX743lDxpHNaawPhTz/fihAKVBy/sVJx2YgfSOejV7ku7VRGoucKlkP2aRA/+m1LcOxTR5pBnNWbc++BX6CK8psLVn3XMssTioGOaxrJS7pW9jzDONOxUf0O6zT7MGA4Lj2YmWuMfCe58D/0LNC6GiQpSfeV061M4xXML6zR4Z0cZAdOzZjBmeCFbkN0SKGDKnLI++Sn/KtOJGSSJwnM2fQ3Bxv7BglGTlmVbghKSwU6AQsnZNb6jpLVSam39dga82QHzSiSi29lXNmFmSTOsSR+vSSk9C8EnYIs2DSqPS0UCzR/YmZw+CYOUT1lAbQgxcYPKUBfOEpHhy0IGBIPXzgEtjlYeINatNhD4Li5kT2LkAiTvfgmYxAM3vLU6HyLXI83+rPVEiwL2AOpQ81iX/+9Sh7SXPQYvXjqtVfDJgyJePIiaTbT7ShrQKDWFBL0t6JoKzb2Qg58pxSx6XUWPYAuNQPgemVCfT4KjvXehWS/12DBviutA0mR3iahqkwxcmHbFG66IZuy/r7RfhBLkLyGPWMg0xtDK4T5epxocYwsAds0XvUbMoNmVs1lwNZmyzHtJFBiDdmTkJfbWPHAJZqxAdY4ZjQjH5nRoNtrfaCkZ56+E0jjR2WJfxAuBdD6I7dt9eifY57TyODmLFLfBGTlUfogvo/UutjDhJzZtyN+wuBeDETNvtBE8tJEmAPLzfOfX9G1XbyTuEcxqx+mVn2mG9iyU97AlNRt46E4rEoc0Bgz5hSLtLFDrN4Jls3YHbRJPy29D7o+2C8+dErCw4RMVNETVAHtxJ1DTGeEWlcQKeUgZOfpv5XlAFkG52p9gmOFIefn3tio2D/CwBr4WatW761jbZTcQAFzczdkhzlAdLoeboKdBcKlnh/OtSpfCwiRXQnK3GFyhShaWvYT9IQ62M6zOUI/K9x2vXj7xbs5b9F2w9bWvP9eFFK+YPD3cpVAXc9qQNfTZquhCemphjDe9I3uM3RjTc/aPOF6+QkLr8qBdZ5yzr51XxHUXxl8M6PHP2XTvbxUfA59APVS0GE5TXnkakzQdSsd5ji48RldLThWdORbOnd/WSh632Dfoe8/27IZedB4Wx77hhucNwoLiWKT1peRbhzZ2zF1BMuj51UTr/a8puSHLAc3je/CMh1de+mFq9mqVRsFCRNLIuTfjSDBnM+1VBIE5iDoeTO4chkSSlHxcCNPzfvfi/ja7ewqxR7EZlbMOr9zu8kN2ik+26Yl4LmqkndezyxJ6p0LXt0sUm831RCCEn4ZOObAIkwZCv7lp4iUmNlfBFQGdnOWnzqNtqlvnYjvy/DHWX6nMnTeUyxFXfGPgYt+oHa+AwIcmo3/Uuyy3KYeo9UeKCt8H31VzyMKaUshbPJSMp80Sn+e5PsPaxklcWhXa8P1Vg3f7GooTF4jar++K3OJiVg8RLdu8O0jdDUimL3fcZYaWjRYUOMFbR1f4XkzJGuIse/udlCf+tux+vWy2Q7Zf5W+7jWWeeHQqdvUyuIwHtp7sIRzxVWU4+yaTK3i6uP6DNgz5DU6u8gpbx0T+NCE9pIVoBZGEhUp9rtg1i2TI9svCpgQt7BtjMHZG8Sg4rQft5jx4eclbdUB51FKhcxuM44BENWlJ1Hka2lgMEIY8Y2LFW5s+1AFzH/9JKryKaLIujs7XR0S9Km6+6qLOzD/z0KcYz8kOer9m/j+9zO3ytsgcdstxAfwD3hGmo9l4Y2VXhZHOFAOflcdJGAhyPrgRo05mU77kFU8UdDGXIVD001AWuvTBTaGPnsoZo70dgv0mUSSt7c9V57WyU48DwXY6mWerZ3jv4+1INdVcERrVxbXDSaqNg5Bic+ULZDbGKU/yvh3f2thOdjQcH+q6ojaUglFNCiUy/fd7MEHzu15XUfjEpGy6Vxuhy2oTJK5fUGVx1GxI9nk8lCzha7OUprJRNWaxyq2UgtIkskwUn79fIEe0MooUDNdkUZclgGuqJyIRNEP9VE9yFOIAZkVePgH27MMvzKHPxoChii1xqFLpRXjdViRPPgtXz1r4ZVCCk4hBHcaNCfqF585e4F5Dl79Fg3Qv8V17Wi1zxlp+K1SyW2BUHaT4h0kbl9pm11ZtpoCJJ+XN6sWibvDStNiTWTJfWdT+T/rLo7N05n8dKqhO0K6rM43ot11s0T+8PRHFiZdGWyXUZ1vZXdt8PZyAHMXTmLiblpSItlreBlD0GBw91yhA8Q0TqpmIG39dewVSzOrp4/s8RZN/Tu3K7gOweEuoFjC7Sapax3XgzAWoiYs8t5N+zmS5Rgo38Uk/dojpLC2v664kgziK+A6cfXyqwXmjsFpUgJn3G9Png1LgCn0nTY83Ou8Fe1mt0XaXqyCFnZiKrMxo7FMFCzDavQcFiNWDV8fhENaV0oPU1efRgK0YjYfGnEU9nZj1TLyXjtcPKnVIdnTUxTE8E3u/kTk2C+Jym4qKyFQpWrF4E7vca55PFy33s9W3iIeMZFo6i6cZIpGjT9UWCZv6KzusZI70EYtYG5sXx6lqJpv17EyAjiRq3Qhb+GnV/sVVC3PYqm0E5nYr+P2xB/QCIOu/OvpUUFGtClYpiNEcR+h6FLcrxkxsVH2Hw0nPfHRx0LND9Yg/TdHXTpxIerHAsSDTwXhq5k17AASL9VktWZG48tovkJc3q7UNp+wRk2oANQViSgFUMayWTn56theXZ4BAGZpdrD2nrtbO2y1/D9RIRBv7IVPT5Y79armPEiXfZKsOa79Gfm5lqjw3irQ3JDBOJet00QXP6lrqm250JI1uCpft46R7LOxDXW6uccOnCTtJJgCNMOqwE3V1o7KVSHWn8emx8BrOarJNdaEdQybjXYXDx3Fyl8TUvkYbDaKaP05T3FS6fIKOa6oZfimXxrl18WZNciOEkywqbpu1cZd8yE8safF56gAXU+xqfMpY6Sp6Wbiqg+pGOKtDMKImfHHIey6/pY3O/AwvP4HS8V34FW+l+TVXIQVGBzMWw0wS02lQiBMnEHC6IxIyYBr8elG4yBwVi4u6eeBIzJUCeZkbrNF3Nq6GLpXf0mJdvcQmgWBVJNsL+q9EzyYE3+NiVno8L78eol/a/JKdv7Q6lefGqf73WPpS2VHvBvbsYt/1duckBihcW+5sKCc7UzNMwyOA6/25kYpRNXcJu8QwH6hJrd1yr/aCLaL8aLw0Tz9dBrxjhYu9x2GRFz7dNAyszY6PnD21BIsAF8Mx6iBheWijz1mgWSpI2+dahNuvXNJIkYgXkLo4gIyk1uM7kWeJCp90s4bMDPUXFCb1o6K2cb5akW0/QMnNh8Cs2LjxJIt53xZiRgE/wNHnTX0Cdm0mwZa64GCpVrKuS+hpvFRIHBKav5eCIGjCxHt/XcpdvOjNu9zhBESGUdURaCweGd4XM5mpqAqyEUB/cogtg7EAzMLzP4TRvkv2dFLqRR+P6XONDqrt09gvP9BfACzr3BEQt0qeRXoIIoEbKu43V3xfpb0=
`pragma protect end_data_block
`pragma protect digest_block
18195551a98d0d3e61f24875f6f80c495a4743f1c94b51f6ae052ed4a4a30595
`pragma protect end_digest_block
`pragma protect end_protected
