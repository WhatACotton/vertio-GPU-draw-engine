`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
ZVpYWct98t3bd+mbSSaSVtpLkVAVico+0KekI3mDzpkZpppWNjSht6cKKj4/DHhzzgKqNSx2dMt+dkU8OWJADoZCuTZR48gYgtZqxLDkHBWkjVnVj2raLQh01U+YVeu+X3/Ct4KRgJtXjMGhN6Z7KhganPnBt2P43pK/4d4I7h7oU4jUF1emTME6tMofbafxiAYRkSuRSM4hvag1JjWq9KwzLCE1KEnpH3RKCXNzvRmNbu7vvFfbCRvlWp5m1/ySt/OgXVXDhJGd1i5XdOA1BLy+YHIHrroPzqlJib8q08jgjjaaSB06EEOiwDWbf7flamdMUiaF85tD72S2wUWVx2kQlzFgY8L2pt2a3cr704IEC6k/SRohEJp0vuAM8UgF8lKNyIujibzPo6ZMv/OtaqLmQRv00JBKQxkFK15ZLFhBlTIBafRR9qdkqiRE9w4DxBdeZ6pEuE+U7scyPctN2ORUO6s4pEwRwtbPpIwDAN4jQ/a1n4w/+GGtFSS9cJsYlNw6fu8gm4IYijBzlYaeAEho0cld02LQuK7ifC0mNPjBFXvO3Vfw8VfJlqtmG4gHi60mSd7Hk1SmNK/p0/DPx8fSU5EtMI8UoSgWbiQzGhYxTEsZfylUUfaxkEXhyzWU7Svo7/tVB9d3cpeg1CuN71LJhH0CEv2DgDvpBB9XZVCuTAbOpjYIoLZVYwMkCvTQP9rf7Qn74Sm+e38mBTgxJ/TmnBQUGXWabyJWyK1oXy6E34tcj8gk9/HLsehCzi3uo26cOP654ZqczkN0wE7k3z9rhuhItv5/FjNuYvThH/P8SzpLMKJh71N6+9UKc1Xxt+FpVfGcblvaPC7TYwsOnW3dteAyZND6B9FfGYd4HshqJ89gahvYWthaQwneYV52+84lFuAMwU3CPw0WkPEkAuOfRTBTiUinze1jHbyyz/SiuLRRJcj+5u7mfM+DfEeZ1PvFFviyFqCP06u1TeaNRjr5MRiZB5A0zgYgfqmqKgwaij+3pgEf4G66vlkHxLIjMwdmWjDjUVI67IIuMpYKqFF6ce3N0JX0Gmmsowskjx+svgH8yu3MuSFkrvBXhOuhqCIlOA9vhF+GPLHMK11EosTsBNxnPTjDTwznqjND4B1m2Enk6+34EqnwwSDDeS5a99/UkVWPjKldC8Kw50ODRPfqh6CeJvJi9R+PLgo1xBMJtVusNpNK/MxCwou8w2llay2dbhoFpFSjl7i2zrF1T8IKL6WrU+mEhBN9JXIvrxSz0FtcoTE4FtY1rh1A0bvtbBfOaw0lov1G/Uy4sPNMFHVC0npeoSlO+SuK6IwJvWRA7hNAZFNI07rTnNM44FZTfQ7I+2ojMhYdcRnFl5V4ubUXD9zD6qHHivmeyHuB7LCBx3YCngG8KZfpmEIXP4g5AQ+zwWWF6egTDZlD9pGL2whUToccGgXQkX8tkZI2ZtkjJocApLJziIHUhp3SKqGigxFyWX+BN6Eb49Oaep7mvuYH49qm4Oceq2Qcu/suVMV09fhALctDYkSd2csYVWquVj5kIGt/bVGVVZROFEKvzh2LYdyDFCGjjpo0OJIBPIiyGwqZfhg0HlE2dkIy5+/f1aSjfEm4CxhCRc4dykxAVkxKY7/onCFp2D3Qau6k9CboTaRA/kBSdrsdKlQU/fEzuzfvnrdv4Nmi1+8RywkSYc1DFXjrrnvZk9sXzMshVOfJqr+DmGAkzIGE7xwKvPFBghhKdF7ksoOZDjie7SdgPDD1r3ZvEDXzYAGU5O54N3B759PrDKL8Fm0mAt4WVgj05Prbl2JGRtvP2GAsmJE28T0f4z3ysiEPdi1zFThKFgFMJKiHFkQkJ2pyX6FRSmtgIMo/bcZr1aj7HN/poNsr0FEHFM9t49k3F3Gv/ORK5SlQHe3g/5I2odAGqs5x/RR2xNU2qq1V4PC1Hm/OAThNU4TAIDCx4kvaVV4kolKUr9kP0wQQ7Y3kln/y5lGq4o2bjQQbQu6sDp5W+L/pgjpl5l+i47kPWM4yFOGlDckZh/xEy3ejIaKytRwC8HAH/XAz/BzAZ1Zyk0tid6pmpw1JZFp+iB0Pup5yXwRDhZc7nM11vqyTviqBxOvfWsi0pbuMS6QC+ln7RWcVDBBPimFhUl4iwR+3lh4MMcr3GCV1YTs+fwYGW+otcRW9FN+T/CDrHdn9RLB4FyPVGzFXqogOhZYgWubXoHwm7MbSwRjyhGJe/bhrC0VCfopM6dg7fhF/bZkq65jJ7XBpac6yH6SjtnV95FjKQeMeBOuhIKPGx7p2B8TFni3NU/fqds+ZAhdb57TeoyQbgy+ZTw6YbWi5XOL5S6pYzIWgJ+1Zvy12riYcM4/OOT5t8NGQzpIWMnae2jPcG38WYk953HTrmJXX0Nu5oYFk0dG273qK2F635JCY3/r3192VVG61eNKcPIeZWv4hzzs0bUXWI5GRZ8pzXcEBvuXkEBF37+wWs3Il7jBff/AWOFkd4y43DkaFcFkLvgRDaolgnMG0FD1CVQy8rShtmiAwa5Joefe1O0wGLgNgDsrrMF7rHalfVhipBqKBDn81mzn7bmFQHcZsr+BNbMzAoh1ViBsTAfgkUGCpnSU+fkwtEjygFF0nN1qL5iYc9OXuQWhm+nA09RNVCd/+ZCX0XnV0Zv9cbotClzM3nZZUNnwb2cT99MQLhNNDu1yV4ER9egy2JEwHEwKaQHabiHC+gxgj9Fk/Fpg0QwlAWFabaqc51XHVX68qYmorZN25NgHe1Pk/vYQ7s2owTacetfmM9koGMW9OQtf7QrCEBoIdfNy+A+VBrmKXbmECk1uZKaBJH+SRi/P9Tnwy1CiW9B+gwudJwnMD9WIdmDM8L1zVXzSh6ZAkpQVOcpuyTqN4UroMz9p1uoYsXNWS1itR6HlnCBA7Q9R+pEWZdxJK7W4k9Kex/BSOT6tbP6JOfoMhYm667g72v1qsWKdIzbdA42In+kRoaEarYUUQbpcjQg+xrGkK9mRFzLk4hhBKdpIdkvNjRnN4yoaWqgW9wUqku4CTVA1tN1dMdJ65l3mcoemkFs/8aCEsRJT9oHCON7Ms7m9cMKdmr+LS09Y9fkJo15FBuA0IKpu+wfxNr9rxMdac8jp/8uKw+9psqhZmH8h6eEpdvvCkHAUDs9O7ZaYbQAxxqOGuQmfJPuPX5iEfuNK/p6rdfqIFDt3SkCn0xRqlTf8sQynmm8EKfOp6f9n+QbLxFa/f52Xw4leYJdH2Tuo6TUjiiWJyN/Q56mLyJgc5BtlEzEZPGBqDqUJJXOak8z9L+Fo4rrFNtC53lJhCbbgm8VmI89tJix+bjdW9yU+nQeWrN5merusdlvPG/R+Qo21rBk+qvdhSntC2X4lqnmEgLW7mFk15z7ZRjwXa15JUzummFdkaIJbvgYxqcIbBTrUkc3SDbA5N1anRw486r6FV986/uTst9r8sclOMHU8w1QlBeyq4iOw37W30gxcoV6KyAGTxALkZ9iTK9rA/QlEBK4856OLBEE9odr6oesCRizGC+ujNPmHnJz4FC6PX4Gu43LTLPytukeCaeTJyCZrEedmhlJuE/P+NNQvDgOKOEqrPd4h/wqfGYkh21teTtdP8hbW5SwEtIW3pe8sc+e4hOsBoQmtHOGElEKM0wm6mqCXYRcCWczNlgjhw6cr7sPCQIzUZy5vQp6Aj6L59v+EjDmEs2y44FRQvnsqMtmRs6WmPDvXP21cHLlGIFhfIO7DUA9TYaGXkaS7IAqlTl4+SUpw2mb2m4act4gYdGBfhVyBxOuPnlt4rBp+WOhSiM4cYzdmOBOmh/kb1wYpngRrDQUXXUYcVABkYyaGKiQ19mJrxwgf4WDY3hWxXfpFehXASrbWrnsbllzOGrEMt2hz0o8/T3kj4MDP1jxU5WakmzsxJFBIySQvYKwTv/sdTSzI/hxAVZ4M6aEJtvEGWqGHgDexEeDJDCPlkv8v+VpyxVe4yvWqmQcXcrA4XXUV4N8s0ahPQx0FOmRp6R9ZBO+fPr7CUyoQTS/45jr7ZiGHv4CpCW3rDr7zSdgEBpRID25QS83gRtf/W/b9LOmxDqhd/CG5DtCCFlA4l/+5hlapy61Oz92cuiAVbQj8ZpEKCayQRaD1NubDQJUBZP5jAHW7H195E6ntq08jm5XjlTz16fZJjC0SXgqjxdxFgRtdPryyV9xftayORHbRUK947nAdwszkVW4oMJOQl+ao3Mq5Ty3vbtnfUE+HT3WE5RoWrplLaRIxpT8hM0uhs2MiKDAuZSxZ/vHfLVhQor5vZglXbM8LT3AceWmmPM3jwmPm64MqKIToY2dG5NDMOBpIx4+eIUCFtDbYKK1GkyMIM+Cv6sfxzibc8e0pd3q9J4VgkUG7NMoAY49N9lL/qTKeXqsXnjHknCh2T2Dfn5z09R/RtVNnFVerkLRV9QiNBX39kixq7WM/nXZ0COUTwFJMuQg7BgY41l2LniYrBmYqdqOQGznekXLzh/bCHQiuPk5RpsWQFqwLEPUd3+k1/ECa6PxZ0/0aci9r9ZqaDgWpTm87Qskym+ENALsbDyhO1M66qc/v+KFuMb8fo6D6mL2H1ksxQDTsg1ScMr7g2eT3ssK+HQvxKZQM6AFTrMtBrhu34r4h7USvyCiKDWkrPcLcQZqit2ZnCk1QduVoPD5HQBAuhVvB8v8eh+Z2OJA/zeVrnd+B2Qm6iOCN4GJJcPwVFYOJKRYRpY7GdWKIgPqfTwBwIEVcm9H39P4gbYUlyCoZoqK4p0j4ygnN5hJnTjPWyMzR9InVZT8Je+cF2MlAA4IlStBEw9sSEYpKh1Lyyj1rC9THjwbTsRueTsUbXjh9sR40csxMwooVQfNK6BPl/NGqEbq/Y2wMD0+6/9t1dvMSYxT8atOcc2aJxRt9JGsFLR7T2qZOjwqgM2FphSOu7kbkKB9bB4fvvflagiT6YR9ibW5tzOaUlgcHJ8oBlUlYeozAlLFV4pG41MOYjzPu1FPBcWX7uVT0pZ0kBgBl2U8ppQo4swWcSABDwxF9yhpy2Uel9kFwaED9i2IMohoLWiO1cDS78ifVCd8n9l4CulWrkOYtft5DKzq1+FitM5lOGdoA+E4rjHVuSmqRxglbrRXeopZG2YVyddB+5MiCsIAxoUcvx4r4UZBMRcR4k8WyTAWgwB8FVT0T0wDwm07wRH/l367wzio/qD0QWc3nkkd4Kluf7ae8eStX2dypRXx+Z310u+maDrZwTTp/gi64SG9ymsjx5Dh0WWgnwbgY548LjNTAqg/MNgXsH8OKMYknk7ildeg5azlbSSWyLNZLCOBzF663eVGf2sIN7Gnc7ZG7LlV3MngEGqxKKcJj/zNr0MwrLH1m8+Z/pdXwA/D4X9ea3ehziSRE3xbJGTAbvuNfhUBfZAQJDEuzVaSvaZK9dw5VwhnMs6wAEicae+jQxrP2r7k5gtmZC1qkfa5OO5DLMnhLzOWMPs5seZcLmgPigMmTY3PX1NADJU5TU+XahJBzBcrlqf44y0gLzpPSNVBDUczGl4GJWUQfcJndoKp04MrCzfzidbfREUGdBp9swxKuSfKwRlH+0s+CTMVL/cDy5pqWYpYMcPIrvqRguFseFwoXwo5QlSR19ISZeGyBVGuAL1l7Ta5TuEhGKr35FYRqNJnJf4QT4Q0emVKofssStH3tuFqCo8DHWDCOFv7rO8hiaVHBIgWNM4TVXuVzAbuM8vvOe21VCWZNmZtNPOD66beqz0kUNitN2+pLLN3DU7jpeSN7uElHeArSJ+BAr40bxOm9PKjQcBQCAu8e9WIgJCQEQrYQ27whlRUQZUl+4O/4u3I1YoylYqVEA1wOWiW6sVzGDLFlwOrjuoJetvXY7sehygJC2QiWTF12+KH0nCeyKFpWD0DuTdLlXqEA0jIIeIJyZqLuk+pnzEI01F0zOtSe90twrP1WCg9Yyeypy8+G1flHntmNVK89BWaU0g3zqr37f6CcqHW/ocyhKm3dGKfY5GxlD8WgCvEmHG+vUiCQ4Q4FY6+tOySxI5cxNsk4r7U68YeNdkMMm6926gqzqvcP66ftwF4baD3KCqXygMuGfcGjdmtmhWczYZNS/VafnIyksekhXbYoXvOziw3eGSaFQdm41v2Sq+S4ODDSquFQJSwl7qTfw2ktAWsqvB+iuG1z0MklTHkdYWut6vqcs3wcPk9+T47VzbgoK9d5J/a7Z86UbK1V/fblkdyJnsjMfeprP+vMtUDEJBKmmHW4MPpEKxuClMCMXrxQ6/asgVfOQJ/YFWxUFRm6aEOf+k5l6Ep+tgFel1o6PhLS+lEGR/OGMNAzvXltGMLfKRADpNoXPbr4J5oJu3JaZvxZJ/CiWP7+7ZSTcezbAyhAyS+jfO21+3bacova1dMAAtr8b2qu/ARw5CASOeQrT8BSZDgcnVik3zZqi4jJiedalYEhObuKea57PUXqnieZV2lvEjabGyGMAK47dTkMGCu8fzmS7Bd9klV9QXtcxXW0pji+ASGvcKBpCHRIi+Mm+1MZkBMDtBq8KlSTfbq5myNM9bhRtXhxlEh+pTuty/iBJvbdPAViCmMVtQxAw5eyixEpdcUFK7Wjdp71l99OZ1+RqPTMfoTl5ypIGVqwjH/wVxu+VNwJafXEW3r2krARi0mkayWz7ynKCcGDrP8DQDXRyv89osQjxaktx3qe0B6VDY2XIQoG1rCgvNNlZxQP9Kbjq4yFHf3Ntr+P7YN6fRul5d9nEu62LeTeuiP5dEFPDz8WHTUY89UcWo/68wuqKkNn3mzo+eQz9GH2s46w0vEPC4NkIMC5pIpaTKWJ/+Ffb+is9v89cSmcyA9G7B/P4j8FXxTDBuui7HjvEZ6PZ1VSHFL3lJ2WlKySN4Ub60liK6i/eyQ7H0OE3zfDwYBJsqIdwu2+HbCZH+uTKAEURQKdBR2kWIJfjkPvTfUsJ9nsXfoMxdU3/fsYbWKXTPJRpSS/V6T/yP0QH9VQOgsGw6IgbrZld22DDZH1LsU1VnvflxCSLd3M/KWU04D4Ht0ufOfexaoZIxmtbYiTWhtRtOYKDFe2WCUwZM+0MqOffc4I2F4I31g7yynt5tVLnlh4CQtmq60q0fsxujszRAjTgcYlGludWXioPSvhEArtWo4fT36EyaMcEUNVx7fDgxWXxvq17gba5kZmimYbC3xxGrNx1OXk1huAc8KW81a3Wlic5QNObirTjqEvSDjnhrwpSGQQhPJnj3Azt1chTTHhr8lSTzNvgefRlQrUuVJAvlBGJdN2dlyYK7u+7N5lHV75IltMT8ZVeDawG7W677VAyyi0/3lX2G3wLCd+n9Qfis/OJyfci//S0yQIaZiPwW7diNUDf+MK1LX3E31Cu48McEjUNBTv+/HKXNYe9FAvz1B8EDh0M4/u7z+Ax4ad6IsQUeVb3MatmnUfoXmthwVTtsUnouFPpIquYHX7Grq/sbJhW12auVedUavrjTpt2YLb+wdYLwaHd6UgSIwL4bM9TSN88WhCyLcsXW4V+PA6BcHN0AYaEM/0n9c8WTJLUa9l5SifE7j80m0TE9bNtnz1fUxQTjSss9R3MrKFGqoscL2yR6np2KP9Pc6lNpGkFLurvZf2js457Hr6nFZTMk0lKAkbbZFfg/dmWBNOuxXEBkb/Ur2kyYXnruQgGpjFajC728/s49cFmfLHYXW06oKTsvLz1Oym+LGzhfCPeWPenn5oMIBErYwJXQ8lALmPO/Ivhv3YciJvPzfRj2dIsp68mK9cDQS+WkZkodKgPQVJ0AQpWGTNflnmifBHrX3bLkI5s6yanzt34N+TWwH29ScOE/gSO/CS0gvqfxOu7JiokwPZy8+pDiRgzTDagMkzqkFJIA3BmgBKKTcyg/dkYD1r51p3o7W97XdNdqMxs67bNq0Ypnwso1mP6j5wpTABUTuL0ssdxjvDQiH7lVPAqiBx3k5rdqZOG9+VMgF5/MbN81m2ldzbXlN5RZbek6FeJYBw80dAPEUyOeYsmicmFZ+N5Q4rDuD6r+sBBh8mXllKRJGjwSFzOl0c13YksfH3T+L3nefzg0/f1REX6QgSDkOnSCEVuLGLXEs+5tZJa8sH+mY2El8dZrC182l31IZ1oAeReL3n/Gjc2jBvOxH4jMOCJ0PEXVmMprQn2aJ2mlmU5wz1HI9u79MG6D2ckeXhtF6LgGvdvaLGg2r3Y+qyPeh+m1orIrUZZIbs2yBS9NFkcs7kY1q21Ny1Os00nJnLcmhIAh3HAxfP/LUgyp0mHqUCwMx8g56jFS15KSV9b1wXwDQdYUxWhWFh+mMQHNCaWhaY/emz/xBZ3Ny516ACZa3GMvzkzh9AmKp8ne2Bghf1NacgGhVa18JZ5NRXZUBZ+yG4m6QcPP+CoxUr+ZTy7/yZtFxkkBafJMEn6PaxWm7Wy9YrY+fgKJpV72naeZBGRtDvTLWTFYzzbNt9GzydsqXb9MfZ4M52LcBXez9sfNVR/DTMzoiDxKqa33SzgXKAatmsgRv5NPdtIa8xX6/RpZAIxrpbTQriRncQyBQ1PN/rGNtwvySn+HMz7svoe/b2dZIaHlwykxUiwsTk2atL4jRo3vHv/NqF8HMcPdmMIUOwgp3red/MgMwiWnuYwPb+eYqyT63iNr24o1jx74q2O68zojHIEXE2QO0T46ANn3NIasU565GsRRpsBCOna5GEWgN9MybnZmUbKroMqosPq1ZfSBnocPske0nVp2+D3vCtYL9bimYzA0A58DQwiQpuu3V7ANNZQScE+gniQoZgwsRTg+nPDzvGQbcWHZfjK5ZRIPvYCGWQUn1V6tEdbp66sEpDE7FYJTIwL9rUg4BBwqRn9qgh8p7dr5KzX3gAmQhq1dsENsMPJwy2sAnNBBHQFTzheKofF5CggZbT2Y+PM3gDpbIqIJ29wu4cQU97iGwTnIfqz2Q+vh0mUto4SO9lFTZxTxNL9zo5lgGq9fda3oYGrV027Y5TGpnokZXqIgV2gwDU9XHzSskzNnlm9nFYqyyByVdxrbQ47plSjmY43V22trTqLeAaireyT+b0S64TnxS2vRo9w99mG9DfrlTtHNX6DwpJjAN1bLQ4lh/0oQLbRWfqtVHunRHAYPWhGQuMqtbgW71rBZ/M2cPsnDQjTBZC2W/D5pz8MMMW9T+fvAgKlh1iI809Co3IbyT5eU/l+RFLcZJ1KoydOcJNehbyrWKQHh6SEwyHWb8Ubn/UR2bfokWs5btREyWnRWXjbZfaDkWQFJsV6OT42vbsSaySAmqe5pNyx0vq2MCvlXaNgYFzmWRtDCPJ8T3VtpeG3lVeOwCloOdnz1Hrk6sDB7vL8gEQOAt4SYRkcSimR9uB0atxqxNsctCaI14eTIbTpUxFbIxsGrYcE8zNztAzFDB9gLyanuqMq8yEY5xSiK5OuxcWfMeeCR/7iRqCLmvHzQGFwpJ29fgqq2TYqRZuLmr1siNrW6Z5Y3WSC9X6FhVpDB9BKuRvnfaFiEo+1/TIyDkEUddyBlq9XuN+6pioeVYDzRB+MEew1zHjFkGTUVYF4RPxutVB+699R+VlPZirMrhWhpTC+6Cz9Rx0jo61ZJFEOaJyXxtp2zrbPM7pN5ihsdNi19jdB4RNY3T0T7cesUBCWV7hiLHEsYdZ+MLkArCaaAycbLFuUl6eUTtoLIfD3yzdJMyx0AN451NUiRWKlWVfznnFrbS9xyZCNxlz76IFcYTVdSQGwV+LgNwvL3n8vtry6hSDIAByl/r0GNjQs1YtNIcNoDCd843tI9NMkskn4lBThqKLrw+pXihi0H5Z+NUAJFY5fxzjeaAPZYMPsKaaYXlkqxPNdTmm9hiruJjPyu+tI4jqGxw+tl0HJGgaJA31aRIhEZnv+DczujDKegAeT4NQe7rJA2PgKs/p4GncrKIN7+JlIlw9apV9M6yV5mcl8/bsuWZI/OU78JNYTRppQt/fORaBRhTy5ReoXZeq6f7spe+O1dcLQXvb+zt2p2IQt0BPgkNrpmsTz7nzbePEZHfRXQRrzh59NDa8RJYn+VpAEdysWAt3uUzbsD2+ayKH/jyddTNIrPQq6rQCcLYsRsi/l9PL/KSxVHlbHaN5rinRTzoRcRXrtfESU3ZLxxiW6iaaRqP3/jIfPEW5nXjHNReIdhcSFRb+O5c3n7oddMsY3IKFzrlJE53YBq0phNlOsDhT/XbRG6iTqWiIPUXmBGllole8ZaEKmJBMmvZ1VBvr+CjK8Yn2AjR5SLAsz8R/+0xgxO00l7INSr7jW3DCrHSFw+KEx8UvCaDrTHs9VNi06Re+7l29FCpo6HQ+6bUhGBndlwtrTB4ujWRQ2rrWi5wZginUHeWwB0ZlahvY01kjT+/awq3u2WR7b2UZPDHbEMDXpyVjLDbH1Mzz+0LBO2JlBkXALopGiuSwxanMVTmI+Dewa+mnYVKRPKQKksdnoNyKneRhg1nUWP15IU7o7ytOPfnt4w6lYPzZ+5Q8jaGpnQcwlafV3CC9G5bARNyuyzL88UZSzU+P9eqKHnjAYTs3tV0Okd98te6HX9RAxlqS8l5yf7gp5fRWlzqQu/qEw80s8bMgMso+cZ3i0hMiaTHPIlW8i5fR604myEiBGHxOHtGusIimP5Ov0X6KPlajOgmeGIqFNZPsCWmLBfTVGWbhjsiAZ66kgP0W6PSVIesNHDWhaJUzz5gL1cOyfIyZYNaU6Cgmnj72iKRo9Ouy5VdMoADJYeXQ0qaIQw/lqMe2OCm40K/B2X5Q8Hd04ttwRwFI20+BvSgSVSrHV35HAtt5TB7BYkpf48SrKvGbF+MFRtJFi9UeOHmqFBD1sMTqxKyGTFjhv2nGy9Xb4r31y2Jysf3LY4bDlUs8zxlEysKGwJ/OH7lH9RVdx/AjPLGSRr8x79t0BWfUWhjshsEMhsQiektUEJdomYJ9hON0wzkiimQ2hlI8h1LqDSYJpu9RsIfU202LtgaltrCQW9+2odi9qYgCT5cglzp4zFP0aR1kEzhUBg1KlETAAb1Tfj4G1c9FbI30W4WckBOIneU9fD30gsa+c/ebDdmjrXyHmqRssmjxLoL27ixYP7NssfsZr+Vihvq2tgqgBaSSENgZ9Ff+CLk2fDb/8lyA3C3Bn/hOJnd1OjRRsHWJdWg2NN0TgKQs/jbdXhSUF3WyRA2Fliqn6tSbaIlrRRUKcsG07XQjBgTX9451y3p/6Qzktco9voJi6xf4LLAxtqPzDlMT8DUamulUcepsiw5iDhhWc6giv+Hmfe+VLxxKUz1hgq8GEsf13urNIQsRavnxIc1gcPvSypVO3cku8nydT5a4d+5K1sprixoq0qKsIMU+7hSh0uVMX/yWAO1KskEG9KEsZ/2Qr9+Q/a/GjNtUnDWVnAnsCyIWFudGuBkGGIlMTz4cxmh+4d+d+1H6Hts9qp2WfEwbv0gZ5ZxSXBUP3iuiR9U9lqRKOKOO2g09uth2LwdWx9ZPDHJPS2AtaE2zx1uRRGpq5lFRFOKrZ/kRQLX40ebVKE8Qivt6Tj7v0LQZcxQ/FgvKx0q7aqC8wFe83pXk8+yKg4hWinJnbr5gFcoU9CLvc/uqQmvL6ggdwQnKEZxK0550uJdF5zAdol/6BcOMqZlTjh3rinMy76ChnmtH6DNek9mKJzPZCP5bJX3zpCGejuKzZ8eVH8lbjZTBRy+kayDIuaffSPZboispDujymZLb/EqqyeRl1HE0IAl5gx7tYSubWLbehRMrcPywmNqZ35Ri+i419KmY3t5aY1rouOW1U+cKtoiz5XivcfpQlo57knFoWjKK2rEeCsWSYSVxRhZ06tMXYZEkDJ9kM1fIEJ3woZUrjQE7aL/xi/7t1igh/gjQvSppqSzIBJ+F2S4C/ppQEp/fyiRcRPwRpZ9j+lJ9SgGPY7FPRfgNAyIkAywy/2teN9kcLedC4CGnq704F98nPse9pKMvB668uDrTUXf56yrrhRc4YS9J8oyidGgufyekB6Ou9Y8xnIFFbPvRmu0aLCro2Db+nc0pPEdEwiER5JC+lJLEGA4I40lhD24LF9SNvDsWj33P9H3Dg5RuIfjlzlXrxvUUKYI7lrWVPKhSaECKOiDfkQFXGaWUBPGz+AEmVI503Bx3v5xBTNuvpo8TSsxB8OU3yLoQzFvsvCmjss/txA1oocmRy8WbERDCvx7+fBpj2h+39eNRvJTx7GP7GXgnAISIFE/cePsk8dXt+ukvSSoPdfHjV3pAVcLUgRm/t7h1dfxOnv3IleRuH7donW8CaCqjEN0xOwlFqJlBI07JFnNj/JnmyzpGw1K12umRikX4j7J2uj24gwlsjUlAzd1hOQVe86UC+LR70pU4Tt6jslTWzUZp8GaMNApY6tAhX/sMSjKSJNsRGvfgpAL3XrUJiZRC5ZiDi/JhuxghujrpheC4dx93klpUL+MZQfq7+zg5BaD0i93tx1Ga0WLwP9WaU2E5G2+OOIz48exW3AHLAI/xv63pdcUjhRwzouFDliKVWbi1T5zKXJ0NDjay7abMObeHpGBcoxqOrT/g+YS0OEpo7TAvBIUGrop/vunT7tslcNQZZB7XdfcJYx/tCZ5V7Fk1ORpjRQbeKMjJuqYD7AlnCthivnm9AvnJbix6Fs5MVORNg0C6ukW85ag+V5pyZ7MZ0cEN3CvsZW+cSpqjy++Edxh0PRi7EajjsZnFPAiRKKRJmtg5bLIWUG8UqSqjsfnWYmna9Gh2A3m9vriCrLORmaL5NJDRH1OkuwYRXw3HchnCfu0LqZCFPCes6VsXslwWx3HDc69DAZsO0bcRTj6hBdm3NdKWWR11hS1HsrDtIgmqKByzWWnIMslkjFGt9nUJIKRudWjHfOuB+B9vfbgy42qoiZu/ak+eMsHzDNoEn32XBhLipEnULGNsMmVlBbS+VF1SlFFlq4Nwe6ayCCNM1iGsBwDsVdGK5gHKnyXOMvTNhqbe1F0CwLFy1CrP8u9xrsSpzf0WCQFdc1hV3Rdn3w92XI6fwwDJiXjda4xAFXexTTNUd5kOCxkIw5rKqEEd4TxEsNtQcH6NOt4cpExSg2TkycHAGDwxXIbSuflp9WCfd5SEdsQjtpki+BQKML1Qx3rFyYKHg8q0b3NuRso2oW3COMeTOi0nrg+ZmpnP/u0vDSvzPQsbcDgB5Ufz/emQLVJmzSAu89pcVHZdgLpBct5nfwElnKi5a4OvIggQuLFUpt0M1GIoFPt2M2fx2qajyHyLgOu1VNTpTWAQdDA/9F0h47bPWOUO9teu2xnujd48pjq080BSpF4zaAnbwRGXPggmckuIOkFdxVrYYy1XUYMDIKmN13U1znzYD42yNpL9btV7B0DAmDqgLhwg/bnjh5WGZ52kxLE0zBG1VUjAOjnAw+HFBl4kQO0TA9oXG1vNJ7FqYQ1Udeb4knr2nI+i69HcILbfJi4HclPKEVfsmxPee6AMRqW72MuzRXbhJzVlJRKv0ys1XtBiFMRYdvLcqQo/1AsQwtoE5GXYdBRmsjKcaok2x0dbZCWUJE0JbBiJ9/L18SF6VTksyXsz/fTcgIfLL+nO895k5ciHVvh0od7nQphB44wp8vKipLrnPBBv/W70S5DzZZJGTVTJlQYzLrzw0MyoBhyHABp8lelhjSMLbRGaui8nNMaorQFx3aFxYwwV3aokaKTIIwWjJQO5ZNAJZA7bRH64psgMRsapBpSfC+JzAlGwm+45B3pKmLU9XHbCfc9bCc1MhzDE0Ep7ryruae+sFwsoPPAUmG4iTYG62ooElij4jwzC5nfbu61sjWbVHrr/4hluShFmBhyPR/vL28FuVLG+qkeMHFnt4EOdHkVowhKD5qYhKu9NPldZsUenXfK01MtTdGfOEKA9OP0KAW2Xi3MGISQyj86m5m2MnIxfZhNHRut0X6KDAeh9AJ0DNO0ilxnwxI0dn+Wm3X+CHXEupxZHSguASiRYn2/vdZZSVIWoQnnEzmtDVGr9NB64NkT005KZtDuj1+ne1JNTnDZ1lmqA9i5y5RARC8ylpM9Ql4Ku7EdIqRfQ8UzfctxOW80bhf54fMepqzBs1UtsDpiAImJwjJAgy84dJbCFtM4kigwb0OPPLM+U5V2Q55o4PnF8KrFupcr9mwTwzWYh4GRhoEBxxU9wIngkfh/fROfAFF4DyBy4CP3WAGAZD+kt7sMSYIGNV+7sd5QZOCk9ShgKXtbnGDGH6C0AI1HGq5N5FDcu2zg83BDyxKbDVp7uzNegjETjbnia0mzkcICP41WX/NhtERSvENplXSr5yEV6ZcIEauz3komCBKfvl5aKssqh78jBXgZ9UUzJ7SWDyscg4lfqaJoKqEEIWSAyQc5yF37RvWiZpo+ntkFoTIIjuXbTn5EcuUsowg/zLoXK2bMFEK2ZMrw0oZ2t1pe+IP/38wZ75+3jDTp507uvXPJuDm1JXJ7xaMMWPMuzwiTUXaPIt7OzQSeZUgBjQygiLxakTFAJdDU0ETmJ44YWUNJe95cX4PjqABh3WDfSqrhJfJVDSW2Op/yTMbVxg9C1KZBDy0BNsDbGIptICMMaz8kCn2qYjtG2FePxbjNEiZmbFVoXYrMn7UkcKBS+/lO5hX6WKrNmt4f5iNaHgD+eAZNJhNbHdJ1XVHuUSynUbwpix7qKZ8SubjbKwtkHcoxpsvI1wf1cMQpnSBxnyELgB07Hi/Hq1PQvM78kA5QxaUKGHGOq9MEqIavLmcMmgd3ZHXtIkrtnx8R2SGxvYSJv4L29JATCxLXv15EqIEGSRAxVfVJhIKIxn9dhKle9EMaI2z3dQi2SJqy8eTTy6pJ0dk9vul+RYkjsfYj0mXr17A/ohl5W9W+GhaucB0NfMHB/DybzRGQdfWBuXBoOS17QcnWH/gBeMQtKYYs1KPNBx3WvIC3L0a1qFXsMOkbp4GDCebFXcRX8ybPNi9tIxfGahL4gTqYhS/tuS289sSxPMNMfsq+py5PqPldRn5qMlh7CFk73bOOJTvi2Kj986kHcZ2LS75E5Qfep8d1EFen89qxQk6zbfqDB292QTttVB5UX9puxbGUgJ3mwf0/MaDCJp2BZZ3kpAPGb5dTJuxViCTwh5Fuf2IRCjldZUWfd69yE73mFAKaRpmz9GlwedPw==
`pragma protect end_data_block
`pragma protect digest_block
9c6da9dadfac7c5531c2496ac3024d3cb5088b200f9fe97c1826719f8964a567
`pragma protect end_digest_block
`pragma protect end_protected
