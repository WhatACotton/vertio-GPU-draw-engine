`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
HjEydGfFXntv840YOq55PtFRUzZQ3Z7FUv9EZQAQVqE+X8ll25hGOO7XwYQdVaRcmpy1N7aPvo2XqQ+akO90wvx7dNASCY9O/M9nu3+9fMLazJf4xOwGcOSV4KfzeDCtcVG1Euwc0LPXvNYhNoKOq3Xb5wc6G0BaDpvc+X+Bxncug/9A/oDl3yPrw83JdeCptENseT/zskjjS9drhDPDhmbCJfmRDg4iU9yPfW4ti/09ugN11p4BmD9evLpFgWq3gguptEttAZ8ypoo/3J2CQoPuEkRKSY8/zCJdI7E9cqf/YUz+W+e9/gVW8WFvC8KHiYsVFNlaU4DtY/Cts/XGAq3oEfNqiXg4/Qcw76IuEkuzPturfjazJQW3y8U0yod7GmhFZyHAJYnyW0oIXGwi4R6EBAQU4QA4I6+GRsBCLcGp4/M9J7MKAkCBInC77TQKYcJ/I/A1FGjdXQzub8jRu5eSwv7jGueQZ7FfWC50hBoYZ987OxfWHwkvqcYxMy5brr7d4eSWm0VN5i6YlLvSQuxyB4/ldBIXvrog9vGdtqmAshO47iL5OP5RPqYAnDD7c66JStnd6uFxmES7MU2nMgcpWI3oqEtMc7pG068obvwNkUEuX68YIsRzwZ7tfXyMFKpypLH/082Hyo46G78kYv7HBzY4+ouXBiK6+e6ogzbxQDH5WdaAxCtVrBLF9UanlQT1513IAkMvaPoXfaaIRKLhSaTtHRLOX1pcDzsRbO3N8LjufO+Zfa/mvfLRYZ6O1hCY2g+z25Mb+bN1ewkweb4t3055yxVZTWdVXY7wXu9NB/pYthEPc0mR/5VkqHfbVibGPAAqNnVJcqrvMAWlebrNpK+Ii0cJxXL8MfaOlVaMIvIcaLW97rSFw6Pw4Pbdgmhx464FiTsrbfPYyJZnLaJq7UBOm1RZXnT9SQe3aRNCXuP1s03i3ojDeLxwgGlWJPzZ2876J/WJYWv+o/oEqvsbtB/au2fwdL6/0yJrgUaj2r+ilP+Ae1cgUlf4LGX9ktqIYLEzMyCfPAGyEPsWmTqffFmxfRUYWZnvepjp5dIwYZG+bU2dv5FsRkiPNFVeAF4IMM1MzU/k/M9kkKwl/v2sxAxx/8bt8htErzp6SOwXhYCnFlh5mPb9Ib6XR/oG+oVEyGoXq8fVYgZZLUlYo3rlfgZ30JEcMvfMQeJ12Vv/CIikFmStioAAs6Z+gb48hEBYAHxTTYLsDCmQdzjx4hXw8rtWFRuRoniNfkGVYgLpegKxnDuNlU6HEXevLZI37XItA5fcMwXRBw+O3+JqwAJBAPvCr4vrS0CnpqFUB1iahYGH+nV5y31Lxcol91wiQ9exZQUAVqU/gf8vPQcqb8PJBEwXZELijW4Kii62Dt6N6vRmE60SwnMNm0Kjci7Fw/sPgmHct2A/A3Zfazm6xLABMkn+VnQTTyUjdOW5WLrNQgIen60JBpnumNVaHAwcl92ALcZ6JhLMVwHrIkrepkZx81XGOMFxLNWfN36WQHqLrcoZeBy0q62u4OZn3TiKaqnvAEMUdXSPVFKDRvrY2EVu8Imi7wd6fuq6gHLJzCtMcTlcf7SroQOnsoy/Wee/nKToS6kVTD+2shLAE4v1INTfSUWeyClqyGLUUGnOUD53bNnGAWmQrYNcfq6p8GyKyloHRw96jQbLbd/XBCmN7I8pE+ScO6702wB4RPnyFSvOtmnN47a5yLa498rRJGxc8qM5uWpsQq47CFlT/GJdcFckylbZxEALOIXJhjvXyna3GEaGZJPblGrx4gGXSX9T6Qlr7lrGiLZ6CurbJ+KFCMyyeYDEVo5WF3LOqtDDGDdlxREnqn3o61vCQl6eL8ROonv+7Dl8Zrp03N1iDR0zeHvRtANKjyMcetln0/0uXPQ9hPJn0yyYReF4sgNbV315uRgHharm5ekqYpgYTg4abpKtOYDCSGeJSWxGpNSaBBEBelpKYYYpa1dfFzCzlzGMpB6FNu6zfFSMjLa5dcGoPCXclMGi3Sair6B86vFG6DoAVoKHISFQ4Apb4IMEDpQmrtokPNEgUNfh+9Q7e9JSkVZ2xiIaSIIKpCo9A+0yl1vvNd30nrmOnFzGvPLcLcdGHJOt0CKOHVM1tQhkinJse5FbickbDShXkXfWfj0nCIBHbF1HzBq3b2xb1mOt7eHTiANx5LrpYAHzj4f62Gscy7kJb+FGrt0gxlN/oVuvcbtT2owEFDXIsgzIOHePERC4OtwJerdBeUS9vrr4E84xydoMR6teSnPnel4sK6LNDthpqy/NqTEZMSsIqXLfUZk426IQ2CfTdFWI0eN3ua3JU2mb0NHRRiXAz9jFOZwUBGGk+y9MxIiOsSnKt0ZIKzJU5y4zfKstQbxJj7BpGazRTH4RatThfytAnNzhZvRXk/fZvNpAqZ20GNJXLMNjuQQdIXLiOEvyDZXBNUUtItwLZxHwI7nJC/kEfaTaBBdJ65vVk8tGKROqjIEzQV6cA2pwq2obHuxF5D/wL49LtadfVlipzxcN3sykMPhWM2nuSnnHLJ6psymSAaE3MjESxZnxm3qHWllwVnSeIA9tmTZpvrYCYzajLM3GGUvHNV3LbywRjpOWFefkOCyQpL3SP8GEnrCfcEL6kD+9f9nLc8jfYRmZq1Jy4d4FCG9IYP+zlhzhRF4q9yNID+1xVJOeusZrCdEeoZ2AY6cmzE5UhuhYln5BIZF/9PvD6kWceGMgzCqG3IXfPFPRxib92nFA/hxS5VQo1dbXrWYcbJXqRm9Xcd15YBWIQJvxk+i1bu9IZDvNbLBoOHP2by1BBDN8CFJzpvw9Ji4OXHU4MHNueZfk0VUEB8DmT9ErOw43nJttADotkaUTy81LXkzx1ElCutTorv8SytiKsGt41Y2dcCKMQSDqPA3nJwqn/gbnXkwm/xqWbPPNIrJ6BYOz1rlypa6zGj1eicFwnMXGYmAawxx2+72HbXCjXzHmUgI5zvmrB+kgYzMYBi8FdP+UvBlM/ZL+Jh153Vy5jYUPlf/5lNpwmGicbHS9uj7CjxVKeyxoE8rTQgEPdh+HO6xJdu03jdYX+zAA5zq5DEnbqwNM3bEjkAf5Am5CNEYln0FQGmgPViiuydAn3uR6seVmkvGjjZ/B7paVpzRKcBfSmTXRDTOfN/GokWhFYZIv7TZ3V5T4r7Qtek4dZceQIrpQfGpk/fh8rPvUBdz4rksw7BayuPSYNkvo3mHLVz6iWM9PsmqqWXmIdlu5jSaGCcuBQgRfmzeZjjqJf4TO3CDubvcYzW2/RyaqdJ3BpK1ZTQPJaEJIwZ2QDr+rhuMSlTZ73lOs79HvkHkc1vptJXaQQt2ub+l/M6q6CJ23araLyyx+/4VG4p7OjuDdICKrAJcNpluvVf5w1p1hZeRPya9gu+jKJJWm8kkk1G/4ZQYY5hIG8pLBHevutG5Bxr8DrCXUtSpHKPKRSZDECo0Ic6n7A3PTwAajYBcHY2T9c1FybSchbLZEqOKrEd/YYY4VR/ThOXMh9lAWsqv5i6rLmAKBdiguh3pH6f1IEd9wm8EYyjuDeL4AOMKHVjvD8eP97ygbmOvAWsrQX/ua40Ds0Ji/xtfuodg7BmK+Ae28QsRHcYZmoQQXOEitTFcBRikFPuELL54vWp9xuTER/NXMcFnKFWk/EJfnvYvb9OFW86eXTx4isUwjECVyJkr0sJ8kQ18ghJOyzXyfMVaL5/B4SGEzOni29v1/XIjTQmqTY54EqR3gxjVDMQxx4sAOVgx5Z0T5Fl7iTSFL1BM2jpPJ4P6TFZTHqp8krH7X7txqJidTD6zz69kIONlEETti0OjWy0BUr0eQIOs2wNFWnfvcvmwiYmO4wZAKa6Wwy55OiVdjbDnwnOVqyr2IsaEW3fKlPxUBDDXJdjIoakryuxBvKkTbw0EffmNR/4T3SDs8fTGcF5m/jF9VVYgFVdOjXGeV2VymDxRfPLUF4DR6nGbpkFvjpHHG2nWDzCFPFYYdpWhL9IG79taLQ7ZmA0AskAMujaJ4nGiVkP/IaBDw8G/SpZjp+eoT+vMIH03q/4/O/D+uIhT/cPyM0cmiGtO8CQtRyqATQy0TntZGAIsbaVADjFZ/Tj8DdXNCGYjs1+aU6SdYe8sSaAL/TgLSQNi16ZS93nFrJ5KGiO/A3Upw73NNthKmp0bbOB7LxIl+RwFDDFqW626kqsnEhE6xuBKONW8vCqnB+2Huf9E2Q6dLxYfjThH6+1dtiSI+17NvPbEnnXgTkmpulczh8nwCi08yrCpePY83tW82D/16W4fJdgFX3puNuxf4O5wiwPKfHbn/kW5keAqHDoMmXRggStyTIUw2/zz32vyBL7BsXqoMIw7T+Jx5giewfSC4loQhqmUiqLQnw4QIjyDlacp5/7CWYoxdI3z/Nm53syaqbEfZH5v3z1mMQF0uxzNfRACdkMRZ27JSYhCWfQVANCoabJTZsv52VQi/0fswX1axAoncB2bfgQ/BEMq/rZ/yYEGgqE9RkzWtrpd6ogAz9xz9rr7HyI84+1itzsRZulSpBoV/M6DTY2+k97WwUQTOtq1dUxdk2tL6/ikdG6GMdXYyxrl+WMoLZGPzoPw1ALPZII2SdeAKLJTVocl73samIlU8i3lHLV+lxGGNFl/NYot7+2kme5WvJfT7wItLQCK/IyGkIog52bKvQRhwP0p1Gf+iKz2QO1xiWKQnrO7Pc030Aw6gUUKcuuyfKTD+FsASVu8/en7GnAN8iKWL+/QRj05t5RUOC4GLC/7fqZvasC7qfiIi7EgH0Mr8pKF4TDZ30NLqgv5rSestWYRVjPd76eQoOU+6ROYasCWhYuc+3TLaHRC7ypTtXzzpsAUB1h54LGPs8vN/PP7N1EGju2XYGO/+kt36Y9mV6ggEbEZk8F9/xYrm/tImjthiEFaa4korCuFGdf6FFMCvWVwvxCxDAGVA3a+j1MhLu96ulr9CwL/AFDKe8GotOwQR+fIXkYrcBcoViD6mviqxbuyLjaKPVJSLQVzg6d9v0AKf3S0dhigRqbw3Y6N38VkIquNYjU2FImb66vhVnnZdMc2QrvLvkt+VnrAC42TJb7GSV2zIXcGzgrJxBI8ieQBXWCuZ4GU7yRuiKPAtz6r22CmBqE/mNBlYFJja+3F3ZcMDtIClWDklZYBn5TBQHq4S78NfiHiVbL5TVMGgLovKSDPnhIIJ26jX8u7abU9GQ5BGWlmm6Woxw1A7/NUd0YxZGU0XWjac+lDe07R1erUmRtTWBoYtAQPYgS8M9disP8bq6U+X9UOJWvlazfHygt3S1jukY+o52dyumezRFk9eUAFqWTKErR71LEUKFvRQXd+3uvwqaZM+Ab27mqztuBfEOBTTRbzmvTDpqseGtS1wi8QTuOfMIEr4P/fEvRCdwpKAk9gFksM2VuzeTA+REEX1Xi9aSMKTGBdMIpDPlJtDiRjsHtrqJoPP0e6oXBXszD7T7t62F4M6tR93M0biu79uj2LFLARVKEWOWmfpKbFLYU4JBO2l+I7kpo7qpdfijs16bVmwM/ZEBBZjjXnn2guiM+URIjU4o4BvfOAA4w3eN72UP19VLfU2ZDWQWk646hAq7L9WpHltjiZRmpWn6/2H59tRVQ7t4eS/854V0xt+wpIcOW/LulpWjUNmg1zsfK3ztH6u4KWIiiVIZRivN1xmEg+FP8u766PgGnoySMt4Ksry8uwtovN6/TnKQsdbbtvd6ss8hmAQwrJxxqj++h0AVMLUJ15LBURhSD7gTj8e/kVpDC1Mt/PzIGbRz8uhUEiV8Q0NVSd7fNmeWbyP7y4R5nJpvh1LB+iDbc8PpTdPQwMiHK4+Qbn5t9pMIlDY+tPo9sliWlnl0/xLuBr2MMaP96PXZj1JOzoBLZViSX/VGFeVilSaExTyrBe0+XqF8nCS4G6keTMFhMz7y19T49m239RQOeyUL4VhHhNUs+O183+9PM5UVjRA5kQa3FyRLn0IQNryvNdMXGaLjPts8bcTisbJz9ce6My+3vKu9IbtmdtodKPFet7BjSiiIpqVV0hbaMiyszz2wt4JFNPqWX/iR83n+5tIiaeNiyyF76L6VTEAclQFqR9YK04+WYuHcnDvxqO8zQNmuOZHYGQC1Kg0QvFcQjKy1kzT70qPM6T0XYQxvbdzvXDQAz6OKY/pZbSkrD96BtGlwC9PzoqvegQB4YRlYmd4YjH90ZA3VTWFAcDq7nZNG1IiEA8fQVxPACkN1DqkrogfsWUd8lC5fNzzD09VoKCJ/Q7Ge389t6YPu55CiFUr6dkP0VQk/IOta8gkdOMxs9rKCvYp/rcpaiqCZyQAV51uR4UyQUynv3C6XFhRItAUT4aNeMFEJyYHRuNRQ0hzlctm3MmSoXcIbe0Hpn3yhFWjLJcVI+rZM5e6CvRM56N83th3O7mztQogXNmeb9qblusp2FAHGG39HtNaqUO6ZIBF65drgM6mxwA3V+U6AG/ePAH27xBdMVPahG3ryz+Vtklk715rtEQfjleqzPUAY3YYWNkdjvopq4GjrXAcN/mJ9/cyVOWT8DmdVUkt2xXYOyBjlJjz9n+tBRfB/teyA6HQmnRmUyCyEMSNcJF6HEb3Cs8pCnG+6MyUNhQXxTcBAYyiHTuN1zWOjJM9PEZ3S4eBuJbx9yQsq6ze+3wqlDp5EfZpQAMRvw3BckTHl4Q34uQ3NwY6HZjHmJrnrw0wBUZyOXekIfESA607i239jLjrlkT3w7SVl34Cm8g7J+JGBlW1luWJkCDfUI0efwnCi81oq9c2tsF43WSuaanvy/6l830KkAxhhrU3f4kkC9o649hrILF9mwOmR/y5mLDD44h8xUWimudDWo9rlv5c9ZPtK99S3AG7xPyIXUbGduBLh/HpSqsnvnFpEEzKMEpXvNMNLLHDTHKp12l0Kk39QhyBXoyLFILhR1ChS7ynCOMhYxwJeP45yQMRz2gfdniyhksMXCMKYyYYg3/bhP/qoQb35EU2am5pdjPRFFnqZ6X5ph6XJjxT4bFR1R3wPFdoqkiq5c6NuSMI0hewvNChw91ueUMvglCC+aWi3BSMhJbaHPfMZqX9BiAANIIiSwgJ4YTbuDGce0CrAMGtyeuaf9au1Y7Az0gpMiIzMeEMF91HglKDm8OSRqHUKZwbNe6j58HVUdaMunuqLT68CCITpRasEDfqmAKUv2aPWk9mdQjAgBm1LccR1igscEBojYok7b93ZlogCyplkMOuP1XB5PjscgRjZZ5cv1ghDApU+cfoTVKZhm8OHGB4JLKZ9EWjdYNU0lIdq3zvv6eKMl0PSgtsbkKpx0grXE0JGvxPTRvgjo8pJqMcxn6cV+4UD80yuEox0pgfLouyIG56r58OJRb3dzy225VofrXWnWHUxapVI95Tat4zdX/TP2rVHuPzsq5NQvKyp33LMfvUprulX+gPfhq3105QY1WnbCnwQbXuPZBTIKDexwS8tfdBEmkfoaxWWXuILkY0BMZJS3dCzKWQF5ca/c9tQAFZTQ9IsmaWO/0cbRNHlRYI+ZcCC5BTv+Q3cWCU1A7Pk/ilDG5kgG1bDyJAICUuD26u6g1yyKMn/mDHm9CIT+EYh5WDcbDBwjvnlq6Nd/eXwhvHULBgYmBrDPyB34O5LpR3w00h//Mgwkl+RlKx1KDU3ypaZ4pJ3Cv4yU84541ggIT85gE1fzwdRBtsIrOM27zT1k5+Wd/4fLIEEU+Pwqq7WM1Y4jR0d+dr4d6PyxKf/mmFTL7A4sfaHvq84nQXyjFZRrIYQKZqbwf+j3x/oS+mPeCd8A27KsU7Y9Oah7wIIJBtOL3xqtMAWPc3F/xehLNJwFaOnUw3+5NmgkL/eAjKtzjWXkE5yFTDwKMxwSMqVbsS15Ydod2SeT545Cf6+6M7V/sA37CJQjAk2z1wqL+gvNDj2feBOpvSDAr0zVJA36JWAI8XI3HZh8aGo+vVIb4YDAZ3U13gqTkAcoVDQkv7s0an7LDB1CH3MuDduEsq796OLrgAuozEb+Ttolso4G3wg3Yp/IaBeRdv2wUqh92wjCws31f4/px3PRD2db7pLeQ14m+bsK922f0XipAQXgd6t3qJwvzS3YDOaW84OlZmeqKdQ0YDnTs8z/XsFdW/dIdtwU8g8TiRKtMtT7T1LA/wexWD/A9BWqFdkksPyPa0GVFjOHBUxghLtRuEcRZAbklrVrr4LjTN0a3LOAo/GEU+WkVx+CloPFMX6FZkGpDHq9ZwhZbZXr66dpCw3l49UdfM7FzUQ4ilOHE144V2UiNQQCt0gaiCiCoUVxuyyMJUQs+vbQ6sDrS8Hj8vkm4xMoi1pO6lUt8iEDp5aJSiSp+ZXf/l8fBj6LvDYSbTHFYo5RFN4jQSBy2pefiDlIXwLzVqXj5v1WP7L6xrPqwcmd8n6FKU0QlAjOanpdbnDaEnGrPlDCF4Kc+50830hFpja9N/pv6LL1HykClDvPY77mtMBTIzjwo04rtMKR+i2JgL2kVzUZBZw/dEGvMok/1r0FVeKb7KXdybTv2jse05KinI3BneX7D37Bq0K7Lyh+BP93xFp5eCvGbTBlov+xib/lNyZyCvlM53c0fX+S9mxms6D3bbYgf7ro++NqPjZPcQcKQYkHPrXMLVyp7C0To1Xgj6s5FN/XYtijXMhdFiAnDv/FfbVMYE+MI0SvoVdIlRElhvllFGQ1dgqG+vJLxDEFI0Uzs8BgW3LIEymjYrbEf1YYkdyLKFBxmGzsyneA8KH6ZwLlov3nIzSzMSobjpaoBq2MKJoWxLUrkvaiNyAAqpjx1w4jOy/BJGe19dMwFrS2XLcG7VoZB2Jzs6jf3ImM8zP+3zYTpRCQ7kWBZtLOaIhAcZJSgcBkaxxFhmzEcqpdilHgKy1xi7uNFurZfYNEUsvTqSFdAZNdYT+JHQyNZBHxBWRKZIjfsrdmGY6jna0oape5EmN+JP97Gn0+2KJNk0RUB+3XUn21F24pvhteg72jpOSgIWLJDRj5/JpfPRsPFQbeXDUsoIlE39DXxiJ+f071acJsOmdktuznsxTKej147cnjL1TdSEmzit0iF9WBsnLM0yn6tj2ijFMXDHqBisuYvT6BXrh2VesbSaV0W33nwMLEDYSL6BV+5d9qpsNztEkEl6ZgyYg6r3YZg4T+J/PxSzjZI9H5iETrHND+a+OEYrFwivEKdQiai8oJUyy2NT/XnidjcvDal9SBPKkb5VKaae/oIUlxkBAqSWM41RPHVekp9YKBSXcSf9c8E0u/U0BzuB/W5igoG6FcGS5/81ButH8zozzoFbyijolAqTNRyf/zZBngKqzGqS7sbtp++mV0B7a4uYpPU6J/E7orHMPDHONQN9FkmYUHrvNtpcucicsSsILt1uPh/AFRtpewBSNoqFpqSXDORpkgiIXSl7HomQrVrh/DMSiVZ2fmy2nrcxlz8yRB5Jo+knCgsTGQ6eErsLOuHQX3yxiQyQOb7uTh10kXZzkvq998WswZZmQ0lP+Fx681bco3GpFIRZKHmAvrDNvUnp/veiRh5DKA1z7RP4iZl8hwILUXXjA46S9Msgqhqh/LsVyvmV0H3gFOVFdSzQCWp8XCuYKxG+RWG92amk8yIz9zOnvJb2XDJ2hSVRkXZ8Kg39WLb6hj5FVnwUujb8cadjRTX2sEXk+dv4UGA1T0KRjR3aX/0B946keuvVJsobbJi4bp2kFk02WX1aXhz0wYIqmtwoRNow9LA+UICM4eCXLlzkx8MZbq4lhW6eQxG4jULfDQD/Huk5lhMVuKpHYeY1zvbz/rTxK+DUAe6G/9rhJjxzV7Em80lhVuo0H2K8idhsNWwpGlkqnHcaMqBwAP8IACc8Hcl/8/84Eg1TKhVu2zUx6QHgBh0JzvN5oWQfxOBrWmXvBHeT+rkdi8YwaXZz9vpw5xFNEY4A94vhM4hQSK5VmapSPqJ+QmEtIPBKq8i7/nW4/WImUdx64LQ89rCElURZIcdXggKMrhOAmypk110QjdXXgDdw2Po11NDW9LFJ5I3ahYldmjRtc/M3gWrgG/VkQec39mMd1IynJcuvM+1oUlGPMj7ZUZIuRu9uLhr3TIp5sKKuDtAAVsy9yrnSWlBsEHSC52SeP425JSyBNeA9MAU4Q0CQFShM2tM1dbN0zLnOXWAamQgcM7NCzlM2nbRKtVhPb571Oc0SpPREfcJTbRMd5uKUKK9nZv4X3nTmtuvwpsRQL6SBC6r5h9o2rD3/5lj9E7ewY0ua83ieLCJytGRTvy+nYMnj2IJSTFk8giCPWVSr/P3R0ww0EVzsD8HNHD3KH4i3OWW5osAFy/Uy4JlYH8r54cb0E4CeKFnmwOnP9iXaMyk6oltWXnC+eXX6rnhVdDe4Q/PnDEUMLfQBNwUorzpAOfZFDyQfHao9kBXuzq/BpL2hgui+Wf/Zr4MzjhsBczSfhF9iL/6o9BGysMeci6iPjicJB3iS7419ZCssjRGd5HCVPnCffKFRkMGpkcuJn9C/5ba9ClAX9oi93xJH1wp0lO5e8vSxeE7d2TysdSclHSWWP5n0YEG7RI4kiugWbxvwpsNdF6MZo7DpkjKz5M3l9/2jqdbza68sElJBlFzrd1NEHlQ/mmWOi9wITVO7fL9W/g3IW0JWTBNLhHfwuYMXvqSiQbH++gYyVlG7tno4WxSbub2JBpwv7kGcDEe5AgYcJHNZHW5/HNY5QNZgsDFpGUdiU8RApWPVlfJyuFfa1ISnylkSsI1sVbqKaFnqufMzcziP3J/Ntx1AVT+f/4JcMZMhsVCbJukMJJpOOIaCf++kjM+CqrCzuGpxf3UjsL5x6F7TGiL2wyyW1nvj1PEIHq+5yLwcIYwmAvqAhJCczsyoZTGHOVXytih2fgBBLx41te7Ii38cP3Q9FSgH38sUxneo3IPNcQ8n+f4+wl5CRoOkIDkIl4c/Wnwo9CSNj9fdIpVQqIR237kSh3PnCkwK9xevT72/dXgIg66KQLy6UweQjDpUDVFBLDq4rXJTr13S2sdg45MT8ADIx3L8ucYnZqrD+lRtHVFMdFOaIDw3f+dyw2x9ql7G2U9HQsd0mZr2QQ2e8bpPNKIBJmjzEwx0qELf3uig8t/DPYZ8I8iQ6+A9ACIPPNmM9dvBFHI2KZvplcDkrxUVXMoGuXu6whBx+rykNTnysOGTAa0AFVXNN2GrBSqSRbuth8rzjoumRvp14BkIaRjw9UBYjHEmsfM5RllBZB7sPgmOnFftsezLzbKkVfR80JjOHqsOfX1iBGnlkkx/olLs3D41eww5a3uimU9bznQqctG96IHk7OpR5MyBaQhQoQiOKBkiOrxEZ26OwMPNYLFVzUIrFHHNmCHK9/kNfqUOPVfTpnt9rLHmoR2BwW3kuKbO+53gRS150SLlJ1plb+VFuyGbKe1GqoLnYa7clRHhZb/+Xo2fCKpCMJUlQHjrkLo5Rv0qKaDJkVQqL1+tqROJduw2PqawVp4HjeYnTWqRePMcBi17BkRvzwJLieluyj1Lw+RkTKjv6TE7B8ed8GkL6SmuqltbWm3rNQ/pUkW7lvkMlfJEYirWfOuNnB0jJH2fl840gLrN3nbNQWrcnXgiATiU2Vz0xOfXTkL1fnLIXCT7s6b2enfbYRJcQVcmqdfWGSKSyD766WfcJEu5lCtbjGWxqfe09aECEqT+Hvxcopdh+Og/FvJ3IruDuv+Dw0PszMQ/iwaNK0JPm7G9Qquqec5gGMQ/4WnkAXlb6tcJydNcmTCOP/HMbgdowvR8rr8+qRbmyBQSFaAoxNhbbdaw0dVIN94XeJpxUrcBsyX1Y5g7egNxLWmb84neKBO471hsOb0dzXuhvpIIw0vwxmfwuFbHEmS31x57MevPXZJ8sbLuT4PcH4X/BR0831nXiyx8ZVXd2iVO2aO/deG1U5Bc2Ikc/XV81/p5tqqXMB2Mw99vRFc1SkwKG63h+i6IIbLiXh50DjxSrygTjPGsfGSYxUVylM5gnosGX82OHgWuvKK2OAb279VJWSVkD9SjfLpcno/lfYWuZsJdwnN0UMcoFDPiTQ3jam+RNqYvLLxjIYbSkF/m4Ftm82N+Yyzyq+ytq1eR3XJHcQ2jB2WlERWTFNPJFfHQzOMRsbZmkeN06CH4GxPoIrPW9HyFz8fKOx9oPjlN1F/VrrIQeE/r0UW9wSTVaRH7Hxnj/B0vgs7fVcXXE6gUpajPC34JCVYASPE+c5sIMqUdalaZUBF6Wby5WufWy0zAzucOt6rWC/t+3VjgAuwE9QdrrgB2xSnl1oDblgru9haBvzT5hGA4v38EbUkVzrea7nOseDLsmX5a6k1JSUgMXnRmpN5c1atXJdHRmN0NWia3zy+soY31YWRkQdni9yHUZpFWIbO/sm0wnH1AOKga1nkL9dmNDrBj8ByPTP6lIGcO17IusJqKFzUvbT6a4Z040FDvGLHdQvk+eDwZu5CUSa8vkXmpgPKPTTuItwdffxLr5tSvNh0Vfv4tkf5Gy8DWDnV9su0Zv3a0Mze1JWylkMcVKhOwoEQd2asIDgcPOfqTsmWfvAx8RzOrlm8I6lQhTxkpLvjy3JVTaXjsI6yfepBR5F66B7DtydvXazOTfRjveIIF9gHKbiT6KeblK4He6kC80SMYKakFpbf+95RcrKjSp6UPwwiZeYAYWo580VvLi4B46ly8L3vCDAFCmrAKeexPzm+FKGshxK45v6iADcNutwQYV7Nm6XIEUoT+eJNM81fnh32W39EwvogiiqUgR5567Wdz5TUL/+0vmjaO0oMr08/hoMzIymw5Vz0Hb8RwxAVMbJ4h6FcloUJLtl2uy0iCYet52jrm2qfbI/zlIlJwZS/Jl9BfS1ONNL5aBu2TU+7j70UCnLT7NxM+pHH2P9tBdnl7etdNKUgayLLUVZhdDUrd8dIQw3xfPEjunU53oidGdK6PQQ4AlW/lyplVms9mYX6fJOrcgv4/fKkfDhXgcpfbQJiG4BV8p6ud7ntC8YhSufnGC20YIy/qrX/lSSQLMG1lgcVwsWMyKWsTGv7cICulZy2vbnauWgzUNefZRyKKHQGvJNCkWpqXyWOle7tmD3S8CN6mBmhi5mHgy9KcyILMT4BgI48Rb4JnUf1g8+p5GI6FIy8QbvVIuWtyhgfSFeKrcZnGZpS4cmSU0jBXNEu6NNPFT3FsNL7ONHQDoSBjp4h27afAHgdm4u+lg/D+JPXS+6Viy5Kz3hwF3kWOpvfem9Elu2EHZiSqEwmvEeW4Xhq51kwjd1nZEkRuNQn5cYdbjIUBVFYgsVFPA1SxDFqPkw8zUnnMjnqOY7kophojlDTZjaP+875nBlgJwet31ags1w0/lphyVMPi1putK/p5HQtTgSsADz5C3d77N46i+RkcXoFepbj9zT2S6x13amfQK1b1XHYuTVu9qxYLNl2msNDxTUr7V0pKcdzJe2wEfnhU738Rc/RE8sjznZTSF2gn/sln8FP3S/A0cs+9v0NugZbqFevHpba9nAsVOYTLQkwAoBJFPI0frDYaUVzlpd6MNY8uGYbvDeK6l7liKWgVLTafNU9l7yiUiP36Royq3QGFg5AUVLdKcVoRI36IPl292QbLU5wKHteqclTssoV4Z5IycFLjLlP6ic6U3eeYpvwL5ahDG7vQxMwUuXOxQIL0pNNQ0kSxlMuV7zO8ev45sd5c8UCnqUHpkazvuxjAMnI3924bnGw7WKDKlqpXixehtc1dG/KI0jkDUjjZKtoYdokO5n1Isq7JEwkfRHHQRIqFlw55NdnjRMO+YtUXH9/Fh+g6uN8XM/y5pFgozbytWprOiOfuyIBNnYTPlZDJMp/MCAPgN2V5Y9LG+YvAkHscctX96gJ4CTc7uiYXJMjejGTLTUwLnQkfWQAFJ3hFi1QwOqcoEKy6JhjZi7VKP2TWfSA+Qlc07OUt4+4w0USYhORIOdy2HkpWtNEOi/ck2Lh+ss69fyxLe477+dXN03+qHGW1RfYiDRaYPgJ1fV7l2gItnS5InnMuH5Z7HC0qh8IsCaCE2pCojeycraIc76kkM9dnNQ/+5+6LIoBDVh5xYxmza4Hbor85+19UzjX9cq25vY8RuaK0i2L4AsYXDCoMkiCxiTG4NsDs8t12G5PJuNJ6t1w53QGb3OnuOpV12vozlRSVAUgR5B2mpUT5LfqT95NXzCudMKdddJ6/965RkxP6dZ9gPYZ087V1pTrmlVK0FEXr7SY3hjYsJ2gdSm5gRHNxTFU5GrLmZVA7IK0gZnmtPJkuCKeHieIbDwM8Sw8pDnZN8epz3AaOzkgEwU0ijGWmKwPUo8/aaruY5n/k0js2SuKvcWEr1TaidfjLPC23Htg+ijlnpReBTyWD9tWwNvH1/sfs46UNf74TmTiDlbi9WCrFm/PqvBau9g5KWfzn+OvF5p7GHd3wbmEEgS6vxnFW8evAdzIP5iGbOfMId9PxfoIdzMsVl1aiZnH0opqJJSOL8tCHq8Y4XIXWebRrtcEZljh9CEHcIEds1iQpGZ93eRQC18wE79sH2tMH3Fn5XoxT7u9hcCA2UmFRiuwKsiwRtRKDblUigJNUIjwU0XKY3p03tLKhgBvhbzuYYpQAJUjIEWl9RvGkivzujuGMZTLw0lWdJ+LCqT/zQXpQlPOeZo4SvEeVYLQ/LWPL3a2XF5DvdZ8v00gNS0FQ6xKxqgg1uXZBMUWLsItF61ytC3TVg/W5jwUuCWKBBNzJPltUjcGfjyGTGjl83fnBm1o8SLGQT6ypcnlbclXWT1WDDIMEplAFYkuv834n8If3xdW6h0aHzrdZenBYHJcKHfxHAJXcUUezVmcXGnQyo4r8qXMkbuebeEm2sycw6nYwFBHERXgfh3nlmu+IcQ4dN81yOiEkjmUrprRUN7qn2r3E7Ob2BtJ9KmBiuH0pUvGMy8a8ZxUPwezRRHgutxryIodC1KWZL/QGw5v3POocpnAyK7HJIiYvklXh+Xrg9uYDRS8XL6fG/TQfYQV4wCJMZ8ie8CIeN41izuE8TsYWfisRpKg/7LdfIcGiYffKiGg0EpljG6N0InxQUXs7rNdgNqmub6mIxuxAfBI6GXnes9JRR49a8sk52kHQZe3wTciKhbaeJ7W5Tw==
`pragma protect end_data_block
`pragma protect digest_block
e0aecb5f74f8e43b39b27bf858b0e904a3459110052f28ce6af0a7e6f75cc84e
`pragma protect end_digest_block
`pragma protect end_protected
