`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
l60AeIGvufHAdfm7LvyS0Jnpokflz5rBrKPzaviEJYckL/M4gWYrBqt6nMvna//jIK1bOLtDE62a/NS6OVq0wSn3HbOhNwrwo+l3AEX+K3tSotbDW3rGzsP0XlUsrYvsxjx+Uc+ohDbhCS1O2fliHIMgFCzw5GP8guK0V7xpShORXp+D3oDDk2nPgd72/j620rta1cWWIeXVzO2BM1eTjQPXXjZR0V5NBXh97CA4PIUhQPev6fY+QD01I3ARgxsLAhjahG8FodWSf4S1qtu9D2Tw6LCh1QpmV/gRiEQ0LX58m/uXQzztjWQnJ6ubWJZEzfY2lRyD9AP0yJ+o5/Wl9ntqh8wmSS2WgKZ8cyt3zy2P5Nl9O5cnKGyMihucf/gDWD7noCUj79p5jyLOJidHr/aUi0kP6oTnSxgafAlMHdGfnv67oGR3HGnXbbN2yT0uVA6XvLgZpacAEjDPCagUASg6Nlz24B0msezU0s9ywsrxX88HfUaWxQEFpLWxhGeoP+LN89zbpSPtkBERpIlrQsADUPvUU4tpqznMdt9jJzAysBDWPxW0MkUl5twmPSS56cB3hkSfXbagQbqf9SgzLDZumg9StKc6XQ2a+c3C9B4goDMpzzY2ivnzC4k6VtdZNY/JW4hJkuEcs8bLy6ZUuKS5Nst+59VyMrEGJLKtyNNMFJjxJzdrDcQU9a9ocxUoMzWLHG8N6fQrOU5OHErOdvFfJombRhV9z5uQRK3+vjkW86XtF55N8qw/mThaToIp+ff8n8qc1T+KEoEheP+XE+4Qfhd3OJq8Cxz2rYgvR8kP6WAdClckPdxnHutesa9vn+AFxhMuj5zIjBe5Z0m1rrZ5MzFNo1MGTjPeq6VYQSSFDWVY4b0PkLyILi8USwkefIQO3Ln3oD7vTU9991fK26VMfcNMihfJ9qAMMdy7FVvPOGMLLl4rrVeXhVPhN83/Abm72am/kIkIZyoWhS43FhX6b0e+H8C8jIVV4C5R91ikaPXFtcij9CjPCfFE/TgHNDuIuz9wSp+iolfae5t0JHS1oD3/i/ZKqluku/JsdTIyz3BE9kopSeb3j4jEVC7AmNKPShRsWI6apa0ZcFWRpyauL4wdpWxi1RhRY/EGxppZ/MwQmageeOWKHiOEZO/4ryjl7jGjCeU60WsZE7UBt/K1VijfhqsjbCc+MJRBvR7ogIujDKlIjVzW4cmPodF8HPrrStRj6UrMB5ei7rqnxymbKVIWQmUg+9hn+aBbBpcV1r8q9waCuam74lD89uNB1dzTbBaWrG0F73i7fTzX1Xt2uW5DqXTwzsqTCCwUx4RME40X2CNEPO+4qKPxFxloO5YuMOzwtX4rR2AHPpI+q2rZoJOf/cdDvGcsRAYD9UOj+/iLO2bgVJAkkI2w5kuEWM+jHYswyQ2JWelWRyqxiL0lP7AYb9PbDwRpS5PjNwI=
`pragma protect end_data_block
`pragma protect digest_block
98d7f0859b089e5f62775d2867f2b69ca3427693f962b718b156fd4cf7497033
`pragma protect end_digest_block
`pragma protect end_protected
