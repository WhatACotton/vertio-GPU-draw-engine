`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
xau4FKkIKevZSncMPeUPkPmbMr3QDSX9m13VBsih55j7wPPGwGrf1fE6sMXWgounV7YxTEJiml7Dx9AjB+JV0rDNByNmoapnUG920yc48AgCDQ8MhIZwOyrSyN8dmKmf6+0qM9hnMFTDVDi0bz76f/Q23i2CkNXlDS+YD7ZRH1a6HNJXpo0j1a+kHsr11R60EJQYtefhbuO0a4Kj8Rx1Ik9ctL1CH0XH6wDD0Tb5mb+RlCIVQ9AxNPsYBP7tOS4Sv86bT13RctUngVBLMgXOcPc7krnM9x2NiVGlB5X5442OWTh3IYBixpp/MEsBQwVY6CnZdIyXl/qxYtri/NVVHTJ7sL6JDlbohdDOcg8G2PM+Woih0sGKXTQ5KEWbJaiOLAFeF6ej372+PejFGyENPIv6+FGZOIHfplvCAIX1hKo9eTctQkO2rx5P9L95fMfQzCxNgq6Zu+X7J9tj4OraEPkUK31LDYjsyyH7/kxtCdR+MdjlNfCrRjfqnCG1dQFZ4IdyWInRwMmasz8SkIepptOFaNkg6/swXTRTtisbpTZKmZC6ANTXOFYWD9ddQwdGmlktX9LLFd1k52mcDfezlZX/WQcwWy2CtxzUkOkRHfMSfY8jA7NS3dxgrNC6Wc52+LOVntAoq6vMK2gQWFE628Uy8WdWJQbCp8HY8TEFVB7+YLrWW5Tmrc4BIfDzxBvOqhjvA2rWS+TTvHm9QeFch7+HMBn0zOCgEPurq5HXvjruai142Mi1ioMz/98tvxypNZZYzyApsCQucUS+UbEp1GCl1q+zqG0G1TNuI+ewMWTSwfnihBci4LZbDd0DXjXwCpfYNMdnBvjArOD88jBRXyI8Za4f/NRFj6jgDj0xbgDZyfA0vVXqcuL0ik+7kbEsZ8SGz3pT/ruTwJ9uyF9j20IJaFq7/roQhAQNA8l9AMb9Y3ZBs8TDK4B7UYroDt5m+YWzl+49PoKa/IR/Xc0enD0BLyTm7K7VED3KP2p3v7IfQCs2db1epadI6PGqVN/OZAYK21Y8Cj3VQ9KzX803ahSghTNgZtdfaAhufZK45qYVTZQp7WGekpvUFr03EPGH2SjSmk4P+lHzsBH8O2lttAkHNs259BK8IkTb7uQqHXE64WW+BlknvB4QARZGqgsGSeyGJxTaazl9amDB8H2NNMZUVEX0GzTIDTzQl1PHcf84lpNAC9h1hmipn4a1LXDM+XS/CYL9pakPWMv1i3zVbWqqKh1BLxvhxR5kMOR/E6QqwQJZusixGotvHkWIL38ZlDAhjKDGAV5pvLanBaKB82yjkaFEmbj19NchwgVZcfj+0ZpW7yim0naMRKccbFQN5l7FLveaHA69cZW0jPdiRM5IV2HiIHoTQXQ9GP27um5OLOb1+oy2MlfdHiBYTnv2hMf3jIrOedJMIEXjELUzce4DQCmWYxYhiQCyaKFJ7BnP5awdk2OW6GiIpy8WDF8whkUnKc7GJJWeOaG+Z0PJ0W1BeoTLprZ9xOxUD1EfXCLa/fo4y31B2ciPHKenYd9o7EtWhBiB4UdDRXDG6dDCWP+fpAe5XhOjEynlD+DNMxjdgvyEMSJrZJh1jO+Qt5vHYU95WWDm7o09zLicXnvAC5HrsRNFDkmPLYZlHPIZcDreGoTjNsJc2elfxYQqNCkuTnF2EViV69dHP8sbXf+hwOag0fPPXc/1o2Y8DMoVuTfj/qo5EM+AncvwPS+voBYuj1DBiCrEOc51XWz6WoiCdTNUfC9W2kQQhR6ROVNPg7Y9tbyKIUY9nkMlfg0wcKK7beIwNwswuhOGFqX2kR70AlubQJIUI7amfC4JtRwdQz5u7g9gHOxZGclIbRnAcx+sq3776v2EJcASCuYGjg3Jc3nHZtTPds6CDymZ5RXzgJtMty0btjFExMprnsxSJvXwalK+ZgZn+iqsJDrYLJGG1PS2+RORgkI8V1t4C9qFOkl7IjD2OAM86mSFwahC+7o3W1qRD3lfABuvTRHY3uSSpWQF5OgoL985dcpvo6ooiiRyIGR/GGe9tRELaid+WVw0kytRm+BISbtdYW/VkK9hBXSgmuu1o9voPBvdE9aKK3kZQiRYrQTFU+JACrjNpZWZ+DOsnWUhWOvgvxQ3PmSvrledUuw9KeOx20FDQjHvLQSOSZfDU5LoqPA187CUaVxoE0OK6FIm6Nr3A8W+EqpC8Lewb6atYStDlfZJqfxQkhE0G0/U0Etyux1Wd7vEhmJPC1BoflG5CIFMGrgFMjrGcsckFI6LmNBiPOAwi7sW6Q8vfoHOmMM5sgXqaiabwm3+lWQ2u8QgeGYPMSQlmfCiDvvrVZNWJ8OSR5wmYMfgLCCefbai+YsThLBQehMIJ1Zx96QlwV3y4yKjwvnwJ0HC0OHNPexMDlDO/189j8fJ3pXel7UGfyIsm/d2DBUZoZoQFurP3yJ734iGeCHeMgIj03dJfMIybNSLELVHrBsb9m/0RPzHBHCulA+kVnzR545K8xQu5FJ2YqfqLEYddhYxtCJrKKRfpH2vxOeVOwlU4pzg/HRjt6i4JX49zSkxNTNg91jAjqARe2vV3Fi8GlSu6F8oDKOJUp5sDLjFZwQOSBlNNixYdqLHTMXaR8IPeFqmqdPqFCA031B73exvh+316GAc7evHVAHJs9SxQD3I7nPZ0zdFTIi/LtvajTrAYwppK2tWor+FlnY18e/qVsK9D5aONhB/p2/0Hr00ypAsqMCxEDCM4aXm+PGOVrtZLaAh3kg0atxhJVZhT4hjGJ/lC+CpGromPz1CaAs9x0LImPAm6EM2XZhsW5S9dQS0P6rcM9LKNnuh70jEpdyHEn7XX181bXePDIEuHtBrW63+GW5AU1Np355MeEXxpWb3047MplzPZpmc5vaDAVeBSC7cbqiz9LWZ1Mf8xXM9EzSC/zSImO+hdBYr9H5bvYzRG9IiIoyn9XGv7jg4OqsczDUO/q4DQWmKE/42sW5IP+D7ZDlf2UC2w8Sjbx9piZ/Zvp4MHqC9G7EYRixeXmithKX4rQitxNlvin5yE4HgrdiqL7OLHza+hjxCwosvtZVS0uJX1ew/0KL9+69MWXPPDBnpICAuxXWIwcp57IhMSSMuzsZja79HC4dc15DTHOqD3taIk7HKCHXO/4/+LcMF/7pgrPhRslZ+teyXkS/NF209a02v47LOsi2oGaGeeO1yqwg5KT0adP5jpdOVfv1qsqYgcckF5WTclQYN/hzZYDYxFi+L9XDCcsWp7CMKavTTzff+RiBQ7xlznQoRhwsmQuA+U3O2Un75Dw4XbcQ/vGCOOA6ymm/sKnQ5PzGKv40E/1pplxtRwd29U5z/benq4jJMoAX1JmcYRRIH3//CHtNKBpg6yhaM7P/YYQLAUrbBR8iWd75a6nHBTp7CrFkqZdw4hLt9hEAu8iXXhun9lXQPj7PWmBxIFrdLIyaDGde2NVTo7MedUKau/dt9mVrwQgYmkvuR8nS7t/3kNaW/NMCPOPNcPxMZa8B6/7iC+OKFYuUBUonhIKK97FiZAz8jaK6/L4aEA80xrQWNSJ97nhwXSWHa/3Hm8fca4dYrzgQVJiF8EWh2msM6JewTUzAJbvPRx9YFXxH45wq6Z53Sh/KQCT/KrxD6rMr0tsQxvsaW0Gqew2fto0L1Q4gRsZCy0qegQvcTqoUjEHJKZf+dSQfsjJWeg5FKGRMIU064dQyRLAGZfPpo7xqjk+0j6jfdX9JYHP+ZsCA3HG2od8lwaufwoX9ip6tuuwsHIM2vfnrG1e8C8ml5A+z7az5X9VGF91dJZ2jDQ6oiuTfPY1mecg2voLYJ8GIJQCxOFFhLm5pGC/A5O1P4+NeyXN1x8Nv4nwo8YrL6PP/r3JsLYxXTJcXl9TRoJJ6bMAMIzj/xB5UwC7UxSAxNFIoakpL0WI/PNpaJbeR8tIL6Ci+FeEl+mjs1EUY2HVG8BijXojlwQMA0ZxeeQnHMdoWO5dNWJC+0n/AusDIGVcYR2hx9lmsaCqtGman587zboiRvWa0re4HgiTLwZWQpkCQEDh8pK5OeX+IZE1DJJw47Dkf/igLjd3HfcDZXg9othfd3LeaRb0EmPa91xxtRq0z92le44KlTZllCk1La5JiWc+hDjXw/sovgWI2ZlRcXLUIhnkuoMDmKpPcMl5Z7e4cjgNXIIUr8EKiW4D0hcend+OIs+oiDVqb6zWRUGxH+QXbiL54Ehs1k/wp7l1hFbsJJ8OO9F9+sC9B+iMXM4mAhdSB+Df4M9vDB71iaNEPgAjT5rN+Kz5DQhE/vJ48w+7UEoxfo1d45Ka96SIO4SgnTp50ATw8gA+v80Ts6DiaQevIqJEIm7FDN8aJM0BHiWm7nBFS7Uf6ZrAjYaW6j4OAmRCWS4uQjbxTkqQK6S1WWstzX8wj2HfDLNIJW5R/bVNhljM0B5v13/7GVRc85pU0xqATjDnCAjzwgwS4K7Xm+HB1UWy8WAY3vUrucasnNs3lvGkWdObE8LBrsM3CUXTKfHRBJ2oJMf4fsdYLLWQD9D2V8+SwCvnjXz767vi7iDO+9UFFbSwcinjzRmUd1gfhVQyLqKDtCG5m8rIlIzsInk3FtpSPV+R1EAjpVlluI5ZgT210uxEsTbF0U2IdZ894tWMY+iVyAtNig6ECS+WA8y9uVatTkcQoIQZlmZW95QTjJUpwcLwmOb722vdHWgThTNZAJVGmMwF0KNqi7TGShsyhXASZVfWzN4K+JvDm0ar0+t92q8eDL3xNd9W7m8heOX32V+mdHMfogAxMDDkm1eM/AyfNu9aQ83Vjk/QVqynjHztmccNwaRW1+pP3s3fgaa5rgIZBhnexCcHW9vA7/YqwNF3y7SYRXKDSH8kg8D9UpZukqv1acZn2mSkfgOozK54gPqvS0K15buS3ex5ohIG/dSgZcMEq8s1D9411npum18i1lLna3+x0Dwuq/FDnFYtSb/tA3S2mmZVnOvnW0k3a01nid0fe31kNBykMbPClG1uDfn5U6d4Kjm0wxSQO+eq/S3cJbowSjmuqDvoQE6abpPLwrvozTUZyKnFb+a1T6BY4ve8xTz9z38Muv2/LG1v4G11WMCc9NWBVGWocA3IuOnNK86FdcQaNSWAciU2yZMMeED8yOnW+gm7uUYwY+9qgSaDX4FmfXmTsou5FuWgnWbTQeaBWDh14DCNeGZHrviO2K/E1LfHpE92ICwCJEz9YpVtGmeNW+bAdpdl5I7+Z2U6vLAXPMsCsgkA/8nl4SnxBXrVVfLUQRH1OHvwUYy6KIeDivWZSWI18I1T1HRq3of/h9oPniJttaa1GQinH0nqFqkCMO9nFG/p23FbXGUOSPN9t+omWGlms6agsFYUUDn7bT7KQMEtqtLgy6Si1YCB164J/6Qr08LNtw981wOVtymftJ+z0vQta2CsnCk7/NuuT2Un/Ni+gCUYEmnim3jzeibigsqK+9wwM6fbnU9kuiMq9zwMCZg22TSxqxRL07z0cU8ze2binXo/wRrCiw95hulifLU/N7gzJwsY0ecF0OXLt35Dv3Hq7FHCZSKADPvw1ebgpddx8mcwjmD/WvKRivjxoyq9IHeT3QO2Uqsj3yU91oH1iPj082nnrAgfv1Cs2FpKMP1UWzjHtzV+Ylc7qFglkNK4YTwNEIWNH+KQryzjLnO3ZC+ZVmOcFbSs1BPL7EpdTQyrmE8VCHmqYzLXckUxhYNWmMyQu/dilogpuk+j7eMFAcg9iJQ2c1yqQv1DaPHYnPMhIKeAKJzNQs2FspTLivQEUJX1Nw86uSUhUuCEQ5G+6wvnpl9mSY2PxV+VLT/L17DXYsdacjAHmgxMaviB3H7bO1r3j9kpxlENooamBZrOaI3CtSFHLUEZsI+wdI12OJjzhNBrmmc2LGG7zUvBZ7cHGeAt97BIPP3z75rrQTLTWGD8DlI6YP4+3Wd2CP66PjGxYD1Igcq6kS4zUZQVecgReo5Tb5rNc7KXipftLq0AkU/IiDtztqoLDiYONFOgo2cKGpWMy191W5YNEl+21/6i/MU51/n50w0rZ8Oe3TYhUDnB0xShELCwZn8osbElG5xLdQ14SVN4uAkl5hDxUCGiierNYqzpzwmGn56bawvA8/iK3RO3iwUN1jltCHVFdtzY6+uBZCzhLDI25w4gxiI+M5jUhDoYzn8nyAJ1pn8XWjL0Mg2PMrKPB1q8ZpxLg8pRdVJxotVujwi9aih7qlIEQwYKuYN/dg5Zb+Ku0WK3o0wSgRD49D9lIaPBKEQxC+sboCkljQFvhM8fajXywZTtFAG4jdbj3cReImxGR7VSb5ddRVu6FNBbo3Rkpy/e7SK7pLYbzplddnIR/pxJoiSeboFWdB1dsBPSpSkA0NvQw4ITmwsqsbX6uPkS+IpDu1v17Bsa/nPJQ/y/It6kxZgKngeLPHtuVmmlUNcpalI5K9WYcePlVJQ0v5nD1ML98h/rrt+LcPZbZApZHSsoM7EsaQQLh8XTPdQCYrhFzJY4Rbfq4pSuOPEgLl/afCwSUt0yxSLS9i0Do2naGafTLnDY3TtTqoDx27rwN/sn45YWTUX8a8mQfyio9+IpZEBt+PuUmHfyZu4auwyG4xCpyMfK99yQY8fqYd2Y31OF+3EDmP3zSsD3+hhF8Zzkh8yL4fUeg+uEhnMmZ5lKI/DZuK+oy6vQApvRtt4P0AQvBsp3kz7COqnrJ72LrddrnYrfJitrg3oI2jqzomToreAMhqa/eKfMNZl4TKbGOz2jTcfTTUcPpt/kCb1IIqigCS1i+kVOYRYqYLsp/1LcBkYbVZTU3tANXNYmk912GHCO0iHFDGm2Ej9qyWSvhXy22Usa5S2gNe3zSHTJK4gHjmWUtkSCNDJv9wYruXrTvLNr3Jbi8Q/vSZk8NF1OvNMpJC88zDvXgq+gO2n99JRTi/tDGWs/jifNuN8PLCvIPtgQotqMKtPynnx4XH5ztWKmG5ss1uD24QkzsXJayj/UjTXL1HwwxxuS0TuIvACJGMEQtw8kw8122BVrJVC4MwxAXdZONOP1ZTzXnRKBaKAV+dKgLKQGuhjeJyLboWyO8OSNNH3DRTse/im71c42L8LNMYSAu6Ki2aMH3jz5J+XNGta7188hh1Q+zIe5Cx+ddl1HGKOJ1WJg7IsK3coHTSbbDm7+h+b4tvQ8P88Hkf5iCIN4CbrDrEmajB13OIHM/8RCEXscJKe0RkhdBPt5iQrj6xOoyFYGDM2UC4OyktsL9sPA9/4meMFQI3vWpwinevo3Zyy2n43rMo9v8n1VeM3N1eLQz4IokOrw3yIr9AOpsqBpMyKH7o2j/u9ueB394/2Gp9UWTFTOAbn85mR1myu6JauW8/zJsTlYSjSyp9ur7NmiwldSDuP2K2CgkoZPqsJSYNuwmJnVfCaCHnkbjNYPyO2Lp7m5497w4mIdnoFgk/QMUdfg8xrMYtRSDQhBPK/fCWklmigQruAk7jRwl0y4E89Wta3IgKiS/Zy5AcDQ1uY86szyaG6arVYD1peXM6pEh8AKuMGrKh6g80GnXIa94wH+yFNZStwxMCrC/DCyZO9PK6adCHo0NFNb4G0SJ1cH6V+r81jf6W7+UFhY8onIzCiHr5Eii9vAHLoCV3EGXQOTqnW9clZvn2wV8gCfsjSQAsB+PhKECemwIrJqe4rXnoiAHbKUz98y7ZlN/ivKhFpsNvmvOZyHesR2bpWE17Z1LWyufQ4XJj9PuiDj+8H1U1VxVVpHLE3OM8MB4ig4Cc02RpiRwMER0+aH2nuusCgmDYkm2PLEovtO9ePgnpwHlmfhcth5FBYp2nsR6uie61RSwMVqeJ5RndOs+GgQpaQs/QfTJhu1zUGBQLsFDuYVSfikWTlpsc27BAthq+gCMVGZa7g1EKTcRk+6vLPwDwz8sIiCsCOknX8UyYgJaQecooT/b+KevzZNRPW4MW4dCegEZEf7xseGkboze1/BO/0xIFSFdF37YiOhoSuUaZwt2RV8uf5bMiAsclwWjDnxaQdbJqodSF9QYN/2gf0SpQYOL+/mXo/YjGRAqHdX//AQZQ9oMyEsTj47FyyqQDWP4I7eKj194D8IbpKq+NU5USWTr4vjK/5JRHxGe/ThDzA+1PEvPj/n0keKmi8UM7K0a9VekojliZC4wIOTkilZWhH4/kxf3HPGzuR5c7zQIBuYmnpRLsrYHKpVHSqrHcguJ1twOMYBxgFmA1TK7Ct8BejwhNWqmpsmLz1sWrBpOH+jhRz90dqTVwrCENimTLqn6Mtx7yiseTzWPOrMw67zrI9aediXeFdKYCfvIaeJbxSNw1Cuyip/fwo+mspoByFUK/AXk3WZlWY71VJ9bQgZ/63eNo0Mz7xDCbFYqY/Nxmt7Ut/K5Prw3jGhA0K/FRIAggXovb03lHpw6oOT0u7af/T/kYyNpr/7x8k+6xTLuHFaIGK/tS02sSJ6f1ZMcmk3uztdPjiBNCwa+vbw2daFahRLYXSp+ezb/hForuP2LGdbqikd4ZbBTmc9UOHXjt4mKneOEQmJthJtpBVpgXzyS9x6x99rh2QWNggTWp3u4ZKmF8t57ojbhgHszujN5A52UvbANLJliVVpeeIV6CTW/uQIzSeIjaiLRvwavSz+6r5xp080ocQ1Er+7DSZ7TEeTGecJFI8Ad9ajCyTuyj6Md14ibcac6nQkkC2KkWpBzUEwITvGj+sQ43D/lgrn+DVZfP3Mgtm+vj0h5BzDIfEMtcDt4tRXaVCdEmc3/R7Ou+M1ytFXI+AJdUBeKsifEi2Ie+IH3Dw+4XlcDooFBW9QDTJTHXg1KpaPs1ofQQsNUXqGicgKLdqeC5VGet9131qOpBjUkozvVdPMfLdXpGkqdrYOhPofR+f/Y04pHhc18pf1P2cD3/PvvAs1Nbgq2mmntfD/oLIHINVbN/G/q9lmSdM8Aoy6G9UUFypF5ZhQzqBswoDIYLZTxwPyW6nBYTgZzUoF5Z7WAKzvQYLZ5ShZiSThnGQ+5db9uHJSgkIhkSF7FWtLQz6uPCIfJiwntgPRiPo7nh9uFyQlDZ87f9plUWKdDXge+PeOs/czR3xR/RTkepS+NPx9KCO0HFPjF3M/QdJWLRkXfpaMiCxyiZBfiEfquZZdCv4hv22qBDJis9SXgGngy+SceJXpHV4B7fuc9q7RjKmiFy3aIoORNaIdUof//1bt42KKCYZQZVRKXYLi5nwwTqn2CX7ocuR1o7T8O1wm4lyXCZz/T5F2TjSFY0k3vyD6makdr7aOvg+X6I3ejVXAhWCU6b4I0DynRRle60fWb8FPZddpHTFhN/eYiM4V0Rl0qwb46n/VjiqNrHCRXTm4Jh+RulhzyiSkdcvHfSuQ67k7aPfTqDdaILEhLuh8GShJWjvue+PfJfd0cLB+GPyuB05WhdQy0ou5ktxEyaeTZ0Ubg7n+F0+ZI1seODiDda6CDogtJIVQCRFI4CZHA1ej4N3amVi8M7oFm/x6YIVLz7WYseGxR+jjBvb4WFkp3mrSt8u1Qbkoo34/8TX4bjxBXOW2wz+HrQZtW0RttFqnegOuIkD0mAdFw0mgnI+PqUuG0X501q1zVQJqX8XpwqRGVQ6JXTq9N/c+rTle8XwfCjud3awwt58VCJwptgmk05ccoCub21LVmrqrA0i0PMe0W6nQrO00m0UaSIaXg+omj8VVr92nzT9OyEISEDvP4XA7jRxIHcI9egePb+6ZjCYtFYJy8uIpstWmDmEmR1lvMhv12e/uyxescFz8uduRjwv8GvAUEI8IiLcZjmEpJSxMN0cGfHwllEmQXGTEczvPYqC7szO0dAMMIK0oNXG4HbbQHPg5SaSjhHmODg6rb6bWc8U0p9O4DpAYXJVPuveDlerYB55LbaOm28B3eobsWBGGpHs35pGY46KE1ZskE4uA6C6JZlz7Yw2FgLBHRoXBatCwYwAG7sqYOjQ/yfFpvU6tX19lujOzjfbCtMUMGVfRHRSEFWVI8NcZBtBlow89VyFLxc2k+u3gxDhJPNcbF9xnw1KYAXNULygkJw3CZ/gShjXgptKRhP/a3cAHvI6beo7NNkckkS+th4IrbsBknUxonqnAOIijgf9AKaZm8B7xa6FCqSX5GMh2EH19txAe2OJh5L/NqBceAO8oCGSG+B8YmCMYMdahvdFmbDupvhp5WPtH1TUOy4qjWTOliwktDxpe2pfBc/a9zkmLuF4vdU0sHZPo6kh48ALaZD9ewZtqsLewIm1tnsXq4dasHH7gC7IxDDGvd+ITBZbJ1jMxYRxsDouNv5JWiQEX9fJWnY8YGRccQWLEZICmzFQ+9EDC4zmx464qMoOpq6vJy+kPjh2BFDnU/xgbV2Dku6Gz3oExCYzc4eo2ZC1i5Hq6YNNiiejMozXXQgsvYckLgSvvWfOKcM62REiilxo5yiqlvzotOLu7VJVao2LtxS12vMM0Zi6vrOqTlzBmE/OjzudU9Du+/mevwHi08gq8EyYZWulGWv49wFWrmS+IjrtgFdFSNzwHxVzG4umv2JP6jhUMq++JJh6JKWHEXSzFaiDTK4f6cPHcoFZhLIChHSKl0NvaaQnaVNuPblr5Rq0cP11CpaSYt992OmZHiWyviZ0Z6G7TduXpJtZXfm4ejiQo+C8EW9nXo0PLsE0OwUSnq4TvvnjT4o60/NecMqIsipJ7C2JtJh6rcRGsttLJxqRhdx7gmzVsojsop1G2TUqWu/IfC/rjz7WnsHYsim8hyYGyNqA+SMxK9vdSKCiEu7wHeaVpFaGOM/6jOO1wf7fo1AQQ0xVHZr5oNC3SMaRre/8KmmZhficqOCbvJZzAJIn8+wB4OXFbonOKAQ7BlpQWxzMCsBNj1m6TswlxG6XusDhr5Ag+pR+VleeMUc9Hph8lsjylsi8mWO+S+p4l7XB64jeVDVmfEsW7whXwhlr2LnsyJNNykC/1MEjzI9wbHWrxplXgCi/JdZ95VFvXYz8lFQDYbnXqqv4QRft1pLxGTekckVkcDz6hNjkjL+2kazem6TMhTTt351uTfPdE1nxpdW1YNHzs+uEV5D9im8PhFFyBgfODePlmei3yXkLxlBxX/f2Pxp8mill0WM0jXa4XI++y7fH4EmMOVsbMgVFq5d9E8o5XkgYPkhusfPJiQkdl5/9z55/VZRHEnCklnc7djpDSOJi6/CxhzzbvrxaFebMcJKU+9zxR4eihzUndzoeKoQB4Xuu81eAnKPsuspWpPJ9YznVRWUzLsBXLelFkVVLFfWJaTgYxIxEY7XUB1/0x7tTwPKZnvFJvR6FL5kJMzuNYtp/Hbp65PTURmn4hT/wEK1LKvHpZDlAG+pgUWzV2ODmETy3H+xln34+mcK8Bet+wsCQaLJEwcj1yYurvokaQt9ZGsUptPQ7jftgeV7AcCNFTli0AEEnFBvOdGmnNaX+pu8uF7OJnvSp0h4BXwIM0z8ket6SGL2m1cuc5gTR0Qz2Mi7yk26M0iWOkKoIKGde8JsZ/EPUfWsOwkAeT3ae5a3QJZiPsxsXhkSERVmwYEvoomGPfYO6ClcYmyiLX/qEEd5zC+6udmPC2Zx4ib5mVweRcfz6/IazYVhX8E0iUgSEa6FwawqyiDdytNw7G99cXXCjIEA/yHCgNeEnICnbEZS06LeMILBMdj96sKTNk7OYrrQLPrayjPqlBlGE1KItWvcJ0eFcPRDM4wG697lRgbf2J+rAK+xQMVbZo5T9AphBB4vzzirjsVE2XRreB2z0pDny4r8DJOpEoO7HtduriSe4k/dwDPWN71l4c9BR9N3mnDHMK36okVodLmKc7yvXWopB3/zYap/AGXPcnaIc/qGDjPkj2WoeQy5xO/jeboCzGXQJZoyYFdPy8pexTmOBPG8SHJtjcpXRWL4M+KO+IfY+W+xzb4Q4KjfKZBlhvIeyoR8/xiBRS0t+CM/vj82gaXwig/ynQYxKhQtKDKLCpLjyhIksHuZjSkrFd4ihoLBygbz9CveqBExgWgM8BPWlBAjP/a5+SqQDxMz6S/wB9c/1pCg/wmAr9PfkSJ93A8h3Ekt8Jqi54ExoefJqicv88yM+dioIzZJM4veaLMDDIaXBOMiIdCYA/E4FDnBZcY47xTy5j2VZwP2BbiuGHI6snDTsId2gq6JCm7U7GIgOS60uyvZ01cUurM8H0C9EwQojgqby2ZP/Nqv/c+NcDtbiiOQ593+FKyh70I8YIRlAns6kICzr6cEAOB/Fp8TfFtCsOeFu6Ondth81h1gVTjpHlAaWUCie3HCyaMbj5JDqAOEOEkXDGuOz8hOFIJ9aJ/eY0RES7g0gLtxxJtEXYdkWTFqUJgHvxvfzIz5sHEZm8Ynadiu7J8CS1IQOpe58bzxgtThmpZ0Usp23/JjX65c37RbKoWyo6FYNKcwx/4uXSomaA0Cy+mfuSyht68Iaj4mHyNjVfCFvXwMvUXsmx7B5r7KrHjRt2WCXPoomV3rqWvoCyYzA3cG/pr4bjT37NIFTlTWTwZoatAq+J0SRORZyVrRDA/dNNQqQYFcCUlvTiShVDCWU8zUyHPKAPGFcGoB9e8eN6QjiGjhej0DmqIFBsbCyaPqvZqYdqHVnXKpUQjG5hL+uhXwEXOx1MWBkF6h+iIa9EbI4hvMM+vVl3Gz36su6L1vU5FP2iqqRMEkpBcdbPqe38pmXRUhX5Z3+O1/e/VBSBQe/PyeXdl5orceEESBySaak/1cWtxhDFc+g/16cUdnWcOvZHNE4WzkFrHhJHE99BO531kUJaGOsQoBqVyy0Q1/JuigZe7qZ96c2L4H5pcdBUfrWUzZFu2cjLrHRpqQwqtButSx9ofFWg2sZsY8adEoJulGVs3BuhGn/k3tA99SM8WnMn3yH/X9XhBI/qFmPLkEHrfxKsOhI5WaPNm64L2Qxsk8dJ48kIedR4JI8xTECkf7dSoP0KRLXlqht5vvlM2+rEPYO1K8MlJMgLjkZtklzKL4x0hW8KEmTJjZUAMeHvncNzXIgh8aXHKKvvIpui5eHmTwzFxRBHwIwHxW61ndyUJR0kGM/X3LCDNo9NIYGqwr7YVAWwRWT1uvFeJsNJxEHuC9hznfhRS5EjjC7KVioBZs2VK/dehbEqUUaVw1Euzknqu7po3A47N8ltJJziF1YudXhsjGfEQbWjY9sgZRqNc0fC+azm6oSuJVwqGffMvgVaBCSaFFHlD+0za8+csJ2QiiY/WmUB6nFxe4UFLu/pXTMC5/jz4NkUojcJZXmkWM4AIUFbM94RuJtF9cSq5zj7kaTvxYWlgr10aeQKdJooJ0PmpQDGwiY/LcnaQyszn8/TPD2+3UMjgLZyfskdofT8zmpWyp5tdySx6M4UVuwexvdBCz/+uJlB8OvHfQxDkkBHvdleIRqbsZ56kMR810Opw1LFXWSOwq6K0sxaxfmvHT9gWAda/U4HZQZz9ElfabEKgKXl/PomVKQ57t7SxZq+nbVgXoi31Nqcdd+v2OJy7a2kDkMs3yrYM8/6p3lC6PVPPlKl3mC3V2iDL072HK5jT3HVx8MntF5PtYKxY5SrVb05DYyZSo30Hrn0PC8UVHLvtnk/UekF/XEp3xkGLIYWePeN6dLq+WjtQ0LcJddF40eGijguamNlc/oqpy0txU/vIKo0hOftygqzogakC81/V2JxOspSSbl2t/lxU6zeOLvWp33kG5xadEVD4QXlI9SW3U6Zu4nudTpqJ5RbXAgyzUQUU0stQCQJhe5cWRTG/+rObSd2XF+ch9YiJcUp3fq2aW3m2e7zxvkb68ST/1JjkWwvdRDl4bf50HGh0UYoL8U8NEYaAJ2g9KMfSDYy8QWKSMsbpR5FGcWTjmdkg5weEt8PToTRjC8qePRHn4TRMiSgAfJFS3Znfahou+MHB8rwaiMFsjb0+IB2m2Gxp+otAZZzpolXJ2Iuq0EJ7HKqeLw7wliNLAkVdMoVorAydyQ8fstGbHT2pImBea9PzueN4Qak8LXYiYCZOLueML5o9GWzJHdUY04Miy6woCpGyAclyOipWO9IsiRTM5nnigXsGTx0YERO7BiLY25qelgodBTAnFSp+meGrTqe4SmoW3COD3k7Sz6x/3xqppiYotT0OgEod71BDoUoDO7eKQ1rLn69EHdRdtY/kk4pOc+eVsLIPXtZb0yE4CUPeCHn4Jz/LkAGjV4kmV6imziOMI17qtZhSk78LOvTNhjdpyTEPKkXd4KgtY+9mbQxUspHrSDfFauCTjs3NzALVdjoITx+RXxj65yCk76OHpPOmNuY2PtN+vvLFNMvp32p4u227vt76yKGUV/8RdfMKHkkiGxJTM2a4AtYI1ctjcdBNKIU+gvR+8XaenR+gocynBqblGrwGtaTYHgSSxa0BIrvpsKIWFXx/EEREYVCVkjbvYK11S3axlF25a9w0l6/fjZcFLOQFggAohdNP2AI5XugCKartgOs/rIA9n4EClV1xuC05xbkRU5uy6LTVAFHwbqvnBwedt2E2maswnvd4H/sdQCTvgMt+q+BSYnrZreeuhkWqBT0xsJp3l+yKjuQyO141uo+oduO1+7X4TKNkDtL2hiFQjL9t9utvhH2oBp4Y81PsGTzQ4e7kZswSwOCA7rtvz3MX1XGxWO47d1+Tfl+wFMt4r0+TlPi0RO/KD2h/mQ2H3Sh9CpJgts9jaK4EL9FXfiBp12RP4QpPG5nXae42fvECHP9ltUBp/iMVliuTFaUAIok0Xxd5oJIWlpm97gewzQkOswxW1aDnmK5Of1KsvUjhR2tY+e1x75I/SS2V+BLPzJhEwpaHGqRHxVxFZMmmaH9Gs1IbEWrL9/Q5oQ1diXPV1Vg5sjdNpWCPoIWYBgmvd5nVnH++jsF4AvxCnRv4BpknGwaa1XkaoGHujnpJalwEtKsqhsEfRr96bABClWACj2yhjZ6oZggIbkvypp6YDrpmjqztfGEL64G7wpdmkwGrL5fXjHiz3x66rzUlEwJLOm32QHH7bKOhksKuppaLNHM6cFXR2d/c7ptxxXyLCjBCwbqgXEUNBaotHIqWXsnwl9j46ThlPdmeWWZXyFrkK5eFjTRFehPFMfX0Yasy6YJ7zWiKlQ6yYo0/dRRYi0lDX3bCOwI9LbU08S7ixjUclGPPTnDvSx9VbV/gNYdzstY698O4JniotTRy1uEl7q75Oeh/9Byb7QIux99WW7oRf21X1o6ZjSmPUhgNzC1GMcWpQpBkH4QIWmznysAS1iEjfR9+s7kWPgsjYsGQ6gn5dN6GHl0W1ZQas+jO58XsbJv5FggfWRBVbp4MsRWWtjl8+g1nunelmNzDh/xqF743nVPTGuvW8RMxsvq4+FVo1zuOnypxT63RXLM2J33sfxSYBow/QWs+8rY9TW10YR0AgTd6FBxX70Vm24cr+OBpB+jLBw7mTSDpPz1Ex+WE40P9zANZsOjnNrrIU8U4YzOgEYfUyKGvOSDrEEtWUdCuOPHrXCHivUVvQPClq5aOUlzQ3quvA7yjpnVCeMoeQKPbUdmcpKMN4dr2on2iTu9Ey1TGvG3sHMgG+/3GIVemIIJNDJjEFiXA69TtcKHUJ2CrvM8qkCAAI7Xv997VQ+34hXVutDwnR4FFI9X01mw1O540TbcEJeHLEeF6TEaDL3YLv3XqX1PvAecgFsB8K5T8odST1jtfr48Dlpk08kJ37w1HiX2BLwwo95SeWsqAmvHK4p3EhnU4fl3qWLxLdg6KzskdyAGzFnnCI9F83y3RJmIO4CzOKqQAn/BvYPFre3vsandSQ/YvYEuV1cShGnkP09UKnszu+DG/4x+OomIckPEM+wcALRr4Q3eajUiDVWqw2Vsin5ow1rW1PwrtC5DyWKA9XU/erRdfgMmhPEyCJ60tV5zbuEf4QPJFn8RITr0lN/6cVDbtRwCbUno1J0QV92pzkWDAabmQqU9sWeT1XeIK1s5jQo8xenP39t8h6JxoZ77opAgSTcpY0bCdhi2XHJYT1cxwheUwpwVnXIZzq3rw/HRTOkcPQ6cIpk3Nq2JjDT42HzJyk8M9CbXjZxWU8RGd0WGTEdve3kGC3BfaoIxEw3qR3e7SJYEF6seaimo20Zd9IpCqqr5KNV27Fe2mPcwrMjyieKsjL37o6B58mx1nZoQuZvDSrQJ+qaJkieQdb4G2Lk7PSSt3YXvJ4+00p366/BvRhfexeNYtPxegBfxhe6RXHbleDqnDsNRHQLl2hrnhipAGmMpEM3wFl9l3Kfh1LdY/uoTrRBetLIRXF5wxUNvB8c41AkDJa/VXv5zCYRPbkMIWVbCwJFxJgqlo9dVRiPJIYIe7W5nM4FF4Xv5ocxVi+Jx6SVGBEkk7SgD2DaRfUc28d8AmcchFYo/r3gzMjespGVuLdjSCgI+P4lYX+ltj+yaRlPG0VrVtGYx+ZNNEFWz2xX0V/REZuig3FpqZbrs5WnxwEb4P9QeHPEyIb19VH1LlvWckgXdqk+OZk84ileMYpZsoJ2to5aKIw9oIw7Vs1qpRe4ZKQdqR/cfXHXOsAwurMuhGJvvkzLbfdht8b/zWByPBFa42wqtSGtHRdJYsJmFnElB0tTclh8rNVOhiiJhkN+W39NiixAsoQIrkxUwVk5vfa1UxFvUP7Ol6m3+MZS3DN017gSSdSkpccpqgbfOWSmD36tmpJLMPqCHvcfNDuSBF71paMyDr7RwZGPfCxr77KLGtavkuTQiDRzi8rrdAdktExin/yUBRQuT9CT8C/oJgAkTSARO8C9rrO/F9EQjCInHkhmt2/Qa8cxDcHs5KK+b/sypa57is8rkJso8P35f104OUjp4THCcWygZU7m1QVQFE8kvPRbdD7fTqMXKt1uoGIWBi32J/Q+uzflQD+B8VGyeAhFw0Jwr8QIbL0btj/HFCE8dByKNzqgVXhBYMFE5+xT5cyUlkt90RpaiVzE6BlAgcMD+dmiO4J7CVp9nhwObkEcrwz/4j09QSb8kb06j+KmNSr2QzBypjwyj3l1cSa7NtFhvWypxy8TmQ24cNAITwfvCDAJ7tvFMNHld06XGv/gOffPWwvpEhp1jwqhDG/gKHwB0U/2rNWQN8kL43Q9QzzFDtozzIwzn0FaHsTBDFhI94OxwS3Kg6F/ALyWS4A/zIM+TqBPX4XKfSYdG7FHNKe/b6+mVgWPeJZDiyU1aL1JxTm5sYN8vhzydJ79NASPGcwA3HB79xQQC+bQFGkfonxZ5EDpwgh6wUBHuYtH0Kp03CNutMH29TD1bpx3BtKCmJavvulZwicZmp8m1sDfiZy1oQkvMpsb/xBBGCsuxZSTWjPF/1pPlJNj5gHwT0yOIOMvGj9/60Wj9yOpyvjewXjDTAHaYK2GIL2UqKcF3KvdPKeCNUa5gNemrKshuoGeHZGGj4swyVzBTR2sMTeAMMyewHkmAqAllQofF88WdzLVL+Aq7aGIqJ17Qn/iJTa0ahtQKz6Fv13pstk74pPPJc+X1KwLkNPr61SB+RyPks5y37IFrRVII+UC2mJ4Qat6mi/vUuckhoZQKqkkXsYsrmSlK50iBaXIzN9+2at2nb3xgtX38kEOVCPG7V3ts4huv7DrF+jdezRcM2We8t0hHimJZKGStDwxxo3m8NbRFLjHdmT8OsIT+WWiVk5aQlWjrJ/5Nds7cya2KCClZv7HCEXyAVqPax9g/cAtl5ii7KXpLe5GieoxQgutHlLCE+CgBUDNotA25Xsf8FD1MONgGGUygvjzytPokfpN8seC3jsOYp++sYwMRNCvei0YJ9BQn0eU6voAAXyQzZc+UkxgcN3+5/UwLJNGqRQJYKV5R7hMA8Q5TfkoPAEegjRs7tr+m/mGCvtyqcmNEYXpFrUiiN5eP9jReEBFn+LqKGjvnPi51eFjDcl6VzUzEKBxAcpk2lSMSc2i+fW924GqdJV/Q/r/CXdBb9cqOyV2SHYH5Ik8+x7i0G7KdaNxEpIcThZDaqLyS87jg/eqWLOnlXg59UWF6kGyPqYNlatR1AD/suanYp2Vy/3h1ktHGoimni1LxZ/QxDwcMBr1a25v5+U8doPDPEarFuIm+qkI3/F8Tcn5xxQ89WOhFjqCpdHaVDQYf9jlsI7I1wWZd1PElybxreaXgOcr/qhxTdm1K3qNnOsBtf8P4LCsHgD70xWOMOu3RNxgHTGCH1B7CKQJyIM5Xt81W+suuGvNCuEH4EVI95aA0FHp108IyOAqBKgA81CcLVaM6oOXtEttvfM/MRxZ5df7pZ7Uj1GyEg/JnIAWDmSho5Lil/FMYC+G9A75XNHP1UlrASR39Z1j+wD+Po5DRVmQ08tPeYBCsaFo5N5QbVW1Ju7MYdVTVW6Be1tZNKPKZvGi4Sh0aiXmUccLupAdgSQayAmPaFMnvTJ+LttI3KegtDuyUfGtYMXDDqjdWe/6r4PRNfirhoMK0o/WezBdTwYMfS6XYZQaDgk4NVeMBRBx7gZWgNHJF1qObR9Wbytra9gg4EpxMYW/is30frybFYCG7bG+vd1n6KKuKd7D/lxOdPn+XfhsMFbzElaJUScwC5cGpffxzOmKqE4oRkxDh8Su5Yqgg7+fKZLYlpKp02WYY0BNBDSPubpw2yg9Pt/w5d/dT2mxQCszzknW2T+aGZMja5zy5smnylfojCuDMNR8ACUW7ZKiGfRXPYY9+TkZToOGBVW2FzVDo6MuIUulQttuLzJUieylAYwiDzinbOXrwpzzTBcVVAUEG2+TwUnp9i4zWxiP6jEimL/QvAp/Ol9FqKrBiT2bX5u/DRuj1jWz/f+nw4YEKhOzH/56ASqaz+h1ZzfVl37etpc7HxKbxtT7GZ9TwIioMCn+pur7GQWEQH5NbHieRuMYyovPLUyy10AWfZ0o/g+UCmIOk4OtjYD/3vWnbC0/T9lJ4F4oNBibnoD/DLZkpVLzPnSLHZXybMaHEYLu5RvbatEzeyIFJHMDM53TXyivPDqlzc9hoXv0HCiK6AXRdr026nFdAUV9ZmmaqQnKgifPo1vJNd0fwoFVWcF3R52Nl0wtCwEU08z27Lp2e0mETi4HsIaT178P7IR/t+tfi8iOah1TnQvKcdviHHLPZVViW/cERnkMqui/Dy2xM0on739DODjF1xEuRKGc5MaY29QsPbyq6H8zW07HezNEEHCkitgaWF7DOvmnMRnKOQedZq7c3fB21ookrKo0+LZOFD3fpvxAf77j11hczpcEEukZcQkQRgDDWWv/0rbOfFlh920vRHs9XcINS0cos8ZfN/H6LChdO15t9shc4vV/re2yU4eYiEXTUX0+XDer4YBm6el6BxwtMBvz1IONQKoR63ejva5R9iNsYY7vhWwZHqcoXjLpfWtnXEMJwKLB/GXpXZHS9cBrxKGuUYfy4Jphlmrea3eVr80f1vNiAqOfhuV9s4rluAWPsEVeVzx2OMB7xQjg4T7i9DMxGCvHMI2dkrOKdislf0lLYls9fqrOkzv2Sg+f7uZinFGNOKu1HOnADN+JxndoIS14YTfTR0TCrODTGVKp6eWALYtq8DID+vmtuzni5pXYLHhYDtaV6peWNdUDq/9r2fXOrRmc2s6grlf68eT7xZ/xPEpCHiIM9FKnJyssKTvP3M7KplzBflSQzNsvnCAiNuzpLn9nRZtCsau+yjCOe1FpsKsUscwzS3wSBg8PtDoSs+WPBKWimQAumGj0xmNks8PIQTy9ZeYYcQgP8PrdVXsTbUflaKgJ0Bdoj2wGZfvXd7ZhBjPgOFjxV1CrrSK1q41OZN3nkjzYru3zkXzTnm9uM9TZXX4y/cjIHP3Mt4pQLAIexR55Bj9sSOy74KznPnU7WelINdEGd/qLy8+57RHauPpEWGU9aulf7DdqeX3GGIIkuPSwSrZNiOwiCryY24LmaVHeYm3qVy4dsa0Bgjo9PWZybQ1UUTShGPXFUfsioJoJg7kBkNShtGhvrYtWYHUmNPLNypyfs2flH8aLnnC3txoEGqduv3KpkYzAjz7h5kOYKguh43VXham0UGQvYyXYBWqE4EMzkWIKg65RiaC4kSg5Lq2YW5XXFFgF0AT1hO2giOfeToW/gzicvfkqQlvs6fZul3WaYwCukidjKET8/6QVYvxzq0QLxw+FqNwMJG2mssdHPtxWKKZ0PeKVy1o3RVJndfYiTv13ER2Du2qoqCsSvyp/TnNzj7l4GBLwGm9VudSj/DUCmhtytTArZrHoLjEr6TVUsYy4vtAl5qRFEl79dRXnOx/Jr2cJeisZeM5sbmgaogsIW3/W0ZSe/T3CfsprtMfJVNEy4LCbITbWVvJGwb89yT4Y7VpjoJJhaDekK4PfsENdI7OTbxibv/zmL9YQQLhRIQCAv5JNWX1kaPqR7nFa31vbP3U7ClmDtk6OvszWj0id+YqxVg3PtgDmRVXpXrVToGM51b6FaC0uqVXyLXePSeC6iRCpmL2F757jEQ7SApAy02YhEm4AMArqcURF2+02VyM8qj3KUE0Zx5Nj0xpOu6jNFS6/qtgJTYrwVgMBsRSpyf3k1seTTsAy7ZglcQJBtufGY24Sexh0eG0SiEZFyBrKgoK5ss3PwmyOLQP9PCideqCAj9ToKQuHrIa8g0ImBk=
`pragma protect end_data_block
`pragma protect digest_block
4e89a8e20a029697571a55564480f3a642d920552b1a90a3e599e5a16c53b1c8
`pragma protect end_digest_block
`pragma protect end_protected
