`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
0d/qSIMV6bNyzY6VGOAy2oMWzB8hog41u+vrBQNlFsIBMZTL2IJGiMl8dqHe7UCKKSRwDg2eL+KOkBBMVdIzX+ncbiAF0/FxQu+dMABAhckb4mjN3dXoSwldntqk5RL1zMdaiP8YGP8cMyuU5ieM+mrm32dwjuvotlTzNTALbiTgjPwy0HIhhFfbJaPauqFB5ZYRUG6BvMRnTgW4BaOiB2OaX8rziOQrJTg9KPvujr9a9k12tlrcpmsZfin8Wjq7YwS5AFnOii1uXHiFzsXzHH/ylOU/XMnVns2Rv4QSytn9iZXs4+vDjyjdtM/YiroK9rTpmH3VeMQegPcxercJooAP9n1wvYjAlT2OvittoKcxIBRcPWZ8jIprKZsidhplrcxXqmKmaM712FKv6OGIdWwzxMVae03X7HaWZ14rpdZA8LqPiY92RYBopO26/clsD4Y+8KkJnl3Zo/RI7d80ZaBztD7kF314vsNiOzDKnpBgTDLBYIrVVIvWZrwPF+H9sc4SrFITxFrmxy7bzq8875Qi8fKtfcjcz8deLW6eBTMarZYmD5uD2NGVGOm3Xs/6fuAMmqp0R5F2jWWLLL9X1Z1Krt4PocfiKBkGeisKX2YMEpz88iECTy5L9ETGg2naqR3/6oCABPC/lVx5oTJggxLup+cdVGCrP3LbBTX/hGWXg4FYD+NZFCtW08ggWfAyjLqUpVy58JW8eB1HHRxe3UWAMn6XldCU8C+8VoBRhP6sFWvz1ji884BqU1BAr218RqEhxWPbtjXzqxuHephW8LTplgFaevvIlBaJHP0vX7hPqU0jAJxkn3jz0CywNpNPRfDYr22F9rZvFeWRrjK5U36TpzNnyv6t2t80pgjV6cjYEHpjoA7M4ysqeN/NOF/qd4hYYABGvlhg/wSYEMk/cUQbGu9hV0ulHdxr3CQJr/tXi7fM5+X/g2gdA0T8Qu1BgZBOTafunWNmx7ZXiOjBwanNUjpSBY7UEuDkJ2k3vIVmre31vwqbkQAnnc2hVO0TKZo0QaHvEPy+opIkwH6ohshug4RNtdFjbs7YGgL0b6dEP9AKXE+kXER/4M4x9TFyxoViJ1i6COzX6N56DCj1gDSH0bXCAvx0D2uYsNWvfTsya94EVIvjgToqZYZ4aOaJenEdnN1YkijyeXkiBOTufG5+Wlmm+LGf5XUBOp7NdS5wQAhGlos35Oa6qRfmTDrT1DM4rU9fYLYg5QmHhavlYTB9pxtvxltTGLNMc5iSHqMSv8P1ccxpvEIc5Ywvb9K8iGuWSyr7uZ92xmnpv7cH5Pe25NFew0qem6HGKicP1uXAqgRD+WPjvsFsBgSjJYNghug7h3kKAsNxOduUgUWYc3aIUVLA+A39CYoBjTTGkOO3qpdRUjZTKpebvc03o2y5JOjgmUwwA+PQDClLJzynW/H0HIhp1jcr/sM8zuepo7AusGh92VVb0olbxNmXrCaUAODrWdXSpg7jmqXUrUpboRqvXt2Olq7k9ZyXnBVTD3IFs/lRFtQ1P65oMJ/kLAN5SKK0xigTUi+1J5fk/kqWE169mjf/lYfC1YmgEdrFymyRJURZcB7pgoNIv6QrSB1xaKkCPqGVU+GwP5k92aj3NUkpoUfSlAbg03bS7YPpi+405g3jyIIVah6t6AxIXyenKDYRtaLgPP7QxeQ/tgLJRdddz+aCioNTW2A/OMWUnalbKr1u415oV/8TydHLcki4N3/8rbvmHOul3ti6B+A2cEJT2AJ0ECFxaBfjpDmv1FQxLJwEzbYFR5MhA/YXQpG9vrhVNA3RJCcVw6/uj+AekKfgLX/IYqwYOlec4nJ+ZhK12jlSJ/Pi4gD3s0DhNIY78xlxoGAIrUSU1WyHTumFx46UZy97vsyaT4/RikV51+mihqGLzc5NMRYVSIPzjXn/HuB4rUTuR0EeyppVy+Y7KnzplbKZFewGxiiXnKMdDVNU94Hu1jNd6d489L9vZ6NpjDIltGd+YDwaCAuaou8w/3Yws2RcYbhJn/E7gvjla70WuepO3hXH3tMC+pEmIKIg+Tsqzpeny6ci1jVTctwOYgr4wrwZ3vsSFnWlWImHTYtGxbzuIcCRq1WpZsHA/ALL2KorcTfDvLN9pd9ohq/MhHjuRxDxg41z4hvhebg9prSudE0NjYlxReLBaHnntxCv/b84bFTCmOrELk2wvuitK87m+kkn9jtHwDz+DeYKX0eZ05zfcXkhu/By2qOBBdH32eziIXg+Dt/fcDnfcN32pP7fK+4CezU8w/7Xv1OHRKX4bL8+mE3Hxkes4yN9uWO0CHVSNpzKmWoIqgrxZXh5zcfJliynqHbYQfF4GmJPqUF/O2rGDSPGtKWg4elKcQnCOxwAD8+CnyrVXS/8rAuI+GI3TOfGCwBbAelp3flKt/DPkjCspiXsX/ayaUKOefAEiOCDQlqdS0T7Q/qmpDCeOR8TaNUy9sbIjxOYct5ertxm6FGmj3mJsWvjzGlaA7Dw/yYPPTMniYuXq6R8S3fztBJEtVW3mxRaDwbOKj3LKqyhgef8/kebcZDDWkT52eF+l7dejIg0gP/K05TLvUY8EJnp/ft1pTnzU3+T3zTKocBQIR4gSaNRTtrm14Y4c/iY6GFUv0JHKZcCmFec0jOk4X+MoxHBI6tcA15wulUQYmbNt/fxXcFTgLuN74Tvci8DO8o9DcDAHCWM2IyBkcANop+J8chNQJmshykeAa29RUMAcMNGHGp66DtuYAf0cv9Ldc2+ta+xTm2BG9o1FKI4huLz7G3B68wj5w1rgfAW487wzTgi+56yEX3YSHdt2fvAZ5Bxn6nXyq8WFC2iIJa7FDyCVywLOGbB6kuLwSTCkYhr4QwIDvL2QEwLer2FzTTVoWlLN2dWFVznDeMzLNT45V5dYSzWtrkG8nxASntWIK+ffL0CGnD6feHHmSWNkx+a9NKsPO+0zvuHDRJ2UHOLVT/xg9gRVTZOaVgpJLZsu8CgSTKh6cH00cVs1jjjEA5fzlQLgJxxABRWK5TEgEdtl9pyeiEN7jNvGiA6YCSr94Z427Mn+NqRz9G4gPsSgO3Ul5+tcMr6XRLj+MGxqOJSbC9vfoyhinaBR/hNoGnUxbyvBEDbA6FkBJ95Un7NNc491wj8rFpa7dwFCe2OZS8yHpjHTPu9evP0914EEyB0PF/krvnhesNOaCAfwWRpW56wcJDyOc48M02sPMiBvheXQSb4wqFmZnlpfSFrO2ospPHaxBIjRdUEY2r8n+GD2ZGf8RZO0bmYAeJDScB2hbEQn/63m/swSvNsWMEEHXh4XLZoO+qvnvcZnNnc8RWxQ3+8crSNPNTuvQmpQt82XXpyi/knOZlksQloTE1FgBxlUvlHrdJpi8nKD8FhbE2eFBLLCYnDIAqRM0oRh3JBtWl+UeZzFcNV7tXnMLyD5jMH9+JD1RvhBoP3+ttabpIOZdFNRvBMc6RJVl2Is1FQ0dJG0s2MGpQIEKElynASE3xN/lkcLK+QYzB0VrorwUUxjunvEnw8NtyZ/ZLATgP6PZW8e4eBV/CeoldfjMCdN8c4qjvKPIxCC2MrKpiODRPwaBTwYaLtnwncgUi7cT/A5eC5mOXNyuewRd3zR4Ta5uLaM7rx7ucXdTiGhiCy3sp19XuYmGTzNu8XbmVKZaYO9qS1J3h6kaM3+y6Vw4ZzGklCS2tTOwxRH/K01ENnheZ5WUIDst1zmFetmKyY1F0RhlJf/rd7b/pL+kGO9q94H/UYibp8hBYJobKRR56jgVXs5N1n0qTKaxzmhLcgpa0KD0Wgm1nLyl1UD/w13pl64qJTcDxZfVTNhxQYgT6ln83mzUlPYkSg/v0aviBTm9oUk1NaRFMIecJUvnpM6j1VejFuGpwXs82W1Bd7B7FCcO1itRwXbtarOTFyghI+sOz780zoCTHepVISGJl0HCkjBmfFJoXYVGQxVJG59AQHwkX04EoikuvKYdz7XA59C/KuFkM0d67ykVxYWAu+9pNChPSf9+Rwwt50K7OK1urcoTXnjlZOkkeQ1o9xlk6o2+zVEO3ZM+7jWnK8YS4V/ye3CQA7gNVdiEsJIKYxObm1IxBhPaR1AmmeKjYbTRJMsIotD+HM2J9W4NVYgkVVnbZvcvcLfDl7Y+Pt0toDoqPwhPod+z1SdtMDSZyZf+QJKwh8MpucUrDhCeMsi0FxHzDM7wP3CJR0RrJxD/FGur9qwHnOtX+BlSchbTGyLn8l9DQBVQgbcVG5coqU3worxJpMaHZmcpnb+owvJH8dgbsBV320OT8Z883uE1MpSOZUbnmMDjSXJj+0/zzY9Wz2Br4ipPT0GQJ0hUC5ahaHu4/HOOuoJ3xZCm7NeBYszM4VvFjjIUMFI+4IQTWoThhuK0CrEfD6IanO6/J9UGWzdlTZ5OwhEfi0WVWHdpNxDf+bYPEOuVyHnH3OTUoRLHwZpUj4ioeHSE9Vw01TwvmGxGoYCiuANetcBY5+Ham8L7t7kfcJ/LBAb6kmEhlIDkueJDuS1rQbb932JwWTOJrd1yYlsDVmvK2M+VpML0sp0pKUm471lauozQpQjSS4Y9i9xHN63ou+Ns/rN74ANGwURPf6MX8vTKUXoNgXKXcnsxVZzWtr0QYASjE5w/L/Aa7Ysc127E1wKj6iCwPmETmpdZ4yQqnermX5Omsva56Ch3g7/BopMY+nwVv5iJ43RboeyXWQLYHXpXylC5FhXJElmoMIiFniV3CHga+wbC8OHIVXEfIGrb+dZFT/fe4TA2KB+7Fdn2QHE/1tNVLLN/GrNKgieJepPeAoZwZcsso0s7q9+Xt8WKkTRHQcSiuDSRY8gN9Li3MYK20cNtU8Y1cCTBzBKi60hQn0xRlzpN1Msdv6ww4rMDVBkXH+K7lXjtLokc2fmxC/WveDXjRjDRvaFnQDeFx7HUzlUF8wG4zez0ohUc+WFvc69NDp5iN4EITCP1RhaT1GmUDFq7DiKLW4jN4j8yIadhFJ3xAjljfYe7w0WkG9pxx5Tl9F7JBgONcH00K+6u6Pd/o4h97iFj9MWjrIPu2Q30VfddiAkHJ9CUh1gnApXrDiqj/eHqwjDWwq9MO3FdvF6gw+DEPIqJtEqinhT2vwECUJ64JUFEsILTPbfoyjXr4TOws7OVcF4WWBE60C+BqQQ22oXCwF1y2snsVDaV2M/D1HKiNoJ8PgbAi5DYU0OaQD/IUgyZ45eSzb4t6lK5eyB4NzA4lKFgqutGZI9uBslUS8bniVdNTDbJW0pn6oPwQttbn5qdipSF9tm+rcqyQn/+bcAyj6P8WVjvn7XuKafSYJIkhSTDuNEYA9u57f9smt69yj27TxMromGdFNbxEl7DfHi52HXBJkxMWw6TAXAS4NhLed1M1wzsqlYEoQlgKY5hgnBaCQEzzU2ykDeppKmkulrpzGLH+XVAQv5tD3xJQ61SJ8uxNef5+kuxqYEH/HMhGiGNYCFTTm3xxA4a0pQMr/Vwmi19CjyZ7pMmWDCLe+evmOONX3weDLOnbpmWIshZ62+zULlWr0urFuOksvbND+uZ9fBv5DACJReFZrT+a7YQ1d2lnAS++AVdtJY3odLjSCYSzAiYfpCzyGzuS4vlwHYoAQESsz5+w6T3jJRKFN7Y1/KzQedcCCqdmbJalihHufrBiweoBz0/XFy6zq0Pq8V1v+0YgBz4I2xjHOlCP2ZIkqatNtqsth3XDhTMOEyPavc9zTioXrgsS+8FWmsRR+V3i3+EkiSsqVydDDrCU2qHLmqoCx8KE3reW7F2LN0/wj9bDff4QxTgWTLAhrWV11cKdxd8gH4RpegHMuM1xHhu6WQr5tfWVhjglf6jBIemJNRkF9nu5X7V7zu3geVH0unfo9KHHvVOwXlk2Ofzff33GccGZVQResYvCz9GcZQUOsBKXZ2bJFhkFLvCSIPHMF/H0OfIH49wIhdam60zA3YHv9oZqi8jWrUAqJxIswUf/HAfw4ik3MPSDCLI7ClGItPSfCsgz0DFksH/5fkGR8PEgYT2nT3Wvz3B4+Wr9/nAS/lq6A+s+G/q+pQoWq/lvwIL8YUqA3D3oOsxEk+PaJ26Adn+aX9g+ZA5rQIUT14DmYCdfMZaR1s40HlSuYhQ8T+fnZ5sZRh+RemcsWvObBT5Ad3AL+KvMtQiVyEjdn/F4p9rNDEdPM0DlXVhPuppC3DSyCCuPmBYvD8qN74GXKbn/Qw/Z2z9KU0Fx3j5mu+BR59/mZK39Cw0dGx44Oyd3b8NPYv5FnpAFIh0a1kLZQpwT3XU3HK4uj3z9Z/oP63qG8g9MEwMKbSI36JBIlyk42Ccn86bEdF74Uaa9SNIuq6Xli3mMaliz908w01rk7cp7HAl8Krxr29NAv352ttpVHLAq7lODQdBhKbshXadVTEp8F5yNpVhKrABPoEv3PmmsRR3OZIe287omOO2U8msy8pSTYm3/Gq2hPDRL47rAfPCTLaPuedHnbRndomyMTGYOX7jD27ENZBrRMUrC0bZRfEwkw+u3I3lYR8Qr6+zZqunAqz12H7W4y5amZmCVNPUEQeE3EAybUR8SdbSCmnvWQNuZBeA5rUyZael9+J1Tk0jJlF6G7rsJm/BKVPy5jNYggqFIE+ckd5Q672sW3l9NnKoDyxhtNvtxfEWjW98/gqWMAidXTVOh9w6RdhUcpQY3LW0i7xA+8IJxnNHlk7IIGVEbJseD+dOkAIJYd+K/6gR1WHt6+FFzE98MLUDQNmHzhPbxASYQb+mOtLAy45+HARlIZqu7c2b8GYOTQfbYvh2S4GLyJmhsUs+wFp/4eDRSGN2B12/39D5bGdjl66CiowEoQjMVNxU/0aaFAb+huglcOvw/t+E5DehUgGJYVrzxjGcjCKaHRu9OjBOR2a4J2Mj8IhEE3hLdkMTwqRxmmqDx+pq8ghDzc6T4+e1WvlKN5puAHECQAwWW+b5YzMqVW4aeUFhdxciB493XSOHPaZmSpJk8Xey1z9+1Qh4/rtXl1yu1WEbGNIgmd+bqBx6AoUnGhj+I8qmFLU7RKxpDkeV8Fb/erwQZ9lfb4n3HLSfrYky6L9yhIss6KRuDWnUU0OXUlfo8qZgZSXKTYP7AmAjpLohcK/U9k+wPJWEEKZz+Dmq3JKRWHUXa77Lwv9Og4FBYGxQiQNYajuC83V65RS+vUJWfIvG0NNYMz82xoi94y1In/vykn2q6hjlqr2rXUzrtNo+sy9HnGIoBbB5gGU5OV6xwlPtHz4FaU5/ZHS6QbVc6CFZj0EM5VWJ5K+jdoDxfv4LrdoodaX5RrK7n4S5/juqcmR2knaDLGa+yy4K7VbPPqKcrbH94BwxcoyfzJg2rlX713n1f2BbW6RqNmRywdyUCEcNzI8u0fI5LRPYSZjiU73LDTYbzwe8WV33xr9ZFzUqtuRg754hQuDLog2cHjD5ToIJelMfAX85FUWcAzzJZTqCVPPadi3WFJkF5xTQcSzy6VpgJB63PTKCdAijEAe2Pn8mOuKgHQFtdeK1ifoTUtMJiayiXPCxfHrgkOCF6GiUGPLeb2HdRUnk1J5Q1C7T3RJ02t1t3B5yuVit8QidQ4D3Vs9dbc4STJSIZzf8xFmsXiyM1hwjw9aEvwVhsSaBQa2l65HwFKQT/KAY7jjXZQ/y6r8hhk8i0oeibdCpiVWG38ATfd6NwIBxqoyOoKxppsDdLhxDForDoZOTJzMLTEGyd22MvolSCfNpZgFwsv8N7U4dAri9e0v+eNv1KBMVc409UdiL+kHOXl8fOHaThgDIy3btnpCR7Z+sldajy00mhsb+DBFVYeONolF3GKYm+a3UoShqrQnOlTSTCd5u4pymgdVZlcSDqw+SERw/EKJ1J+dP1tYC9zbisgstcfZLALHMOmbHW1nbr9QDX3ZEki6ciTexGg8pDtz4NOH1O2iWOFT7TXJMZTMe84Ur6KKG3PyazS7/vF87AmmtiW1YII+kKUbYCdW74nx4ts90v1F/KUSh9O2LwBbTuk4dlPJ/1jOuR0HHGAcIGYQEIO9isIs03nczzY09Z4dav3u2QsPC1zvbPtSFo7E3Z8xiHwni9y8wqEwA/AWP7bpL7OewQC5iAoKEQNno3jsQQqVUZUP0jruIdTT9KHe3tvN12I827i9xymIRr2AlJstXbI6vAqAiPX9m4F3ka2LQTLSX/bhQ5NzCx3F3EP6B4gJbf5C3/i9eMK5RZxhaB73OoKbV6CZ4J8jT7Zlcl3fjD8ekjsCyf5LvQVdWdHSCjVc0OL8Lq8qLfMSjxLthQg4Xv2fu6ogLKlujv4mr5HL/QsGw3WKe/rwrSB2jcWFaeIriDIcOgLAcoe+MYDTOv+BorjmHCXc1jskfF18pxGdNRRFc/7tmXDi7pJ+cYIC9njZsN6RSBiiE9ok3fSMD6SDrXvzJqYjUbyT3JB46tjfephG53cc7AYb0q4hKyYJoxfNxwtNItudslemt2a5CbiafNQF2It7eY09mh0BC9sPpY+nUYBqmvKqz2VW8jVglEesGxtUignd365HLbDhLE4rXXkr8wv0tGomTYpUnuKjxiJjcO28hce5BTIjNf9/AbAJvV9tSA6TNRq2YtpABTc8BWu7oQQuKpCvqpekSGYevm+qG18MqLFkqpeGt6TNyGcNMe30+L5ohMq2XKUppPC8B8mkYXjI892suT8aITtUxjxtYNjyII5/AB/0r2XsAPR+pHZAPBz9OuhRqbD4i5U6CNnLzmqPI9u0ZAlAQXrrLN97NRb0QvRcxEzm9N7SX8sBNcXS9HbOgj8/MRc+GnNp5Xz69AtjDE/ubF0YTtqc3QAHonBxA839GUsNfZYWhHCyGijBAXVyO27SbyMJd8jMnYkzR1FraAXMXvL2B1+U2q1pCdzBr7FcS09Lp6ED9D6ulXRiO7Mf6BvFoBnkgLW3t+5+P5+KYkkeWf7EpMPuYar1fBvH3ee0x39H8jF+Bnt7dbosuVZYn7ZPKi9AwNz1vGtqI4C/3MPLO1bzoAheW8yvSqOuIKWITqvDWmRhDxvLF7EtIEhfYAH5lBLXo+0Fd/6p7WcAuI/jn7nX0cH4H2ptsE5Z5sYxVo2rB4Al70dFoavmvwod/SUlDEYe0K26I385TJIwajoaKTfwFkKJpCJjr7Wc8h8PEdPab4J7h+F2xQP2I0lLPL15as3U+x7UlMveY7Foc/zNjEXK4WCglFk0zJ/WM5r0tWeQF892BdkEMogb9NOY2itT083dkUmXgQucbktTGyWxcdf+yVQMxZOhzcy2pxc/DXPKF8anZXnORCpnBUQUvdAEW84dde8yUcTlZOdflbawhO2oEZQZFIQ2vZixKebegn+WZcLY89btOOZ0I5AbKYWC4lAji7ei6MnCgOpDiGueeMA9fLDMpESA5rTh8j3455nYZo6mwYwLNVo6O6Px4XkNIz9k2vjd3917Ou/Uh0C+KYKPZLIw79Rp3DJk5OJjQpdiSVecbaWEu9hjxKhiqDMwMkJJceQQjpTzKrXiJQMUQ2A6Om4LBXqMOsxCyAVtud75l67+d98QKHjnKKghOzou1OuLAZk/hlu6L3sgRsHidsj055aG6SQrn4zEjkFOog6Zt689GFfqjnDfkUt68SRA6Hp7ztaxjlYwOPvxZIAy/JLuWIbaIN26bDfh5mAZnSEqLgD1EcEl/H8FszpQEL7DpSKwypHoscp43jzcwNV/CnDMnvBgNdMHheRRxSvjo1fwMO+zRed6iI5eIc/XDWTzRsS0VbRJH3mTEqUzmP7+RA5IbmSEnXBGefpf4jjNgzyk6u0RaETLWxOFPizjD9SAvvcAq9qd7cs9OMtCLuxrdKTsGg0edezRf6qAu3i2AsvARCoFoOextJgYRGUUzX8TwwZQhrDpPWYNscWhN4A9mJIbFaJDfe5NlbmFDWXGmaLI9m7UepKPO5DJCyBcpN1irBuFivXNP8pdzuvYrkjbsVmgh9062q7vDRlJHv3wkzLxFxTdVVqm2IjctjyQnp/538jQysOgyJUG/JL1QpnoGsG5zmcAEIH/P12TuVL79yur/NcB26Y/jPN69ENiYGaZGNWfaJWmF1g8cSdVXBiLa5sqzs7j7FmRtMBuu+nGRe6U/H9sIB3PWB1iE6PmL8J2d1BymTjPeEcGInbv5jIfaOogtgAwJlyOR8UnGrZkFHjf7So/gjZjrjwCn2RIbjurZjgrQ46wdi5fsLPBtvnbTqktKO0VdBOnGeheQCCheBcVZp5ZVGolBww09KHJdP/j7N8xJABXDPNu5nGGkAnvUhLyDifwEK8vZlaFoiVtzilsaf9My07FTKkVyWLtUQSOLK2PdVYmzKNVWbrg6wNWE3hz3YOlD+7sqHfY76U1TCyN6BKv5HX+zH1ziHrFAGxM4zmgtQqG1NJvCA3iZyg8SBSl2gIr0X8DpeUB01G0yOlhJ/I1gWwQt8FotlPCdUDfRF8Ym38mq8WWJYXevO3E9LCQnhGdaox57JC49eJnGuvLd3Ucgne87/2d1pVn6ABkF7L54fkEQNDFGvJnkQSBdIqvuYkL4LOkEjAqzrX3zQ9dI4VwJua7+BtVNV3w31L4+GYakwgCoZCeK2uh2mx/2EIhtFaqGWbtw8+7s2lmdNV6Q4TYYYRaEHZqg2TyLrhIyktWlnnx/Rdyy93KJjfmL0k3JGEhdr5bhWXGrjh9zAIEoeFijH8pr+VLmksXmijPcm+B+UpWDdfAPP/TSsEPVQ5mEmba0GXCj/bHUnGCsORXEqEbxrQbEE7N+XfgkDujabGnFA2KwgzR5/zU54KJ2yU0tgaDTAPTkJ+jDhA1LZb/Cs37cyoH1FBBeb6MmEPp2h0w/ytJNmZfud9BF/qlTumRf3ym017avpTx0wtct+IBuxFjIc0xbk7R9m7HZyx7qpXhQzZ+uNSr5Wo1/uAoKcbn/TfqjZCWPjvVL2VCewlc7ExpUS+SbdQTjkM2e9U1w9RNzIoErPNYHYScfz3lDfUGubLSwZGRPm9RccXkbABmYQ7jUhBomcAH9TzhrdSoMz0Z+OyBZE9ofvBqY9mVIJXrEoqSiEoikjdCFUAkJ/cgo8NxqKaVYBRQTGWdSTQHK3cgwNsg4ULjJfAzRQTQDpgmja4YGIyKWu6hHbmjVvWGdWHExUKx3n+lcRctXzyuswmsTZ/yFaq2K258wMEcCaFeZh3IzvIrBoJy/vvj/SPWR1EW31HFH1tLpI0C8f5+/XmP1C0NX08O84lHZRftGKi4BI9KHNU6VXi4N8OwqgTxlr/XWrFvA1JKGw4ucWok8pBNtrpW7e1HjM9A+Zti7CFjyNgxAzp2EdlyCcRwxAf+yH2JSyZEPSo9M1xwnJg8iliAzW7AQW1GJY8JM2s1WXpW1IQnTMXeQSYG6ieL/WTus3m84kTRoeVeS6Hk2DOuvIjWKU8264eJErIK0p7fLu5z/aXW8lUJ9VKzyzxCHvoIvG+Dz97iaqRU3PSMcIHnBC2unx/OWJvMR7y1IAda+0sGR58fKPnYZMh0SmQugI0fZPeYhG3DiYXKmnooFXRUnVfzNqIh1FYRuAhgZvH3dmXXPT2tSSP/pwMk7FrY/7LzduNsceYTmJMD7EvGfla8kRGp7XV3tjF9d9KcgeINjGqVAgCQb7iz6+4N/oXtjN0M7Ht9M/Avg7/E33R9U/MzKw7vVcOJnjSabsIyQr7tc0KUzv9VIFMbOSB6QN5cEj4PUfuUyqi3XBqZXGKnuMsSYFevwMeaOsMCTpC9TlSoEVabO/IWPfjsOMGznunKVgdkzPg+BdpYKs+VXPIb9ZSw8nGM83bZxZXQZQhKnRCyy6Mnv0qOKOXmtPxTi3U5TJKx5a1mazGNPMisSRtDStsJ1VHU2cpKSgbsc7SM0VteLj+SUu4hJRLnbFfcGrlJXb65QQWXdldK7mFMNQC2oSrIhn/W4JDyZu5ahVjIuA7z54r8L6WPrAYciSqpG0RD/ZE1h2+NjdZOI2N4Sbl62Twmr5GKKHArL+fTHSAOq5RYFfV5qBbq2NPlpJbz3VLU/OsP5PoahvWfX4TcnoRayXOH+K6KoO+Cv5bArONwBC+EOQXFPEHTPghiSqtjsExmOHM/tSAbohPCWmw6cPZwxg7qkxNRcxoHkmlUX88X5BnSTBqkv9rfV1dNhBXVWbtY0OzQGmv/Yl4YLW5MiiRLzR88i9DxazUSY6JzWCG6Yy/XZCjeIM9Bl/fHV1kitsdFwC4s1vtgy1XPYGcZ7omWkoyiyxbCeehb76x1L12+0OYSVWIjdugcYtLnOdhzhT1vLw6jSUEEeLhPRLrBet68MfmlefwchfzzeAXcJjXAojuVmIMgTcInAAHyQXGBPsYYx5HlU7XTm6PZBnZlJl341ieRpFvV7m2rxSskmLXXLUr9UGyhhI7mngsbDCf3Y313mSorJG1yIZ6t153H3hJkH56ECUU5ouFRTHdcawJULOF3cO2ZIfIj5ayLCH71JoxGkfe7F0s2VXvns3voGgwz1wJRRaxhjI2/lLq6GEk5jWnj023F7Iy+fpzjmWHWptUA45D2tppeRsqA0HhQMhQihQa++i3ylHZapvfdTFLBhXAKhyc1shhewXhZvn8Obf/bGMuLWHoMHw4wbqslAO0nHujdrqixUELIb0mXr4cPiFwVF7cqSd0fX/FXYDdwjwSKH9Q4r1o+tJXAOMmm+b0J7wYiT7FYd6lbBOBWurh2/rgqHbIxb7KPsaoYb0NMTHRKEk+p6tLB/FAsfL9JwS1Kyc3pUWuHOkpSZOApnpGwDH+Md/2LYdhncTyFiZpytVPaevqApNdgO5nOfQqvPmTfUUfpBeSyjM2RW1kyakTodm6XUwh6T8YMnwoMaAIBmz8qAup+F1SnJa4KMt7gEPhmT9FNO8OQrKp2fTCV38AUw6r6jjRNxSCVNCD5N8TfoE1Ke0RsLtHkcN+3l5vy4Z7/xuqi34JNmlRTqklFMDPojKHq0qtOTwIsx61gPXnLlARKJsAINMlAsSdoXvYAA1az5pC5G2HtZ8u2G6IuC2ZtRm10IFc5ZAqjQoYkG7SrJT7TrmKcJ4MICu1CZVgjEPgempcOfHsNShX2lQWOb4qAxkSyu7bNNMqpYc15L+nPsVtMThMXzOqVri+YIqv0SkZ9t0FgwDwWiBaD5O6j7jP7Lu6z1LjRl/FNTSJfQwdo2HriKqRfLnqg/VhYOt+HbCprWhYF/yC0XPLPAO7PXTi73cZi3jA2MDkUBIkjEOBS1Gxgdu3rgn//nD1jA1+TdgvOM4IjjtVEXL2P3Qr1NjEx7vO4G0tC+iSSnGRiU9ETpeVqujc0PWI5VwcIRGlS0L7yX6XEB/4xbDEKcilAr774WEPzxDa9n404eYeSPF3AcaQSkiLVGczq7bRv4gmTwpCKIu46EgtD9cgD+pfUsNQ7zNSzMtZu6K1neTcoUDZFp291dA96qXcmccMLfM/FU18PkcvX6pCGAvkdovwaubKcLNIZWUr6XUh0HNMHaQG1k0yOkSBovsnkPim2tLoJ3ND69VaKIzTfKEUnOwgS+ah6e0fCQzbiOd0/vTXcb8+M+sHbqa0jmDQb8s1eLsoSXmJ0xx7xaRst2lzxtxPQLt/dsvw8G7s6McXZI8SgFl8yi7vHPK91pTMevyeZiJuVfTUZmBFe4lrBX9UqNVAdrKuRF2GlAzdZWKm47KnaZ/wdqLIAkc2qtlOOUm0MpYl/FmU5KElGwdS2+Sci0cP6xF+jVCr0UifMCVNGxHqMeXtGp2ch3eHiLCRpqTK6o3ZMS+5vZEO8JLarcb7WorXgoW1VPTSOy69G41aADpfgPPeNtc39pOq1qt5+2uOqnUHaoYQ5qj7M38XsduRSZTeRGFBbhRfhzBrovpSHGxH9gkXLwJJACa380NHYDAzJ1wKFT1UJWx2x1mL0r5Ic7NVW2YCTUTWQYs22P3BdWpcnvxMXOjBcN8o1sKpgG1sVRItHGUuaIGBpIGbOi+zcN37hnZbmZdVvisNId509+1IynGHjqBqNbek2qOAtnFbzGJAMZyeL3Fi1KAxljdYIGYiNKeKVtONKI20I/PLnJ3dt8G5r5vi/gl0WZxcPOfZZGXwh2HNsJzBGVn855SnEckQ6Xfg0Pdtn9A/EeTderAmmZCcpMWMImP572n97QWhEg+eMnJeKmafi7ezT3QCN2BiSYa+ZE8XiKGY2Wwx4ThR3bWllO1TedmIf6WhApsZl57kkHZ03AzixSFUtfAJj2Krkn1OqGHV3ylH5UWWGevEbFWSY3I769Q43Uj5xkyj/rWJexv/NO3IL1W0WJGtFsflx2LR5e9ipfMTJwy2E4ysk1hs0Eb167hbAHBtGWQB6D36JdYVZh3zaEfSpqHvZUujjWrdbML5RWjdlAUM5WevBBfAKU4oHFrNjIQYtiErWIkx3pp/GCq1/rjv0OSIXLUbGWiD3U66MtsPUJ4Y3nmtEeuTVVf7kfDLhi3sL4nKbW7pxR+xEdd7EcPxgMLpiqmAtnVw40MhwLZHbAlbI1jwem2HFFdqiPxKxXUPeXXjNO/+84BwgjYdSgjbu66nGL2EUChPSaFn2Wv5LxCduTpv2Jvy6pEojMdkwLP8nOmTOm0FoPNFBSEfqOhbwWrE9dH5xkMYl/ZSo/1alrT4aaOw3uyBYmv6N1XyzNv8bykKrURoAdV070b78a3Qf90c7Ue7LTumtFTks9RIA5iHcbsZKE8lOtvXniJVZz/8vyWFdwb1IhCfsNKyq22yGBFtRIbZrHDQrhhR4vI8XOIWoboW6r4Q2wQ7tGsaYS9uJ0MVgfgBuYrEzuODN8p5nTiHeHMSYmQjSaTqhtAZ2NOlBzSUAOLSCvz3YErK9hg3U4JLiMdjaA6FAoLbNGwquYsMRhvq+XIYYl8AdLJAVWhFWDjZyPZCGGB81FqO86RhDpAJoyjfPxlJwLzhieem0cpbCOqelGddlK4BDwESa+HNlcT2fy/2PKxVAtLXunj0WmVRkZAyEUp97WpA9GsbkzDoJuEHNiBiplm2zfORr+L8RE+oKgJXYD948dWnvMXHHEIkHglUJGAbppKNvu5OaCtazAl8BIejHQcvDxNIoGvDLWVkEUcin2kHq3BzP1gi/qR0Iz4/kspca56Ljns3xowvbQ==
`pragma protect end_data_block
`pragma protect digest_block
2bf76875e21a25239bb4497aecef7b12c191d5306d59b65df80943582f335629
`pragma protect end_digest_block
`pragma protect end_protected
