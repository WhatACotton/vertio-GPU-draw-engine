`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
XMrX6lMEnOO1pg2I0Vdjo1uXYKY3M62VT/swv7WqeNexz4FEdFFWwC82ZV5VsFb5Om6sPWyY2cxe/0GDA0QeA9KKoK647NLdFsicjWQ5b9VTnIN4qJ2rRPO7dCzYNao58B16Yhg3/5ymXhlPnJ/Y2HxW6Ih9caCiS3K/f/cKB6RqYIa8cwNvp6JvqRoZhWLaayeM2VzOSckBZQy3JTnF+EFHNReRL89Sb2knvUJD/Ym1yZo2xxjLNACT9zCA6yepOn61vBVhdkwnXxTMBekZ3WDYq83Pl0sQx1gNVN0Mi5O30LdmGbr+0muXZiTlUd6rua67WkhcSzY/V4c8MenKZHMTUAfcabC9OuNBQulC+9DFSn1JiRygeXvtDmXb/Gz/4YRsyOkpZ2r96njom4CjjEpMlWCUna1mcd7BnHDIEJrZkNErxM9TtE+7n8xM/3ej/DOn4RGqZ0QQcd70K0gTsoV+lbFtp3wjIGiJhcLpQvZTPFa8d7rUsbLX4kZvKFLodTaYHacRFZu0C5R0g3iuLfO8smqhcJb+KZ2W+UmuWyESx3Fy4oFZPsr4YNAsJTnVEoSgzEsBMIpMuiQi69XnruimXzpJ5QS4J/1bJX2XDI31RTd+9NdXUjM9lhU7r5UVdVSw9Nzr1AhqCvgi3sabKcKtiUO/rz+auuLRuxRdzXdaETrrwyxW5j7GJdvEU2lt6JdGxCh/LQU8Xr095c7gU2nwOJbL3bQDkc3REYt5q9IRTa4p5hH6OT25IfpYOXbjLtOopOkqx6Z0e+JO8DhNNGLXOqDrIsSaBrCsa83ovAYuTqKmF4c3hZH7FcRXxFGx6035etvDPVPmcXE6Wd6zC826AnoGHWhVBAUAvtsYiVoeVSL0uYAtIZOPmscD6tB9DTTuPJaPXetNcVDresr3RLcAAv6caJx9h/EpWpivK3Zr1LeCMTDGuXJ711PYgHGdBZCCV3By7IB4wcL6PVBb1rAFHj8x439lEu3m41BxI71KQoIsN+kydApAYy4uK9SWiW1kXSsU4vssjMcNuSTwkH1vVujEzlxPP1lNIjj8QIC4PtJn0lBslwGjT1nsc6WlP1XBlh9L45MInZLBLxwYhkbyQV9f5nS8ZdKZY+yQnmCUXEeo6UaLQzi4NPQATfSBmhnwqBdSBI2KN7x511pIk31vZJAyi7YO5YQNzbbtKn9nhycpnYj7hgEzRUi08I4rQ2cOJ3w4QS3Z/y0DAZ+eZZsPJtvxTJJV2oeU4/cwZKEj82oID4t5vzKiA63ZBMMotlMfXTldCXs/uqJNrvR/XeAMNIWfhY1f85FXHlnMICAWZkgz+J2N5V/aPE/YvnK1RtJL38EQYI2IoCt/hWY3KgHOtqyHS1APrAu5hL/Rp2HfmLl4/nGErGz+DE0fl4a4gXQ8T8AKRLb4Ja/uHQsTJ1oB4CKNIcku+dVU4K2bq5EpswC84XvgPEF7P7nDeh1cE5OT+dZ5QbYHR3BNEQObWG01q+GQk0NV790t3mkvYVeHh0U5WT+b18AHIXP+dNJsiWY4J+2P7+l4FkkaVRL0h8PzUXEyWRtgrEW3QR9XBUrSiS0IDhCrtEN2cMol0HXd9iObNoCN/hPfEDgBR/iV0D5wZtk5eFIjBqGVZTdJPGZK0RcMpWRYxTkT7gIS4OMz9gUO4YxLNXgBc/XCenkgOe1j0Gbx+f7QCBQLgGdInbSVkEJQ2HQHNBkh2kG/bUXlqWJ81RwnLJ7wlRNMsc4rju0bcSgAeWgK4ghvsUc4Ep5BqQylc7H+NAkSKX2AnxZS696Bab1AmuJQDiiX7FAX/sBtmZyyRxc6eZnIk2Fpj6S3TbzfjuJlqSdmWN/DN0ZDABIvyRcBSvgJyn7pYdyrloq9t9by72cBLgHz2DWHhQ8IpT7RwhWc7InxZxIDbiFcY++xHUPjmanbvxhbMc1eA2bdmidszP8OPfn893kDJcQoflPXhdB5l/g185K690M5SRjrvGlNvHVOrH4a2WTOXNID/z1ki5M/lTR5je69bpUHo3uLN6Dq9/L2oscmVg+fCVWa82aoqFH0aSTXusbatnOWgo4EKMabtiGbAZczVu3svuS7MGDiFlZkcuiM2QkhJartADjn48mLDEA/O7UqhNnzb+FKY0iUX7A13p+f5PHdNUYbc82qVkp51Ekl1acGJ3OhTeeK5u9o7vmOze5c4u+g8Is9uD7/eWBNOhxkF3yr7fGwBFq20gq1QS6bh7TR2qcgb3wuDIZ1Jy9TZb1kc1byVgElmZEXRYsrQgJywpLOuyK7U6H3d5e1YvwZ2Rw/CwT9pNEEq3bb/DIDgXXzJwzIS/epoirw3WWNX172W+OrEn2RIj7FODaqsx9sBnor3LCy6+vOMoriS/k5HBftopjStPsl8S6Zpy+qlsWgkUWgOI215h7wC6byM+oqP+UjSgohYnxrvAjjSt7AKMd+yXCuBdHnl0bpjgnGuyhRV+3QkZaycH+xPXi3vLEDRSKmnU9cqUZk5R/7rIw9HgDzwau735d6NL7eXyp49nJeZEA9yvk68ARral5C5zh8xWheO0CubJk+FrdNGpHyf9V+UNSXDU8PL/DGswjNTDeMExRR/3c5w0C3Gm33rDoGutAIDI9WSpuItJgYO0bnUp8dqPc2jdQERPMoBybSjo23mZS5DHdcdJFeOSYS0jxEbsdy3W3UKYtUMOAbKRFVDqTlZR/p8mH8GNq4bc6e0UDyxvri51BF5uQugboncJkr1bBRfXuz2+vDI/KQdIvffc+gsbSkaz8XwMaRfIX7zhpWmIjX++3mtHunnnXds24X+mDt/107yerjmiXGsg1Hf9sTZPlV0k3MxHhlXTIqEprMcJcX6dEBzaTUweTDNl/w/V4jYuZDcgJ56g52yygk2y3mn17rpACLe5Ut8k5Mi0kf0TWfQQMyWq7QVWg3DuuoextxAjWkCqnygibSBSuL3s0z/rl0yojXqF38jCG4uJFlmS/i4V4d2czqZwHA1XoF71OVwfLQcS1GwVhNk531dPgl8524f5TpFSVZj50oFw8x1IulLdolPMyHe4ziBfjroJYaiQ9pjHRvxJe1SRuM4MNLG04Zs9ot6esa4a+mZnW2Io3XhP1lwMSSm01GoJpFsAJJ6Id5IzH5QpEM1v0EGxgx1o+XRQdSRH8sVefjXmZv0hYPhpPnkj8CCvICnVlQXS8fjNtG4s0MkqbRwto737b0Ru1E5F96JWW5GsKhu8H/S6pzNKsvDhzfETozkN8FPUuBAMFvVTrw9ixDplWAZrNP97g/fgJjjRNyY3tJbdqxdwUqTovUGtFHv+lq7sqbcBbReFtS2z/2qjOqjuVLuOy64o+w/pjqLL811irKBA1mTfLi9XiQvSi3SPi65iYdxO3M8EOfSR8nvj+nlXw+xj0ykc93b+gheuenpFtD0j9CKvPWdFm5Xe4nNPJhV/V+0h7NqCmwGrGknTUMDJg8eMfN5yJrhLnP0SHwNd+KwSbPlc8yAU3/6n9MavLBhkqSspnzkhLlkcgv8BZTIkbVZIBfwZ9GMCq8zcRS4ZH2omW8uOl4cS3PNMDBhRlYI1jHurfMm3fB5S4pL79Jhv2aru6ZITxOMnWixn8Id+qljfjbjmTYLowmiwz9+IpqyMN+RhTVYZpda7pw25ozBla4FSmVyN+sTH4k1FsZyTu9VLLC1aEz1r63jPJxeHGVOXr++uhW071+fxhW9K5+slV6sS+7hfLhCbVu5yDJoU2LPEEB0Yq23R5R0U84FTS95FtRkD9L474kafnYWUIj/KSY/EQOYqfMoEzHLrD+YndsAF9ZXnWbvC5suIgu9OMlIS9qmNJ6YXzp9ugYFMHqfmV77kBnQJc50rAA/f085Ff0ePXMd3cQn1Kl+ofLWva4w4QpdWcpILiLo7D3yiSwLMM8ttvHohr3Ix9m9952qgIPHA+tiMzYP6y2rx4qr9tQ78PZvgphtfsX2ubw5GhnTgwtln0ZoLMBksw5bYCMlXCg2HqPavCyiuN9HN0WrMjnQfRb/1DexRt9D7uwHw2na6qdGNS/vM5qRuehnulpuFTLH5FnWl3nCAUaeVCudNQkErODURBo60GKhrkvAJUPZ4MY0fFGUGJyyGkwblc7lfdrPYugoZ3FvArP2Q9RYxNMTvznknlj4NX/zq/p+7eVhY/H/XSIq73b8p9x3OUnCvI72EUxtK9PcPDZarLe9mzurzd93DpUD/YGVkKZT3yCjbnqZM5AFP14vz76TyjFD1PNwJCAJE1P6nmJ+jXB5o7kfY1zJvRWXPJixGSBq9C4Ah5HqaY5WnfvEB4rkuTdbku/bNOlp48Gv/pL7xoc1y5Lv5ZxzyuWMkx/HzIY7xHY+GosmwlofZuhJXfFnRqJHksApFHFdiUaUZ+yE1CkM6Fr8lYamlq0EcQnpgtS30zbZNjlbyrzWkxWadYeumwU7zAeP9X91KwNHz3NVL4FZDUa+fgR/egnzdBs601wbrsrhNF5jbVC2R8yopfqHblzNf7mD1qVh/6HlvgAisavU65CEYPMZ8z5uZR5uYa9gyMlUmSGl81ryp12DkYA9ARDaTi1YawEwVrsQGsaLAcX2VguuyalWTzTiYNyjrSRzzI/BVdZiubjwEIy2FxRsc6D2HPkawJWyZEFMHOwH1W5bR2NwjXI6lKLC8zokyfMxAdFy47xJvsuyQUfl7oO2YK2EFhVh15nCloQb/8tByGVVwIHoLt0tBVaK+OaVkSDs3wfPLl0KFkIpAxYOgxPDj5j4kYV6C/TQskd4f4M4QiEsoxQPCTZWsU/vCu5WG3fMkYeFhG/bbIU22t1u9simE5OwN9ouN+4rDyfCL/nWYuTNO05MSNGTkCPkms1BAbrgfTkH2iG8pWvkK5f+vdb1WHOaN7wShC8M147wCEkyEGJQE5bnlDXBSz3pe4xqVA9kT/WaPtbrzunBQi+ymJ0oHBG5XFsE9mo71HplxrozoOUPYTD+vdarBMatSl6hoEuTA6CPypUcBB8ZpAMCnM06RKq1Q9G4nqYJkOEQO77itkSsRnLlhXxXVCipJt1ULUFTxq/ka9/ehkMKr9LpGoXiRcfbziZfqf4VTIEXzNsQWrb3oZgEmPVI/v3Uo8S4AJeYbOpCz1GYMseUB3wXHwckaoXPHRQupS5TuVuPAsDa9bd3ZU9gty8H5Bd6ceaFpNH8gzrF/AyYkJ0fWwreRBmoOtFsX/08YBtf9ueCg/sb4KHobmS2UOWMEWrjFOsORVLg8GhqJ/Bq4IfUJHfzpMQbsoO7/UeJwRg7V7n1ZzrUQiGfRONuQInsqYyliBd+cPZtwz/REqCQmUoIuVcQ3cyPPqOoj6hkpVvwhz57OZmakLkekX9RfVX+Y5IVu4LGGtKLnK0+6O3mfmQ731mUCT/Pq2PY4RocRQB7VmusBnFsgILFxVy72XbnSvbbEwWVUhZZCPOqK5TmXVBxh03VKPmLF7M1AeeE+OqeNMj2wjoMYrEocOyZymqCHYD4nJSCa2W+rvqGqGwY4fxqSD/Bt0XcK/a43mNcqvkyBu49//9Yglk1aCsSScNpajajnWW8vXM/3uSiKsq7JU+/6o0vCu9aT7MQqURpq5020boaBJqmvCpe66ZaVCN9mJ3Qg16s7GyG5kW6do77yzy4udGRAntSYu6oAqSFhDrLnMN6IbtdMaE5V+7vhPJB9TBCNFseGxKFrk9DI1olq6++QJCA+vtQ2B9fnbgJW416+1VMeze18LB1RJsWLXbu5qS2ukSH/0c//2XfnzpBNtfoO8TRpMbtZbo62zhfUbX48kqhTyDrv7RySHnlFy1WO7I6CNAaM/PewjBrbQzMqFqoA4uaDW5HE6KDYXzPgZ/1/IVBzlxCRGfZPauOJEjEi+uXGLlo4bUzWNcfo2ml4dTVkPAavE+4BQ9XIGT0a2bk5gSASOY6PNqr0XDiqGAuKPiB/hNuFQd7hoFd+laSauApWKkbylU/otOSshwCucEmfx71nb/X1RQSrVgulUfOa4LJTyOgPavY9am+o8N2TjxluhITJYUy7h2j/mvJYfFnAKfBvRfXCTwr7MAoGjpbf1sTvqR31TEkti/pmvV2ByS/+EIbLTq+ItpHBIDEXpmGOMZAT5CxbzwaUhtkRrFpmtssbvjzZkK61hn+WJzxPu0Ox2ZzLtEkrRth0vnMKpRrEyEh2s0dEtTZ2RYa3CkvWTV2qyP98g3TftkcaXT2rWmXOVrJzENNX1T3kw2KvwYmVfREBUKfDZtqLt6OYkDeD8alHSnYi4k+eGqgFFzrhkELcOIJooj7H0hv6QBc3/XAtmSvRjSzhvunoRpbeh9QzsSCx0q/UKP5m3vbV6zfKR4mXbdON1jSZG+XNkXJv/z3yxiIiDjVMsgurmlxN89sfr0l5E/jAuirbyENxnKlLZUquJ+EZY3mPAUY0mVFmVop/w2csyMNwQZe/X78eieh2MTTxXWsSw00kmttl8xtNF2/tUykh0yCq8sJ3O4C7gwcJ6LKOuUPSh7W2Yf8aNUeonNb9XLMTbgPBrLXCxl0z8LUhwnOvUTSJ28tszE2+t1uaKGb4CdlAB0V8RmAHP/ISNxrcb7bTknu3szXS0cEfXZnkRXpGiGVHY5lTx8MTmnE3D2z4ONEUrb3k0PlY0omjWJ2BORYTDe4hrMJhDIZGAHsi+WNrYZGtjgTqcqCuXfAOROvGCfxi120Y43kJShCUegu8M9u3xymiWQ1PIrsSayDdFSMALJqjiRVLqwyKbXiaSAaDptn0/mt3YOVIynAx3M9HNjRDFCfa8yz0yGe4YK6b1+uwN7nPg3bMndx2Uh87W4EQagGV+lkSBcJh3hXNFIK4kEFwGPuuYkKTD91dJoiRriOr0dO8ZYvSIqFuSphfxpayv5iM3Sqa2gGQtIiQEBBoEl7T3YHgkP8suX99yz4I8A9S88Bmo2TG4iWn4niv48w7qEAQZ74Hy2isw0eEIDQYBcvKU/UEtm9pWcHvsdEzHp6uyVJoTbOFhzhRVBX391hBZb0yNhGcC3eAPVAf2Nplc+fZSS752TLXGbug9/DlX+g0SYXXz6Xu9pV5+vVx9V/VlTwOO9PynaUYe1zxHHhvOJzWmtIsuxmUMWd1I/VZIoKDHHog2D+o+qsTeLUveTPmJTD7FrP5PE3q8RGvDm76z6T56MAdFjjVo689L3weBBPFQ7S4wWzK4jUV5mGLS5mmSaBnrgJ3eJldZM9dFEA5xfBNg9n3UQNR91x4Z/maURIwhIe6m1Ged2NL5xX7+yAZAuP3XG1NDJMqDWwG+4msaAhVZQMn62XN9usK3Bx4YbWYwWAPc0OSNnn83ADH9ElkcXBp1SNJNXxGcu7LJmjBMomOtPiNO2LB5OLusZ1eVTVHtT5cKzYK/oTFiO9fN2Mec39qBX6xfgXgjdb+Of7qSichHmA0qqceYXfkCSSSVECTP8Ide8QDPSlFEEql3WxR3H3kWqtRoQ7XQxS8ExvtRnxQsvW54nKnwGpM7BSUNKFSDvmc82OaaiHt2eoFRslSJvigk3c4cMXPG5blsrcSjudgmL/BCW38M39b4tBZNVIwXwtTdj9ock1Bpz2ftsOkhn3U7hyg/OAsVpuA3ieCCSqubJiQoGJMHOXQOTQgAyGunYMSjODeKS8bCYoj6fQK9GkOz430opMl+HDPuHjt3OPrYf+4DA+ehCgkelPMJ0EZniH+zeil6uIQVdWk2ipIajE84zFoUMbPmXAPyu5ZSxjbZg1CVS16PhzBB0bW0f0j5ozbYI7WkVC0p7U5Pr6siGprQzRPHvhY5BvZxittQeYhcNK8+PvoN0tV2RnSviEl7AzZpNFEA5Oqsc/U5sQUxnX/YLoRHj5xg1l/70M2F+Bj5AQGUWpdcW8qt8tKg+Ipv1qnjUIWB4jbaAkG6KLeMr0jp1J2E/daHGcY6KRUHE+nNW7WakTzuYDEhqnLwwAKOiPvsTZxKgI3AXGVVgJHdKdmIBEC1MxnGeJAV4R+M2/jq+aozYki+eDX7DVWzjDprk0t17m6zQyx6UlbiFGTfdy/ORVm8coTtMhwzxFb5rZz41EL3ayPrToguDqhBrsWMjTIUPC82EXshZWxh6Pg9T5I+833dWTl5JEcZ1zNQ5asnhreCynQW4+qIFCnpntdhSsRyc/HtTMpL03w8v0tc5sfDQRPYTar6hwTE00aegqj2T09wEGSg7FUc/EuDgtYseyHxUguBEIBMhusr5ko+mS8lBiCOBgsM9dDoWURWX9YFkWwL5UcbVCFPrtkGcvSogtqwggCrdSZ8Jd0oRduCmYuyKz278CtwSbgrH0FAoC9NVYdA9He9bHrQJArxYqcln2LMqnqYlRxK3LgmC6HW827Le35Lv3hIeZ0dM8b2me0XcUCYlS0RyGjIN+BmfCMdnR5urZJYWjuOiHkEdf8+BkBWWdQLYQ5P8hmYhQg6WPv+NVZHzZNkAvmbciBfy51qj4xEdKeDhMF0ksThD087j0FOiWJh/IHPrmdxypVeSJL8qWO6LTNFwScQObuByFZv/S0aZErQkv9rdHsuuEFQStONpbHWMSnt/tebOuVvhFDyIgndCko2KnmYukgCvGK7F5YrrTKo6wxchQEkwOcgaeP730mdR4/pHfQXYGhC9DUoxb3p9GX3JtGVyNrOTXlQ2qJSbEk+G7rtW+sbgCsenNlrqf2xZJiBtdLJeNTmp5x1kqK4AUWXI+BvnCgMbbgHGRdZ6DNKpJfIgqszNLbYZKCQCNMhp6Fird4+fZv7wPyCxfohxaygkWWayBMkfPknF9hPt9eft/KAGkUh8CZ1hqGJm2HHqe+aGUX61f6sOreXdazIeGAmjIp5j22GH5eJfMGa9XBKVAofFhVu8S45ark+7oCHkoSYCEt3IcR1MoWDKu2sd9iaBUDdU7KlahIcHUKy6Oz8trMtMn0Ob7o+BLm30I1Ur8YlMT3mF7xjrpy12f2kgQPigpVZLA1y/sK8KGOQoC6EixvdxotStwteH+IDec5nAl0wFGGAQZ68eTLJL2pS0O5y/U5iHt91NOdBXDKX+8Uw/maJIiOW2/C86qPkgHmzCgiltegTEgno3bYJgotUZDRnb5alKlU5de+0+TaTOyCP5SNWAN11/xybhEsAarNh2DZ7eyBa3hWvFPGHq8p1SgIyaXDWlpzjbFXkOHufg8ccGjGwC8aLFylTdn3GlAARXoJfgxOnIEq/Uua1v3g4qMZrGA6Ia3yOgw7LAHfj2pPDPoQ9fKiFHnC459moYFzfUgp487YFsUYNzaT+rzzwhHr0imZrBl5ikFdCj8lOdu2YFMplCDPdEaqBQ6jtlczvdlNzjqSMHosqgou9FndmWKeW/K5pLLy1Jekqj4K/07wz4VxIvNYeuXeIoLyWIXoJcC8cQw5qZFDLzjoc/kaPOLM3sSvd9yPSM3ZEZtFTEQycWYFAOm1wivM8laDSr1aJTYMJWCJmPJHmq6WB9ExnyoTELRGcPmDtXNqY+Acjmwnw1dbpl78n9LKOBFyOwuIQ8gwpwBGHV8NdMBM0pj2XLFdJwl9/QE++P9XLBltm8y1ixzMMFAH0aR/4UcN2xBy+hmpwpdcG+epYMh4MHpxRqZf65WXB4Q5QCb/sIoQ6D/plYq49QFnUFwugvD03+wDQ0ZKB1SiGKEh4T6DdZRY8jXqu3qCpIn9wrcjxUpFS+cdGPfr5olbd2+Wh8zN1i4g13WTQgmbK2nWzKodRZrrlVfKrBiFkupBNIymYBHn2Cocvy+8hNBjqvqUGiYwUCfi1oNf/l9B5RPVuXpmLw4WaGJpKVsO+AbHxeo6Eh9tPbER/n3Xaqz8VMmdP6hAnAlIXQHI+4xqT5dDNRuKUvs6dNwrQ+a5xRiTndpIxAxG8iIPhWCGNPvBkIww9vMvfPzLvL7sbK8Leqqpy4PlgLRFE6HlVI3/IueYw+4PDZPR7pjjFKR8uu0OM=
`pragma protect end_data_block
`pragma protect digest_block
f579a82d7adbdd2198c90ffb9537e66a506b207353fee52bb6671ce1be2a539f
`pragma protect end_digest_block
`pragma protect end_protected
