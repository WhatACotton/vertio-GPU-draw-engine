`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
S8pAblQCVela0Rsko+MPCfY8N7FfA3zCm2yBJ5zzT9kfcOJHptDgfcMe7MGRvpWuM6SEWHWYBn/mbUByfvXCR1NBqwlwT43/afeTXo8rqxao/ZB/fsDAsU2xADLIg+/Mj39RpTSfWgbxPVv5TSm0znKY9Xxue8wUvnQoR7gnLcjYCbuNcfXEYWwANoj3V5XGkvw5dcqkBAMvFO6jX+3JvwU4EtzNL5AHj9q/AlCTUmMQCx7IwKlc8IqV6CMJsOkg0I8rz3Vt8mnE/ikhvIPst88enVxv8naz0vTSqrZgMx2HgIR16G1dQ5G1WbsGZYfknm2wWOP+h7xvBi0V/aIXxY7rRk9ghFO3qlcEFX82KjH17Vyn56wZ2BwQ+j9NqA4LPvgPLq9x90GoovxnumAm0KVVWRQklhV3L2ZzarFD3C2onjefOU/cDPPoRfDdyF6ls5Yf19h4D2ggOoCMcKe994Ix4kU5ZD22jhJbM0NAjJuxQuV0xs5D2B3vDDvqM0npmoYB+1nD3NSRPpKVXNLPUT9/COZingUSGsPrvI+kcEfGpoxtvjakhrsXWgqsmnDmYvOwDcnTrt32fUHKXiEi16JkTxdP2JZR82ntFEkuPH7lBRGdHILGI15MA7puS0SaSt0kCGj+6qnoZMUauf/1SED49qS5EI4MzJCGtiym23WX6D7d1sUJvhi480h/TP3rzgGiSpS55U01PW6T84+amGabNHFPQwAykVjrES6iKaMUsWhKYa+h13wCoKtzjQdP29mTvKHj+hQOwiEqmxNnqljJwSe6I3LYJi45g9m+HAGpuR5xsOKXTKLXPT3uPG7nKq+i+DDIb45f392N2ZuMOIRim1zml4UpQpvF2Zzv1myPfQJMUNxwOlb74u9TucbRmuMQmHVlEHNxBlIGu5XEB6c2hbOgECPr0zzTGe7rH9DAbT7zemem/wPa3We2IR/xEnBvI4FZh/XlYt7TTdZL+3kUZRDBaTlUzZO27lHQvsXHZAZ3LO92REDZ5jiukh8cS1AFo5p/4DlMFy6gUDb7t9Z0uqr8a/ZmuAN5ZHyS1k8nUdDRYvYxLlwURn/h3MdmPWoSa1v6qXfdItlPsIw/JYsSV4+WdmVTKcgp7wWVlGRKipE10WUhuL+oATggFDAU/9xDA9rOhpTp0mLDyLCZwZqOga1Xyvj++lTAelYCvWcWG4cOSKQzl2k1YRO8XBXDyI6DKwi9Y92aYhIYD6k2gq07ove531pmm37NAriOiMg4oGHSu93Oz2RyQRU2GJUGIC9clCEXIChXJIi2Q7OoSX5/7h25B1XwvyzGiP8xToAJ0U3EyWEJXG4Zw1D4OmxFi54WCMs6yqd5ubRWG/NkMxoQXeY88fz1iCY7Y1Mgl7UYBMdc9cj1GUVNLki2XxIYLprNKGdj27jQ2DNkupJ3pNAyZOknpTd/+OIbtXridUt9Uf8ojoV9uQ5qiUWnUWh5SwXkHTyk+lG664Omo1KIRpV1CdzRwagAHONqv+supjx0LbUCEbqnbXDxnVZN8a1Da7V0RLTPkYAuFUS3neVT4B96KVSrcitnqKmg+yQUy2o36qZahtZOaftbKC0TuqDzNNmsr/wFWw3cHHB4BKvi4TOeN6Z3JjfCrEWtNjn/OoJU6S1ZwyaUwQq84CdyVRyJ80f3vWeaae28W2XSD/o03LxJep4paRJGmyvhFS6CxRvdZc5fU2NHbeBFc9VThHW26WRPog/ig415069m+DRZRLg5RlMUZ7L6lxEvV6Z7S37chXGoCye0nwQvUeXNMSS9eG3hXbOnejXwB3g2vSMxTxtdkFVdYtWSGTUSMk6EMU8z641sTBl5Nlk0Mx05ufpLsIy2e4No+FSnwhIf+tpxC4pWnpJv40Nn/Su+uDVAH9RsUGOuM7RM2PUiXGdFw28WITPUen7ufr3hwJ1DWDCZtD9gXfABSMj/nQfdfHvSf408ldNx02izvbCPQd2mLsnnKkFNOaApGucu9o7f7jAXUbXGB4MqtP+FbATySOJ3jCpoSwyW6MjRTIIcBuv7OGhfFeYp413EFAxTKHXIZaE5RnzvqvEEePE+1/s0n9MxDcyxJ6n6d0anp5Yemz3tuvX76551sfz5YETs6Ajl8Yb3aT6qXPZWg0cDN/7o5vgqgF/vq8WddutrbzH1kW8I5pgV8/EipfPxn1C3zYdpc228Yop05rTCaL0O66N3tuLgx+a2O52ng6jj34UwogDA/sq6WxQ6hCB0VskTcCaiqim6mdYTxnU8IZozyDHIPi1KecK6FGxOdN/2u7B4XBoWEXJQGEGMJL6SpAZFkGfzPhmSdVM/9eUSXhKROVqpXaNEM5BHiWH2QU7aktZAkswQge7D3A8UZxeAQpybKFDfFpYOszNHbL6C5R6WwKAu5BCGrcMZxJvjx1JNy+04f7zRf65n4V7ognEGvef3dndSdNq4SgeV85aIQJJ6PJazUXZ51AGLDJyHQD8nyzaD2VwVJPGKNRlodokywoipML9975c895jTOppfFsHn9axsIkxfsi6v4i0+1+pq2nkpDmv+n7kqFfx6hgvne0y5KA3SsFKRAx6P1HWfWXaAmvjU4qxdLLNJUrbxkGjz7odhLUGJje1+lcvDpyqaIICMwAkDOk8xG3yJRGtX9/bKwrEiHhL6Bh48qy4yr9RtMdeOYihC9ShL0R/BPRIG3FjCbsAelT/57Sb6vpfMtqRuyzO0qUWIhENYzCCeUo1+fV8LRJxXSBWDwMJUhpefgtf7yfxHyqm0XNAqGHkH2DOe9AR1Y2UH347wtuXg1xueSbTFu0715DG7nQ064BHXMcZhsrUmgzKwXv+sStCgVJ7OOYG0cvnqB5tQH+2fERQa4R9V4GFR+kW+T9vyezJRt2CnZGk7/hvZgaLZ7njFYn4jUo/KAwQAdszAJE8O5COYhLg+xUIcE5CSQRRPn/bv9PoomYQfgxrilMoR0/mKPzQBN9oAdZJk/c3hsjaoa7/CWieIZkkUuG8IS4juY3vDeMba0h12eQw8I5b/akMPy+5XhvoJSpbJQV4/W0tB7Boj7YN+pncgzOR8f2WcNVijDZpQovYohTMnjuk7ZXTEs9Xpx1Xo7k6GTIdOsRdLbvOZkPNi5fajAJZSnQmdykdBmL/e88xxFmjXbQnNIIJhmQsV5bmdtUHQ4W+QXZfLfvQlRmDzcO0SaVi+6WAEPJmfkoM3NXjHvcYq7UQ10zg5JPhipJ1weZEkMfHYBm6YuBSkQo+N0QWpql8BQoAu8mJsxViBxTc4GZi0Gc8j2hIAy+y8CUrzqI7PvAMMi/lOUgM3lYvc9OL+JkxyjYUmHeRTi50QNrhwDvKhmBjXtT5W5P2+hgPwd3M+pwN8Vi05S56zy2jFSg/lQHbd4B4izQEUm1HCdcruTSQObGu3ZAUjxZbixzATPHVq/0uLz7X3PJygsxMBrTUcLbebpJ6wbPKEDfj8IjODnlSerPH7gWECAsIraAI1LCybek3Y+En1IE+NcKRLoLbXZAtdGwWMSbUHa7Pea1glkBk45SH0QldCWJjIvQ45TjOh0kmeOLaOBD3dYDf+zh6SmxqIMFWTYrNU2BFDOTRhms/AfmJio0q4NraWBpbwAGqeFVuQweapXHiD3pACIjS0Az/vICn3gcFQVQHJY/RIe7fpeJaOTx3XdzkZ+fZaDTP/Y2xyAigOyUH87IG8mhOYjXHhCNHgET4k1u/I+fwmHNMY+csPsDuWud+d6P+5g90V+qI66GhHkfye3pnRd9hjHjJDr/0It0YrjzfdPINeFjbPFY3v5UjswRXmFU0/8AJ43mRZQMK/OXvYGGsaHFgKfUBcULK+fiWRO9KMQKfh5iq6K7YWd51CwV6V+TgSPCc8ouOu2qKYfVpOjQNrR0Guug4aHHps6xip3JSnxyAXIdnA8p2gHIQKG3jyByBD4EzAUuq0On3wvWo8F0wgliIkVB5I0TWsUbY4Qb0bwNPnOcjX1b5fEy0B+m8FCp/eMXoBM5W3HqGvavi9uY3MEvidFo/QPL++3p4qh4qn86odD6Jwms+0OGL5WGwFMun4c7qh2kwL7g9AXeKs7Rk0G/6IzqRfZOibIdQ4qxKLy+jkdl9E43HYZL0Nejjv8K1nKhQ48atvncfMtvGgOITargOewl51zg13G0fwz7Z8+gyzPL/c5x2xBxDMK4CMsTEVLKEfj9+HFVwZmOj2d7B49ovYuQH66ZElfgs/LvLM/3RNtF/VdIgVA+AcX5WkGZusfJXLzL8iSUdWJHHeUQtaW9/YBsvgm2K4Uy8E+qYgmxtoDE4KaONSMvRyo0OUiuJ7NSYHDPFzA4F0rWAouoCDZxbuNdh5HGb/FM1GCo5+KDdwf4L5wSJzzPzHGi+0Pzp6+F3U8D13MlawP+vkLlZJmxHr8REOQN7ZxonWmW4SDaaBjHumo0t9imo9vSUc1yFvniTmU5pW7YlK1Ulj1jOt0ngw/IMVIW62ZiUdFcGMAuINHYHbbeGnsF2esZGBMbGmZMhJ198Dps8P0/iC4fl0XoW/P0zcU/U3QWPCCw0ulDxx52/RzrbgJlNr/CtEt425YsdYvcu2XcZF7+36lM9ow0U4BUG39NRac+iRRTCYaMHikRmeQlr0bK61toIkYATis8mj8UQ0ANxbWZerE/EgFDjaH2EEx/3LYfgNxRMV7sDkxCKIuKMrMFBKgjCHxMFxTM/5Ptgm7+EaB3DqA0tDd8Im2jLo0XjYL67THsDbdcrV0ji9A0/qnBgQWwZctNEMrpHQ+8BlCBDUhqgMygiUQILF5FQW2EXto++Fv/CthiSpZP/828rmKvu+a/hOAulb1SS9yPTe4H8cv5sAIpwWIWwkQ8ZuMd7+pi1M/XcZ8P0BSt40cn5/R7Vm4mJsqTfj93jW31+MzwLoYmTELSCS9GUcEYDsHkpa6HBX0vPIqEV6cWBzG4a6c5yisjMRHja6LOTBV721E8EsMHQkYMNf7NuQ+9iZKw4j3k23cG1i6pqSH+DNQLOAue1TOhLfodh0C6Icn3/tpwIx0Kn3hVl3w3B0PmLvECV3dSOnQmIyl9YMsKqcfIEI5dCPLaeNsWdi4DJ2E6Hmz9gQSrT7h8P+cvlCOAVzlFhaP8Nu+UUBeclv0H9ojxsMWqXTSGsz4T1Olcn0z9YBaYTW6JNzMVspeED86mp4fIg9h/gvKscuuW2Y7PtceRn4rycbYFWr+50Ia85rLgK5w2QqDCP/t4NNj0tolCOuRT34y1g804FDut9xcp/0cqbCT/bohJUdzizNqs2NowhXKqCO5whlbOCjT678tlQL/bXNNXN1VZUQF0vYrikQImfr4nU6fz3JM2TcYi2JpIwxzZU78dNYWQR/r2sKC7isRQR4OJruKIXnuWn9hye5oeNpOdGj1Qmgkz5kgxpgMWCM2DqzFp0aWM8M8sK55gSiYcJdx5Sxi5ynejrDZbpYZ6ucjlzDHFUkoSJT61cg3IdJ5JFweTNwGz7wnDtvCadUDOKXJNrLWxmQ37Az1ctdmYuzhkyh/Di1LDEdvad44SBUzpNLH3Xfs6evPPhCajPVHvPMyxhGmh3LcF9EnGiS2e0VqED+kpCWbNiS3/gxl2fBHb+RbP9YaodHXPg0eLBBQ9LU57eh6tT26W+qRka4AQW7vDln0OHqKLtwv/8rdUG45NIn4gkL+tkTNDAYd1vzQRJtym1nsShNKvKweiQp03LDllh1zuv+Qz34XXUdCd/JxNbui9M2+UUtg6YAHLZ6FLWHWccH6oqUpkLTDQJhZKSa7woN41MyD/VKeqBwTTLQCkeq7TT9IrS7uLe0uUTsY1LHSqwp0afhyRjHjUCZHmSUtQ3o8pFPcBw5W15BsYppjwgagko9bbFO8U/MmEt5V3sQZYXwo4K3qMBhRUy+JsyMMlj6Q4P8LbVR1Y9HIuRxCDD9BJw88halytt2G8RVxiV9sKdKUIvKETJPqS6zkCxC+XrgH61951k3I0SdDgopUznRYZs6xUyMc+ftmGFj28gCD/LCVDCP0sh1wSoAkpXl+r/MxNqrk+z0ZPMIP014DqmCudXMnEZ6PvA0T987njpAolY4/d4VtxUxGRejU+uhFlii5WXoXF9pYgjaVLIvupMEYp0p99LqTqFxXcJ16+65h3XSrpbUYeiU66labhEjjUxpIemWX7OPRGtT+KiQdtOddO1UHOi55nNPV2L8gKd1hdD3dNQTSiLcSc0moju6NJ/wHFX5kOJjd5/y+5jmZ7mcB4OErt/CQeMAVkVSKDZ5Y/+vpGWMK5m9D5u9727gEjrlkR0StMkj6xR3M+NQ/YjpURQfMu72OyGp4dIz7rfF0RS/+RQ436ju6oqspLxRvNTI1pb9dH3z+Sbx7E0VXvJGuHUI5S9J6UqChqu5LEoSMxUxGVRpnEoUF/z0Tg5wGSJ4rr65LxjsV8DdPT0K+0DZ2UQdtosgK1OOww6TCg84JYtQTMJ8ygIn0p6HMYWiW/IRfN54v5Ly2BeBOQoYzrBNOTrlV1tRlnVBq1ICbiuwquSS2qjPmYz4/7DMomPJ6z7DtMf38AYR9r08TVvFld3jDvAw01NphSrPhF/QNBsQrijnvrYoKpc1GpnnunyWBEVsLz6pICEMhewkiOykiZ2FKQiBsewUXbALr0yKmMdAJUu2qybbusHUplGvrhabiFSrMzNl3IlZN+X5O+n4sJjgaCjQpP2XT4sAQRNXOnVu3Z6vzQastvoNoeK9dt/jZkI8sEQUZD9tTf8wOrnMNhYVb2vTJvQbVZntj1S8agCGIfrntbO1umlL87aXKqaXlGMK/vZ6/8dJwhtgPhetGfD2eKHyHaE7XwXITDk2D52lqe5It+LO0pheyR4pA2t5AY923nLCioWUtcmH0bXejn56shmX731INtnIqlt7zHCuW4fazv4C/zNGDDn50fs/IBAV44Zoz+Gy4ij1LSXXyazSx19D8f1TTEWKfqz5XKnT/Ajc9zL8AJTfQPB4BiTJk9q0hOreh8gY0X6fjyqHbHSYf6CGpPvjLwmnwNDJYhlIAIO3U8wQkoLMfbz5V2qT9plwXuzbOJLPOkVrZzuKnn72w/eaJOSW3+BFGZnSq/k+jkDQxABk+X4EUd0mF/m8YBqionIZvIp0oe6zB5eReduOIGaDvE4Ik7pc0qfS/qg4FYAzVrcv2f5Da2gOquHzzY35eDPd748nm5utTeTSeweMsQ+3zcVvI25hvujXuEXdOMRsCbk2pi8mcbo7hIwThPvfVdCf4hZ1kXW0Bee2a8Em7arrwSkXnLVM9VPFkK/PbtwuX3iMJRRq/2kaOH5FnAZd1Le9mD0GaQE8BfoNl/P9nlb9zOEl48czoI3f0l9kvAiYnRsS8DASefJQ4fK2vp/XwKrisL5FcElIeXeHbwl8eGtHwPPA8Svnl1m/O1ti+FCXmseukkxmN0Fo4UQEJS53NBT29T42AfCYeVcxudH3j7p+nwNvi8LoKdgv4Md/05dTj2ksj9XmWwhbslmYxh9y7Lfw8plurlo9gxoC6+Gl27VbYieNK22prUnFp07o29OpsfEbpNKT0P6vLzLaML2Uu3mOyalmyna1IUbYY+e/oPHX/Zkcjh6EW533fXfEoJq2SnNBPg/EmgqjisqlA9TpAew2sDkszGVQDPMU/SUynMB8+6kSxhoym7mrkK1XOc+6vFZjA08g50+FYjEDEhW4MTyaMidgm4gmGKAwoI7huZzqynapKr/aRWazvKvvI+hC7mkfuBTnjUsIhK3KXmI+LLVck9lUer3Nlq4llKtvAbg38ID/zcXIe8NClc+gNGP47ahgtYcpnZWltE+ZpNxZd/rANMZ7igett4SqOo8aSNR/7gTQ2szqJX3cWoue4UfX1qYPnnoYCgu84t9W+U9FmT82Ylf5afnjW99IdpMsLoKxfXT1q67rlbZ50V3PcsF4BUvbRJzG3t4sUUUbf97Dsq5CCBjwHwVvZ2JWoh2lRM1iCxWFQw9PMTSR+fnDzhbxQmlpWtBneFLUZXa2dYxaFCBHVRTFX703eTtJ8hoEZIAoRRycwQlNqh17VwreZkYFEAYoLnP+Pl1/q2EW/0JSvA870eD5dV2usZlZ+6D6pqB680qRhEunQiDg+t19mpOF1yobSALFjxANTY/dzy8y7r+ukRS85418bU3mXtLJpZNYQLHzqiJWlmHJAAzp5YXnYLb/VSE9WN1CvwW/uEm8uGKoEOpJjwb/pzlAOHgfFgtB4PRXGWd5drECqdNwTge5HrlFouHnREhXPTZ7LGBRczWKL1TYaPO9iULZjHbG841rTpX64pnRN4m7PMQMtAD0a4I3YFjyjoxtyB8KNgC9/ym/lPs2DkRAoPGz2mOaO97bzUyTRPvgi2sykKruTLkkCObDyvprjw3D8DqEtPoQc+5fB8LiEjJ8vs9AuWqfwU3shyO/jk5iPOKJwALpxDkHBCYs3RcEL1zlTZAcc/Eabu164xGGkEWsdELq9d1lOpZAtvWnB4azRmkKFrTR8Mo2Nfx/Q9GPA2rEupgdnBB1oTTZ4uAI60KpFJGES6gtoUWfN1ijL/IJ8fmhieV2ytE61IYe7IH2yaEfrrLSe7+C/bDDAmo5xjp3vOxeyI2btnPzUuVoxFU9IJ428nYNopn/GoKt/kvRrJJnaVI1hkRm6p3mRzT4e4kCfFLBJYQnbG3AGcWCp9d0wEn+3Ak+DRv1IOaOKZR2X+AIxVeNbcel5JJtU11J+OBqSld9iDik5ppL8jjT0w8Z+g+LJ/+KvJ+RTg8g3cmbBp6txXSkbt7xQYGirUbZ8n/5L7zEhLJBSq0XeUtKLNqoCrfZJh53oFDXy3MNbqeyzA6U55VgpLGjt66jEIUO6a/UutRwgfHpOGXF2oZ+HFY6okKSs4vOMaQP9BisUsyRipa7yrpY3TP9ElUDiXVEEQpNMLdnw2AbJ+7rcodCsckjcprS8ytRlACP+oV9KoN7miIAUbwkR6VRymLwJ5KYRyoE/WAjGnQqHMKFTEAHNKcaCKRQiSYpgotT4B1jNX9LsXhy/Sd25dYsvnl8XHbPB5xFG0N1D8iv6C17UhMX+AbyujdpoLEOwYpQTw+bBV5ociw8cAn1H8iIOKPguISLaFe0eQVl5qIZbYgCLQ1zm95s/RV59YqfKy2audycmjidWM0kXzDKf2o/PPPifrWZIYF6INBjcERk2Hj7TparQB/yVLvEBkBsst8ZnqyDlz3V30wTyGjGziSG4MP3YiXaaxHZmRiYegaqhnd+3YQzMGJ3bs3s14oFfcYP6p41m64Bv3dxpVFG3bptfs9A7zbUh927nyLUhAA5ztBTD/sVDKwywLWQ3sBxzmQM6HJqRE0UKwO4aywg5bNLO+LtXqLXMRyAETbYzCIE2LQEIZM73oafgQVflaph04G119F4GeNEq+af/ZF3wtyhEG7XxFc8FLaM9xtBYVdMkPHknJ1Bd1I5lYGRSwbzkXwgubBstkblG069ByC385YuHVZLk/xmMKDFQ0ithSBdQTFFFmD32rc0rkFdu9nOmFn9+jPWsOi7sDaes1iEJENGAVvsuo5ATh8ZmL/BIHLTaku4XHLbdlhlNN4Y6PKEBYd6xOof82AXpWotKTl/XGomVdyYqaQPh7vAwxSJMoplc3Yb3ZMDB86VDTGwV1gVxMrqkxQ3z9b2b7SK5E79BbQq6JFsstyenVVNqnSuAfcP1nkbudequGUiMnAQxiSJnkK7MBwOoO8GOSBNwMTuV/gV7YOr1i5z4YKA0y2wkw7xaF5BJzaVRqIBtfP6cM9bDE1OdBTYTGfN2FA4v9GZ07S1jOZ4VspsIfcwBmBNtFzJ5DvUsBkn/HkCiU0++QsUph+F//JO+GDl5G6fco5iGS4nl2OdecO9lBNly8UX8YO6qiDVb9csj0wLv4GiZmm2snHKjMXOORSW7xWMIVJGJxKGGRPO+Vy8Z7aBIP0Mxz+4Z1CHO2BpNnj/mdC+seklujYNNsza+kQbJy1MbcD5p2a9Nl/r/DfpB/Rf2lJkGdLp7TKYRlUMhgDiOodCPbEheMBte/JDUZN58872/EBCIj0WBCSC8fFB6+Cznd2fBzutrV8FkXG7CGkS61TrW3uDI869ah1E6xE6smuBGRllJbehL3tHriX4A0lVjgmRAV5ZwwuBPLgJFVB6x4AGexli/0LDCOkhS5oEYz+DrcSv94dv6dVzA9zuc/RZa14qTRnm87NpX7kUegJgQM1niEGzX7qQrFHHBan2ZnFGusXBZeMTycnwpl2JDRnc3YCsyxbJGUKWbtALbMwroOL0j95Hvk2U7tMkozi4FgsQueYP05NrCh0inqXqkW1PrGACUtg6EQJnqVLoPU+tKh1FtmeZir9jW5BE2upce2ZlqMsO88cLtSL7JUhN/xhhyPEC4nCvYAs66aaKBGPRc3iUAolr5I1UemaEKXRH59J9tAqocy//nh2nm5wRGPl1Sp/VA56nEDHJc7eiWgq4VcuH+PFUN/TXSYsHlCGFW+6c6dc5GTaJdhwngXoCjBJpliURcZ9lk+oRl4SY5u03FKqZUE5VaVELYRjE9SJdhPCzG7LZPkal9ceZ5z9A7UYUGjw1yoU2W72P6C6AS1UK4ZXJTtKODNJgXj0ssDGGJixim3LYcT9Qw8GWkmzAGHq86qpMqxb17OO58ybfY1AXCYkRDoQnYqwOfjdh1G0cgwJ6FoinbvAsP9Uq4JVbJtqiEJKpgOI29hnxLHImtJiqonsYry/qcCHWLvGvY8iNuogfztbMN9KGAaLGpWwVtUVz3+55sQu36k6wVHd7VcMthprJM4yOeCJd+Pb/WtetgGXf5Fh4p4jPYlSu/6TxNTvVGpTac8rD3NkixUS/5KV1YyovYptUkend7x3UahWfWFnk6Xx2SoYilLjHZ5aRpnDZGhRpKa7VnW7rhOnEEao7jSfkSTlMK2eL6Ps75SnzNpNJAXpOFw8pXMpQEI6P0RRup4+HfEr1J+QHDYqFaTvvkhdxvGIZ+6B+pCvclV7Km4wxC/T4F03u37SBYuVeJ5YQWgiRlBS+/WJ5NVP+pT/JdGTgougaMB+MLB1LKG0lSom+eNu8ViD9KTVWzePuDTylqSE2qdHX0+OWzFgSJoLw6uD2ixowwZuA6kltdILvNfHFFGgVojUMErZnCXgvo5YfpQ326B6sF7M3AJHcUf47Fm1bURXTAy42GP2D/Q2ZVsCLJCyaGVkIJ8o0ryyUgOkDDeOke7fdkCCMiv+vqcfbIC5SBhIUz9nJT77UNxiX89I59ZhCTPPN+a08wA0OnH/pSf/rpCqltcXFTjHjFzO8YHoR8/oh6dS2C/IedQxtK144FBQ7wqbHMMn4A8qb/by0EJ/d3EGXO/fzD79fO34EhuyeF6xN0gIlUwlt4uyfv5l5ctvFOR6XaAm7x6G4xmzH+Mwon9Giy42qCrnDGnPWxAHB3w+rs7MWqz16xodNAcY2nqiJJ9xJmGuuEIq+rypxuowfl1FH5t1ieDo7O0uNRxQUIsm9W5ibF9izqrDWmQCd2wWCHumBXMaRC/98yGV6OdF0CGPeo/ncxTNusBvsyLV+C6SBxELgK0B6lNEpByHR4Nzl0EE0NxA4fgMetYnPUuISXkQ0OrkQ7UQtwmGRR8VhE5gcWWC7G/Ata1YQ347SVZr60BMKkifUyoScCMqthwI8hyQ6c18wpKqp99PNBnGh+LHtIV4nZ7G9I+0RE7q+bb2+T1DKGHszPOiQYywCiZgN8kFaibrSlC4jdJSW38ySHBdUTZL1FRCJ5wC8LXwYPt4tywOxODBjPhouDrAgrccvlTbqfe97edADl2MJBh7S696hj3eE+WVhE4x9QjWTgc3Q00TyOT3zqt2T9dGnJmb3rCGYm1r2m1I4uL+VYKw24KoZpqDwI+DWaIcCoqALzVEFGHOkKpDYQj94HLQHRxF+LZEp+CtEpkhauNO0RQpREmuD+n+V0oMpYPHqhT3lCXGyM+qj9m85xxdXyuR1E9buyXCFhXa3Hs46oVEP1umvMGKVg5Q8q1Mfam5BLpQGR8EK2hPxs0014iY4oVBoIudvaQI2DNNSw4GCPF6xaTBP9MLWD96VjcKfNdk5CTs91kXH2grgh4ay4AWtlZ7bfn8EX3yWgNKQNyBonOpFL6Oq1kNZqwXK8CWqOTyPVoxEVRR5UmdF3nAgeVQgGUYLg6RCxCWb64/kcHugBN9ZzSwrR1VpxQNXTsXurJWeFHwk0kAveJwGBcsf/v5etnaTlru4ge7Fs9dCemKOIxQxQMonR4erdKpJGD0m/q4UqwHwLMB470QQr4WwGjGHScaHlxFhm9iyPMYGeAt2NZvYL6yuAQEHfkDhuHFbaz5N6Cs5fJBdEfzQy6qwjlmc7tgidxwCMJ5CkGQ2svaOVEFIny0BuuCZFbTodVbxGXxaLaDKreg5Ll7Qefg4k3mBMFJojE0w6L0zx1Xqj9EbaSdLWsgXA59IpzYyH4ERdRG2/wREa/qQaUZ0ftK2iaAPei5L7e5ohbyKKVC+MS+tu2LOeu1YsyacRak4Xx2BaGGRg5Z8utmnfLcuS+BjVpAjDRpxcpXqGZEO0zr0oc0ymaorKP/V4ES2QrVgpWmOQipsovIQQLBe9mygV0IZamAnPAWeAo2LL3XpbouMf3qf1yzwMmjUIKSPCz/0rWub6jWSvfxuM5un3dKXQKhffxLwWpyfX/pEePd44CCKVSUWkDEmjkr6CaagexP7s1OW62DGcCvmZOLReY1hZ/22qpBnyMYxZkC/HxJHcXR7cPAeBXhpKgOlNIPAJPcI3bud92qvT9UaAeARzgvW2Qa0bE06OFil8n52dY8mrvWqMyC2mWtBGWXdlNPjKdIyhAGu+YO2Kf4bpAIHyLbmtoONaWot3zESabQ0KlmeyoXDSimGN+jcnflXb6k5nNe0VhhvFl7WRRR/TRI0sAjsW1CQPFmnSR+GNKrGDp5RN3kxo8ubcDmNTPOkpkCuVeAcRTCZW2o3rlrJyYsSbydnFzsf4RNZX1P30mTESfxugsBSvWb/e9tygr8cspDSxVoJMAA+TRzuDS4WQKwWeYRxR39kWVrU0KF/mUGtQYdyI0C03rd2EOMmbFURpDHP3InS7Pr90CYWeRxQSFukYxLYPRXBwP205BhvRs6/891+47T7nWb2FvjP5YhN5hExN1UNsIpKf6XfF41s3Is5nFiqoZnZL5zPBvBRqB47Cf8eoBtgqjXM9qTRx4mfjyQFlW7LoyiK7PaBKaVRITytpKiZUHMMaAby9SUHyCkrvARTLEK+UMBOqPwFPoLwb2Tc4ZBj11Radkm/QGgMvozbwJMfb++uT+HD0nsshfYrBshet3GJBtfNNBAcK2czm8wzpjq1wZl3BeULMPL6TXFpQ1ywoeFU3D7Ow3vTGiwtYBR2GJvPoNUXLfQfrGB/JBr24XYrM64VwD193LBD6fQ828Qt78EM2bpmjDr7sjNbybGIiEP1fBBdHldl7nEdzr8Er59aY6JdDAA+ovycqh8HXgpbOiVKhKJzO8DyQMe0BuG2aRsfUp5G58AOxdkDSzUNCu3lGIjJ4WIgRPiQOngQUqxNa+snhGRDxyU5+P9G/DtzKCdL81KcaUChgpywv20S6awQAtJ9TgoxKEOcABZY11ssUZd3LgHecVrWh7eIteVJ1hR15LJYLdYuTszE4XHHBmVwejbMr9cHuuyctA+rQ1uFGgzsWmtoycxjcygHwfdLZ2Wbfo1JztT6GmmTpKoXTulLBb1TWMG53fSLwfMJdyGEU8i4z4NkV0yg5DXysuxBKouJr3SzDZDkTIoNz5I9gvYl0Kdpr+T2zVkyJLu1Q3UO6kYX5jzUpUXsPYyEy0pDVMwK2dORn4sVAFNcJsPU9yz/Z7L4LOv6z9rr2RHCMv9aRneYZFNefyEq0vdFbI1yGuBFBHr5OGVIV/GVoWCw4giYTBbohv83vPQgT9RuH49KgDkzGxIly7PMvJ/1DE9e7YtLu6oLvejh+0NAl4ylG7jTBwKeIoWhyIHIJR3yOVAvpqT9i34FrzlobssWtcsYnDzT9I8zCosvSpWW7mpBHaTewZ8qSVVODPVB4S8kDULjJFKlLuksnFR5KHthi9oJ65z8lYHxmmd72n9DBphSX5OEfXBF8Afv4yhoT5WFkm2hEJ0hxefghtxgU611msLA8mwIkSC2/y6jnjpqLmG7t/XcTWV3XhTEeRQTD0Jd2u6PiiP7qJWx7qPl4pyG2tLoMGep7aKSv1iRLt3gDAtRa9VePJgKZtCZRUZDVdHJgApypnFvpqqf5he2JQQtKxiojBtZNr5MlSsvMHQE1kF/63CCnmO/NoPrW0x2PaWus/D8GQM8pwsi89SF6Es3Y0Zj75F08n5RTBn/amLR1OywL51oi2fMopTavd08miCYj879dsRKZ1y9slHBwOH+ZyYXruwsHxgElhSHSHE08VnVh3MHmIUoKg3oMgzt/T87QY8UONru+C9Bi6kRTG+fGL2IukEWhXsybRXzR3dT3GkoMAv4m2b7trKc18SVcYBJRLmWChEAyKJPOyoVc9mh4y/SiK5WtAXSo70Sgrj1/UVFjLMDfyfJpo8iT0K8gmXQdN26tjvhL46Uaj6OF7YTIUc7BaYANy1x96xZO8ELC3kPaPNNtWsMta7vKnmJkHnSMj1Ml9LZclHTEExTgktNMVqsbZGiHN68ZBVlKdz/Y7aVJDPFryh0Qgz6ha4TdhNm2xLAGoy2W40D73HX3lwQR6Z2CknPq73eJ0TxXT7R0c1u3hpSR97Z/lgMUx2sv9zUoi39kIiSodDLfyOqdSDIqd1CBSWijA6kBQgif43fxtpUNprqytv8LGBRQrec+15PfnhN5faCHhbc1LijVaxHZYUGuOTSnvwTMRsY0YEyvZCiKUhzEijAk6lWrLlMH0fwRjLoS3QlXCHJEd5K+dtdR77GPEH4d1+cCtHqs9bUUnG7mQtIrPNYmI2pzHP45wJQUgwlVBvtaNOuWXMQSMBJz7QnC7gF9Ew8KJYjwhjJWSbTxo1Qo7tr4ZTMmK1ocY4cy+Padsqb06O54fNPWQR9tWPRdQ1C2Yu7xrqg2ME0J1Xt+EBdo+0Cv4XQBOiZwy7E8B0WhaaHPU6Qt32xSNSA5heGbEzYo7XiXzqcOlk/TKXqNfBURl+wCXNiGv716yOWjBQF7X8lm2E95u4UF9JzunmbxsxzRRW0hOSgJELBS7lyhfFL9xjDqg4YFJBoTf2a6MNzKNmB55R7zmeRobzgLHy7w75YkxZAVrCmQlVW
`pragma protect end_data_block
`pragma protect digest_block
d5450d2f901c6d499aecff562e848b29206b336b71816ecaeb85d6774b7584c9
`pragma protect end_digest_block
`pragma protect end_protected
