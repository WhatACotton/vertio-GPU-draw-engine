`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
d00yRNu2/qDzxZI84XtiHeRZUwUvSGmvAfMHdqrnz97ry/YPBlCx9VtuHRFtC0AU9JOzMr4yNq+W1OlDt1T09M4A8L7MsexqgUmgtmLBPSXaFWRjb7v3EAbpr7YHiiyXR+BNOUvqZ1CtyTiKeVsBAgVrRKTDioSa8DqSvynLTAnQvE92AexXDzNbDvlYAHmjLcVspVEfeI7TpMct/BZIcVYwF5vIcW6oHmg3rGWvHEPxqKy6cbbBGk7PNpVxHZPXH3CdWxPOqNpRpTRPbCiBbPdTG0h0KKAWknbtVtLkFHdhT7tWFo98D0jyza6N5ZKp6g7WZSuF1fy5mkERUd+BpuMhZYluVZB4jpkMgIzOG+UqdzEGO4uXTMJmlVe9ftCgAL7P35Z5M0hRv1lY9P+/E9pFI4YA6Ejq9ekTBiGYnnvXDuOKt95j9LgsRjH4PJeoXXFF40oMof8auE5nU9tUVP7MNnTnSeNxEbgctAvIwFfiUJyoe+mmoukXCfhcLMkEdTPgB74p1jKAFJ4QylFHHbv2JAA75hNWeMIMRBLV2CpNdCkVFjTI+8iMme2LlfaYWFFusA3HjJTn8Y5vV/sGGNio5W5Q6IZxSOWvvrQJnl+Yr4UJB1Q7s+x9sesaLFuJRO4Kcdjf92Mc0yLegHVVTDkiKlMowzoGy2Rj1u6cuQ3TjlBwFXLpA2AmBt3vEjvMrK+PLXBaP/JWE/GRO1esqlN4EgveUzv3+q6WlHAF1oNyxUD5ShJITSSsiXuhaX3OxgrtegoJmC1U1LCmMdDsSOIGCHR3jVsQE1vFeWCvzwjMSUkxrJ4Dptl/63Akn0WWG7EP0hMLVCDRn0fAi/smqSQWgzihsy6nJ8Zh0oUsflOvQcK4L9l00T/HdPcxYYT1KszNkMcASs4tkI2R++TELpHJydvNsAr0EPeYKw9psBRMQAlPzZOKM7kvBrEu7yXVnyw3+hzFRNjffB62OF9VR80vOMhinahjVBiRlFEYEp1GdNG3INEf6OTShG+HMzlqYEMtts/bUU+tdFKjcUpeSmlImGBD0WDzFEZDsVLD37/jKCjwmerQwT2qUh3ul4LLhXDFz1lwbkgOHBAUsewQrw6+cmI468K+iIPYSxjS8A6HzQVfWeirxZBzqnVzIRTOgYU79DpVYXV+FH6OlEu+axPSt/r6QWQRrAoD8LBvhozeGFxmGx2quQPc/BrsEyTnCkJfaOqzX2Ctj+720Ajbw9Mj1aAFz5L6B3E2RUngO/IPP/uFfraA2y816WuciacXtn85lh2sccAZrsdvcfcnaVRhGxqpi3JdoVfMFqExf22bqpBsWVprd9BHql8U+yrLeka6S3u8XFpA3hlUoeY6NNvmLo7RUUtJF9XwCYZQXkaRwQkP+GzA97goAaHKk8vGRivU1lf5GxsKY/UWo7Nner/oMo4TQznVH/SQMzkb88W74mkNSsc5ypIEaKzUksu2PAzmVbpOtZKda7fJMQWeEia1YROKhWRn4wC1b6aXC85jJLqC/93SxRzHrkjNuvv/5i8VeDFhQGldIB5HJGsL4lOQMus2aXMoQzkTHOGOiLyOBVZw43l9dO00Q+sUBWmoFwv3uFJur/QZ2I/EREUA5erGkP0ddLbbj9awi/9MC9G/L1cycpe64uhWyi0v+587kjgwiBCuuGzWIKy0Ib2Tza9571/36CA/0N+7bTV5F3pQqF7BXBxKeg4efnOtN0ylxLPbhx11rnjq2WKYI6nn41pU0wN5PywWb8GTWYKcYoG+i3bev7dQcOGO9i9CzAiI5W/Eu2SYL1Fuyi3jmL29UjDI4KQX8v+MPyZJyf9ZMRk9g7aUvUu3wm3dzTLaFrTFsBKlnG0vfw5pfe3FAF5G3GlbAvKx3RS+1qbJ5yHM0PC9IvDnTm+Dj0DdkqnlUOvnTT8hxM0VWS/Z/I8J1/scH29bOKKp6bQEDhz1ivLA1OaLOa7arHef+WReXm+uHnaYhCx7wRKa1aPw4Ne1WqM15ds5rgAZUcyuL8Ig4Hh+d7VI8zJfdlZEBU2wfaBCIyY0kGL4cgbyskfu0Ax+g5lHUBMD0leUvsTZnbW0Hex8EhBIX9UiNxldBl5aVmbWQHkEaTvkDu6XGvCYve48MfhhVGj8vuqKtXslFHMpgqq0jmCFWOUqJyV3msYwc0dN3KZ4xslKvFys55RZOSTSKJQBOsDP4rpULXnB2StCZe8/NP+VeBzL9y2nUhayVv3jDiWjbVkYYQyX3bOka+nFltiO/iGsbmpM6+sfd2soyVv+TnkQ1WKKD3X0Py86NXo2vVTYzrjQy48NPEoERXhdY7sTpCtal3ip5ybWepw6HKUy724dqEiYc+z6zNUIGlZVQReBjBOBogVX0F8kVWigcqqzBlCdf35uCWJoIhqdc2HX+qS6RWXthJsVU0hias/2AvSJr5PDGU1AEwUxXLF1UbyG45FDFb9bhZDN9e1SHwoVP/3RB2Vk75qcWpUv3I/9ixgkI9RavAyKsbHdmXMFKgvDf5bCYQoEL5PyfwTzzZy9yK9Y0gp5nNrvZG59K4sQ6gu3jY26LAQbS1Sm8SXknDx9jBoAlai/GO8HjGTqFyyo40slqEwPndPV7FNPexA7tHBI+IJafjqvwiVOEOw21zZ2PCWgblXZ2hQ3+IGYJcK5mb3v1/XXA1Dh7viOkYOf2KOmLBxEe59kbysUFAozh0YLqZz1mYnOZeVT7r2elx3NFWNyBW4IIe7K3bGrb/NwkE9ZqsTvlwlIr09/UoeDmBjs8gnnlKr39ewUd9AJWJLl6HXUR9ojyJfMccy1Wg6rVQUXetMPmtVi2jxo5/9EFvGBv7MGEEi8mu+mnVkqYmF34IPQtdY3vTStyTWUATm5QREvMt4ZIbPTzvuvS69V/k2sLtacgl5fT2shAf9w16i1qFJB3MDdYT9uRIBjFoV3xoHqVWi7qLUtZNcskEc0Osd2PQZwZl+qjl4iovj9mTQkGPLZxCIpzaj6cpKc317Up4tQYxdE8n+Ao76Vu6L25kwJUlG4l5z2aiaczKyTZ/uySDVwv5pEKIfPZoLu660s3fgnz3gfGon0rNN8BCvO5fxGCpnQtTacGZUamEbkyXTVIwUg/0BJn71brVL2qh58h0MmM1Lo+CIWWhkx7uIArubFTlYgpn4j57AnHgrcRNiN8ySmL4/341DZaom1WRLcTa1ChPVFpBt4ebYpXZ+c20on1Ma7/mtYIUkG0Br6k7gqblMvWxHTEUPTKjGG+zgOi2fZhw0R9+9A7jrSk5NwlaJp7vx2f6um/Oiyo64yHBgG2g09nK8T6YlRBMVhicgg/EV4M97TZCUGAafEbsxVSKNzkjDcCt6Q0IMdc6gzjklYLnL6PQXlsqdrQDy5hUMfYw4mc5NCIoaQF76Jdp+v0UPFZ2qY6HGVd9Ut4ggfdU/ICkLhLB4gFaG2a3MLl8Yk67fMfrpwQTrbFd3ikPxSoihdhifDnBbXeXX2Rj1B9ZhA818km+fI8cA2M/Ntw7l2JkydFfTJ46ciCbjGRonc9wEQ4H3lIFW7s1pB77GZQspZFqezYvpjM1LI9TA6NRn3O/MWLN57FKkJomMOu7ZE5rby+TfcLxvbRrefY+piN302P8MGuXZ5ID18YLWgV2gz7hwh+CZDIaem0DM0Nxk2DObIloF2gS4vs4qRrbIcireh54n8/4orhSBE1jvy5jA8juhMnxKwFoG5QfKwNbQQHSKi4OUTMc13qCoZrPjlz3XhlbmYW40/8iZoonjRNh9F23vWyPIszsxiYHsFJFC1w0uGAEg4I68eUoPDgQJecensk1EQRmfHG5Z6lqSe+K8G0dkGLTonPjdRjeKHAlTeJYjJ85h1wW9sx5fV1fHePpvKMnNj6ctkTwigZBDdqjhM5SxzTVhFS4qNgbs3ZOuH8xglC51agRRTteS3K5Fy0bibJ5OvDPxpkfAP9wlOSEtk2FXxTUZCHrl8vvjNcjNu4Z32Du0sAPWKZ9hRkjOCluAL+yW6fr6iV9eCPUaSAr9mROPx9emmGP1660Z1nGewnGSsiqnsFVS9gsCTAXH5krK44QbFi5GfhtMxDCrk4QIa/aZeEJwnx5bWgWCYbeXOGYYyhsukLCULgzKHFUIDaKKwu3c9DVbUlcV5Ql2KZK5rn8acrjyydoKV0hoW/GsHwwzSCzcYL4zgTRDAfA6hgMrjBrsiHtsT6pMRfz7kTP/3+3LMBnKl7SLYSPs0knncWBvyEXKTqI5StYuOt+ClYyyVYfF0YT6Pspb9YtkrG/bN54Bc78O/R8YS3SCDieCuIUzZKVoD4tbb9hrk4DgzxXjf+cOzUffUaQyAR4pYeqnmj9y0MeNwfs7wVFI1OfIaXxbTlRnWheX7tw/K73s0lM4bxpCXsBNN6rZk+Mk5XDTpgxAcX2djzdQ4jlks3soPKTJQZyAUZIAauZcrI+wKVJzU6+1cjilu/HHtt7otp8iTAaeZvaNukRkVWQwb+16wIM2AWMzkqoISIyNVIOyEJDI8hCOLqls0s3DYVq+HlUfL/ZxfBDSCf4HeeXAFWVLy4h/UsNRiXmHABxnaQoz2S+OWxzMeAvI/CfwzjS6tFlnpD4DPev8+ZGAT8IKVItYoC9XuvDOxf2ygmU0xd8dawsl6c1PYYwgavkHHEPpqQwX0NCj/fX2kyRobBRRRWknWh1iNqrorK8w98y00VPXw1o/78qwVVMV1QOhfgJ/IC/co2+/0I9c0eoi7jpEqQAgOTXHklsIQZWMO1+fxPV1nprHxBQFT80HFqL3jFH0UnJENQ5weDUgaQw2PgfZz0IBZClAfYoNOgFpPn8M+gc4JWt4JW2QpFH+i1CYSC5sA5M6783elI5ACgSnBrtVvOvW1sJS22N1cmGfy2KYhM//qEOdDdxjLWqHHstnLzmJIx9D8AxUm8/OheenKvd0kv8Yz0goAsiC2THw9SvUXAO6Whwjcrg16IrJ4jSVNqp+VgXiz4xPCuSVdk2xwb766sVbZmyZQhksU+cjj1NmaE42YFVa0fbESbFKADTAhIouubQItfNjHiwREFZzRwsX4kxfGC1P9zL7PBM6vGw91YS0Pa2woG6URjOpLt4hcaChceC8sWi956bBaNEbsux2Nr+Nt358KyYXYeReRGeYTSfz91UV1CYW9JLemgVl5FzOzl+oUVS1zBFNY0mnqHMbNFyCJbtr5mdjEiJj4kq6QhinvM9zV25YtIpNoVUZjQTZjzMXXXyVpkOoLcFbaIj29RUq3N2KTmEnlADLWKXDbUiQnp8NMayWcrWPP46cCD4MAl0jZuq0LCNZ8G2id/nqtWRGlCQXjb66VdojCZmGKAPHAfoChFkOmdA+3oGDlilhcUctuu31Wes/UVRoWMpqFpMqok8Nj59c1EI2TcZPexZUX/ELfQYRTgeLLncL+llTSbk8P6rTIZG1kJISZETSeTVap1mx9ntuc7FAruFdpnG6A8hs0KoyH6ldMqjYFb1F5WvloCsqPYYeaPrx02fmDB0A295ZeKx5WerjfRsmkHGpeNHccZQZzj7Mv2MYHOjhq1OQwehFyodiI8NKtwcab6ghvO4uq3I8McPO1RkizwMdVq8RrO2XSFmIGztRDghxEpSW2fGHGOO4CvMQp2t3XBm16cIg7O9jXEo6VgpUriuAx4KRGJIshoce06tl3hgKxsqn7iNqpXKZnfqxKkZaIXNAdu8U3v4WH1CwSaB4Y32Qz1bOhhwmDi0MQXetM5fWrYlqRcpBWCf1aKCQlYISYvDuB7HG//wou3umYl8bBOq9vC8tygj5YUyfGXSg51GPPkehEzZHIAmIjDukT2LpgMAJ5g01xihl3ID5fAWC7spKFCEC0PtzDUfjivB0rTgUceW3aMMm4I+6XbbhnuGr/jRmF768usV24AR3jMp4tm7ekvUd+0msiyukrHMGOIEg1aSV23W019nx17YkM2r1BRDD+q18Y8t2GF63pHmzDpdzJpLDuoxwh05k8jjFb5gbqD35udWQhh3/OYbWHT8BZix4Wvb91XghwRQtTnxBnlSkCRj27kkEZDH7hpOYrF6u0kY+Qg3QZW0mewhAE0fIIMc2IJkiXsPxpGGEsiQmsyui60mDPv391i3ccwVxQtfno8zON2a+0yHdMxNDaVyLld1VFqDbyiThry/XrpKvUialTnRIq0z0OkFPGA5zssutPd5CoOz1Khhjai0/ZLQ2lFwdLr4otRVwJM5010d4thXAk/Ck5m5pV2ZHOZHo62QXBpF0emBGDScIXOVytF8uO8p1O62DeXU2SUVYcrGRleCcBuy/cumYShReuk2rsEP9NqkDZXXBOT4EZZlba0ypX+vgt7/6bE04O2nQf3J5h24ip20RZXfWGP8tB75wVj6Cl7eKKUYbKEfJjBXubhx7U364dVQB2wTEfS8yPHb9bI4oOk/aKbagZttu0casjnGbxsJCRkd+ew+iciZ8vAS/zjK2HYNEApujghyPBY4hK7y7G9N9a/BZV8pvVgkEX7ABnEBKc09oSbE9NTmxnK6IcGv0b8lvkow8U3CCld9IeT4/63VO4ODQGlicib/iXld8DANao0o3GIamrekAafWz2ZRlb5SyxxETRbCIjsANuODqsFP8E2KDHh4a3N2ppxPpKWGrbX1At/NmJ9fh+Bw12qGD4XsJ1cBUXStqX2CQhG6tcFMZ3frfPuG/DjpGOY8OCqaU3SsGDDf+cMgJ41TKdXqJcgC2O017vhzghlcV2T7PCESvY2jLkvxa0q06g0qSEiCSwh6Cza3ZijiNcwpsTOepZiKD1W1vI449JtzHkYlF4LMMsmV060MvxveWvmDRdMb6a9TUCRxZ/LX5cb2qOCCQx8X+qaHE2m4d36aD/82ZJnFJ7adojeh2iy4dVHfHBNIUrsUYv7UNvZaMMglaE0rXK0g4z0HawjtkRYKbbBH42cEOE/LPwZph8i4MGOL31koV+oGEyQGbg262nCpCMQD0NH2Oh4pcKeNx6OBQgezaDsOwoWuy+fw8bvatkPgELwACXyN82sHLtfkEa0cEVyrLUV1eXMyoNTlJFuDjlxYUQ1vUNx9u07p3LyYzzn2q7t07qPFKMOHBqt21VYXRphCA9nbocJM1MDTShDKBTl1Et8Mp7IYiQ1bDVVs0z8hgfLkqRP9jU0elHceI2ZnYjprI3qULT9pfr9khvmyQMA4jR1PgZuEBUW9HtSq5JDOCzw1MCc0Rq3SL8bPoNz8BAybCXfB5RMb7D6F1QDjNG9dmqmEnX9fCjYqxeJGqy19Xg/XpdjzMw/4h9DlFnjx5dE9XOJ0MRODiUe/GKTxHc1v0zf7K16Nn6WiVucYQCCvBqqe2gM257ti/2vKZPWZ4p4+pujvIWme5wbF3Tsdr52eE+g9PCf59QNC22CB7o9I52eFDdldLlnyOKUna++kSyKmSNVeeIigjuxTV6CIX4oqYo2uBOZwsAKN8RG49htFBoe0g3HOU/N/wRmbBAD2CTk3oQFprghoEDHXH4kw9lYuUA5Wey2NPM7GKIwroJv1xUujX81kgPyF5vx+RuctblQ2dML3uIISyWioRkRn4cee6XDVCxpwYPag+SR+K0u4CB/vOB2aC7lawqzPK0SjDCx41Xr8ScgiMGjpqo6eO8x+WsOmpytt0ANRp4LcHUlLMEtSk0j55nXNQeIiHowJfPmkEUJjjmA+kXY1cM7wcdp3/OGs+I1dYJHL4oC8d1gljzEerEeybQ8ZGVOmy4n4+U85rU6oElnf+rrkxgXdltN31bjh0gRNgIJ0pmvuVLWLH/1fUHUEhM0A/hNrZxrPF2M4kAU2ZKBYWIT73HCrIAnZWf+k/m+z/cQ30Vs16ALYKdharexCn7+6mh7GFLL2hZQedZVPyuw2o9PzAEC6UwEDkU9/dKGih+ipQZ5zt6KXVtVSZMJkpx+iAcMZ/MRrCe9V3bDsaxuGdzMsxMSjzD5DeC1/mhfTRzGQHjkYilETwRg6+VBj1F8rS/pqvlZRDSa5aM7hj3JFo2BQ1f6lj/vLyD8K0VZ/m1tKRTuj0UJzaj6Wd7zmQRNaBcYlzn7ruLPtAZwyOIqEOnBBmZb+4KyItGEk6KQm+V8O3/mJ+OZnuMUoM+rsOlI3/CjtJmzbfaNC4qf4OZva+MpV64tsS7jjz7SyfK7lnLKdH5mNvHslTdhrUFTfuMRhGW5XQjhdLlk1o1jozdeTRq6DN4Lx+L9zNdfcHdcOO1xVbwZ8QKlJ/xQO26PLkKr6Hn+AxvhCYJaYMDMGOQkJp5P1GrMnneQ15aDNJO4lbCJpvvxNhe7aAVt/TnJvh6H3PSFZ/X2hIOq2TuUd8dP7gPArM5VOUuo8JozF+o0fXYrFmwVKm5vD2eqqwf8SFUb84xZuk/1r0rKDa0bSaXr4PYGH8Z15A8OUtbUSuRP2z9PL8AgnYZxfOHDhk5MnijqSFpk7CFpj4h/QOYXttQ7VTadtrSKrVO1KoBhAIdpdIa3hYnbrqE+PypFQcnpI9uyssq+JKGeWmeJezgNSIQ67Vl1YhZk+U+o0SaofLIv5cQIrEuQTwxS8rrDBj5SwDbx2ZtdM7AxTLvnG9VeUUzVo6FOc4zsaAVb+G5JTxS+qcxCj14XflPKOQC3E6JjyrPzkn/bthKyHZaPwTGAliNQEQEeDnIi0gAsBBy/5DyH7ZGF1dSJyEJlgGbcOPNLuFR8DF9fCCuatSksv8h1pfeRDUbqwn+iY59/mMMB4AY+CZXwWtBWyL+OttYBlivUdyo8WYXFI3OADziULIFoxUd/gIVhzIp9rnPytMwIpIKUosESS0uVsTjEnM6la/cooJYLTS737ImeOwKsj2YCUlTNEPaSo8XrGo3ktEQAmrqbeapbkupW1NPU/3idcUUXb1QUffnFodZcNpW8dPHIM+CLwhwp1e5OuSPILtSiZO+t+X7+cjUDZxiEmw66eCNNhJyROOwTLMoTv9sNWZJYrERdeV9VoDVpDz7dhsrdM25M4JZGAW8g2GFBg1i91sOO9XuLPbny338u9Dxa/snW26p3XT6iMsIxk7GP4hTV+aaiD5itwJ29T/pO8ru/3zykZC/RxSqrIeb70pbKSpFkYu9nI+d46rRX6m8iOnSnQ6yTyQmzUTlugnBW2pkfXcoMWqNAaI9arABCNf+LDKEKGvmOL6rGqDFpE3lJ/j/CRTSR0ql8UEPtqQGkH75x8ilcDUC4GEo/nKwOuF0weDfRlPNDuMcTgC4UVTKNJEkvpUSs0OXiTH9N4IZxfzpVHL7Qog1wp01Yu413mzgQsJvEcs/HkFGOwNco6sH0YnqPVT+DwclvgEAMWzZPPn2ZObNSLqpToTBHMQgAYii3jmLM+ubAXPtR9VXMHXuMnqcJqQo3SyTcpokDThSLnJFQP6siutHbWqM/U9Hd0IILdJVb8t4LtTY1DpENpKGphWQyw/WcttNBqGd2zjq4GetdPzexS4KO/wyn34FKWKcrBIAJMwrE7hIvi9d8qYpz4Baf4ByA6E8XA5QZkunv42sMCIdIzSI/BHvMPhAtvkPCXSYskRfQeDOf9S8wtd0WY+3+HdfD0tX3Xui27Cz4Eu/QltR5kYz3y3acOqaOBXHS1l4OAqcfyqxDZdYZc9/iLTEPoxUa4CfsAcjd8TItW59YrF1+VBEugD46XDi2pT9SGg3OO7pteixfUSHhsAjOgPIVVQflm4rqwamps4xOSnTjSw6f8yk0v7wAXI59B5AOYqWM6iUE61vhdPiHy5SPFg9w1JasRAVfRQcRPQVZGxK8SMglhmrds2KAQXxl+U4WkjjahJtdv3g8SKeuPYw7a4c5R7Bx5sUC5NXUK8vmMkeNl2vOli4wwm2xrZuyz37Iwl+KPlmV5B6inc0FP4KZkZIlzuI37ZGE59EwMVD+sRWDiIT/xG1g6M8RJ1Bg5bi4htLesFy/9WBsQXB1NjqQKzjPq9OBancLPaKMpHHS+dMFzCXihtocAsZn3LNIGRAWMb+8nALOE0Gj5LRwIW07+TwnOe/OGRnjlDfGnITjXxxzdExhz5yJw9AGjGgTAFvgv+GH6TpjrtbiV1R8BDqSR++iHVZ0huxsf6UbqYXQqQ5BYLflX040HkGQ09wqjSD3lUFqhlb0tZIZeeafhtaqoIOpxdlM7M039zynTNEStdleRMNk1IhrcQW3MPTjTvXDWougFe42Z/P9knks0zlP7U2D/ygILe+SARNWy3KZANDw+Iy5zZsk4ed1ppfoyaqjKHBcQydHTLvQ2jKqHGQazqUgzc3AgcZuCs3xhOK4PnICsRPYf0aNUV2cQrpn3mU665/YW50Ir8S7E5kOfPE0miOGeslDC7yK9YBckzjHqvIHN6m4Z8piTWMD6I6eFL0e9gC53vf5WbKLbXssImDvoffoSRmXVL62bktn9GAmRMcXiJz9CTi06k0gGysaSrprYC3QSJgb9X87uDN+1nTP2dfHl+ed/FxdPhHr0IBYSPXkfcE9CV1p2tBqE1Okbh8aLHNT7064oZMiV7bX/LeLFm3AgHqf5EJxjkqFwGltHwa6xoemLSdNDbQUaGPXY+DCJdBbK06m2qvYwM4ImfNMNyENh8F18CQjN0hhxrgl3gcy80ThnQ8KbUkzpCO00Ak5+eZKr03Gjm5u5SnY1KgKrgMlAl4/PTQ+jBAdsTHCnnEx6Bgz9Cpsyy8KcOd/9CgAp+MlnTEYl1PABK/A/zTAQumKxSlfPmfiXmxkWH9BMKhIzOtekCL5HnWeEtOCElMH0vjNNixZRNXnX6/bgg75O/YxPhLjltTk0+wlL53vR/Ps369FuKy+t7TC9XimhUwrQ6DjcNRPPOBfiC18mxbX3vSYXa0woZxsF/V73THe3BwstosPv+0SwGBAyXUXf4e//jtWp9FQWq9gby0oM6B47Yy2sDRsqZGmfiW3wCtaFqReLXZLvjG0zucLl2tgrkg8DE+xfV4oKzGqbJNJJMTCb1PxhJ+IcHM055ce6WSS/HvWWi7PDsqZG+PKjZSus1d6YJUlk3b4nnEdm3VhEwsvAmlk/o2DsdMHEHmNX+XMPrOt50iWlvkWcmEuFT4rK5ckMcSdD00A0wXv7EDFdF/MVJJMuFyDIa1EAcXOMCgLb8pl7zSEi2UNX1dD+9WiMPqVYA+OL3++IbVnA0AJba6quiZVw3nvQik8CuPb3XP4Lo88Ld6XbKF7MipBsDCkbeQbQ3bPpsFDCGiAWltDpmwqLCDGA4Sxde8RvF8moeMAdBFNZsCNU+g+jM/uZ7+2JuktQ6eQtxrJHmjCizqgMF6B5D3z6LknnUVJFmHeLwBYLHilGfSPVlpi6fm/mIDHzveC2dKLwZ2/tBti7qtavJDaZ+U/yG5i9sHONxzxslifbtuAJnMcgXvDVWN0cA2a+2HHEOe5wzYLpNcmVXYK1dOUmw5V0e5mztj8RuuPUhCudMyF8De2acigfBHOUHPbk9b56YFv33qX7c80kZPHI5k6PV/tb3XGx679OXoHnBD5VrW+CKVKMHzf3n9+7tKj1Cti+nitGWOzkWkBOILbfmlqo9tbMe89yPZv3qlGJ00uiDLLxoZPEhrlE9o/RzT7CtOYtADrBrU6mr6gYR0E/GC9JFMykABMqXQGfWYs33O+3A5kWwIrF/dBjJUZ7+7OS4ln5AA6M0h5idYA4l3n2/f9mLYioBSbz2CAv+tM5YWhdhjhIiDxyFr92c5AQKP2YvsuxujgW/lfO1Dc6p+3jfoKo+BCa+ZDr3z/0zBa/aNWmPqikS9wgR/AqNx5Ebms0VW9FxfdMAL8D4azLASW8zx1oKLn52WzdE1C4JzvBE0vsnY36Swp0pz7rt9RxV5G3s/VF5qxeHc2aWvfIAJLBCW+Ax3Y6GkuxxCN528Th27zehi0G2ItS14up7+lFIyi9hSqwcYvS3lTtaq0wH24Iub2+5kOQQWQdWq0fSZC8L8yu+KlXz1mZUuTbYgJ4kSlsCKOiZp14Qs2cB6AEun+o2JphuKr+e1IBF/ZTvMhqH/2XNR2k1Kwp9g10ZIsJ55pYNlL8MVSiHuPzURgUnYKT99wzPPpRUB7k/gtjlF8zGMqMRdiWTpRpgSuSSc68GinFdMKJIoHRz/G7BdaMApKVIzTqfUFOXAWm299y0YpxxSvJc8Ipi5dQ9k9NPZtIgcGNt7ub+VvMGwHxYyBz34DRA5pbdiIdAtcHa1h2Ljk2r24zC4E8z5Oc6ujBjHx44CNOkIkzZ9vQB5nsquXHDODptY4mfcy/K5V9Dg9WtxqlCkAS1N0I82e5Ioj7L5hQ9mmlJlT4ohwZAunGIP2s8OcLcds9KKSBMcmCtaExYxjDj+FtJEDyK5+RURoMV4nwvEsJPx6njpZ+BcG7M3FJ0e3nrSSqcALrq6izhuJf8TOsaR+bufodtw1rbfr6xTzEWFDDCUVgyWJPFDq3YSLdFI2YECwXqA7GuTpQ/fgGPSeh39NVuQ/kh3WTW+uLloAL2T9lMw3YLn3N9tg0Jji0Fhmoh7MDk6/clM4TRD6m7LFmlZhSs7vZGY/Cwmkoq6utNSAqJ4SOC2s9g1sBDqDeAuzhnBiXCfELKCIwP0jwZFdEN+RtwDz6QWaGOeIldxnKJztiqsX6tdlse7EM+kgxCVxbjra8/iesSp0DlqFSEck1vf4D2vaHFDCLWIYnYBtHz+ZBw+eYy0Z20+cHUyuqQps9a5g3rBQ8EC2AwIopU9Cy3pUzLCB+gPLJIhbg6EF06xMeSv/nunRUuwXbjU9SsFEO6798DoN9cjucXDZQVbFxyw6gCl3LLWBGZTkovUC2wQcw1EpmxjK3nknqekNIt6nLkB3E/Q1eeAPuwvZ5rIcQVWez2vxAzb+0dHNzOXx2cxI+rQO9Gn3XJ6aHrVB5XLew+9SgV7v4rXuCwg2azd2NrNi84aKJSvpXDMJbis2eW26u8MTmArjccNniv56nJ67gyY/bbdIoDMacJXBNAH60ZWwORVQ5RULzKnB8R4gwis5kBXQ0/0VwWWVAroRvtKqp02GwU77vin/QepNYv9KK4FyxQmy15nvQPLAPlZE5Ib8UHw/l1XoUBfd7oEDW4+lZZaokOC0BRpU1/tesLKdfLlHZ9nF+SjtI/fz+TMHYmT57WMWVQ85AH++6oa21LKa7hhnXVgDcyMkprCm+qA/bl2aPnzvyb4m2Je6f1Tpgx8bPsKzZqcXXQI8OZwJCxXqWGlrmy7rXFXbGEgZBSd3uvdm1yBetwCEj3358Y7UgHTdWSDqcn4pZ3ZIKzdMgQAtszAekpB7SuBLjOWxHiAwSv+OQREqubk0A5pFDaFGRc1qP41/ulFiMVaTMiBlsRUYMavoIjOD6HjIbRcGjN+G3jrXM2iA+iQ/d7x02+xaMce0ZNbe8xjqvTn6uuLWMQL8AGp0/jKaq458P6l02L9L21ubLDGWfnd8ydrDrlm7ZKJI8ouw9rO94u0L7ucmirio02C2nbtysPw8jbCRjypX4/uC9AmoJ069Eh33FD8mE9Nx8f2qXcIxlMMuTLb7n5FWzET3F1JlN9AwyaM/j9Zhj5BSH1BE1979R/ZJ3KMiH11c+KKS69RmuVl3AVqTTjQ99CwGlLwaAEOL8e3s4JPycJdK0GhLGaV9/hK7t/TMVmnr4NaaUHFcxf/ConIrVoDEftSqBT4r/vEnEZ3kr/nYwllvuAcZsW8eInjCDNI6ZFf0YUfjf61c/mvMcYqlcvUPQ8/LUfuEMmgSWBc3zPShUe7g4NdBajie2HRv6B74h5ZCvbCXXY0VSI7d1Xgp+mv3EEZlJhoRnPAKiHmdLa3aNdLBhNM+4DP/zR7JxvxC5S/qvf3Gl8wq6ZQ9bSVbPhrpxvnxIFVFkbnZTLjVhB6olpBOmppBE9zjpI1ohML0n9VQQyr9K+Nz1eVQSaF7GmWWHbr2yZhqoVf7wTYVFSL2DMafYvHv/VAgqOiulLmUdlIV4GJv1X+hiiuIbPVi1pKoc5Zu+uMqpYRuyZGbEmbpcixQb26VjzAG5zvtX+K/KML9ODtc/Wi72lQ/cF49fscRI5XsKM1HsWPaSQvS/1NT3FSjZ7VqLhadzR1X1XM7Ll7LwAnq6q0bqJYAz3pEHRCozPWwlPkmTR2KCgWzQgx56RJZioMmLuWqLVctHT2mL4H0U2+sdR643c8fIvu5NyF8v3JX98aSOdvj1S/cXSqaAl4SipK6v5tyEcDXSueU36tthygwCQwH6P9mudfxUIs+4cLdS2OFT+4oF79XmrXA/3kid6A1eFrA2B4C6smtPTwl5m6DdWRNXsTYoCjKep4EIIDKBqprRRhsP9PT15XAYsnDjverzwipkbWZsim/rrhidOcaihj9mMjXNd+2/KytJTtUEkIrc5wDUfShGlZXKKWHZO7KxdLlxZpuFm5+Vg7aM9ml/AI0zqltLdJDhymefmNDa3+rh48veMSjz5zuaVcAffbXdswzP9lbdvxl35WrCIYR83VqTkRdASja16ucseC23r6obE3vnj9mF61IxdQr0ya+RUnIF26xER4moHmPOMFWTKHFVHv5zU447ceKTVFnGHYMpl8hN9Ngn6ZoR1OEXzGPILHw2nFhpu9WcL3FbKDN54guZyOOMqjRVdBsXT46V+Fplo+kEQZRexq7ifNusK99dglkI+oZGT4WndlKtJZQwePQt9i7VSSNCNpFJ0saGwlc1T5ysIPuUxgISOkFG6fqwzslSu7F4DfjEeB+QBa+5eMAvCKUXVDY54jwLPjWrMSkn0R5k6s5y4RXnVX5OzSvs9qohF2Hi7XJ9oklH8gUvkaofFCgJuLGLxJyJBt6L5KdQkikqbgl4fiIrTFhFuBP22JflrQSpIB9xStdna4+fMRIHA5lt2+pZoiyLMBUchgcFAzTsl474yUiN75MrLc97YTIxJA6VkW5HGPJSq2moi59uqmTs2k69ICDJRv61q00Auqij9O6vxbvLUOn+PtjphVJdy/KIlsfWl0nPguPva4D7ni1P1IXJWLGLh/Tjt01jJEsyuEKGPMxtUPfAU/cmUZOwmpV7E63dMVYvJcuAr8L98SmX7161cFgz45PCd/b0NqAOTu3Frfy7uCq1CiBAqadoA1I2SttTSzrj8917SbocwCsZgTU6Z5G4vOT7b4kWcQZ5qXAIic/gSP+oK/4Xa1Vo1huF0rvoaGi+LRTYfLfLN2K7wElPS0P0SFoL20Q8JfWUdMVvqtsgy0meX9bLIMHXScLAwlQz+s05cnQ4nDk+3SWbng0q8HyhNoG4atLANfnHNbaDN3FmLvwMdvDc6dI6wh2ojhglV0xEWg7cR4JqdW34UvjmdELmPH9AM6qFPKs5ooFLkiDjqfmPSx5UCaIsxWKe6K9+TJhSoRYWIADucf/JN8ViAAc7kx6GFsNvq6GepPo7UYjPGhYiTcHQCgfK0KVTRvTcmjFApRGk+qZDwUtWnUZeO67j0ox71H8dEw9AQ16uI0wHQ/pUqlSiCV2QnTr7wEsJtsdhYtVRHQWNn1dnP/GD9Cm1IvOBU3koMW65BsJTxsp8dSdWiVqjgMdRdBdFQZM+2JJaclI7NOAU6heICAmG68v7sJh970OnVYk37gwLuGwsTGTyGMNBFdeneyYpACQGfIv7jQFAAnFNpofXIXPmj1jZ8+yVmBpn1Wx5GLWXcrXsz1RM0CY/IHk32GtXSPqBdiY7M1TmmUNylQW8cDtgw1FM1jhrB4OFDKGWw=
`pragma protect end_data_block
`pragma protect digest_block
31d29968d7d92d7fdd4740e64bb12cebc5c9e5ceb1c999b3a97734aac1cae55b
`pragma protect end_digest_block
`pragma protect end_protected
