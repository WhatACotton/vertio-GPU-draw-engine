`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
Y7IjyYssstxbYRf57/BkiUBFCoyz6VsFUhwFbRaqrDIVOPbvnZ04fZ/44T0fsuaKYQ0S2g+ozcb5q/z4ajmwqjtCC0DUwU/H1DxL8a6n9AewXxG3bVGdwcWapZHG0Rp0zHLReZ/f+1eJFpLq/o0UZAm94YWLUUjspEwLyj8ueS3ZW7xDJLVslSZyLaXyJgHyfgXlfy3OD8c1IHrz69d9MVjlgy13xeWJ890na90pMTlFkmMy2a7uNMjXiY0uPJEselpwuLGPRnruVkBczl3BAkKcIc4baNKj+2a+s+ul4ifpHMEpjIMzxu8nfnJE4+5URdqF6ZNdsXadp0LfHRK4xylawSKDUk6+Cj7X5bZpovdP7S+CVk72SpmHhAHmzF9KwlT8DF0eJ+BHf1nklCwdpuDJSzWMnZwrjTVVausuBGvPi4NLzhYAzNSqnprfbMLTwcW2QPqlmv5LZHa4EDDp6grpFo1PK/6Yn4EX5+L00LNwFHTQ+Vyz9F4udM/J3daiMaoItKQO9N/QMEcVOCZ+FrTRUQ+J148q8nxk1WVIRu/2ekHcNeFGKX9PT3lLawMvBuCuJEs3KBWjf0RCpFVOcmVrKXyRJPt0nwCISKjyyUZgFuY33KX+r/XfGsL5KGstzB5vC/v53oivz5GK0AkeK5JcwOrzXZM+pqJ9Y00r1m/+NmhZ0uM9zOylrcs7ALcdRbb1q4PKPJrYNSLmVXCIw7uBv0Vmw21TXqRweNSwTU6rLsvvuoi/ksD1B/MPniS6SmpWnwufcqjQPRUo3aAtf6Krf2b4dK381Xyq7ruth5Tdv+XkIBhTTPMaofJoKEQuNKz04Al5uyAnfAok8y5T+R3E0Rr18eCHuABdDtNF06IeLPecz718J+ZsDuQr0UmshSgfX4ND0iBF5wtdqToTiaUZd3Trl0dfIlfB8Dv6a/snwckwbhLXz2ymWuKoGgXFdbhmwHnkO7faGKBiCDYGGXNuJpFpjNJ+eDWrtJ+1J1mbhU0RGbzK1MCM51o39W6GYUuqz+BlWz3im179euNHugcoLWOJWmF7vMQtzfk4qYnEqeG4tcV3o2l0msAL5z1HFxpBnGDcKQE2VkFCns2yYHe+D0VJo7IHyuSVKQ7S/j03/tzNWhcpj09tf7R1vYKbiCzCVCZ2KaVmQ4C0O4WTmSIAyVRhAyyONkTCBrIuWc8LBCXdfyp7VcjjMQiV6dkwXZSn4Rt6tAIVZmSg2d0Q2V3uBW0w+PADUo/aGTPM+SXgfpG92zShKdoPoKD5XzGbgq67uwhiA9QqfpIAmiEBSM6nuO7FmwppwTwacQDnOPAyJxExvNLwdsK6gaC73igU1ctBPLAh8VYyQTDgCS56QnDtrYRH2t0mS5KVXD50w/rX0K8G5oRU1Fw1nF9d10WQifhADRsKFXZEtyzt5kSyc4RnE5eEJsIFRFCYIERu7Nr9YxXw1YAKgfEk7W2NRxVnteQG1Rrf+znlf1HpJoBrOaC4NLODbhuOLCXak9m21GmUwNqhxheRnxPK4j8zpn3IrQeScXSDdkdA3iO1xpsf6NHZQogv+7qe3j6qUqQ8wQlq4CGijxzIaWTBvgWW6IVJ66C5vKE22aHEj045ZbBamwa2kcL99R/u3KeJ6SsraM9OYIMwE0dKggc75O8siKHupKabqMbxyyWvCHwu/Kqqx7fZQK7XgcdMAFArErP2+IXDO6d2yfJuGhicv3wLIAR2tfzjRXZqtM5EpVJ38dHc1+RtdpQhhJKzeWCNx8HHa/5cEIV0qQpyKFsePwMtJnHtU5o3SdFIPUSpKxAyEpWsQuyJ9g7QBl/7YRPc++as6zdExl7XmUJfxxD9yeXUGXZJnTavD21zjTRPVaCIILKwG4aJebrqE3H6hNqiky2PTQQaqKPpvuCrTO8+HMtYwCGLpkw6r6zEHGijSWxdCdiQlUjN4wrbIiFf75eUZ70ru5DHEwxhJpNMYka/z1cPuXJTxGVRsscAGJSbsbo55xwsEexdXrU33qOP4cVDYVY6B/ON+4hMdqmAVmO82hfE2MxFBS+sSIPa+zVhhYPBgljv7//SMvGy5DcPVw/MY4AyJ6WqwxOOlO5X5FkyDV5nwVceYOI1XXgKlL3HE11+8AGdIO8ToO3oDLM0DrlMp/t6zKEjJHbnSSdHgwDSLEOeoIC0Voz/+0PsAeBBdh59S4zG1nFq+AM9sPZaUI2jhiqp+5oSxwqqSD7Xm4AjNE1hWsVvrZ1a8Hy8Uj/mmzr19muXA6tPpzAa2gj7DplJfzROrcyPlkWbHbTOFlw2Q5jbMQF/7vF4RxxR2axmhhRNhOb8flY3Aj+7jO0Q9kO5cW601WF4f0qfoBbfyw5BRhSxOhD9Wm+qekExYJtSRuYX7Kx2RMjhB/Lph5vBkdkDAy3XUL9w59frAEB9Bb8ge7kQTDX33MU/a8rFXXmdkpoqQU4a2KKnejOPWyV1SQzA5NqvZZICBQEYhLGYyDAXci03JPXpvldypdQw6AI06EQua4c7g8zf3jai2rxqjGHmKjDcK0QJ5QQIbXGr83XtX17emNZnWuKnimznIEaRA7OE8Y9tq31M6ub8Fpj+uNdZeH6DD5zYQhPMajLy8LiMrOBc3qTeoqNLJadrlP+5GptrH1/eVCyratJQIXKrI50F1Adew+Z8O3xUNyEpmjl5lFB7gkOjUpCl2LNEk1F8GQjut0QEtXZklAxxdEgy5uET7X/Z1FyU/ThoZx0PcbrQNhXVaAFWPglwEjQ+RmHjaU3e3H7lxRYYInDhJjFXI8z4Ak5BQgm4y693IeokvO2H5gOCnMhDBPVPmaJspUxvhcWVlaIg/LiElh8JNsSjU1+UtDB1I26DLlmmTRdg8RX2K2pE2Egk9uCNvKtp9WjOL7Nj4t0a1M+duF3xyJrKiotTKeUzMskrT9jR1Q7O4dv8GzVLHglNIU8JVXJecKQqVgRdwniEP1ZP9tMgKpOuYy62us8B6/wO8W6eAo5Vx2MUQ6R3MSo10TT6gcPVfw631Vkh9Qt8r7wzQpY30J+dw5rdqSV4Xp6QgQk7teSN5fB9K8hRv9dhQ6ZfHb1WVk6OsGyzFz/wR2vMFSy+uibnzOwXvO5CtEL12jJ3NzapYkHYZe/j/QwXXcEHywgRbMX8ge9HRo4rfWc8wpuLr1IZUsgNO7+A1IdHGatsLUYQ2oQkRNTrcveeI3LdruKGpcpBb45oqBB9OGDdATb/2GzJZRn1uz/2fVcgCikQw9snz81mi2VcUjk0GLNdmjtgBE4OQFORMIVsr7psxOg5AVcNfw/pMQ5QU8RaOQaHzcYN5vMDhfBuqRpndTlniHcQdpfKTXKHXSlMfH55RG7VAj88SWFT+em/H/M6Momp07kdTsoxyl69FgmHY/w3seR+AYx8nUM3NLosq7T8mALUaCa4Oaa1GqPc692YPD0mWAzvqE3Z5vMK8usVCClFjHIX8r584Byg7Hqp7uFKTOCPGwW3OAOL4tDNM3Ba1d28hxdpY/tQo9yegXhKXyr9VgU/nFHOEj03VMo9GNOcOkklh/gVWlAYvVEhmTCkI0ISkHJ9ae6nxm9C10/7bppIVUEy/fEGziEtr4VEsWTF4C/7/xO5zCzHEFlJGv2V6F8SDa6cBpM/pWFGy+rjwGX6i3mHwKq3XJEoMziYMbAEfHJsqpjMC46R3X4slO+pK+3NL3ZqRtBcjV0oqnb3mFWKpeKY3NNNNqBvSpUa8hMWoJl7WVzAT4LmFcPGhK/xXkoRQPpCwghWZ/HndhGEXmeVPBHUtHenpJfyYVXH5f9M6MzydMaXabqQcymt9DnCxWpD28wmmfMn4lAp+dT6r4WZFeMO7oNmr8tvufkYmwv1gB8FxSPmcIIcBKzSpQkWf7khaqg3PUBl37s79SFlSlkE1GKU8Gj/ppHjg7hArW2t9ixoMWvYnnO6LTv1b8VfA6N9WQLqoKiilsLkNhhxCx0g+TrjEF6EMs07H53IOmAoPLnec333Dg58+es3ppdsRplR4NRnXKPKyj8gkF/mE5f7ARIBAnbz0mrcBC4vx52UzBYkpUpnxSvw7eE2N+K351RMluhE/IiBR/0Yi9M5Ar7SV484IQPF1x3Fh3qXOBBCDC2fkz0xuqcCpn9Pmat099lbvi9XIwjPkogTF5vXekWpZMjLMFabewdu2zqH1YeVu4e3ogOMiYnz4x9PwQD5WBDEgwwnYlBT9DCCwU0KEaeZHK+fB33r1pEZsu7bdKE7789Zijst/Q8inlDDjpJmKgnV9z2/Zbpwjn8LxLaGBv/V6TDGfNArNZ77ON7VCIkoHvi6txPjtVoQyp7pPRDRpP4n3owbzFb3x745VGA/pNg1NzkYp594mC7e/YjBqf+VtNTFmWWnyaIlsZQ47AcHR58xA396eKl7LIdwVK+hXoIGiSvOmI8Cg9vdBGkNv/bIQxWD6uSvSidqjyLHPzajUbkTBFUQVZebrWe29EOpuwKPkBCo/gTMjWJz+Uqb3+nDsli225g2bBVAaIFBjvL7YILr6x3lr6OEg36DCF+FzV7zKKcm6iZDTSv45GCU2Ynz7xh9fkzyu/9bz/A+7wPqy2kYhI1DgyBwwPsxdJtTjracAvG5KFI/QcZS02M4cstPM6WPoe3oJWKsBR72rREELPmrTE9NAEbLACdpVNVUVkEYKz1SKqvV4MMVfyyCWxOu8tY9WB44lrZsjVRFvyy+3G+PWgvLrEDqQ9mK6i9hM1RdqoNcdv7GWg4dcrZwGaKuA9gzlOl31ODiW6IVi9R6d1UNnaMiFfh49x5am6EF2S1uPTfRX9qU8CAUJ6+ch13jcrWM2ZMvnTFQrSgGEsHIOXpRbyIoId0MgvhcdjJSJQie3anyeiQS9Ig+sjX+hDKBiiN+53o4r0TeC7XNmxYqkwGAGT/24b330DKQDZkwIpT8pyofKfh0uctLhrxRodaCg1hmBft44nBb2Wpr/gwFhH9F90PczSpwi0+dtpfMq0jfU4NNDWmzD7bcd+UL+q2RYOGQSSQTzmTaDeAXTBfWzZmQOfcEuzfKfH5dv0zMND9oAygnjqRGDVbv4zubi714K0QpysvCFF8OyqmMEalpGGYs5wUSqf1ePTRgaFEheobYf83yvDMm/N1yq0AEeKLJNkb3cMIdHwcMt1DQQLyI4S6lAJHO9qYoU5c/TqswrKmnWAdHg69R0hai6qg++hSj/7O80MA3yCHY2bKFIwOFiARl48Tx7WFvJY23up/WjAmwKNa1oMPnUK1FpLqGd0+qi+T8RKfKPVTwrApsH/bhg9jK73ISD+yoCIXXWBPl/rwRsQy1u1S3XDFMNWsqUVafvYuzcwGeqBO11HgK3iGQWwUsZBBY9WdjncKNV9Uax9k2jGHRAuTAO3jOEqwLmj6UJeQWnSdVJUx7VN25Eg7HOMKWSu3IXY1426wPYPzGZX1AEo5Owu4oLhrJvGilabGNa36F63mlndqdlNiisRLwGMq7QRnjnXvBTTfUoMixB/BqERFg9DZPW3Mml8X1nSPVQE6V1xlqwlISa0DC+kXvz6sEP/u+Ue5lwl3iUHa/G1SZTHFD1ig0esBQhCKHrjS2GgyYUvcDsBw47OMGV830x8TgQGJpU9s7xxUVS6UosTe+PKiP4V7dqvcwKjYhqVc9g7TCbC7DWVYr+azFk41ANdWwcOP5o304hd+0gI4JnbWpDG4+qjC5wKtKjw7HMk6I+6brs8jnBx+Dj2EaHn/kojpyIMNeZVfsoU2EmqmGvwIkAnq7hdWO22nazolOgSR7+scojyD0ohRkVqzuC8nYM1/gpZachekSraYROxuvfJYFV/2I1SzuPSyvPIJCpzYPDAgj/7zSmSt8qGo2yMB507FvBgXOWuezQSZODK2qlYczqDzXlAKJLLxn2mTH7no4MVNp24uHOV3WbVezWyc+LClJueibcjYpwUEf3M8ZEOYs7V2hH9g4P2Io1bXZi86jFX7Bup19WqMcKibgmaoe1yKFKszQIvrZ9AmPgfY21JCHI8pwisp29NpTrD60L4+alv/wmDoA1iTmjxJt+ruemkVkmX3k8qvf6dlrlV56RgvjXyhm6y48AI0PYoBHVF2BRq9KyQArBBlob/hf8ACIevU+tofDgUfiO4sJ/2NCBz5thG3q7Bvu82qcxkRBkrbU/9fwCLm4WEKF4iS9Z7mBbQbWAw0ro/orNeNAe5FnEI9Kx3kOTZ7uytXmqpcsULTJgGtrQlPKiq4rp3ToF3xa+edgY3hN2MB5oX3OqQ6TBZrVqrEzodGmcNdK7u9oJY6aC2rIDj1fUWoWktvG7U7itl8T1qkbK9mnrcnGhEboYSedTK9+zNji0PKHuhe0jnjSyuAbdKFMxAvnHtq/NzM1Be1q+MKVAI6WBIochCst0hfj0SCMfPygmf0KZ/BqIYfXKNQAXBUa3Hq7l2b4hZSXdy7lqsGjqmcZBhYVEhX/fSJzc6PM3ykNSvW15qTZ+KZzPwsQwBpOa2MlQPt3KOKMvxBVYWM4Z/CJyGklLIAZj1FsnDcWmGvIArXKk//1OJJehuXd7nxqU5aKg+jL2R+tLjW6ZrkyHKFHX5If2JlybS7WG3fuHxasyv2DXdhCoDgvAcJ5AK5n/k8dBcsxPayiS262fo0hAMzqM1z5gmYpb+XE6EtazgCKSnZNtSsW1k4DWZiwLbBB9TbcJyVc6U+a0cPXeGq/h53PJepa266VKyiJQ7OZLHg/RK0iFEjtqalz2bOwsK+OihajE+H+AIKe7pVkr/jke3oKvIHLT35mZ5HLmxmy4UDD6d322enhSjyIZ2aPiz0dxYCIL9yOueO6P0U0kkdFKyonRBkpilwDSqTwbGUyrHd19wlYV+NgmzPAeaAh87/3Av4BEyZX5GGNLalE9yYfmPlXDyXeOWDyhJ11JvL92azHT3ZMLM+5Y9EVWdP/qWaqogIyKMC8nD0B1PxzilGaHqtqDYTaJ/YaaMdIW2DnVTcVGR6c3W0xmTXpbd4zuHfs3/0rKM9KXpNGGGjJdZHXX2vXhUJt/DqdAmd2COCPFKtnJ/uIVcZ+hW7GSMUEA/Zw5fT5AfmwBgl4wIofNwk0+qPuKiLxco0ODmo6TUsMF3rVA/GrG3pQcxMEapRb8Gr6R7sqgNlROaPO19HDVHIWWwBjthXTc9z/iqWKc3Wq67TFKig/x5l1yaAIuKqpHhyqx59YTdIpcH8GwMhbiucNyGaMeNNR4CYd7e1okTl7ECMzffoXyUOdGggwpY6lHpmuU9qJ07iIzVrNzTfmSoFllDAbUzvPW5uv/rxJFnp8s2AqZCJwhQLHWrSQMG3Ct2NyOSraJ1dJUU1/WMYDmuFw4PEnq74YV452/xoUU3CNOU/t5IsC8WZH7rwszY6DXPOGar6jFUU/kdJeEhFCk2mwO5xBxE4ITOL2/4QUPx+qPOAmryCQKeF/Q9HZQ3OMDzmq6g67+8/0aG5756xX3JW4IQbURL0UZTf7b5m3WAEjxloiQLEPkHSzaPbmMtkoRaNr78/fSmaJ8Bl2VsiuPfwVjM4pXnnJVlR+jmEmet6N5FwpzA+M2NZhnErkhoL/306nuDzU6B96uU2exO8s3mL80IntrbtOBwR4yLUzrdMipLJRHPum82cHphlALw8zVc8y2HrwKhiAHKT7ALZqxYqtSmyQ9559N8GY0YeRXnOKxO09GOkmIgqKAu/wrdeHX5VU4ma8Q7C38jcSk1uIEU0K4NDQTt9uvS5ShkCxCn6zQj8Vvo171KPXZ2sInge7bRJhEuffltIBaBpYC+vrKGlq35ZabYWSWMs4Rqu6JUnpcjlKGPHHS0aS3UMgMORkySTft53ce9upsstBc6PzuzJ0/eb/flFfxkbYbOTY928bBMA6djEg9yo379eavnVvJt1LhtwqvocaUClNRXz8gE1sy6MfC2HQdj2M6FysMDZWEWCiiJjQNzwdV0COQNYZ1sxNX0qZH4rRxw1bWL0zQY6pkFjkOeWShq69HXNQkOMiww71958psgedL6qTZA0imwP+G0O/CejB8uv5C4ORrTiFkDA45M1bXHjOn/0B2NFAY3hLmJC/X7RjyP71Brx9+ckb/GTHQAYPHolZ1LNQzH7mQ5yb8FXpKBEau2lbNXnRNq8gpfXrk0Bag09m8ncuZOLcW9MIVN4Kv60SJy8WS3nlt17WgYztFilQAWLk0XnZLXUPGC3t8xgWWyQLCn0bN3KPxZ+Y8ryFksMwbRV6enA3bzIf2sKR/dV9QtLBpM0RMJk+XvXa/7o09FpnA1clwPVL9tEdUEArvhbQ82N5WeyzFLhQojjJETVhEjKqaruugPBq4N04aC6B8yfd2cI5YSmbT6nflWjP4cEmTtd0X2OE2YhbZef8CGZmaGAvZX4lXRBEc43JyAL475jXNwBf6uB3ANysXCXi3hzvAqNr2Hj0GQ22DCjexHsHp2dFMJZ8+ozrTEI5T7wP+m2yAxactLe9uJs3f2HSfLHjH3thG1V9ksiFqyuNmQzcIbUMmNpAn1llCH02CzCVl45+uAnhK1PIBiKJrpXt/xFzcNh3JevL4c/QVp+Z2kgYqEAwhhI+4iXGYjmnuNroltnUn00AnZHXQ8azvhU8heOnmb+32bEmOEQWxcW/ZTDxEhmmV8XvLQiqSw/ab0chLGMOpzHH+kxjU3iLiJZRRdG5sS9Pas6ekPe/H33jYY7TC19qVY4wRi/lnl+rYhHdDory2hHJfRyrDiE4189Dfq/SQiqJqLHbzhjXxzx9hgz0b5zwmo37ElfQbeYoSjrOsUI3FjWcNrVKyEOZbZtNWEecZ7NSDGeNp82Hk9iJa8MWMgsQBG1v3iQ5DAO/DVTVTYJT9Dmn0sz/ZBGu4rtJG7v6uD3Z66ZWDdf3MjFJ+aa7lHtBMpoxyOX2Y1hPgho+AnfZh+etUm3mf5gapLaxyv+vPIcJ9znEtWFE5fLkeTgUPajEj2G/qAlcu+Mebzz6vRO64mvT5UklzWeKKhe+BxskMmm0k12p0sozSwLdWqxTk6kSjnOPznn+MrcfG90SWWgFhyL1kVt2jUm1S9slRAIP1K5pKSpN8BdDPjHZNmaBkdEkofW/wWzXp6VtZpcB5CQeVWnUPcOc9iUztm+EUU130L+BFrx2z5gdB5X09IfR3foj7uwOAzi7U2KVxQvJzHMl4Fx+uUbn4v2PiNiXnFLdLZhGioHIDME8bhzdm72wOaT2mbOUnYPZpB2KQL7WxX0MtIQv53Vw3Z2M+HN3p0aI+O6e8ocEZAO3E16Q60cbCKQ114Vch+z+I6zTefgwuhsrtDcYot7CpBBFN95yOcoYQCnCAVJR9ouOGzEPeCkd94+ps1rdrcBfs/yZBh0gWQjBz38xmUofHX/Qja76wc6kUzRcjGgT4+rhwYJhUhP3w04a1D3o4JKj4fzwBeRvNlun91DFsVHOXeHiMA4CTxhtlXk+g91eBG50K5Wzfq+c/Z0Hx3vMPGBjpF5b5fRcdmGJzV1yASVmqulI0W1V6VJY5dZdrYuewPG1Uh1xlcGPcJqQKtNnheP2ySQy93M0mO/EJ302rxbN/aLhdhGMGwZLdUz/Qz3cVzA9W/gimDTnF1jB+SJ6LfFo/X4g0o8d3Z5TroGeEYH9F9SjuntuaxcubI/e9Lbp426gLwAGB6ziXbL0Me6vPP44PUO1gdIC7ln1DDPmNuuQyWfhDNP/minmdvpI7v1QvcK295yid637H8Axa6A4QJH7R02olYzVQ5V+V8Zn6l/s6h6SNbwn0WbrixAGv1ps/2n2g/IjU8BADtZKDuF3YUZIhrZjEnGmWDIEbyoeWbzigFN9kzFCa9pdMi4hE2Val4/nESehuE7V63jV/t7de8zd8pWIouu0Bk/2dKmaU7ZnxQCdn+7Bbi4/7S8swj1OS9TnoKjdGvfKzNqadjZt5IQoA66bipUMZNOgLi3Mx1dcWfydKtP3mPi+/DkSNeWbZw1YAqaieIRBnGCihwnLhQQVpLfdu0v6doRx+gMDwIWfeXtjRfJ/ADRXOjG5KZPKxj6UQ2hhgIGvM+fkYRe6uflMwRS6Ey7b3lm5lRPqunYeW3MQdzJnOq9SCJtSwpCr411R05BXm7Igp4uM/DbhK9lp0AsmocwZibl61D6RMlJGuPBlv02m4FuXdX+5MGmg6xEzTVWjYCNDgaxGpqQNRTWb4KR5JB4L6qkFK9QWs9+m+clfelNt+RAA7Otal80oU7BWiG4MVn8dor/VoV2hrISW+Hy5buOYtzzNdrzwVVjIXyQh2xQ22+uexsIe0voILLO6D4BFgXuhNAftIbfeChZo+gKQba3x1S4eyVSPZFkrRrGttrFpT9Dbbkp5NGiytgBYNdiPEbr4j+aYqi15jkBYvGfsGLqwHqR0EUz8G3NJVF5FSYISzsOV54+IQCCU66simq2EYIBrUKlpYfipp2xbykhpZfq55/Sb3Tm0hNTpLKN8MfcqAX4XJbrNCRaeH+kMS0894BjKrsr/e4AmrkN6MinDP4Oj1aUs5Ro0Mc/GyMZUV7LTtjxpjL/S6KqQXlaguMGsVg2Ik1kZW1o0o8vGWTwu+pbIEg4QHIWFmXSWFe29ZAMJ6r+D6NmfXQ06oWiVcPYBtvTOwswvquc4o0Y1wHcYff5yTHZNCJp48aF4KMKILgwXJRb18OOgggDOy0L3/R6vfU1rHBbhD8pq9hCxZpAxYY1pHSA42T+0vEmaFCbcn2wyG+BZKx9dwEgd2bD1lQyGLYOmZuUaRdOfr1uXJfTkpPCw1LwwwnEWmyTeicX8uOECw4392VCzvE0BOVR5LlVRG/xetujP9XpNgdzZm7kawmseNre4NuWi3gWkSLPKBg9g/QA4J0vRr8rk5o4rDi+et3bvrvfJGim9id5/3XwNIHfxbh7dbm2M3N/U6+WvR/CSaAOTvGTBsavp7g2t6/c8UyXIfsw0R+tcYkrosTozVFEOHGBk7BEJSQTnrgwI8nBSPRGGTMID/uzfTb68WJnuz9EGYmRdNooR2DUxN66ebMyWk233DkLgTy+vS4C3fniqela81yvP6ITXsXz1o7bH3YO+0rdQFs+zEj3JVUbDMRnqmq2EFBuztv2MPleHEpLg4qoMtdcsa8rVsvrnHQvQ3QcOj0/iK9KL8FUqmQqXlGeR0cQgFg4lpg22qWLJZNob00y4hZc917/PtwLt3lADXAiARmM+dukiucv3z5IG+Jmm37HIj4scWDz8vfEkxxe+sYVQPhvPIxdapnjFEaBIPbCszeoyXbOCcWqVrqsiGY8IT/aJq8HAG+DZwDCBoIdAG9nGEnLQD61rBp2QFK0s1YNrdbboBAQPMl7TLRHwxUm3IhXjucl7kc0XsgqhoR+QveSbbTDj1Hwjd+0QmWBciqpki04SEUIR+PKfBgmqWnQSAu6xvLFEAkn2dgUbrf/q7Pb9CkOnTtGL8vHk1z/P21n2yzD+kJ/6vsfWT2+5xweeSXR+9iRwNR11gyHjGRSaHsJ79djeMSN+PFpCmidVGnYENX7PZcIROhoelclbzPKeTcE1ycDKTjiwLHuwdvw0HZ871NHWXAJu1lAm1JhVmLue8tW5RzYU/vGoNkbziFh9onb0u3b0IeEJEYvh/i6y5w6FBoTMp94yfajzfWt7NQXE2Bc1OwBywhCUueYuTBSDY3hqNbnKnKqWJINo0EcpiYdIJiVb49BSSxRinQ7GUYOJZ9TGC7qFn1wnXxvmEkEMHRFXfne8CJNeY/4ScM4ocbWKwlz5GIOouACoZ1uikGz8KE0SgMHzrOXpZb6viII+2jyoRvRyhisFRDB943wIQw99oXoNcKzgWgExqmGR5rUKIXX0PfehO6hzCfRz1VNbPw/zshHHVOC+TexWDq8+sK6S0W2hSh2B75mYTOSIiyuhg1QAVkyuY8LkG+UGU2EJ0TW3VEBTK7pkWsNFbDf+IgMyYhZIajThmsHQc934elTUmgxmlwJ1xIWb4jYqR97O7uCkx/EG1diztWWp+fwBQRhqpTyFdh/RbxO/mrAHOJYzNMnhAKPEB4OrowvjXsstgXPVoPWaDHzb2OaSXJ9pIjCYVl0LgtdWoJppTatl2Kvqor3IEPPfL9lrdUVc4gcUAYHNYvLe6PhvEqH/anxaj0Y99N1IFO7L2hk2ZA16XBA8zfr6w1aFVb3a/mVCfnSW3w0yjdfydkFuvX0Pbfr9L8t34CSWz9JacEUyhJmX+Q2eTTq4aRad0U5BBGKIpAICrEHrswUjRezddTtvGH3xqGZdO+vHt6CGAfUloBqwZGSOTI1OAvRwzlxNC9a+tGVCbe8Xj/8v6BPJOekuuMx+N7FUDf4qVRvnN/9lm094Tt4Dcz8qAdixmfxsPekNQTJrpt6ZpsF0q97W4t4UoZs9p/b8z0ESlVbdF4qiiIITzYpT1/05U67JN1BeYatPeoXUUZx1TuFn4m2WEBjxPwsovd7RwJBJK+4lVLMLUjQUcHPtcltLEcuUCxTBBSkbw7rLmpaGE8lGjTxKvt3MZYjp7ASAH9iWc9vqCVit8gekUTVlbsLbyuxM3WCXJRD3eYwlsrhso5+Sr1Vmdx1tbA85Xt715H9fVBaFxRHyUPPAjWGQjPAZpw+xiQ91OytmJxtc+hgpznXTXJdl+TiDuo7julh4WNR88FX3JP1yO9M0GQBHDBwwxiRVpiMLtbzFWiXaQgMq9UM421ZJbM1TF/s/S2muyi1fDNz8/UhRuYRhTG5NOzR243TCAa+15GfzEdHI+IEvF5Sngj04FjyS78cPsyzNOBzDFzNVKFKDP7I9a8TZGfGw3wXUXDJwU8jFNNx4A6WZ60AGw5X/Mus0oe6vJcWPa9RlYfEAQKh5lzWF1WvUSlsGeEE+ntBLOcQ3wNiKtEkT03OiNF2xqBrVjSQweoCGseDzGP/StSykZ42112iwxQlwy2l+QuOpABqXmJfCHL4lWAwcADA/Ho3lmm6G498p/AcCezZ/WHGDGwleSg9RB4ajgVoH8MTQWziue6BTh0tXDeLm6SKV4DGddPBzEhJbWyTXaXKzvOGhNJ1Gw3KkZb0fpVwHKObVtOBSK6qtfsrqARN2/mt6Un7LDpAeaF4UTQhIkD2doteZlW8zjxFHb1hkWzYnAZvHeJi7zbXv0MwXYS68SlHYexSBR2BLHv/qrZ3DNFrpK5k2k5S9J0reAUJNlYMqEetWbkzFTZVjgCh9Wj/nImm+KsYVUGjbFtmkJ07/8n2UZbbv5NQsHXvAW7OyQw1KptdJ2ct2AY+8x9Nt6dreU07cm61nCrGR7hZ4bQuToKoc46excyGuebfKtdZRh7H/FylNeEL3qr/eVeVlZrNFI6zqSklqMFXAGmFIfPMEyLlLAU9ZdxxoJv6pSZi9/iw0/7nO/pKX3M2+1U3M0bokLg6uzK3DFizJ4/Whdxxy16fV3OpATwTyZFh0wqnQUpESRMaYV24JkK9X7abSuJ3+mjM2gHNP5g/FzxdxA/q5hyIdwEm2wKTuTv2ZvL7DcJm0wJ/n8qW63EEacZwDCnno+uwLEjA8Nu/JD/bgD+sRQFvh/tt78hQU/7BzLhicALRlTl1l+8ovioBO+u8wHYMLDkhQTHmiLTRAXMEbCNdr7kMJT7iyK6Dz5bWiy805Vh7OBFDdXNHlJazEytEAaAiuUM4p/K8pacmmFE00GMvMeNr3Zrk/BpUrx6qCuYAx/je1I/ursDGFn7nvaKrqqolUW8UxXsEiYuw8nM0faI2XPhEXuHNU3I9hv05p4pY7zUIpZl8x8YWJpSrUkptFUQr1kKTI8/rmkT5Np4g3KTkTVDLgwQQS0V6rS0EW08QzVTYWZi+HscsG8VCEITroLK+I7EGDlO3QSyHn2k2MwS/wJGfY9Ub8AVV8u3TMe8LJQNDdID6hcXsYdT+loGgcFcn+mV+9z1dgdZOLil1emYDfMQ6YRuDcBCrTPqw4IwXvY76lJZhuxkAci6NyGanQK591IWrggFhEhVA+gr+Sd81KL9xFZ1qfWSMhp1jpKxr6xzUWEWHk3szEjUE/+BMEMA8/EpUYyFO+7tl6lCnb9XGN0Kr5TUIyPRPPW51oLQbed4Z+G/R7DxiDXS+baLXLo6HRoxRKIy1dzdfYgbo1EqB/Sv8GXPpwKEzqD4FxmBeNDCSb+z5ULL7pMAd4WOnmoBNliYiv9EA+W/OZXZHbq42EFoGXvhu+da4FuaqWmAp/2HNdssGToWYrO/vL2hGYd1+GeSBurUi6osabmqbmSNdNRTqDODAzzntLC8BE0MX8mHObKhmXvDn5W+njprd8grdLKCRH133igY4BbepmH9P/020Mo47Tq9NTxUJ24LjuyC3vxw9d2qLNZblyQ43i65/rqUT3qMmsHMlLxbVdufJm3AO7JbD2hXBKlnrpGfzFE5nBmvWTO9fzxfLR7aSPFK1qI5PTtZkLyHlf/By4izPspT9drszU3rxZpjOLVN0IANdeFpJW8+PE2EtyAvokyFf3WmgMWqo9d1WW4b54/EUUls7/7NmspbfLIGOH9uJF6i7CsWyI6eVj6yIMsZ6EqyCsk48wJ4kJUoQqQQZgYT4G8tLRZdQGkZ154v5jk43k3wDSD/ueCJv+VlnQesUYxPnOC2Z1ZMvOYYIfS12cUFgB8Ds/87x/rxrks/KWinIMHiftCgCiCwcLqjMONZj1lOL2uUb50eVNf//ypTWAf2v0lpdKAqBB4ftuGt1+58K6s5YUQem1NKbhBfG6CH59RqH05b0B0o4Syr7LiPmBRnEx0G73IOLzXsIuVW7AspotZOFRiIOvyE6iGChU+isVuJiiA6fa4H8i3epXlEs3NVK9JjittpbjYPvATLDZViHpb/zYs0J5sZYEwv27P7kE8KJ3mViv107no/pvkd8dHwmgKyLia2z0E/seSXvt0Dku0rUzSlqf8+u+lyQElObEzzHQ8dpntl9SFYP8H6x0hWLinNiO23yoT53GWT3jEkfNg3BoQNyI0AFlpA62mxzNPgC9G3iOj+DfJiwLvz3Be4BuowD8qGMD7oc2OysOI8DzHeULYoXCkduGYVCFtTPokW77l4w1lVEMSvPPzDDkdiOCGJR20XOhwcQnfeqqeAXROUz+s33KSzv5NzirpN2q0iJLwjmkI2AmC9zy6/GiF773vZTGI1KsT2p9Jkya6XFU0wzsbLzK0xb/BVghmGA6Z0vbi/yqEPtV7/XuEC09GnH2wyZb3bE+KeswhdT7kO8LgZV+n7d7+12lhLS2AJibWsh8R/0N6zU0LLl3qkwpWV6ECtc3l/FTFuy7jMuK
`pragma protect end_data_block
`pragma protect digest_block
2bc33b2d8841e56092a10695c3d9f63e23c5bbd8eeaf2363aa7db80b2ac66cae
`pragma protect end_digest_block
`pragma protect end_protected
