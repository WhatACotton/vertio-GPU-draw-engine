`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
cWsuMS0Dnsmxm8zoUkH+HTptA8zVb5SJX3e7zKXAfN5Kb12ms/qglOXg3X6E9cztlUPiQywDnsx/QYBL+BOL7YVOGEA4IZjaW3/NYs0qRHrpajPqLwzbzgwMMU5iWtqd3ORF0cwrSNucGsHCyKa7pi9557etlj9ZCvn07Vdfer4g/f3f57N8AIjnnT6WYCAgtCTqTitDLdE3CaEWfEMP8UqNv6dbrmDOK4rCcSwIixrKoUwUrr2YeL7vQvv4N5Lp7LIIUMmBp/J5+3zyGGRUGHdFYXQeNxn0WgpWCmp69vcy1WNwNFQcp8LOLqs4rGZfip3SvmeqtOAxjY4HzG1p25uw+9OcDYOFxmRUQjgU51WtXXH+l8wBg5c5H28EpvijOF0eo3MvOwHJJuiDHLAFG60HFuUuNMQGZMk7aIUnV6V0KTaYrwQVRvj+JrbdsQu5a0tVFkabbU2Cwv7MHo+r1TCrYBphpclybuCc0BAD/2XRGD2ZbUZozaNezwgXmRA7H/WX/WzPpJ8weyzt4u9zzTH8bbJCO+eTE4XOcAwO0oIuuRO+iL+XZiBpo+9hiFzXBD165s7PXQW8qJvjxKtFgbnKfwcg5kkOrRMtJzf4AI+TYsFZmN1/NEeKuTPOgX7zeBmwySKXFaxOgh7Z7Wxd9x9YjhhAWjKfRlsCwH5PjIEmOJwRR+rpySwJ42t3kulj55NqFyYUEdJUu1ZEK7xe3tqJE4438+pjeAvtDIgBwq1ZxHRgZD6sy/LAQfQ0GP9YpXujXRi0+V0j7bM4mDg+m6q51I9PxJAQ27UmNb57QxkH1Tn+QwFYO/2BZL0c6s7TPGh+oJzrl0NFzvwPV6MCJHNvixxg826yu9YEGL3a/QHZsdm0fnRrmPJQ/CUHtBRYNIcmPzGz9/fCXLKZ06TT83LSmGbMtPmzs70SeJsnKp5yNzIxcLImR0We+GmlaKXVC613SGjka6SnT5HsQ57GFn7nKt/5hFh5kxqEBIi8lvOpBnmyT84tSXAKZLl45ZAe0+32GFsSXdchhJskhkp02JsdUwEiFwBF/aLsCn+EQiw/Tu/mFSrBC2l0sWNZ3rbIxaKC6R+1asV47RI+g0IdU9SUALHpqDs4Bl1Uffy8RrlVLmCizqX92XAcELJ5DEn0rJxAwariZrFvAcow6pW6pjufFYLYvMkqsI+QBQNswYsdApm6QxDIpUtG/7tolUZat44+HuQBNW5TstXpGoCClJyCt40Qhbl5KZMU+ycQ7K6GqSLg0MvM2ILDjgmzN/rn0UH19rIQ324+NxuLaPWFK+sTWycfdRjqmMZqQoYDOWARkI5X6Xgb1+TMGjmakEEDGB6oIgq4ExIODxuMDD1X2BhijosE51s5GBM/pcr0VwGBIRiV1MKlqU2Xmo2SytUqqs4t0bRazsa63vX9av7KL/Xuho2oCAmPOF3H96pJ9DrUnWIePjY7Eg9/wlYP2huaC2TjWXIKJgoe6Gjh/qLf0hvNqufBBNTOigvVB1k7MAyFw+hLq1V3KiqdXeIp7PqzZYKlKdKPkQ8BoNUn/nxwRnrk3beiVMPx9vTZtY2BlG7bFL0zdysCm5XUrADQdfpD5Rdhp6E0p9hJEzOSc+3hklVhEACsTcq202cjjotvb5NCucXZ3qPOsqQNi/kyKh855kdZpw+avkf2eemVCH1kT0trEfsCUwNqMoYJcuTEuwNf54esVs8FouB8+1wDWXYW/4EH1S79dqSEAZZAtU54T4koCQtyRIkRqNbyinyMINol6DA5Xyj9M1FovXP/Be67ydxZ2h5WO1uFzabAlNYpIvjTyZ3I4FJlj381hT4O6Ld8Bc+mx4wkF2y+TbwfRkeQ2O2cfKqg955cT3aqlrmsfDNF5NRpIyZtOR0XjNybx2FiVsoQCVn1ujYTsymDhAxQF1Sle8OoSLxO175DXeGfZZe+jGZrsPcxGZkkYA9z7bdn7EnYhqW/XysYuD7xSiEl+EudXvvqh6ougF9cdgtHmx2aZ7MNjs1Snn2Z2+yGWM7P6DCnlv4ldkr5vn/5sGtzLzWgJ38xoOcu1gbUsRV3v//uFjiCqCLTIHsIYy/VOdCHd3uzKc3keEmff6aWPW0VhdJSRVnkCRtPjgli+i5Eo8LrvRI6hE2CefWXlSUoYjvo6QrfV0vV1bDOmamzsn1AN2M72D5FWvZTIE/yZNNNB1GeHzfMzJ1IqRY5+xe+Q20cz5m/cK1HTHclPN070YvGl6sIU+kNqo2HM+2snLhg86I0vgA/e5KmMK2bSqa8QOXUjx/8IHnjJK76E2m8KbHIFlJgt6bpYDBCQZHleoNSP+xPDp8jXkIoTZ4AxPtYxhCiOwCN8xb+JOMGc9bL3Dt2S872tECWsgIK/MpT2lhlSLMlnTxjL6/0xw6Up6ouYz8W3a4yl6gdZzu+tRy0CbAGaRa1p/Z8oGBDkhQbf+fRQaRY06gPcy7hzUucWnFd/8F4yOTRtKUNDSBi05We3HN6mA9fGZDna1V7LQx3Kvk68b54feB0pA8PJcP9nTXO9IFkYh24kRKBKRLfPlMDJI4sDWC/ae6vKed4oz+7L5eZLPF3PaYVcj6gNWHT7++a+XFlE6yy/QnrrpTknKxzmj3iUCQZ2oTpwCjPBcmy8qzcTkuuxBpktR+2Z2+thrGjD3/lSBZbh6o7f7RZJ/0+ZL/bKhgYiS6Bdd/XRpiF8GEfagWRhJizW/MO6uhYe3UapdyGrEbU6s2mXpMqsp7hW+4QfQ0GsQjjSnJWXpHVsApOCaRmgemHOScmUB0iMMw5E8XvERVTSHXOSSzDI6+871ITlllB/86s6AvXfg0mUASHdIUT41tk2As7eSFH0TNYMasHnPr2O7asLjHS3jxmlUQXxUAJcpFMtBVu3gJqzlLx2+r+nbojzH+gX9ZfOcyjH7J3tLZj4LwPlEJZaLtRxG4Tlz4Wq9QGKc7LC/8lmEMMul86fJ4F/qvGhtv4J0Go5t5MGrGZ/kk76Q2BDvXCLQ50DvzVu5ihp9nN4dq87z5BuoNVinNfRoe80X6+TRpVXj5eXPA4Ws9V/fHQecEDiPlPzNoqJBhR7CpjoUzn3t8P1hs0rVX2ATO/7ZKs3ggwfL/lTO2idcx84MaeVnIuVK+y6dvE+YtpHC38fYA2kPuW/ZSvmDW/tEtt8Yj5Ck6e14lZ76PYLjlCUw8mJRhhEn8dtDuutJ2jtOU+8+RCoCIQP8MzDKb5EdWSb+h+hp9CAWFwesfOpYGH1kz0BCf6rbySR2nzyVcevX/mXkUSN9/Au5mLFNhoWLB9FASFMItzJElJKt2Y09cMljs2Rk5IZB4gF6Bia5MhUhKtw8xjmSZKWJa+TKPqDn3YPErwNHyaFPQjQ2vKAVwlXNnl8yMlL5Y8+CXtHdCOM72KWIcLeo0XalPHES31jL0rAjF+Qm0SrDBqzyradBgMqqqTNY6qGnFuVKXVh932HFbVySnMr840DzyCILmYTEYzpsC7fv8/+4xYiurJ7P0ZPSjNGEK6VuKlcMUnOpnLhp+nEtRFWdLDI0dlJWhZKktugCyiiKG0SnZsZtOXPRFU/Dz5846nig3g2dJNWru38hs501HN5WVicVK0fcJOTZXhJVywX1LeT5z1UzWLOJnahEp1JRlgBLiCrx/0IkeVKmbtd4Kgn9nOxjWCMP8hji5yaODTxTNIagrEyYK54gkwmFkwN3ch7AfUyDJM9s5oXrMrvjpDS4BMRYx9msQcsndK3e+SE5QwRRy2oVzS3SYF6D4KPsOTb5hDLt64rUi675+8aR8LwSA4Nq+sDp2XP5xiMQLhXKTRhS12+LyzqDe0X0tbYGqssJ3Z5j7GDWtiGeg15FOAeBUfCNC4ujwYFRlFRQUaWtJNxAdqO/xFeC4TuPmzOAGpf0wuiCzogliCvEcdEN33ERzmOAU/EhvvO49Ls8NcJCLyRPJiEM405roXknKcnkMILZbsFBHWXqIm68WncbBfyskx6JN+JaOuZ2fIGXmlGFoqnOFS0w+P3yTYZ5OnMTurslrAlfZIge4nb1YB3//ClbyYk8fjrLTpnB/kUBhZ4R9bdDwnAUQ09A8teyagJQc+PbqV9aRLjHG/F3ppxOGR0GZOiavkqCXwmxvziVaQSsJBdeACcVoHjK+1X88stZuHzNXYeVXPKgAXVb0+Yvo2vC9EyvE044a5ZGZAnnErq+qpqgy82tkfz/yb/GAWUl1ncJBMFzhk2/RYTMUXX0hnmjDPIVFkYjPehFFudWxtNoyzbvaSRyRuUhZ3sgSRrAwcBd+1xNQHqxVNFzAf6H2YL4ZsDWbb4Ko70S6w4qV/nWsgX1YjwRwLuVKHwgkjx6xgXjU5OKiUo/QLWlZ5qvc0Wg5ZwOdwa6ai7N875Hik2ZE/X0SYyGj9BYffQ3adVsRMIVhkx/z1jXWsb3vrNUUtKWx5n/+BZAjShkt/tPvMdCF2/0hmlzEQxEp7aBJoeOEPW5gHogE68EzSfHzo4wLxl5ug421ZHTy6KURYiwlym2q5TRCucyL1t/jzxUHtjVv5IRMiVS9eWaEfRQyi4K0/dQf4xErRqPj/c1a2Zq6YyKSohd2ff12HjrUGObazBTiOkK+YsF+TL1yCATCx0E6kN7LQ8N2/zyjQ+N9FMwkzZGEJsdtZPWsqOHNTcfj5BxFFECK7Jz7KMQ8mhslvVTA7bkd7D+4r60oUhxdFESMtEpgfa/Dt+L6EnWNjlVU34HUKVB3JzEvuWh9Haz21ILSXbdgVpgLQWZVZqZ9aJSqgkFpSZAE47boGN1xsHSXsIRgEbDms0QJ8t2T2g2qQ6UDYHziRaifkH5ImcYl4jkXxTPtlFDm2KdsLmLCLv5wrUrLbbZDWwmTUQayV0emG/WIuQm5bSZ6sJXkFAKf6iJYsbOfKHiuoA81rkdfnh5KXAh4q0FyFWpX6GnOHb5vgAMokV46XNpnYSy+YE5e90J8A+oxohllr/M0CeVuGy8szdWWQiUc2oEZgpd2jpas9txEjcH4iLfreAKN/U/z4L1aXPBlMmf/AGZ28zSFdMYGvvmzVMrX3hCwJUg22ghFvqbFxq0yJO0hTUeBZpKpoPsYYXm2w5XLRkngHGE1RcvGQb+5ME6nP/hgNaX84Tv4mN7rHzUTXpC1TI6fE0zU5syc5FVQutJ8aBO3xhsc5yxNubDc9qyShGCKOVd/jnuXILpyO33I4ARzSJTNar/PTimc/wLS87xHDKG4763TMo7be6ZvDCoVIYkKAuyMqD3FN4XiMsGdhsq+AZFEMY6px+JoBGC67EaiUIq+Xovut8utswjT3if7yT0kkL1MxGxna+lbzkIAQQnrp15MQDSPGCoswSuUn7qHdICZ5oa6XCJfTeKCNcFAip58mDve4GTBl6CxyMlFQrVR+NT7A4cV+qmCbNnaNqhVLZ4defnf5OloaN3rXW9vlvtU0oNgF8xev22aJgqR5HbbeOPi9XPBBNwpSytDFS40kGtDZdoGvrU+T/wJwt4gGzQsM3NuL6zinc5z9EBnAiQv1gEKSls8B3Y8yU3/QP/ruMKA+XlFHPL0EaQl/ZvXhKOF/wA6VDPOCYD228QXsx3S9+8Ta0oIj+djKqNI+VtLEoxvdrRPR5PvyS6iKgcjR4N7qeNXARyTLKPlcpxNjP7aF7p8yTG3YDz/pzJ7aN/DP7af2nLAJWNtvXVacDKcfbsixaeix0h+mihPHlzdu4CJElxnmZMpgJHLAgmO5fshenF1bx6yKUojwxiMIH2nrnjrg1c46f/k0bYsEja1WuVdmEiDgwXzpRITxFq/0zuC/9d4zQhBRSBRD7F3RBwHmFIe+WeNzUZSBdIJsK7PX94TD85XjxJixpYV3uBXU2erYFiM7+YOTdBlcnVt6bpvJVdVuF4s7F8kgKDqWhI/k8NMb4+7MZS8m8e7jnnBpl7/vGJ6AUQOMhCqQGuN6goXq2BCIHude4Eqf/EL3BWPb36uvHv9NSOfi8h1omo0wP+5aL2qfk4m/uZbYD8JhOyT/bw89o07fgoe3WkpOIchEy6UWgQqoUZD4oOMl9IfSkIg7MCKcWlJAqDMd5xCMxpJXPrUoGJz+HH+z0A7ayBtkW2dYhFsqhyIIz0/5gGHxYp5yXxK8LRC//2TbHux4HMiej9MCLzwSL2jlYwC/vwsFxS0BWbe6Kek87cw0u3TsSoVvJklQRjVKFeae8qtVJb+iyYZMO+gWJewu9e6hO5kjKrJbWKRcT/XgTUYxky2VqFUSFyaDfiTP+xMhZ7Z3Oqxqr8lurDpVMHVKau9E1VkGfit9SQnVBE7g2xQmNz8AL01dz7vLAide/tjypwGIETt2WIBweP/2X5qzUj7UIrdtiV8AlkDTqaydG6kazYWpyCy3fZ3YWl0dd/J5ipcbrpn30GCNFmiBquA079Sdsm4Q2kcJVopMU9hrmHlke/AehPVGro2i0dxHJFbvUijUXPd/1+B/Hz3mj+RsjMqv3uToHv8s8BmfvwRLPsdNh2XjpxPvf5N6uEsn0YO7+FwiCbkdSh2p29EyBWMNXPnK/TwRkTUe6oLkbT9cNGwgRowfybToTjNS8cy+EoVWW6UkLtRnIWqMqSBbVyzOB8WHfSr0cGWJgW6blVFUiyCniuDpumavp9OOGx/w3dxeP/X6pE1iTnx0f8vIc4tv5Scg8XEIpda1VSyz2jN2vjn1WHkZSjF3/63oJ/xPgH7++0atAuUcwmgeMK1q+JZ5eIMMs85LdGf+1IuFv9kulKNOKHuPuc2qgM7/++AUHXojSWOjIveKIDniWdbd41UbGo0ULtBwWxtMq1JL6ZVjwuPt33daGFz0P2/AtDvx7yHgBiuNJRGOGDSypXa+OWqZc/sIZoIKLZk0IhUKZ32pKSTCrAWp//qTbGC4ka72AruvFOJxN8BaTz0GLkrvCE+LpknCq9ynGij6tAt2O5ZcSZ5qhCr/UCV/+yjrIxTY0HJfDwdlqB7Kya8kCwrnqw5UVwEyCiD2EkJe10cJbn+qq+iK1KuZ8CFsQ+7mG4LzQp6GpByoRSnGrb+v+KbTgmN3/ED9NnEBYM17s/jR5ULO53Gr2h0J6idwpd7WlXXP4AVukdJ+wUczBw+VNQM68pm2HM1jnAlfqG3YOUk15HRLMtoP6eItpKhGPxUZivGOAXbUJ2yefljbukvPjdWi3SH48M3LunqF5KNLyEmzMdnglFBzcnNn4jZKdznD7vIT9UwPdeuK6TYO26L1wBmCA9H6zLW9N/hMSpXGNFGgvFLIrjfSCkM8D8yCvAQaAaUqz1knHzc2ONOg4Uc8EB3xxsQGJEKFVj+KySNkWnFFpd4unAuz1lEqtSN13wU5deUpR3+zbK2WqQqEF12ZmykUb4jVnauF0+wVubgiNeKyArhU9JvPa3cFIOMRrVJotoFY65y285jUXeKDpSWLlwShLD6tsetDTDnZvmlHOu/YSZY0b7U92dz2GmYQ0ifZx4gOa3hyAr4a9YWhzCpw2SfjyiroiVBOrZSwlPGvIVi29gcgobPNUMqlpR+ATGCZIlz2WjfEmMN76rx4VWBAx0tiKvPOE13E9ExHR+0vuavAfYWgceLzAJPFrEUc/G7gPjjVkZ4XeeSWbPzEZdmjFO4FWFxbQy+6irCNeA9ch9Xou1cY1CyuSzZQD2Az4ZPVBSBtVaB4wk8JA/b55yDu8QESFqyz4rU6nnVvD1MgkUEKtfhqWnLExynYPq0upoXfQHKT6iEdMn82rbNaFdJvJtse+XKJzM7AaWIBwKvVeqtL+qYN+XlYyOHK9TIs5+T4OUwFHXNKu1L8l0lW+4C8Og6UuehXEMvJwJRr1ruyaRr+XaPULTK2J1MGFgs3jyZHsnHket/7/0ZwxLGbI8St3l63JNf2H2pTqXBnhWPnKuX9POHqMmsId1q0kTMsxo1GPwNCHuOWbsnAchOPGhFpLdV8o1v3zSnGiGC9bk89QvCTTZbaJcvbXote2L1cuE9gRCarIqiEOaecydxN5sJ/cV4S8EwjSyEMEP2AUfVwr/dodacCUpyVMxS355bNqugDH1o+HRnhBYZk6H8h5oqpwS5J2ozqnVf8ivZcGuP1ZpgQlGe1rhaGyKy7WvnFJ/MO1nKBDUA8t4BJrmykTDPYE3B/S17ZQH4VUsnmmAwOT9GdMZQUXvVKhiJAYpnl3iDZkOUYWS2ABiMh367VnZVR5C0HH93KMtA8Xqn7KWnhyyxXJ8ZXo8loWAjZsuF5MPDytqkStq+gwnrGt42Glg5sT3DJVJJDErX5Z6C2eJdgAiZDzDahgHn45fdaOwXhezRphlet0DgvTA2Q30Of36a3+lxDpmEkD5ksJ/YaIAM3MDhgayXAs0Nuh2QOQ3AxTKRViNENSq/vOcZg5GcG3bpY5bO/IIJaKsbjv8HIotqL8KwpTohAHt8mGzTWsSDtUxkb1fjHB1l+e1+Fjd8kkA8tnFz9lFWYxSJMQDxGcUXP/finUY+8Npkaf3H+xyS444twm8pPfMdfwG23QcwhCzKszxsxvbSevkkong1eG/LSnztMNV1K2YrjbVasVytUa+/9S5Gb/TuYpICtog0Qb5T0SxjUgy3WxAFCrZAey+hxJJ1G0Sq2GSlNCOe+tFGeIE7I21Xt8LI8HdL6/vJ5avKuz22tO31xcd9RLkFgNM7qLgSQsd/N/kxkmi+iA5mAgkl0XFs0P8o5UleNgwel3k4l88nl6o03JFWKe+msxqgPD0LvSpzT/3TBPJ9iu7k3efSQ3KqNnvLDuxMONZe9mmo2nHQKX02pvLTD5kg/UFL+LgPryJwdnuvpqGCgN6m33xdi5Oe0y4CxP7FgThjjnLwWRvB80S6avq6pTZIkulFMN14xwKCynk+6DMNRkl5RelZBDN9R3XEboMgMcNqb3n3jQRGKSaBc/mSq6x/irzA3GlAbqrw71dLrAs+xXkj7qTMT3kpATpBGJ9IjwFm4pXKigCwjGvOkG7LJbbwDEvh5j8NqMxXFMvmkTJc/bX7JoM689EuCCimJzWWQcj+W0438+gB4WxrGCcYxWlMrgLQDGKkJVM1vgs+tkGYVjrbWxWqblxzTy/4g2MK1qg3FZ/8BrjOc9M6lBzVHl/E+QgGm4Y/oBCI8RF5ARzpAknTuHpCB2bKNnQH4Y0FNJLXJxUv+R/Di4ZMZyyxhbx/s2KhCFmAuHJgmKfbsNSN0ouDkevIZ3SOFaStmJseBD0p1CMQJOnZD5ITZz3MaH4n+J+Q7UuZCqG9B0q4NZlt637vvfvH0n8MuikrERr+XHr8/i3vs5RFO2iXIg0yF4kI1WjaOBEG43lEuhW+ttBcGgReMWt8uxotUDTpFAHDgI0QPi4r/Xu43Hzpa+kqwfoOeGYQgs7SWnLjvphME8mJNDrg2Eba4d2NlmxVmlVL3P0VGwLsUtnF7x5lFwctuWBY8JFAoNseSqVkycUUrXhNqNXKAu1D5mU4XJaZ5y7NroW4MI8Z8RCRJQWJ0MbSeRO06FYBb4OzxpthRSbNP4p4zYmIcuYim6AmUahIeBcX1bZBrt6vx3/AtitBrTsV69Zoo8swB7YxwN0Op0rO5/KX/ecFgUs4+cEHAwKoDd8tHbvGXobYUF6o22q6Mq5hB6A80eHHG5+BC5wgrVPS3HAidqI4d/BBrz7DB5p/dC5GELcIZKWlZJLU6+HVj/w5zchLtSeJX0Eo3QtNi4PjFMXPgKtyxUOHSvpO1Ggdu0ZWfho3k9bv3xkNM2Arh8ZNKTFlU7BRZ4W0sTlPe/KeYwQ+4zUfXJ3rSgk7mR99k56zfvk6F5sWjaYmgWEB+1WcHF3OPpcg+GEa84rHCNTiTJsgz5+gX3roXq56xQmJ+TY5USCEAkFPbG540798xnMVMCqSnlZNEWi3Y+MeJ5xe0U6T0jMybopnjDVTfQYMHWZ+oUc29cg7DVKQ6EOVsp29IP3LveUBCxRzUdOBAPjolLQ1B3EUhE5kt2PchyyZ+H3uWrAY4Q4hsvsDuaXHRM62VbkvP44rE1iAm3nTaw3t2AtZIJazOdFV6LpSJNchzEnuZXlLgIm3NYgS1Vw/RRWpHunvHxXy8wN0fb7h6MWYrxmvhCFwD2azLO96XSEn0QoF4XBFlYhEXrqAUxK8YhcxLntoSumdQWlPA5zoCdJ5XUfNG5rCC43k0R+li0cf+xeaz17ShpCHbPecmfEI2gmfk7S7T/OX/S/lxsgGAl77NMyOT0sTPK6fisxHVUcWCFkPndmPl9VDuyKjet2EjEOZmStjSeQID37A6uxEPYz/lHGNNcbeFrU5ss6szKsByel/7atTWsSCg93RzRZZfqjDRqxEMloW8Pa3we3m3/1ftYZ7kMNbEhzRww6QQt/hW3X2xrS6TEp5/xlUWx5xYvlPFZQ2CBiKpNxEaNvcmxOhCe8xLU6oKJxCMjUWGC+I+VGxHkFpOkkdgxnOQ97UPQ0Ofg/1X7sYG/etqRBx07gL/Tpe6fBdCGQWeUwYVh5X82gTbdetlMlZ4iNY8hjNSNFtFOq2Se2Wa+3V8d1ETg7bSgEuOC14imaj1uwjHGCr0KiLqbPOzw4TdTrd7ccgJvcnZ6sA6Bi8z0KILQlInr+BXnYwqaPgfsU250Rn0p5J8+tm3vcxk2/xIzOONV4UC7UC5n+R9LOikp3ITKZlw/NeXUoVUo68b7IWCuQV+rtEow42v2W65ScI4zrQ9DEYFsxtU3eesYfNT5H54SJwhQMZK0PU2h5IOHwD5esQ3PoFfzduxmNgeU/wS4PapYtdX6LhefPdInIhthmpTD8yTECm41jWfJU+66VZ1uhDnawsQ/gBbRRlJdgIuEWxIYr9JpDCwcCGMv4Y4frFr1fn+jfVpsyaKFWTHC58lIj/A9Zp380FtyyGQNFXFabZah91UgoXgp6yXbGyKsdtrJ9z0y/04Kk2pLOQu0FouHPCvXx1VMTwuNYz6uAxPYl6A0bYQOaix8S/sQeoSn2gy04gUiuccczqJvTD7HKBpYYhLCUvLbunD75NaHmfKeJVyB/x+/JacLM63LQZM4r8swaN6MxRLz6Dub2aFGbS+iahJjt7ukXj/YdMCnTMKy3hEpdJ8Gauub33yinl55dpq3973s8ujxk5FrVSnvtKOMkI4nomfYw2Fw/rSo009D3IQe1lD0BvQKqlaM9T8SytPx723PDZfsZTNp6trpiiyQAZgvZlIvq05Q/kfgPvf44yH3Z8o14pX27vExaYJxdXgFReFaAjUnOQI1pL6fCAhf93wVPVAU7e8ktcfRBdRObDcNVKrQaQThcEYGMP9AYNHpckJV0JtlWLCxGoAipcikJ+3ajh/krGn2Q5TwEgc0rQflrVZYJ3ucoW0W/M1OIcNmm8j0LHcqzTXYkeFB3WJSqjQfBHSuCe56LBJ5Cg2cl35Y1zkwWG8pqONoPIIlOpGXjviPV1EjRFiUYTTGQRfR/U8GcGHLqY2pHInZmf5uVaMbcQr4hEq1JQAFvq7FHGVYeGZyAOBjujZ5WElNVaE7lb2BQzRrtW9giITYTWov+amp9H2+7GJbuxQddl/V/N8nLL4kcm+bLQiSLSOg6HnQCPNkEdb2QOo/kHSOzzhCY0g+wTKxJ+eu8/7dJT0emsoUJ9Esk28ey+AUEi4FyM/c0AXQyBIE4l1DXDR1+cpqIlZH/7fdiIqRJI22pnrfGWCmj1bUua/ig5iceiVPjYS1VW+JFQZnx03oe5m/Xz1MwpRZwxfoHe1xWGglq6RMJwiNToRD0Abl810QOtMbFPwBWfcVgW/fA7YoLH20jlOhlZmdLO53P9OpqZKh7oDgeqxIZx/aPsHcX3mZ2zZlpxfb6vVzvsjiFgu+V/i5GnnSNJ0pR4iJAfwI9S23yRNawtkYonV2U0SRvKtHhJHsRdgpltG9jwYsSrsmxEcQxA9d7uqAxY6hAnIDpNBbo9CSIMHY1Y2D3rq/ooqhHwEGjo+Oz4uqzvZGK38Ilh1mvcIy/fK8Ff2nXbGyNT6BpkjXVN3nfvkY8DI6VG8NxggkzNcH5JBc6gm23ezyXsa8/PmmraOHbkRkDdnKHps9yODFY6/SjHHIPbmjtrxHXRu84OauR4Zd0WxSPKOHLqmKmfbx7BUiVo2snD5JXx+94KvNjn4a7xGTL6vaq8/45d2LUfwdqvH061vGLrRpfwLbJcgTgnEFXwTeGMwfitwArU3fwy51rh/sYMZvO8S3SlLsyeqe8hR7Pz9lOE3euR0K7Rn6RIdwzkZ2E8eoZ8HqReLC/nkw+KTCX2nZNi5YblD/zTYdDN9IosDCsp8o3NCa0cf1qRMBKek6lCpoTuPYG3AJmxEzLAzJYmmvyWghdw69ybEs+CUz8qR50en1Ggkr5wdBuwGxUCYF9h39uMY9XrIAaPq2v1f3YZtET7jhCJLkg51YRxT6ou73l8G24Mxr3ZtVL2t3t4VgI561T00T6fSr0XaZghatt0DglBPHhkfzoSV4BH+q2kgHrVNWfS4lYKXRalghAyckTJklpB6cxoB7WBkxWCnXkcO/mN2mfSl2Tgnvz1ZuXW+B0PC3MQWlb4DfnYhRpX+Xd2lyOvO/oyc3dIVn9RSUy23F5IQlBu8hxIRnXgqnN79R0WXNok/GegRuS3ZNM5nkVKP+ON8OliyNAdfhWhZseGXaFOl6tz99iNkmHjtrvAEWGP035/tCbuViF5Xc4nW3YFuZoqWnES+Lg4IlpbQ775siDEVSQ2XakrrKgMsH40zfQW76q4EVPJtzs/2Sj9VOs6zEnGjZIEkmUIy9iQYuYLrfHTy+HKwibZq0lt3dfyTFzYxJZkcOO1KkdjtFHPsHAGZgUgXAzK59oV8QdnQPq6u3idhBuaGreKANaLvSlLVMqSufqV7DtRwO41Xmhe8t4BXV50Yt9/XNcQ5iksZkuPIZoewtxVe2bjL6btIyy9egxJfWivJFqLKyO7LEMvOpMhjAIp3ySy0lzyOO+pCwAoIyqAIC3tlaviE0dovzu0+xgsaLguYPvnaIxeGxeJ/EIgnHv30VJbLBP8Jkxp7Xk0HQUO5mG/XqjMGWT0riVg5FS65x3KMuHpmkRFcau8RlMZJwLZOl0BVuBgtL+ZKIzE8+l/GViKNXXkqUHgpwr2/OfO0HwtHO9/e3z6Vz1IHVkqTcbVhXSNrVSIqp6Fo4Z+VCIC3m0KdFuY/FgM821B5hu7lcDxSHwK9jKeS+L9wtKBu54NtytXnIeV4R3+QSr9Ze3MI33ULBX5mEjb7Oq1xPMIgMX57IXt9+f3Unye3nNhlOYx80Z9BvjuRWjCJQ46Q1lqGeACpCsHA5rl/PWyyQlc/OgkU320InBopCCalJ0o0xQ0p2GLYz7yAlOU1Rf/6orT+MS4IodlYTuyJc8cAj/M1GQfC+Zc8IjPBIS2Z+3IJu7bNKQyaspvqRfjftg8myEAYZQbKHBMOlrwevfZljFnB9jrgVVjX9qUtJxFXUKfc9inE18M13M0mGEcpgBN3ofyw65M82/rrvAaw1/2tLtn+ZPx0qzdHDu0oZcCzppWfjHm90D3/S/MPhCrncXNl+PicK4A5oxGPGGIoEF9rCZ/JQKQvFISIJvaN22JZOigU8kwNnQXR7xQZKMuCeeEJ3WgiNlkUs881cp+pRvAtQznlh38BfBAvwxu027mg6s14Q5i5zkVTJ86ATDXIsIlsZADzc43MQbagwpQYSfd93ZyqSHv4JSiHMYqplf6GQbVPEaGewCA8tfBykj9IOQaVdtNqM6/hQsQ/MoX0bTTBo7kAzASmHzzhlk1G9IcYFY/rZJGBVZZh0PM44CMKQs3myoKYYZ1JWVUH66s325znNFttGVz8RFt/1169FIByMu8EpXT+J9e/l4Daj1dHiIIlmlXe+KFyF6oXbCvfjn5AAquOWKlmjpjs7bag+Rj88kgDTZqjNRatb3/aut1wVPC9OP/gt032jCYazi785c4hYXBWxm0MkUI+rk6h+iemiGshf4239WmxI9RYrmsbi0xjs5JQz/vUMbRMd3E7gPdyuinzCNbfk8V2YHdzPpg8UWIGRp3EdBkheEsU0DttT09XhtTFse5Qget2jJMDpbldi0n2LXpepQZ3RyWYddz1TTSnPtpanDY2gk5UELuOyPZLf0Qo7IkTiQ0m4nCxw8zJgUT2DuhMOzrIvfOpruQC1eV7JZ6sJ5hVWCa7ZjJWew0Ase4pgjG+FzL7Cipvw3GpWKcsnnSbs1inqDsoVnvACPW/TUOIVO8+nI/WtYDp3iIOflTgMZLAklmzkDR7WrWb4wwoT0vrSyM51nh6zyDqMJKVieDJAq3Yc478hyOCSWd0B3GTKl7ZSHbNFf25dzEVlk4jqFnGr8K+2shr7MZKpJRIz+W0JMs7LyCPpm4lUwkhseL83c6TYQoHqfyGV5h5SD+Dopke76+dYd9sOFQGxUqfJW4het0rU+RX75s2WMuHeoZeHqDUL9HhPESCpBc9sWc1T7PFZE6Kxzqg8wA8MXgGXA0lqHk5QihQv1UqIG20bWyo04BIgYFNjmI8wG3YP3A22uVTL2QlDEvOSLBkTVJXfgEypQfDOr2cZPUGcUmyP6cLBJvLv9ZryzfeEi6lwHhptLi7/ANypwwZbcRblBNF4G/kcPxxzgetpyzqJNKe399swgaNyBpyxaBeRlAhpulTJKGS6BLjud2yhdxkqSfPCDR+IN0ACbKRbxKrNDZYXuIGKlC3AwDdjw/jv1v6weh1piLH8FyyHZweEYVFYfsDJ+Pa3TwmYzPzpSBWIlXQlltmCV0Nn55vFTTgY3D37cHbMAuXu/UyXMSKgNIO0FsZn7WqOeXSeKCa0XXmWuVvB7UuaqyK+4NRJeCWmuG+MnqbaPUjxGR0KoADowlxLr70JlggC6sl9J0i9XvWcHbK8MSmXT/yLE97MlSlTDTIp4bxhbc+XiuV9a43qO4Yll9uCQhb2LpwT1x2qP6czKvX9GrxCi/cgbUz0MkJC4CE/ip3k0ynaBVdY2hPmIvNhvT2eb7in5geSmpi0ozQlDHnMRQudMO9jjj+YCwX45AqR5anvuO5vbm9bUTp0lrNL0IShWNy4TMErMzGL4ofDDVF5k4zQKWinWMCwBXkn8oxBJJXRTqZH99TIzuhHJSvhZWDlNZRnAde2kOaevv2yYGccXw4AX0C4sE3Iw7ydGT0x9qG3zmRbKYuGY0LsoxRw5yjp83BAxwT3N+gS7FIlvZIXjxk4OK0MQGEnNgdk/2eP8+48lWbLZracszcBaN9YA7njfEA/LMSk2IcUNVM/yFyP4MRCFKI9zYziaz2wf4CZnXTagWOnkxljRBdM568TdU6WK60ElXHFpLprwGCwYbiwW0TCYCIWQoXl3pCbHYBoAd/Sokpx0VvEwb9RYl4agT4s6F+bJVByqmZXlYXf8EkIa/pMH9O6qnp/bYClsNhByOYgaItN0SsnCOjAcfBtcicWV5TNadTHS3T+UNQz/HLQwc4gNd2IGoaZnL+scnAwDuzOWTcdUbNmciYbw4aZThAD9JLv3Kv7++zcY+fLYXM9wnntQZLteLDlfFDRppQu2MRAMqAPeGGNYMCCrIx3PzO08nY3VdVF+FULmujIo3d+nUjw9uTZSqu6DzxaB3OMk3RLi68ILbbLDSsHklbc2dPQxNWlkubJCdu2RvjqVU8+/5zok6DEULPdkkNyJrXAjoB+wIyxI/+eCLxL4RTDzwmJoaykjum63Y9GRacJfRi4byxUH4NC54A1DlGvigZRKREKurHiSIdeXK3GRNlo7f2zp5ie73ZCTmb2N5XM+Zddhz1VQODptjOJN2/9FOlkoFvrSyr3tFigwXl2FkyNOXTTZAXXhn186IkwVJ0ULLzKKnYE60aRvmhgfi5yY2FDOOzZQ8v5I3FiAe2cnUkDNVaMWx3TLkUOw5+CFR/6nCYtJPkedUvIDRFqJC7/PjTlwkVKoimzee0TLre0zFQ6k1brjUktynyly5FCceCySf3wH90M3BsTPvH/tZEf767BNobId9/b3nkNE/8nxCT1HIa7HBHi1nHZAX3sfx+/yfDCWHP7ezmanyCGQ7Nq0HzriGe04DHjUDoEENP9y+lB2m9MmSYM73ymQQXrlNu/zrVUGnGd+81ZQSHSShUUKlR5N1VZ8jMbKEgHgAH/Hbo2NN3xY5XdtNYLYajoFcjaeIsPDhTk1Iu9go4qldFDIRT3m0ZqxPdARO0DyKqlBvDBYzGu3r0JlV9XB685bdpZ7mwxayqbwyjteqs8yMbN0wIlF6pJJTEJiDC+VOrgquOztt7mQqq4g7yQgZj3wqt3V270eV2KKy6NnB3D5wFuaq6Jaz3wVsVZFASLtcv4KHEd3JJsYid0CYeFed5d0IJ5d45TCxFfodmt2Cwiy+Hp3Pd1JN5dWB6ra0BuNkP1c+SXEOyelmgLdIAPOznUp447fw1CoK5hDWZVy5MegsFTsg9rs8CXwgvs3o5xZlP+oaXDpnFum4I5YEnMUEiZffUpfwNmksxdOAvBgxef8EC2DMT2y6qUHahzvRdsklEWk4ziAedbcQnt4QdpLwBH4129Rssq9c0ZbvXlzEC8fjNL4giinZsc+gkr7TSy/IkpMYvJoQzKtHNUTyako2MtTkNGooF1YGFyALtSKRqBCgpen6Z7cf7yU3eTLGbLDBDWkXhHftoagP3V46h07HIB1GQAk77h2D8+1q0CqN08JhsZpG9avrYyqPNtpa3xkVktrJV4kODLULzi5pkGoJTx7+JoKQw4/codWrme9nJnRuLc1f0KAj/fw6+Fwt8at9LuJaMWEhlB3luTlJU/CWxP2m8qIGxTXtOpl+W77sDjvd0sFo5a0oO20ZVtBfc+2tYEkZHS9DyIG8JdNXn0a5XfH+THR7+wLdK1/XOUTJoOLWwT1T7LTYAIV500mcVbR5Mqhy6Gwn1UQsEcHzA5wFaTYyOdF+GfsK9ty0fPvL6IFt/WkMKnN6Jl77CRsgjjWgBWUbETASOcQsWOmISPAb2K308Tsxonw7f4mtlfGtyza8dYX99NowbbZEVdR6PHavkfZEfDGBVhiaepVPwLOuwJ3SkaHTYpMCQYErPLxiJwloRFrHcLVFKM/gkgbq1QCQpZq2cp1f2vqfPkp2kZs+W/Z4WnLkhGGpoKMhEeIS91UP4Yzr9jVTLQiq9UzlLLUqwyhhuYuRrVN2jMebU3oAfeoF0H8PhaaUuVIxMNKipK7CCEzTIgdBwzDpu0isgC0aCQX+XoO6vASxuvBECSQRrs8WZw0AjptBFIZEPVinrzIDDMR5Hz538EX2TzWVXrKvGL+hnJJ9ozuWUZhojKizvuyBnkvMMAGrYFdVY5oDHhXiEreBvYhu4l99VZ8j/JiNsPSw4Om6D0eyM13kP5axCxUiuzmt9y2i1S082XxQFjJHOU4CsJXWy6n78cVNlDp/N32BEKvCgrbIz2s6TA5TSfff5FYez/Uhe60pQti1AOZipynhrP1m0zNJZhkIrLe93JAoW+TGFEO0WuqHtwGTsBrMJNL2YM+R3nXIbUE4nx+bVDonC6r8xHEnFV0WtlwTRhT0bcv7M3r2NsPpni/WaF3BTuzTTKBbqCuFonLDvXxNQNRllWmS6ksZSLkZm7WvE7YXoM7/JogEhqNbdxMs47jJ1Afr1IlPU1FEkdRyHtZhE4Q7TgoCwqi19Gt3CNPoAfvy0wU3VhWm2PY/qi6uyOc/PNXmtR/mL+B/UrPcoKvso2Mv7Hiv3Fs+ZpdQYSRiptxDGIW8QTFDZA7ASwAFQa8xZx4GnLkhznLL3oIgn4i2YWiBsoGr+eeoK9OcxpQcsWVZmHwFPzrTCFeH1W3zSIC9tE1znFEddmtxwIHIzZYV6rMnNPQJ1/fIe0ICajPqXrdfM3zoa7ZIlG3RwdZl52NcjkNI0QiOjTEXIvYL2O1SW3AiT7cELSs+TCR1Bkb2OvQOHhNpG2lelrpBnvfzMvFjaaKDY0wmTHyVWXCIIGj5bnDbj6FwTlSfAW9IU6YFrMjb2FxYZ3GU486glMC4jq/2zRgmXsQ38kz83I2KK73oMQNA1Ah5Vx38EBJRKqqjUipbqX8K5dNkIqek34agcBwnqMHAfdthbAP7mzJz8Z48dyz/vw1YSE6uEgFGuSXcypouJ0RzOXTmWwnThhu1YvAYH27wHOZiZ3FFHIN30kAvuv+y6LHP1+EKvOx9iyMga2OaZID47LJrnNZnkdlcvPi8mNg4CmDgICPqyE7s62Vq39z7Y0MJji8TOdFI77iAgw5kA1mqmD9x0p1cC+2TI0nSxl2IhhSwZFcHLcMbjynMRci42+2B8IjWMe7tGfCvKMAg3dNOnpu1lfBflXYBhoVLPzuIlkFSaIE6licB9FaRZh5FNxjE1KYOkaR+/2Cwf1Lv/0Ucs5wdCl6KeRa43ufX37nUqd4K67kB2+sm9uYpT5DdAAH7D/yZNmz4w3AOV4amcvfGycBvhw9V1ok7UagxHhTRcbi8G4Mm11OMTuvduuGRUPJuAcFS26NPBI+AAhz+sepL7EYJYCD/a5kxF4LOVRHtVDhqW+KZu87mIBHin1Asa4JRVYQyihSHpkcp5sKzVSDbBgXV+y+Pcw9MjdyJpbjZ+NYfflYIl0MCOVzYL8qyqBkyb6glFLQxgz77/Wh2d6yZAMDqp+YxX5oKvm9k7hfTTQ2kZiFx+D956qmCJ+mQbM2lzsGMEIFdcBfDWJIgKcPxlhTow80tpKpG2pBkrL5BD055C2uqC0AGxz3o8PmWTx/jWkJN+ZXosqVYp6Xzj0fK2RjIcQkD4O3mg7Ed9o6n+j6ZQlWld/NcZrRDszDT++P1/jNA+FJzTE+Fwt5togqW/W3OR9KZDonEG49PA4J1MeKxbUSecrgMzmmEOR2s2keR2+3eB1k1EvYg3XuAN73ZI3Ub/mpAWJribqTVGGp63DMnsIAlZFZ49yrlUcK5nmlpwwQ5WKLdIJIItyGHfwFaI2P5OlZz6m9RY2SzYbYhBzhF+OHEc8s1AbZpfG5Nt9GOtdPr8tNC0uLopYVo8T8Bmrv6h6ZBQlNyb1BzoHZ4rTwhr/WXMAg5owBFYTorqSX8xR2w2DjqyGWApGOASU4OMhsA8XQI/eoPQUkaGNXorik0AP8YkSvBP4JxU8NO3UX1WxrQ3QkYTOUCf1Bxe4lUpxbTUh1eEcwUqNK5qnFeJ/PmH6nmvA24CVB2zhSiDy9xxPBVVExJGGRvTDeH/ZrNAImXUoIFD71dJt5X/vxRKDZapeIzwfpLvkLQifRWUfr/1v7UkQEm2x/yw7fbtIn2xhge8YnUteI4V2ciuI7S/Hx9edR329r+xXarVVvPrRWL3e76JHwOQkTZN6Cvd2EasqKziH8dRuO6a70uGBZKkNm2vXj/sA1MNt6KHCYzWb04r+8xjo0/8V7nEokSB8PgmMw/JLfQB2+aHwFy28IRR4TyqYWNtv0A0LOrdQtGWB0DWrxYKqFfDhnEsIl/RSZ7R7h761coKvX0mRyt5yeNOVZnrev1Xrxl1xBr7HKXy7i8dicNn2iKa4OlEeR1hL/7W9AiGoyKVP13eM9HOKoykpPzNfweh4K1bdPvPhMCv8UpWdkzIR0vYqKc4/U6HOsS7p5Zuzw5Qlq5YUSq3S53yaxXkazQTAhOvWNjHPp8iPN3mvp9DWkv/gjQIl4/D/HOvknJ7DRUQI9K4oJYQKSragfA/VJ2n5fC5od51gOih/l9h6K6FaxAnAHtREz3El3slaDg0Do3krGFFbDvu0gSPMRTMseHvdGCpv5jMcPywXTy83JI5weRyM/01RHlwCehre14H5pqPQj2xNcm+7Tv2UCAI60EjZH6Ba2QafavLN2ZsMsze5AOV+AMkdYUMMJEga6qaSChwbnzjKsbWAb5cjc4RzBWfIoYvof6AuRNDv+84E95AYN+r8DqyHI8Yp9jPi/f+rO5s5+SVh6k/kS9S8g8yX6kat+Nllv8lG3pmyVsv1hTRGfBUKpCkbLDTf7KWrVtSsz4JTZwq0+BHMWulbaHAjmc=
`pragma protect end_data_block
`pragma protect digest_block
b6008cf2b477ccca921b2bf0f3ba96e5d13aa28db94f3ecd8fa3f3736c0d3375
`pragma protect end_digest_block
`pragma protect end_protected
