`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
Si/1MyAdtGZd3a9Qwmf0K0M5guFfkH21v/d4Yz59uNWb0gUmRx6AnBapy4FBvswP3+KRa4d5qHFQCVIWACPXy37aHRJNiAYdCbag1Jwspy3tIcmliqLjEFcUTmps3J336a6AZiUs29mnXJI47+u8yvPs5QW/AXrmYP47XnSGV6O1d6ewUhywp2nFTG79oLwAR3Q4wYf7AcrV0O4x1M+k+KsN2MUPYTdC9Xtw2+WyuxYChV0H143MYEQURk6mhIF3AD5qWu7JFdcr/LNApAvOEZ1leWYMVnTeNtLdaS2GJ/MusHaX0ncoJrKJDVc3c3v1TwwxeXPOIJ2xRhjIlnIQ1JfHNoMZRaEc/q1KMa4kGKjryrc3sV0DpXwlRDTT12ux9/RI+732BPt1p2QCc8qK9P56SufJ4tNmaUrqZz9ddmINcQ0Zg1AZYvLK8C3RkJIGbsoKjcbnW09w+SMiyNrqqOv7PGMonIWJlcoQ5jxN25u/zS7URXxDtg65ahki3tVkquDo+7XKotqo+Doy49KBwdNXxiooH50Nbjp5Hg3HCZX8+FFJrQhipReC0ZDedEhW1SyRRz5fVmqPGsMo9/zIiywGwucCb3GlUEzD0LRBovSsdzQlJMB6eLV2uksfO1KsAQ2ku0eCYo5/ttL3O/VcL/4seWyw9ylO8/AOWCeKR4+5lU6/UZqLUtgXRnklyTl2iNEnsaQevuiVHKrG5rZ2mZBbr0zNt9l762+tkcA/g9kJ3h8UNORzLzN9kbg5d2Mb0Iglvu3gaw+bUDf8S3acLHlnrzlo/d0Ytk5KgcQRMSq8zkHTldn1Tw+reZx5X78AHH/4aLvdoCavOA0cXApGVxspqEGYxSP6rys6i0fOViiBRfSUB7XR1GpucOeQZC6Pmu4UxD6Rwv3v7uxcL1gyRWbQtJwlxQTxGNmhabnJZeRG9R85Q+XkWe7A2NE79dy5Sl9/OMa8xNW8mA6nJCfMSNytgdFoz3s3STPHZraln1qzd3qy7fMl2ulFSwH/Zk2MDDZAgYIQ+Z9RcYsKtX5QVw5TAL5AvTo0B5G0wKhOjS0rp2YzOXQPbXGthKgxPLn/zTlR3JM6qncTtd/J1D4vZheRh8kiMcdtSGBt+r3RHBp3nQGXcuC6A/ymJSKIQovFuVXb+mXwZJTSZMGGysb8/U9NrnQF/4hLebXqAM1iOHN39lSOyvzCAPucWX8TSAKpK40wJ18A9q+Rwhbk6Mv8ecxcVsdz9kCjCByGdo5u+ZHxeJhGnRAZzozO8ZuVDTvKUhz4SSN2u7V2yIwLGxEbgI7Vyqub9RQCaeamIsYr7DxJyR9s4QrJ8mrkl60u5k3YeJJYe8/QQZaTopLeBHKp/ULwwUzO7k/M5anX9UtGKhLenvE8gYnzZrDyEM2p82z1yUi2VVwxL0ZSJg3dE/tr5TZu/C8HNMfeqdS4kYQxNlmgwl/mtn1PInH/wqEx34T3C0LVHNS/TVRP7E7Lp42e8LA69ouLte4aTgx692SNQ5s1z96LJwLpB3rJdFlpb5if7LusCnvZmi1d9UNt2Cfb9+YjLNRUyonibGlCRHf9Z1CXzDBiDUT9hS64IZx+ZivWTt9dZ1eAkt5cWLdyj1tQ3lGbHpgRJBIKKFWZxiKlehD0U0lPQN+k7YEzgZ7wEd04ewjvgi4aZOR5cEwKvIYdG55o9BakCiQZt6HPb+X+PCqWBgbVd4ZW5deiMAXUmp6zrMGLEWzvOlhqrNNJMd+P6XsRAUnrjDdP7dixJ3ryQTiQ/yJ1Muw11mFJp1BGkoWWn3vmsWXWxyIQF1ovcf8yN9z/nLWh8lMIGMzaZI70zPjgEfP3mLukYG0jAITlHTmdH8Acn+y5Ejuxa5pjR4oOva92ZyWG5yKx9lKPZXmEo0NyaBPhpXNuDZwqnZ4zPU4yRG3UgXkDawztUgjc5c9R23IcMlf7oxpvmEmXWsEbPS4owYC22VP5DX8sBAUilrJnd5lFZlbnPyYzEsk7zUGdlZu5jtk1bm0bWs/xqrjhq3mVGCGqPRPaNXQjsYYekD51EavCWyFnLB9uf16kEWOz1jncu2yGrLURWt9b8N6h4ODWLMOwaWj5ExT5FpoWjsN7KGmCi8XqO0a4YmuEYZv8zF2VTw86yi/47UL6l/yT4QHEkSD1aj7Pl/2eO51UsHh9cHW7Of7qRWysF7ablXk3ZhO5V3MqPgPioz+rN+X0bnS4mo4ET3TYZoZwKH2txl03l3bcmKytbESevJYVan0wK0wiloUr+wum5CCegk/ibvvg37ai4bdjPragl1rb1l5o2jtFd60kab2dJclRLoxQbNv5zRThx1GvEa7wA0FVBpdVA8dqhHYQ6VSZH9brOdYTE6KZ7gFYsT4Os7IYefP4OwOU9DkkC8iIMggX6ADXc6kVt46MLMG7c7cj8PRJpFZWC/NOBv6Xf0weyG8ZkdoPVvYFRiA8VF4RN4LAHAQLjGk54KAW4Pf8AfGqgO6mhxmJgYn3eK9ju/TCevwl85+6r+WcS8YaIvUF90P/13s1MqR7vSW3JuJrAkFJy0cT5x50ogl+TuXeatqA7tHoZ1dZFE6KdhMcTINF5WduL/3H6xYOK9rXDs+gKHU2Qnrrrt2c6W/ndXLZU1uExfrEaHsXNls2lsJoNuB7mRVTOzdnIbfan8IdHsFpdUgxjFgg33GY2u5Hfq6uVt7xJZy/3J/maTWie3/BDcEHYbIx7nLRTw74n1zjsewRjKSB70JDR/Pdv80h0odsnn5Yo4zi8TJYsgTy9ySJNLrQv3MoXdm3Kjv9W13T5zdSUPIZNvET5a045EGb4fQ0Be/0o0FRwOS+b2LC48NGsI4/Z9jbpCdezUuUeO7hr/tAmfzYuTaX+RAAulodfZUtOH4fTZcTDSmjb7lgCW1HceuLltoEU6yGzgBOos4WuAz9H2rGAgijdRMFfFfHMzQoRTw5zFAkIWhT6lLT/NYoLEyWiMETRWxU1HixLgjcCo9MAOe19+WHX6PJykeUM38YbIldk9h8dM+TRojeoRl+ubjh4uGuWHTuK2/FG5Zw/ByZCms+gya76ix0zPbcmDuBqVdUkIbGYXEYzqtmOLMSKf4M1SQ39eIZiWLxYfWOVKxzDh7K66MrsjGtUxc3QqrcyyjoFDxeJDxERBBa1C/VFP43Y0a/XMdkMe+/YVyZXtvM/Oh0k+ZuhrE1x1Jz/yIm2YIeH2PMSnoGxiT/5ALFqc1CU5fLyOaeP4gCttP8Ni3tCdwEo+aj87XkQ80HWXr+FGmOkmmuWgl84MKpa0sbJFpKOM/YvQzhczibQmz2go/cbDFvl2i90lzu8Php7jj0TL2Rqt6w2TrR8OycdMHlBKh8kW93gOqb8+ox5CnLpTBFtlAAWl8J0Ts07JVwSOyZCSBXp9x8ImovYWg6LOTj2/AEdkBfQ5Eep4okuACt1+SObd9eX3MFGUSVwzgumjYsq4R9WfyvTQovtO+AzgPPesddErCafAFUqXklSGYe26vfcC/VueyHs5kBAfuLzwmgjoMpcJghD/gXseiDmLPYH8L10DseH9VE56UcynPSf5/dF/pdrGRQhUhp9ME8wBskCYgXgpXBEyEteIPTRVJcTj1SsmWtGRpWI2WEsbODFRTzoPT3u79406xBAs/3d2QGVjpNXb9Nxmmd2tcsV37g6ng6TgzPijUVVQXQDKr3EjuU/C9POVbsg4iKYabJCXWMKJnsaqcafETFZ0hpFv9HeCL2HYX6QGoXyhMc4zydfCZiLortZySKQbmGX5yZW5Nk6Kbtycw9ewP/kEbqUMawxqawBAdkNx2vdyplYz6JkKr75eRu03Wbg1S5nlFGe8mkcltOcLcQALKG+rn7WqvkUQ18fwy+cXYkQKc624KXXz8bmTbpCMbPJtgG3wLYXHt21fk6sdaf7H0QKeuhTIvJS5CRJPYjJEjNuUrp3knr4U9OfSDAepXqVjqmYMMQs1benLEvJUXbbT8AmfMLwRaZbH63XfdAiO6pNEGkRw4YBLFc0pS86tnbquxpbyvbHK8ox1pU5ObS3cHYASGgkweWXAMwA+qosVnp2SIVooJ43LVe5Tt/WLYgHK/GeOrtPahTNRwW6kZ0Q0ryIIQbrMed6VAV0AD2QakIT9/O909aQZAD8os/FGDf1BdZdLp7Roc3UfXC/gqp7dgp+NCHNtBnEXGmZJajOp/dQ4B1LzPxuiXtb3DOO6BB5FarYAhBJ9+M2GsA2AWvPBk513Zez1gQgXSb/cNM5ccllUTiEcMSGqOUQa5lboNinhXEjQJA6u/i861wi0VOM6PkKoh21PLp8OreQOwMSu3fkXaYtMmpUVapB84n2bndZjGFCc4oPyrOFfShiUY0d5TkPK5/QOfimn4lblc/yyBkio55wQkIayD+lTjL5W88mEEO160uOv89UmuXL2kbfcZwYUqM3ZKBw6mUPVw47EYybFIdyFBghxF9OG7oYpHq7D1WB1PNuPxW4tdQfcumTJg3ZukymwglUesbO0poUvTz5ZiM7+HIAvC43nXy2pUNW6TPuw4ilZe74RlhRLaEIT5TntZ5Y6Z1PNO7ayUo2cEE/4MkyKzu0qO3Q29YAi9bZ/pfF3HV9mRTcFgfWC01/1bpzn2JPvzEgkt3gqS9gtDWLb8JqoYaAHCxZbS3B7CJowcE7DOwM0ukhZYSdqjQimaXPpAncSOBFu/Hs54za42UgCD0qe0AfviPLwcvhRjwhJrKgSWB/gWGZvwEgoxLyjnWdCyRgmfqyv8yj/0bLmII2/zGToj83og/V0LU8Co79m88mOQvmr3q979sidbSaSfZp/G7DScBIGkVfWLPB26ZM9tuo/c75vCXhabX+YkD2OjZ0gC7ngJt2vhV0vpdmsNMnGzh+1gnkgFiaiuVj0WqZQ02X/Oo8wvwVMeOhv6NJVO1e4opwFj+v81Sn2s88/4WdclEsq5zJAesgx9Ojdww4RQsxLTW0FQK2GZ4lroK5ctFPIQd1ouMA7azVZSX6fxih7wqw/ooS4APL69vZtcJ8x4qqjHs0b4f2g0v0v48vSbHrGCidHRy3Jo04cQmMgoYYWAE/v1tLX8J/LpLauTi/31UvwvC0BlHlquzMXl13IlGjeV7A1fc5EJEaO/+CuiEiGr1M7fmJ6NKRSoUkbu7E8h+arAJbZYb4WcvIBVY1vqoa0vEIw5xtMqpLmZKkQo8u1USzYPN1b069YCjmK4iyvCjJwGQccwNEb1P6zoeXsc8bDwMh7HKasrh58gpWX0oCpRwYTZcLT54jIfHVd8Fm0Z3IYyshIuOGcNuBT65qsrlS9IFQlhTXVPyIvQt/OuuTdRo5xMIPJvxIZNgEZ0MkrG8YUlO41fTZWDOWxbMpCIhB1ZFVrSmb5ZSwhZKXux/KBWUU4BWQk3jeA94dEGcj/68gSmgSguY92qRNEi8mXKTwYVFDffsT70RHPPFt83ubek3u/8Rp9Y+W7jeDB2ci7Ur7c2S9cpVGNcZkt6/MY7rAnpFhXhOGkXehL/qbKNhNK/9OGRcI63hRg2ExKhqZVPMXalqynvrMSrUVwrFQxIaRjprhKav/K3zgWg/yfolR+ArZASvDzD1nqYqo/tosSZBksh0elxUHXjM8R9N8UGGZDclhR8vfSYQDxYXLBHH2L0xkY9nCwEE1MS2RAOZJW4DcJSNP2eKD3nxwiboWWodt9oD4HeOBQ3Ub6eIiMOXvlT2bOeDF6vNsCCkVLEqYn/hym0vBKkk00Nlu6JEyBFXJZ7jbQ5Ll5ojtQfIEEHAglopoioCWhvR1WY4vs+DRkNrYDUQ4ZbrkiN6Gg1gliEt3OvsuhwUOlQXlN/pj+Su9fgU+tHiGOCfekYK7nWIDVEEglzE/b3C/pZDaSjnGgRCIw5LAEjbBEEruc4izht0rujXQfEg9EsbAXEJFBlRUlXmeON/n3SAVw9vgi0GXDCCS5T96VRIMLPpChlihOpkxwRArWZAqCdrr12D2tIU3jvlwSgIU0vadUm60Y5NdU3LOoWNlcUw/xlX8ZTKN8749CWaCEOY3DDr5DR4gTRFtpNHuLMCVxTJwZk+vc4C7q/wCQ3xcia6FSEbcJNos5DqJQcOyuCF3NcwzpX5omYQo8IL7LWNoBwK1QdSyDL9EVIc5S1ho43MqQdtaxubc3CqjETzQtr15HfKRyMRLEGqLMPleoUwPBaHMVa1jbbufFha14CYGil+3yUnmzoq9MULWSxioatWG4lszCoI1SdDsY36BGozp4G/7eU7fQmZ1EXfIsWiIAWd8vJo13D4aumdOaC6iaRBP+opghR9EqwPvvv13TEbDf3R3Eb/5awXZUAXLVvBYHibtsV+qg48PhBEsh7VUT4J5MsD0EzGH+O13MXfLZIhaxCbbPMVlQ+oRV5T85rTyohyt/1+79AZVMLAh+R+twX6wFJL7w722ZxIod7TmhcnAOyFRcGLsnU/Gm3efLvYKSKHLycBH2Wa+zq/cABG0cOC2QWy5FWzX7qXggdjxHXmgudN6p78P+Lz/tQPGTzlz3/D8FXFVHObiYFFXcIsF6g87okVtvQT0QP2VJv3I9qq1EJRzZglP78kssnDRN7vPVYxc4DM+breEoBN+/GwFndxE6g1SCMdq0DSR3rHa4MHFwW03SIp9ZrbkH4+gGQXu/mlYYYdGbXjw6DwHt4MKf0kF5XfykEuUxWJZxqs1gyvcDlsS/XKIF21fW3YCzeNjaoeWFwssRoPIIpI0ihEX6i7JemHbNvvPydysNKtcvlp2j13RtnZmd2rYDinYVGZ1PMQoUCsPXCdqT80Yg43E8tqSdMfJY12wGmpJayhua5gTqtJ+3gTzLkW3RgGfxXi63Ziu0SBlWjFxa5D3MnD06g79pcG3vqDiTqU6O/QD7zWTLqPPyRZKco6KxJqHxpPaPNxXgruN4lJJVdF07cuU3EGuYhSFtYkGfgRlv2FGjVtq+yB6t+7h7qUwmHWGS9gYzeIf69XffanwnrS01kWlgQC8hqUHDqC80UBBKXFKjDlknUqTS36appiWivNJgZrGDi/7g0zk7jPUIsVibWO7Qa0pU8ApZUTB7N+96P2xy4j3mF9IbfgG16njOXXDXih/ht5kf0O4y3iNUZcLmoletdn2cCrq+nV+63AjctL8mH3TGvmEXvfc9JLzpUbeGUk8k3eJWrPLvxahgTtsSC/X3yT5X4BmOniONl5ghDMRlCmokLa5PBEIMKAsqUyA6G1IBuF2ILueLsTBZ+PAeRkn7fD1b871QsxlfRliyCEMFjxvgbh1O43ZLw0AxW0PiSdyk/JHykEqrczTbOcWkZZ53rOeTs7bLSkwXKcXPN1+ZIEXcmBrds8v1Tap9ABkC76AHt/XSY2YknQLhrmRrQcE+stJc/OLI1Ve6XreiEH/hEK3fI5qXMbHIzcptrKlmOnKKtDfGJk2GMAljpwiPptan+U/6yk5CDvPXDlzL/3U7L3NFHzQm2yL9FNNlzdU2orRosGTcMN49RnrQr5H7GYXzuFnoGn1diC+H7CWCjmLLDSn13agSjQq/XZ0qGE5Nzesx2Q03U++JqAC/j+URWCkWMcK4XUDhi53m5GHlU7TxERXhDCf4UsIkofifj9bZOWwJVjnPnlBLA9ttIrUdsVmf32flORkvpCpRXI7CqCLwkTqFZS178RXfTlbZcxoLCl7D4sl4TXGh/GOHqbsqfSGl2hWOlcDRKErjcL/mpmBEtzbZl4icwml1X7Ot5VPwvh4d7TN42RlAGgHayJmG7wT/aw064OoyEoIjfffnzxnt4iKk+18C/12hk7YlK/dOmTtDZrzDy84lgGZZW21mN2rn80gR7pFKTvRUPDMF71PZSK76UvuWbsNn3ybiF9jes0hSaibi6xAiZoIg5nvjYMQQIegvFayfCZMnWw0sVrwB5ebAqUs9cQcC8l56hfnpGKH2+po8bvuYgOIgndrKA69m8nAsK1vz1qQvjMYCCYIHa5Gt7Ck0/ns8GdD7wJORHmiSkjc5XsTZb/lTMAsywPLe/tCxaZK45079ly9ribo1KyBYD5q7UFBc8UJbF4rN/zEDiD4HkwV9FIq0HoZRTYyy+wHFnRnMkXoDHTAExklEhDMSJZN86HQ4iQjIGSK2xqeQAGtZPxOVlWy3M3PuReqVGsBcpub2qiTHEvH3ZVRSmSLZ5W8iVOOnZnq93k58aXhJHqAGhnQkKTAW8O7Ybse4Xur4fkC8TSP2mOw1hyg1edrNve16sMtxKziwkTKW0OyD3Gxu+IqdGoMLHWKGUfLujTwPWrs3mIzZ2NUikDQWv1XtpwmpS7qsD7JliIjEGnfCgQ6CfDMxmCk764GfREgLwDBnHYAUjQCTfhJGHBgNkjA6NC2v07dwyO/gdR0zJMmcydAsksoNA9P29kVyJHLFiUwSn9sCoUC5hvmsVsASjGkvwejvOnq0I/Lxg/5W6z+BpGVo9odIWwQN2jNUiFC3Cxagxv8+biFwmjC3cJQyU/+bAu1F5017oDHXg8pESeNVf3sHyBQM6pHEL2+rmS8k2SYuXhGR2Qq8wg3GGDibMtgMR3EZDtc3LgguBtkxxRhWq4BTnX5/D3rDtI0oWpA4tyZsnI+OsbHmYvOhXF27aqS9crpLItsLHtUGIpFxR7JJHLx6vKSWaW9lbpK60FBCCiXkz65Cyv/LLLCxytkn6XMtX7VMfTfK7OzVYl2jE2hjj7qvkj5Ai8aFnWuT9HPqBDnGLqJIZRJ9iKzY5UX/Qwl6TgyyAOf0LdxLtloZ0pVY7BNfFmZs0Ny5y17y8sl/wCoZOX5ZAZqtVFo8bWglpCtQkFOO29qwUZzbSzAHZg8L2C+ZcUDVE2YDrVrXJMp0ZJRycHetOxEg2rgFDx5PkO8LCQs5M+52yb6RyiWPeW6QNr4QF2NLyFjl5djZbZGintDrOw2iNeUKfYQbQap7FmVSSOrAzogpvKjEhb+PtjTrkgN1ss/8x0lHNNHBvhxqARPD6gSZbscYXeGVdwlPW+OBbqoBBBsuTuwoo6UZiXI7EvAD8Gb5tXBoSJMlbnG/RCMOJtMAzCuo8GAlXk17WNzEwY3Lv4FYxeUsZzY7OPUKO5e+ZcjOpX1sd0s7JBw4HPwL0nfYeDY40mKeUDChR6wSyzPPdFijhZAyQ6xcygS4bdbmngT/IzaATd8rDZuxAA3XTKD8ywtQ/poZfyXRw9nAHlvoXFkTeXF46iCawkbctvfNu1P6Xm8TAGR27WiJ7yQEGusvCM4xBie7pKb0gX+pVHAwshp/6NyCkdTK0vKuGcFnVjz+WIN0TUWcrBu+gKL8AxqjLHlKcMFbs5DsPDq1Ryny1kF7tAi+J91Jxkje5HhJ84JQl2m2aLGey8frHx0wk1yUl/e1fmguiXFeFULFNGcWyGfwBEMc0wsTNMkSFQsT42krJH9FmiA4G14mKbgRx0+iJkja+92wgWi19Ihc5RVnaNgzGjhdY7BQZZ4uZIbStLjv1XFPc6ugavNH05yCu3n6Yn4M63Ra2sVgwSoI2R+qSlwOYx137YhIVGjK9rX9Q6lhJCG2crAMofAydlpUNdVmuDQk7ePZP1ut8rZvqav3WzpeGLDDUSu1fO8yv+EmP/C+wHcP+oaVUlqnz7OgeZ/J53d30K4bS7z8oEYqEir5F/UC8ajgxzyJFXc6W8GIWB3ndVwgvUNMN8tuyXCrXdLfznHCF//x+0+zYBHeOGERrCuKEvMIjc8Wy0OduyGeKV8K6KGb/0JbDir1uosb18rAPaxMJbN/wYU2+Wa2gc0MYim37YTWeAkARSrHf6BtpEflMjpqF10KzFIpcvSSU5XlTtTS8nMaOCSYBvirG5IwH5uyrkss/BO3UntE89PHHGUv/lUcA5HEONPlMuNhCCgEJs4GohVMs2K8QBZGY8cAuDsxsjcDzsahUYnR3g3weKzpspqT6wPZq+C5xpOgWfFwineu58k8z69+8ZT4GUPIGA5+8dCUz0Q7ZXr5nNDWLHSaE9nMMSH+pQvUEjjVmvjPK12f8Y5zKkR6X4JqFegTLu1r9+EvOehJ5oZuJAYB1AitGM2qTqDEjHlEsc1CIktSD4Uo3gkCpoVxBlWYO4CGT73YzvxfLblCNDwMp1+dg8pRaHakPrhYNohZz3v9F75kB+DCfqItCpn4dyiiXvRRqyErR0+sId3mxlySLVlsRwqEATU4p7P47RwilT/UQGIuIFbyDtzrG94ueEJRttuEpts/LZaA7kLyP2+7OxSVTUsFFY7iDLXoJxeup/wxbs0vkTXkOGa5Ert4rKI+2qbN+mSveVoBU4z2zja9d/sqQoJSviplywQn66XFOZ9NttoavFbhF7wnH3Ym1qXED2LUIPkbVTKOmDaByKu5MeBPZBD86/m+AIoXfOSqfx2/TCoq4zfo/ir3KRpkgh8o9QTKuhwN1i4KwDzSVQhrbebavdtRbcdM6fVH13LDv0Too04MBVd0j6fK1+IPnkoiRD9nYeLrBEy9UCUg+J37B3FUsOXtaZQHBPNWuicAM8xlMfOyACCamXFy1ZrblzcKfuXO19eYALKTrce7bAOndAJeZ78Et4vsH1QVU0bY/AJAA4rl8VSJlIezCXSVD9PchzTaIWVf+7wn6B8TdDn/SzIDsDLBxmqLrUGEytqZwqgVKxPn3irfFjRFVp3af1KTNofJNP6jcw9ibhXzjuXXg/grTO8i5o4cP4kvn+S9Xhxd1TpYTxz52YNB6eE0kzpAWYwLE7QMH8obMc/5VQXwItay6UTkl9xVIzuQW4d7vTDDI87f230BBLCYt1NgdEG7UUMXv6EA5zd+g/ojpVmjrpRffo7UOWSY0hzgl+L4kv/GuymeqF/ZdPBvrVZYfDmcPrUuyqoyakJNGm8p+17/mQSmX9edsu+4YhfBoXj6Kwp8nVsc+T5qSpoCh/V2VA57PprkuzJqNzzAvTJ8hPSshYzKkYoHCPLwj12shKGIAwZW0pknDKDQ2pKRQPKObz4lPrHMy4rVhyLaDVl/2LEu11RU+zSFuxtZJKvHfwI1wxOIg2tBv2lqYRkG4ooDBlJwHIYV/Wizyqe/F+mPoCLm4maxI7JVCBVoxd7pxLIk3pmP31+zc9DqE8GAkVgv5rw5muOMHtGB9rqv/6TEdBIJXKczWmGt8bffvTpH7nitn6+qmKmWc507SdZQ1DoMpFN4nZi5CpwsGebVdP3yzMCCKiI7hmsJdaSGgWmOGTO+LnyvbfjaRF+6M7jytuweQ9JU4H5dUXSdwxwIWvUBq81zYnaJ1tHzQZq/brccFVXFcSCJPDBtra8tkaYfktmW8FTMHizTrV7u/eP9UhZx+T/7X2RBD8HMH+Vz4ClUJHjhzw0Ukb52udbvmLOTqLGFv8Rmv5tza2qgmW2xK14BTpfixdN24Rbo5Dz0CM6hn8JN29cCcSMMo7pu9RRhIBBxvVqVSzU2b1kdlWqr7ml8zVsS2Jw+ywEh27y6VkCN/gxAS0YDJEd9KK0d6bT22jzd5u4Kx0O4q2tUGfuhetbCs30f08RU/AVnzeHYhq4C8dfYLehp8e4yXA8asevfn5BNIO/1M5tKlusBX25mRS38GL0j/JPaKV9qVH01/L5NA6VgJunH7iocGXy+irMQR+tXiggKOdp9ZvrQXLEpEa7MXcuWnRs0RH1qHxTRmIBu8FU1EDtJgzYAJokFBL3fWXq6jUs7GgcW3PFwKdxW7AVwZO7otXm07VX1vjTYDOFiD6qCnsOMU3/iPSg9SvtlC79zp9t0qzwyUA8EId36vjvEWYGvzZFCVNsUjXQfcPdiB49Xb4NxuVPb5X8Sy0oJW4YuXPYzCrTIsoRFY3yjC7tSDqWwDKumnLdthzEtDfwZYTVQVx4k8n2RHj4psrTXSw9gkxNIMIuBgGbLRNIS/z7VRBg5gUkSdvxR0tWc1G8N2roNANfKZXqmRkAxmtFseS00Hi+jB9pQn0vixKSWGGvAz9dolWZf9UHblpbMPcwtSPijc/p3djxCm0Vju+mE327FY7UjBviw9z1Jj4OqEhxRs+j0xbVHqRmy40OMVaA0G5+2tOTNEMMrvsKTaUpMxtYob5BxHW0GRLDoYPP7tTtT9OUDF2sE7AUyoR/GNKhYi4oMsrDHTtAyKKPHxMN0JB9HLQ9lTSTFzfLFpd4a9y0zXI8mPrDo9GwlRvvhrXb1a/7Cc1VC0tOGfQy5nFbNdKbTECNhN6EVpDqPt4CBq4OL6vXJ0AN+VXB6/xV7cQVyvNd0QrV04HLZiMZeg4wXI/V5mVPr+YsK+su6hMTvB7bGrfZkVeWO0QVtF3y5/MxU2tk58Fm5utN9S/MZmjfwUW10kYTxIKdLVs4EqBtR5pVbQEhN+Q44XU0HqdYl5jPn2u7iq2ZwQaeDTN5dbsXC4uWGiU3DL6au+t+tn8kAq2/AXyhJ53s12/MGdX2oEUHjKxOHCpwEJByoPi2Y/L4R4qz89noE5O+dQonnSfj6qCjlHwacPLV5YeuMdFmRSBEF1SLvqpYQ8cqrx1PgEj7CLddE39GipKBYCNYPJgJVrqCFBIqG/EOWMG96fl7eS7SN2VQ+CQ/Ux4qKLa/0Hucg0T7FBdRmDvm7xyTimtD9jWcAS0UCE5EZTQaDnxZLNAUxiG2d9z1wL8icnnvgjXh2CHVh9T06+rtwvbpdZ8pLH9FvZWjJ6BhUsgx5oUshrCaHecr/0sJxIM9F3uWkP+w7uaxJVL0SCzL8R5o5GTO1YOhFQU2XwM0KBmR4HZR8rWK0k9czwD8XJuyTE0fVMKZc9VwkvRHvqDSOQditoA5M4ot7mAUrUbkpE9MrlWGrMX3qXiN3HQbSZnwey0aF09CAj2D1ot+06Ovv7OMbcTDtph2ptd9MfOpFadeH6MS/7NT+un9yrSI6BbSK2P5JCJolt+WJJ9g+jlFCjoKIO2Rl/TXUTPLvym/3OfAxU9a77l0su4C21ZZfTVG8vHrUeIIRkCY4k9XYnXfQZVcUFh20uBPk6A4XM0Ndm2jC1GYHf/nbGfjq1uMyNnW6E1XGJo9PlifuULZ9zufzBWuHH8PB0cetQQ+95BB75Vw++4zzfldi5U65s7Q4rcF2OTx2JkGoGN9JfAupe8/zfIoVL8oytKyx2nWOyjHsX6UMVIaFh0dC19NW6KDDkFjjAXmZf5q/G4hRkRDkVqxfsJAViMz0rk+3rRjyEPNH+FhcoB/6rc2mBewJHF4fhqo2OLZODcNewmi50aKmSOzmKc8Qq6BY59qc870d3vhEuPhkkh6OTLTvXp6YQbnxPwHBCBPUylASfrQuf3hsBQjyQTmehAL0f+O1gETbnuA77Z2HuloJQEQ0/85EJBdlZmefLObQEYB9qogZPru9QnpjJWEWZR69VzEvdJ/nB2k0LRQIreAUy5mLB90byzPxWByVqsINf00PHnXzDOhWBg+S+Hxe8RcrYiE6sHYrLbOHTy4r7bLQ2kbRTIkz1tgRRyCp6Lv94IJrL1oMn5j/0mUwP4RWXUY86vdpKd8NJOAjh3yhec5y8KnqfVb1Bd3ZgIt8WE0y4wXELx5kAdm76OXold/FX3DX3oxlxsOrE4DOFdgeWYD3grsRq1W97J5deQF2g7Kvuy7a9Y9AaklxmW3Lp5kbRdRJYclPQVlUZ80l7w51DV6Ae/HaPF/hrKj0EhcW0jzfLGAfCgb1dSLrQ9Nvxz4hPde9F9Hc7Zyj+FUvxtB18Rh1qgAReKGbBtTtrnywiJ94ApCFZsUvb4lkoqW+en9hZbpOguSwTxzfq/LlceNM8MvJM8C5aHAZrMwBaoW8dN+k5wvnX3lk1kPaFHXuB7y9uyZRcv0D0nvabIKS2AAYJkfP/mJAyxCfE6nOAqf7lDg5iIsQ9bzjk8yi4RTJqIlM9jrlH0tBl1jJ9LXb808+etHFAInZjfXJJjEnE3VQIFm0beXA1zlr7VZx15clbMfcFsxv2CkYNqCbm5QOJ7o/qHWXzWpCadDf9TBsro7u5m/MGmZIQI1eyspeNzIyJr9KY5emwwCF+0txUDh4wPWefkNIc+PPKiZoZFR7BvFtnmzt0V8lnKItK9VcyOj2t6BAKY4RzOnTD88r+pfZuEoOS39OOZbuR8Q4Mf/MrN9SHbIfqiy6hwEA2ecAyxlgPQHDiEA3JykECukEppOwHJMnFrsY8Hyxd9WrKdkf1eWqZz1/igGqM6sR5CMqQF189Nlcpr2vv7707aIMHRgwTl15o1Etm3P0LsqJJQYyuZ+2Hj8S5yIXhBs5oMNTc7f6ugt6M6B/5eeU2msQxpLu+4F+IohfLnrcMN4/hM3kLlbZPJq6ZSGtIVxmD4X5HRzNuCmH+kSBA9URv6UM5HtfTMmGBMKvug/bjcrKvNkvnz5agTIoYFuWm7Q8aZlQGIRFDrfxtqUbzH//Cac5mgjHqSEwc3GkiXDRpT92A0LzI2lgiN1jpZm/9Tgx2I4a0PxDSe4PIqxvJVmxxTn9dxWfIPGK81gwULIwdJ7punyievLPBds3xtBGsHEjRiscfmVI5fkNCIEeEXmO7aebbB1zB7dSxw308hUEzt4g/FSF9hzmTAth+Dazymg1Bt7qPIBlqcnPefY5JbQ1qjaPEhSpJUaPB5IIJl8GdB7/GxGTDIveCXE3dkhyXfISmLp4HPtvqGXymL0w/J5WDBEiUt5E1Tn55f7XH/i6LpwK/KTIsI89FUJ27wjvJZSkTCpBgmeTGe1EbLTzRph0iyiwU9kvDszm0E76a4Kg+VV9Vl7shLSjxtVjt5I/BPO4Y+RebdcZXvgpqmisL4NYOKMNy82nL45WbKkG4QlEf4UVpMz9GsA6pcUekIlTqOSVVnFSxiGJcN6XYei/HC1DMsyskNmSZt3JMasX8V+TfjPOVlp+pyro/vCNLH1W3w6SxxLsmRGvRkc3MdT6HtyLNlxC8GQkY/LXwrP7VqGHPvrjF1XAER3wvQtlI/xYqmlT2qRnIuHMxCcvtjVgcPNc1iJSzYr0jIjD5ZPJ1pXBYfnLyjUvP1D7d7brO/87+bhDClkKcOiwZlAN4uDWHXjKCd+iBtLPLqj5awTY3jMmhQajvXbCevatwaCsfZsBpDnqmPhDGh4LOP7pytfQl0dTGCVpaCzxE2lJVj+AQaA2VgcZ9LjKHW/pgM3TLAoE22zB9CjPRE/2nbRloq6qSUSyb0QWC0Z9oKhTJpQXkX+6q2reJZTSJFnBBcryzfxlWJZIWkYN1e3r9xIdC3yQdyJxugbyrNsNNNq/lStwDR2HKLH1mXy9DrwAII9AbikhIV74880drIN67QKHXuR9S9aox/GrM9D0nGH3nEUJJy2rhiO/D+TS7h0aIcw52yl2V6mangTS4PEX8dOzYE9eQk9rCVRkPwbtT40sWfueat43I+v443p235Ue1eey7sac2jMWo82Wr5h0oZA2eYcCVFwrjk5Ms8kmf12bsVS/PR5t4fYYiW+6MUtUZBkHraosEYyPUPXbibyRhL/tAUXaip94kZZdfBaMptlIVKKiilxgYTQCx4MHkjiBdWAsheSKCfCNQMox1VC58q2AWyawA17NoSl9mzh5pmn3inPmuDJYcGhQE8F1ipYH8a9qo52/NkK3k0bdNsicnGE2YBMsY8NR4FuUmQ2k2xfc8Ml71sSYyu5q8SgOwGCBJZKtOr/rwSwTCt+tw803do0pmU2jcrrq7xVnzHCfVWkEf1cUh7gVXZS5Jip7JhF4jNgvxgyg3Hyz1BsJpatNhVnTzGOqPGIRukanUnSHpvXHRzJUartT1MH2XAmY9c0RjHZPmdVoexc1j4TlJTju2z/l9jWtaZYNFxTVDIcSTgAtjjFx5+E8RhXuepopdto5Wkinx47v0H8ha4cJESivkthFSAR00vfIEVdGp0qoGrLF7pVDXqMTVnlqcz5EJzzgxIn3kBN3/I+sSfe9FomVFnl51yDi1pwCN3QNiDPAbHAalMx1MJ9BkekdotaK2EUb5Xbidi+xIsu2mDnLOtffxm9pzlKen8pV7Geb74D0KRYif8CyOYUKqcsKSeb+JpwmuCP7INg7ZP9fiDklAlo3pOm3b/etcO68QiE59mwP0PanOCNvds590KmO4RnUsVihjn/ZsntprM1Ax5ZrIZLEfHnrSzCiVrvnfvVD9a8CrzREmtm1u4ukAswG0SHCpcrEpI60hwdXWhoJgPhi0BiY89VFswRaLbxgtK4irCJoqXEyp9hD0477mh7J1smX743fHHEglhzCT34OvveMcly+pG0T6HWBvq8rSTzcfsLcAhhYSGOqFbgn8EAtRjxLfxiukfa184o/mdU7A5PyUDQ3IuEFRzuBrIGm753mgZtcW4iEIfhUt0ouOdrjWznmcAdMoOyuNig87II1san7VvJ9H0hH2afjj0hDxKrHZfqi3Tk/FhC8rDIROIUytmVMOY2iCh7MHqV/+4Mb3u3EU90gasHYW3B7925grZT/ZhMe9Sc3TQOWt5am7/cOR9b6HqveDS1JSF0AZ2auB/f1ml+WyZ5OfFCvfw8ZpCk7ApfNOB/sZQISETkkghccA2w6YwXp8ZIaHYRpUZRyb66eZJYbZ9wFQgj3h8is7/2O90Q8Y2LdmeeuJ9JYWdWl1m/eB/pHt9wsH+NE7EGViXJn/U133cShIaJ42/7eo0BMNW+lRBsVYj0Hb1hldjSM+woGpCwJFXf9+kMfRRWqlg23lIyCbzvMKZcV7B8+34MCMqZv344UqNcksqVVYTD+hu7S72pnyGTvR4C2uNM8M1u+uZWnF2vJz7uST8Yt420SfncAVhoMr/Vk9Ypm7kEIEAcQO3IsoJLL2RXRIBPHLzIAjV2N+MjeVUXeGKMtKwghf/tRjgN0SoCMIda92WM6MJM3VPs016RDUj+Stsox9R29DSDMaTvtA+b/4Xm5tLE8mQVieRYd3HmbEr8tKOAnS1xTNmrJnGAP38zsJFSR9VEM92bhs3bkb3H7F8buuCOiHUx21ZhPizlrpJOmVEBj5thV1TMftu4kX5WgBq8EJeTQ5G4gyn6v2dBz7LD/OcpH0zQti4SnnTfIfxKVD2PBcvhUW/2DTIz8u3QjyrtPRBr8rTAuj7nt/i1xQ1DrKGxbGQeu8HAimNfMkZmjssxcTJJ6P7C3UEcRcSFhfVejjnVpc4giinVs9KhdhSIT8seO5X1toLIiGhe+SV6fIbKNISAHwg9rLtAkobII7hN4V7W28I2j2+0GeEoIL/0M+1m+iHhlAJbAkG9DPPVGJy3TZe5yy9Lu1LbkrPFDhXEmN9+YNgsRP09CLwK+fqej3Gsj5xcQQkJZtgDT8Uvn3uRScQO8+wK+0adOStG/qaW3ShMihqN5KAtxwV0kju1MZ73zesmpAaOpl8Z79CndqrwjFP5SnNtPCFYQbtGeReYH5fC3O2T86OedCwFd7Bnxk/nPPGix3wtYg/c34B7W9R6q66Hz/KpUxlwiaXGKVdWIJPa96csyuN3xTz1UUuEQJ6lU6vZw9w5B2+HqgPR+jOb9V4/kbIiGxO6Dda4bFXnNAHiPoZdP5NyUTPLTn0+UX89cP5lFZCmx0AXl5kqab4TjI+wto8Y8h4HoCKrNFmluwEAXBJmjWoGF3VX36tuD0LJucv76vON1gLzHYQC7j2OVsnrcauS0sNrarXgvvGSJgThT85BVIJbNqAlqFqXJbYBKDhRUYpwVjhak1RVPzX+IZmA4v+hCHh/p6awVnI/MDxghGCrWcPtO4C8YkwLIwPFsqOnMZimI5A69NGmOF/qhZ/Fen30sT8sx6CG2KxIaf0qt9PEBt3+psTUPf5Sl3359z2gqtiA9enHvYEbMcMDELeAI4FtLJ14wYdOwh/katAcn11HBjmazencD3IoMw8THB7aAFw7j6rxMOAmPa25FuEbT8s7GZqxLZAtem26qEUHjXIy/pS0Zm9ttnJQbyb6xXD4FkDQyVJEOLej8qWmQjENqpBR++vr2OxPJ/+BxDDUzpSDwm6HgDzSac1BnSCiFQit2bfRcB0fXtjjheBg8Qay1+CzkSwOmRvRGHYAqxFfivGBWs9ZlXEA7KKDjnBRIO4su4kZqCw2l1UWtZNwY0s7rUs9yJHHGUwvFh86/+al+U5OLVqdnUN3oZ1hA2fiJCTAvUmwGJWp1cq1WRtWvVZyX9Z+PPYa/7rQN/tVs9tTIjra9Y8UVH3aRc0OW2Xg8W0M7bFJeLlH4pQUMqPAE17H1nLtmO5HFakvoVdguWo9ckEeTotpDNghFlHZrn+IlYEWLtViea5EtmldAeMF+xPbuoZLeTvTcorYmFPw8FoygNIDg8AxFz2Wsa9/eSfLjejHh0+B6Mt7tiwBSeKkDe0gBc9X/v6pVLF85BvHjOyOsOgnKQVFs9nw3JsqAMWkMM7BSpXeLqs/gnIfegMjSPKzbQwkmjM9IWCDvqCSB19MSxA0fC3QjXhA1kcvgvqVCvvXRtM8hdDHeUzPQIvFLMsbF33boma03llPvyPL2DG+mZ6kRTaQsqGVAd4IleMKQh9PqN5ITFG/EYxeRis/TtwpI1oZ0x11wDbYaxhkvaXFL0PTD9MbPQ+3tCWYCyMukJq3yaT254NFhQB62yPS4U1jJ8c5Ijhatg+quFWEZMrjajvJP9A26Ew8q1LmqlBZuKREAIaikpmubqvtTLLQz/oLtRBEzNpcCOo4mkPrO9MqZhidx9vqOKusv1A5qTSYxAPXYf47aDXpJDEgASBxlqx4t1AJnrWRMt1CG/4FMGRqeKS2IQ4ki2loi1AlZQuVpK8QOtpm6CSCJlJNprG/aaVstu/jAemsJnnyzGteX+loJ9zjv5n/WJMQBerg3yaFqbMUowSJpEr6BG/D7bTEWBh3NzulLA0p/EjBg7i2k3xpWEm1up/rLGiU7vClw7A2t/bc3/SptzifAEY7/SPbvH7LUJdkkHNQaNKzaAb1ie5tWhPLQHjgwmrJXhJo1zkOIid0oVVCVa08b/bLIPr1XlTEObONPzo95DzQKHCz02YMuaGqaEFYouD8GiKV/VMNl4SNE54aiKjiAPxQVsOhpq9QjPYyzGw7ITjX0MZrjzlQG+bDnVLo6XcpNSgjQdSevP+6TJ62tzl55Cgkrnv75rU1jh/YjvgUTKmajd+5ZQvz933BQ3kNzch3XMXBDitx74m73SBMiw0BSidWyONRWzM14zERNcD9R8Nvg4y0ojwytv+Afv8KoPfeqO3feSBVh9sn1jFB9PuoxA8b+RATqkxS30OhMTlHQ6e6Is9i/PgnBFeVMnMVqrcN48nxlUEUYqQc8jIs5VNp/lbCKajILwnW8FIhHS5yx+TxXz5Qv9fO4pH+Kg9e3L6vLWI8Dcv5ycBgKSjDvjcmgjJi9U8lv/f2bN7iUdN/AvDtOkHs3N5gag//AelRHXAMRHK1U316hyn4EEBTLE4MT3hFYu2M7FbbTwRtKihELzFUlud+AHYmBoSt8hSgkt3+/puOtM5IZyABDvVveczEEcHi/sblSO9TVTMtUcx8CGlix17SYW8BwyNgx40RZ3iNdnOoOiUB9vOUCwkbCTxLbjNYufInwIvyGHeeRBqjJbxZgp5rrzQaTzUG5k0M+ptizt5CU4w9Lyzbad8NdfRHXXOJoQW3dSeK3DP8/huFu7QZ7XttfCxWRz8xyVUMMV/E4Gz8Znk2fdeFeSx2koIbfGLXXkKK5tvttNRM+9kz0codwS1LX2thegOStiZG0jkZsCj1kIWLgFSwrQiw0a0uUblFhUSIZiNrDiv4wwGZm4Ahf1yeHhXqbt1HEWr4eDAbqDJ195/0GQeEWqR78PkJRFckrRYOKr08S57S9oKQCNvxmcZLNaZjtXzV3+qJ+knXtISGiXbDEp4NhCbOCcipK4PQsU9vxXmfi750OuxsZl8jreH4tg0T5dAD0ta1qw2Dv9xXVxMYPefmeJP5/LMinTTtifGR4HtcDg547MgAGavIvjLpL9LIcB8HPtUb4tZp5wmwqJOvrH9mrVDNB40qep2XmKk1efBe9omo/8PhOdnUbGya2B3IUgdtevj6i5qCjlND6JUpISHyMb9NXmnuhBmeKD4B3Yq0FW1G0VRN3yH7W1sOA5gx3wqIZpnNi+yiq5bu+v1QGIJp2ouo9Gd6bn2WD+1E1RmXYGV7uR1pFwTBqG4u9p8ePUP1xr1j6TFdk9clLDnBUk5yFTYIl/frFrj0dVKPIzomAsiA39tmlLxz8TZ1TlubUtkmxssC4elyJ0gZVPUgHziAvEF/1N+zZ3kUJJTzazqLK06t2YidYzbbO8OWkGboc6/uPNSfdFrIQlAdXUFq4Xmt/bMbWTozBckVBYlOiSvYjENOpCOLf7RRxKU1tAKUSDvejwFTiy3ozrBh1YZdaC8NhgEdMnKEhhegNInbZSzkyUvNxbl4miJo7zh4iJ2rEu467j9jumemesKNTcEV3tFfM61XQcMitTGR9+2u3UJeoAXLxmZwdERU14gLE4ihFM7WZZlBp0vgmUtPIGzcZl5h24kYR3nGL4lVmNgazKWakvdNH1+9vhhWIrNqxLS/WduyVFoqfP4cg8KoHSuRAUxLtOq3nVCPfK1NDIhBotQsJyAWfpN+UkQjiuYg78+8zMryktQvpuReOlK4hZ37KXm5TA4RHiuWHoR19FPm8zZu0hOsaFqm2VxLNB2bIcKohlH4TZQ812y3hlT9JgSloK94ZXJfSduk9VxNliWoTLN4CPKxLR9coIdjEHKm5jOYmjWyabyhFsKt617j0cSCF4yCTebwhcGMaVH+nlK+pXxx3I/k3GGkQdh6N1Pq1Rbhty5DCl4EWXKJLniPYWUi2LzOSzN5Skx72UugG2d+URWxlOSN7oP8oAJu4x1odDT7MWGhCJ4gm0l6T2mqvurRpdDqToGWOKkZQMnpxI0Map45WpyEmSKUTCwymKDQ/rBS4CJw+XB2cFmTr2vZUC+DT6EmiNgk4DV8WpKYdE6eL4ar1Gxj61UlCuq6GFgdsBHEgnJPTn9+pTLZzLfugh+W/S7KTJtCQlL9B/uMkHALoRILzVcOXkIuEysWDLPyr4aJFuIo/7/vfZyiMyxA6YnXwWAfupcqAEh1n9AKG8cXZ58x6GpX8QSDyuwNKCOihWPiMwG8M6Asf7GCfLolx9E7iMMH7aw+qknHxjG7dEu/gpUEHxMn8sAs0LAcVTEFLgh2dRcUelJLoEtci64kpRC9uxpBdnwCP6aNGU5jrBvwgKsqTQ4PiVeeZ8Jk6pWYMaxV23BTzpvHGzUVkoumhotXYYQdJm6fYRTcYE8HZ3ZVPIpXfjPMxBFMmeUjj2rLgiPwb++bZNjrGIphTjbhVO+5tFscwjecxlZvuMyPTabd6zkHwMKpEUMFrb31gWcXUn22vFva/H1frFyTpPoQhtI6N8ASRZpTf6Q8JmVfNDWrtUY3dLtqKxt6TjX2jAhoFi+Y1N4fMciA0OYp4zi2poWRrun4isJmyd6J/02+jBbAGqOAp+YhFnrHh/qQQ6DmqZfzJuexQ41rkvWfq6GMIm/LV2M5/A409Lu7Zk8ANimVCm7AOmU5aCf6PCX/nW/383QusMCTfOZCCyTZfJM96CB8ARznMDJ40VWnoLV/jdFIcr6q45EG5Nssbo2mVx7RhNISWDI7MJRtFbQMMm4hqxb3+MnFjMNUum2rXMRPZM2X/a9vGnBoC+S07BtbBQl/bcQtozGsPsW5YmgtDVD7wYykKc6uDGU+Qu9o/+apLfJBYLKXZS2e1Gt94kwYXsVwH4kSmbZu/cb6oOFw/F9FhaLAXNHgdT0stE7zdx+lVrh5tm6QMpI3mrR7dDepVHAq82I2r/MfYksR8WSryDPQXypcxMHdp/YRekLuz1jgebJ9S1Tj46MCY1mlMO2kKsrKMGeAx8pO7e/RZW6hD43VMSOeCI5USShcCbcZacS9y+ECZApHdoaGhwtL1wK74FLuDW4qDXu6wPiXG7qbBm7h3LPdAUYvUA+nZgtLFYAOzQsAE2S17PDwsFMxTuuz2gIN/7zIUWrxmwJFEm/8WRn/zAtjUeEMpmsmR66B6Z6slB9t/9/amvqFZiCRp5Q8znMi84HiaQsFZNmpIfiey4NmBE7wjY+oY/tw8tPh5VfvHtfuDsvK28JvWPotEnEx0k7Gx+LKwYd0dB+gCN0MElZqGB5ghOawW7Js0I7bcqqdxKnrwBp9x2J0FWupztPdAjssgNhtjlioLbXdDX3j4KbpziO/P018KmjpoFSkn8Q+EeZqnTO+d5HgLfSExClkpQBQadmuQp4kCgSZkPleZm/6TrwMKoHufs2v00FGsW9DuXBDmW6gxc0zorQN9GobTxe7skFU/lbjy9NdQSz4IdNdFmpdRkVBqKC1uy7TNeZaq6OKBXVViEt6mZB1osKQYjfO4eHpmj6X3xIrBfBaAgNA+xT4sLVlgQBNNxjnYawdXv6GhvEPzrJl1ZMEIYithOp3hVcV30ztmCq00CefNkO9CNMX24IlwEdVOjoPC+TtH6/+quZ7r8eJkGtU9s4m5bttel6ri0ZSNYLT3ag6efhIcufzE8677lQd5KmLJp49HjMAstEkAG4OeQ3K1k7IDkC6uQobyEqGBlTBPPIMDIKqiHpuSgtJ+jgVmJPInV6WEFxP1ZEsAqEqQnbyd1l1f6VZZ4lJbRtSqnw02ENzVtRERk4CL8BgvnMsYBFDh5XlkOSeDau0DWizU7nlmCu6keTAHWcKZKoQ0l5hN8w+JlCqofmuDawbgtEdqUZlbmETGRKLUotpw9XJKuNBZL5Ue7S38fEzuAK0U6+DQZ342vZFR8Ucw3ui2L8Ni+hVGjyhaBxu5/hpHVBD7rEEa2X/O0SGdLUGJk3g4m8Wy4iBh1sTuRNJE7IcsE+UXKeGis8hZAT+2LomNgzYVJlFvhnaAT0YnApedQGusJCo7GoOp8oS17doIM2i2ZPuAn0FglONIQDGkwPDm12Fq23Kp7EI5plYwNfeOhad5KUSNV3yN5ElvtqvS2i5SkMXAsIU9/yy19BidrwqOpJQ3DuwR6DwqnarOfUzfQOLrCmtNZUSNGZYCruPPWMdUHji1kJcIpoNbQdmAAmv3lm8+Govb+TzNZvPK+ZFeg9sGcUzP96gGIU5xS/PkIDzNdDzNljIzV9bhsYi/JB+K+hU00yAs/ZTTkCAGKwhi6EOOySYej6cnWQlhxQJ//Gnoj2lbWmmSpFWMjL+un//xwE8D3olFM9PSyGPMwMDKfBKKdbeARRwjX7UDHD3jAEG5SbOHWlqXFVPWKMMK4OPg5nO5RIP+xENUviKTIJjzL1M6WVNo77KEKaURpccq07RYPgjut3TfyDTwdFAfnQpE5rnGgLxCqgqKww4GG1ThLp3WqjGCY6LyDH3eL5bLSi6PkW7hi55LfFkJaZSzbdkhCQxvZlHnQSey3F7uC4TBS8iiwRCEgoUFPUoMB8VNU0Bl0YlJg9HLYgvdxApGdzZYyO8+VHkuXp235OPHhlsf5nsMxNO9ibgNd7EJjlhB/xQdiJl+AoUGPB97P2NCpbPcuJendzDQKPBGxeZo0HWltk98Nj1SAFdzEd0zurph1fSmpOBMEXLQm13yu5AAMmX5VLtPtstlJSAC8tJIoGGqE2RUnJdrE5oMY56th3r2r8+JRlDuooHcmstNgNfNKudvEk3fIb3QCDO/xXYZ7fTJA8fu3/5EMOK6NpQs+Gyksv9CJpFarBaDfjlNmcXwki1BWV7AxXxbEvFuvHLwGUB//8HlzDUlVesqEbBejPPlr7NLoYaDP2eX0SB2jn7mnu2c4eZhIaKWq+vqpMAyWYZroKa08kM/Tw8oEUabEkIDcCQeS13CJHFkwWnYiK4y9qejRIjhbzhjprIKufJ5MQaStI9oHkjT7/FhSnRsbYlxM1AQDFBXsFGv+IW0nuEgXEds+jw5G70+gEeyiWYlVyB3jkDkW/2F2YVPhQ0TwPkD3sNexiPVku0cIXc9WXA4X+JMW7ZvbJuIBSZ2jyg7FuGtBmaOIoZIeY3Xxj25sbGHSAEbtffDGpPuxyxE/1jcSl5XKJ7FXTuJARY/wDYrtBbXQ9rBwPOW347bm1jTXyLc3pqoP8HwPkNE18F8yfwQXXuIxh+ex8/Gbe7+golfwjm9OR6vEd9v+LQyYNnx0/1IyYvomewLMXqFD7OYGsIxG7Oc3lnsGUO2+f+IlrIrEAWFvHDfEHVVhcQD0Ielqx/3d46qimhTPj81mnWnWVoUwuU19hsClTWxTBt4D+pu00+VnZKT+xMy6RVB78GIbgu2tEstGL8CmG7J/qZ2oyTz403Gvu3wVo3m8gcgXsfCGWI7iQvBI+chcOWTtPBMxECOMWbCYJlQOF8mPC/m2fgKSAmg3fZXOA6lQEYoJ8PeqhjdIDmxkprWK6Wt141X7M3cZ46lOeyhWZ+AstYOwjjWFdsPfbzDzWHh+hfFALHXEXVsKRsEltVJP776SkQStet9/InA460bNIBN9jOWmg/44gQrjBKUJXrg0BnoER8ChsCeXpFTgHiJ+vz1+TQy2r4/mCZBD9l86C86PhWU9uankRGM0DGQvKwRz0093qpa0DZ5Xqp1qzA158ETDNNa0cd31ItWDA5mFXdnKjm2g1O07CxpFP8HUJy32LM6S6+LZWOL/A+qVcrmwTuChPl4Xl0VELDBiE9DE7v/pJyXq2ZDVGIVpWLmywUzdOc6WWVH5R/eaQqlGvfW9vHYm5Y25NPKziI1k9uPv066NLjxZJzDx8/1grvr2/GpQbUM7IMrhBhDpw5zhU9Jm32IaUaf9uAFaGLSpnyQo97ptCkhEFMpJrkXZEyoQkGr72++5fyfSyab5c7vIL3wg39l6wyb9rqyxeL88fr/3LLMQXKU1MmRCa9jM0Yffi8xQdartnlpoh3RkfFz9d56eDmOYjkgbVgdxk2EiqSjL5i/45H0SbypPeUGP5T6SC+c0eb2OITYJt3NbCAZ8XSOOJ8NZXZjjd4y9feGZq1fVWuNTJ4JLGRQ2YR7BUW5OfIO+952wEdojRCVH087vxKKPjgYCEd0toCi7KoXX2IrXg97COMIFlNIOp2MN7ZpA6FSDMucnM2quUDqixqSPY07/yAhS6kdMjZUgukutN8/AOeJljGz5vf5Pm46z+wESGAp1ACeQhzTTvM8NDVqBLeEHHG9oAIsD57+EjAikb4SFHmDdmbTedcN9V6tXgjmUZGqfkH6zmZ7ndIDPnTtQ4w17XqOg2OAjg7D/3vkQeQeuX4wGetL3oAfrzZ5i9UytcHFOrRodQ+stjXkps8lXzgioK0SB52kf0C8knXYqMb0xx0MBusmWAEGwXJyYHjmGcSc8lUe+jvHJPaQU5VPQMCsLoWDrrlYxhcuSDQYUuXS8OSeh3FUohHbUXxX38DaAP91qdKsNiUt/IFixIKFWU30aXIK1bGDx7pu7Oi7IzWsmWOcscW9VyieihTJohAzUf5EPeSM968oVm8C09l3u8JcMFiDfHWJr8eMqSraCNBw5agUvx53yuH+mFJW84aGz4lgYVIKUljc110iwGNMPCDTv242/ohmqeM1ml0sjF9ZvEhkcAgH/1T8NA0GlzkRUvIjMV3UJdu7geMbs+xQYxXIp+yQ0mAmVJ5CnEq2DVYyf3/b7KCKafbPi377e34nBNhU1EFCEiaYZjR4aaFoTV3zMy3/+es96V8eYA11CQ2eMAdsCcFkRloNbGJREfLFNwI1T0oeh+t12ddxJDKCXJuv0ylEvhdhyfIWDNtsDo9H6SMJKZcue1JFvclbajEHq+jDI5Mu7a+sQ+SEjZDCntWri27spSmQIA5oZ3ADVpMyPpMKr+5kLjft6x5JatrVklprDf213/HYzneLcOYK0O/H3c4qU7H0ZTX9fFonz1pUzpadvMIJ97mm5BkkZPQWvYeHVrWqDDnbvqFAyQTYULvuEgqLiPRCfVUmgU+ytESNZNefkJzn6ggoQvtPTVowFxS9Rb4n1iscLjgIGMjuOggn8q3/yiMe7D+Kp1ubFS6VDmw1JHlT6oXtPBBZaxKhfz4LEcwQviFCzrWM3j8x71iceFGxjZm2jo7sMZcPZJCDS0PepZPvLpe5H+ITyEpVVuboZcH/Rbj4EnTpswlAqCcHbSLn9oB+syWxqs8yj4hAC8xDTuF9JnWLY4Rwqsw/I0F7dd/LgYbVvNa5JDkO+6/3mucQ7thw0w2o48lg1heyEnKgQ6nsn4aKPSQ/PRmBVKAKh+9zXN3e4H0IxDUr3aTfuAKwzIHFZnVTkelka++tgWAwEzhvuwOTP+zN9tKaI4AHdFMqT228yUZ5lZFY7gA7vM4yBlm9rHGM2/jUwEZJcQh+GlCemyjyb4OG2hc+1BTPupEOlYyV37o9NVXVw1s2fky1uDlZGdPZaH2b9OwlmzS5QczQgh0Tsar5h8+jbeleW6XOMZYoa0U8Ibf3fEeKH9fqqcAIw0SJ7H/MmF+0jxXidevkSgEgFjIsLxy9OZD4rFL3ZXc/ZyYLvim77LFKwHfHd1Hxn8BN7vp2s9A0Mxa7b4HKyKTew16FJmlvA3ARk7WIJRiIFFGHKKYk5VKOt3bScX3V5VgeXOy1NSK6VESFZI7b051sjPCzait8/CFHktfOH1VbhECJLKxKnlq7WaKYsDC32fcXzmPdlvSghfoV8uXMmv6yoIBHJ4nze+O67W1ggSW1BSS14fcPqbP85HmdVL8Oh06tmay0wlTfAsU7ubizcqSOgaVTxpB8/KJi+J+3XsEecxbPrGg20pwRzpZVlDVHreMd6NGGhsPCdwX5xYn/el7iAK5K1wNbUvu+SvgH2bxdHjGU+Y8NI+SXl2yg4Da8XOBFWrO2irBtJ4sT3nLozwLGu3HKjBOXuQ/s27ZoXMpyyL2cI+qmcw434zo5+AmURP+6Sy7mtzMfFwQv1ZJkMJ3x8zTORY4lZlhfBqArLRHDkKrx/rNFTwg3zWizeiOauc8jq3SRCpZ9YV2Cpp61PSkNAtRFTlyLM/ArM/m1GJiwNn5sqe8Zw6l0Y8/7qfF3nU7xiOeLXM5t+aZ+vbNwaE0q1pMBpej3cRbr3yuY9GVvP0W8XReyq48QGt4ed7cMzltkdlzMudNF2jGSyem5n71JvzJ+o7YWSABtTA6sFH+9asAsubIcrZEqx697Y/W7c+Zr8BmZA3kPwgWYUVT0Ye824NPm+d5xrQY2isD5JUfKIDZMMY7jEV9t4fCfTfw7woaLmmls0+lzalzylbeP2k3n/CsQIG6Aees5+WlW4FqCPplPytRy9S1FBt7UL5upvP5R9x4tQmmLtJaj1ntmQ6t6RAlbSqe6AwPpYCU8kNZE9AL71MgNYxA333sTkEqblSQIKHbjS+tox3TeBOSDE+/x6ACOG054TcftXQKWkXjXpzgwTagCe6CVcVS2IeAVuFdjorT3Cv0BPBfUo56xlyadkqHj0nofndz/yCHpfKBFu6w9KBEAU1u1Ow8kKlW2CQq5wdkfFl0Tf8CsRvknQ8DOQ6+bmbbmPHkhrEthc/TLzj4Y2ggyVn1JZepsaqCsdEzZKgR3cAP1HH0XvKvUH2+M8FFyKYGbsimVLQgQ+jpX8LfdfzGqJvOx8h4LcuOR6O5mQheXfxxNOdoeeW9nLHr/b51wqduJfWkTeU/5aiC1B2agazYcmkX9iPVuZajJGt0IjD54iLxUQ9zUgnOQZI89i8UNBf9OK+2vHNW/kKO+HalKT+axGuRoSgwm/HQauuoVrkbVvc+wjb6KiiZAUsgDpmxXfrpjGnQFUFciODtlJX4VXUWYJisFbz8ogtvMv4JdVyivZFfyOtQg7wsb9LDzZRJeVUZg1wGzBNTBccqFs0P3LuWW6yPKJ0XDfUB6V+DHth1Pbg5u7qacFDhLtAQ0+GKPffVXf3NogKxvnJ71yh9qpPTaMKdVEq7qNgEbakobGFXjK9e5Rk8TG7vhf+DdceoEGiiRtNbNuf3UY9JESpZWLufzK66jOPwdqnTUkOxBQgBiD+odZ3oQerpqnsy1QV+j6cruyb50LepdM7zniedBUyEpqmC5njdAXAHHc4w7RwqzACJSiL5FKcS4k8x3LMVB/L113BwGuDXRG3ihNCQyk1J8MfAgc8oKtf2g59/J0+UGSyLsJ4cQgpNLlhIaLfs8QCHRmY+LmJ8v2wfJpaJhaoauTX6F7128oAE5Wvr1/ZpikJl87cx5TOMNvTflv9wxqJ9ZG2NUCe6xkp50bzHogTiOzLvpJ2RrcBcVulliTXpwTuBzIB1t2tg4CJnQRCqKmGAYkWlrRi9sF1HvzUnb8igOT6k9pbc8qlioYY+pWGo4nswzs/Oo9X7+Kk8TZWxB+pnqcKyiRoDURijWKyRsI9TovdpfD1HKSj+Q1v5l5vLh0dHdDqccykcjqce5qV1hkD+vXWTymtw54mjhXxUOXa5IjlnumxNfecnk0Tn4hGddSWeXM+nukTNpCX70Xs9qxFY+i4pwqAj7O2fXxWyajxzSXzrs2rM2pMpshDGJpEP6rHRuk/kp4gE1XeQmm+iM75+xhjq9OGOFhPDKCh2N5BkJNNtvP57FMi3WFJHMJwBFCgevxlwQB+v5jNnV1cT6uCLgPC6/MtiYjUV/45mGexFPs6Pm/0oejLEK4L8KGDDaZFya/wxfjrra4PgUd+40dhjBH5fFMA1mgk6XLoBRWR3ssO96NcXUQY/zWiLl/on8V2PykdbKMqzqPFAFPfAPDCPByRp6SfhT5k++NHa17pv9u70K8Q/SQ2BqI+zRTVNEW+Gne9iTTMwF7227u1d7Y2UOW5sIx09QZQixRmG3ZM1mZcX9dPJiO+l255oY5m7692IRZFBEO+oNhrU30yhLNOh+ugPkIKQ4WqttKtqu08NP9T4Eg1Vihj16mPkpYkekRmTZRd/VDmfICEOvqz6xpOrOF8zj2jN3v2yFi2PD+cgWxCtZnJnNER8drOfAzo5ZaVAoihdqQqh5JgRoZr0G2EuLjtz/S+qkhCgUI/c606a0rL61Nm7ecQDzhXdtU9G3XAHa3KHVbPIeyUTGlWvGZUP4Zef5kZHraS32sopgLLLqny24mdMNKoOq27+DPdQrqd0uFMRrN1Bubuz1YJc8YvpuoMKcdyqQ76ZsHSjTExv1yM8fDJswrqL2dgOytglxonAUONGgbkbk2/9cgKhM57cv/H3mZKYOnh0yBkK6XYTPfB6ALrI01inlXZIJJCzCMyTx2e4x9++Cyu3lH5CnHr13SMWKnz5QJYPrRmYM11xrcM0E6oISDfiFK3+ho3RiUWYhhbwH2wKiR3s0qLVz/+rSYS4fXaMvPbr2LDW6jxaNbBosaSyF9aufw0r0NFUIsZl6uKaWpp6OvuDUNp7V7ufuFXJrZI/Su4CGXCi0pDDue1sElbYZsvEEIPK68dukEAQGFIQiLtzp8gDuzB8QBt53kItCR/48qIy1JsSxBv6wZnENcXVaWX8L7IbnW4ouvvhxom7Lg4A6m33Sslr7f0ePsSqDva3Ncb5yiQt0EjMca8Vr3/fSDVc9u4WnPtP2Hc66we2pKmvCmKeqZOn8emzbVmIoNlPEPK5JzoNIOw6iqptXNFk2RmAGqRQ1xn0118hjyL7SEhkTrWL7kCwVAluYxvkke5fZ4NcLQwvUOvF2QUKyLp4JNsMSzHiIbX1cJx+FQsvuZHmnms5iGpp1C4nR5/Aj9ZVQtDOTn+xY5elaql81WKL4rFVUMcL8EZkmqBCalaIHVWFIa0tPKklMm87dDRap/N1ZUifkFL1AfUVWDe2/fCkqtOxWLt2YyM1DHIkrSyZdoewTPoicKwa3VQTuyn0pcYRFAmuxBM4WW5UnhE2ZMoC/BWG26yZI9g5OODJkHejZe7UFX/727veVzR7utNsrAeBHZ/wZm6UfQ42UX/vT12j3jfHoaRy4wHgYW6q+v17Ezk55jP3euR7KJ5bUKy/Uuvt2LfcHi40sk7XmkDj0ApziTLPq0oAQJvdkciu6s5rqKLzEBZ7PL+vCNHYspJwilnYIy26uSe2mRuhYvyUxdXBqgJP1DDfoGotbHDBCeA4CAcGxntdPet84Og+UkVd6jUcW7M98+HJECy6ow8oqWzpn5Pe4EKvyY1VeAesNdnsAZUDC1Ph/8dLgYBJNXu4BtVkuo8QpSMZVxs3i7Bvq0KGwbPRj1VlBG8EIx4qRGgW5RstMgH/FqirIrsIQdvUxjW8VlDM2d1POBEhNv8xmcCAYFlZ5gL/fOZ7HwW1jUcMmLQS2U3v+1fofFaEkq1PAZErhy959kmwHB7DI25m3NWxOdcZ0kKmILRZ6ehKSual+N1juv4C2FbkY+20XJOTatBi0JP1TarnbN4ov5BGbsXaV+uWEm6iq3BwXQZE8i366GrTJRkC3mjq3LP5v8vz6brNKEfyHDI+qtu3JnfYWfQnJffMUpTFBotwfHyxZuJyw+A69JxoQFv56L+4PKC2+UJP2SPKsogXTE4/lux2d34R7C2jEYTnI0qiwD11jpkkAJtJi+f4grqk5ylK81hhZhxSNj6mzh2MKlelpRqYRqpBZ4VMrmrbYz73GPK6mxfdH7WPS2K8YYDc4W0wxRhQPJn/B9Aky3Eq2V/T0i+SDu1fBiG+hbbf1Uk7q6sbVxVzrWzFPbwzhBduWl2/JqYuVlNWZTsO5u2F2aNeW2HZXfFOMQScxTlsud6Kt/JOYq0jESJYS69fLq4zC5vjBxUrlnGZnU1n68UxARF98xtBv5mZ76RQr+bUVwEkcfT5TF/GVuGjTgpxSMOZu23OPk5Gb6Fazyx/qGYabXSBBL0uaRvPth4sH4sK+LZFpGoJK4ecmdUGnZrZYiO1GY+LSmv0ZXSbdBEv9867EnK4aWMr7T6rta0voE4N5nv6vC7Raq1ErbVX21WduV7AyKgkNQGzuLfMlUvXpfYWGTDxzU2vqlcrBanVD8xIdUGjajDZGA/1LLbStzfbQZAvzud50maXhuXG2CPCNiXpMHkgCJJtbk6DRroxQr1K0WvSHWd5RB5PujUgO8sLlv1gXLYiGaW2cKdFrT8wZtME8Mzd0HyuLd7dj23AEsDNVDX19d38H7Wq7BsNwB8eul+Sthiya2fCpAGLxDZUElVAy1Ttb1GaHB3shDsrOg0WWrEILgPqzx7mCRXbiCKRK9jctKH7lY8e+6kvPM7Nu2e0gwdkmKLInK3XDCPzIupMbdhcAJSwB598bHSI6zplkVjBMcboWy+kHvjMFN0tFd+AM8pq6KlEMgSHhnABsz4Mox4AI2spKYqgkc3dNQUa8kQPoUzeTjnZ/QWGYk00A1BYiJHU44MWeYycnLVfVZ7/YmonGheReRlCo6hPh5aUKjfM+06QGVZqjkmlJulFE2Swy9L1dNqHykfq3ZB/TJl86Fq7SLdJ2An9tJ0boJqKUA0YLOC2Pm442KHnloXXrfmGH+nQCRgPgorx/oWjX2msrcWhDFRKnA82NFTFJ/7D6S/H/YDDLAUx5ZAGQBU3yc4LqW8nKEk5ad9io9MFzNBlobIrDB2dZLEv5Zf79k7HeZwQt4juvnpc5DnqAsoWuKcZ8su266AmrcP2hbq/V7aFarqPy5+p3nkbkhNEvt8r8xt72W1duNtqBoOOMaUSZLspc6P/5LoGQDSQwuDMF08c9cLvdzjpd9S0+EEm5xGhJLMS36bD4h6VBIxNCg+DyS4GdQBzGnuhel5v50EcKOkCg3oL8mzAXYQjtGYv3V3PEE2w+6sIM8//jPSmO0RzRC6Sgll6BDPOIO+kzmeFWg+6XLYARbqTX1fX3hhiQOiOP0TEuS8KCy+i+bGhl92DKOe5vw9UOMiiDZY8mkxaVmrn4i+JzHXtGEqtk+8D3NqFq3Xoe7y5EuAwpMpCeb3ZWVGnKV0r9z/PM8cgFZriiwTlmqFKhkOTXH4dxq+f/EuLGxGkJPcHiNVx0IDyH2p5tegQQjSn082/OId2Q5TOBoIx+UOuVRPmRNmc+PqlxMFpHuDH4NGmu6wuPuqFkUUtWnzfxA2uEkBKsL0GPD8IBq5aq0r7ncNQPhAcQGpQseD9K6mtoe8CJyWB0p/wiFA+i5t0KRz9JPkvM76UCDmP+anOB1rkf4xS2IqdmUYLrGcC7nL6iPLEdcIufaNiVYdUAscEzgDhXKQCiBBRPoTJYbWYd7dNcsuFHpo2OZVkA5l7pNsUYLz6CmvGozh0kLwQsJ0psCTZ5JWoHsa0BmqzcsaS24cAO0l9AX1LWqnZBsiGe3ZjJNLA7mAovsBE+DESNYcotPUJgIuSfgdXYBtYITGXftS+v9nl4nrGyU4PuhLYHMVIevSsmvBc71PROdMB7rgY2ZQa6J0O38WijGjuUFKzdRuxFaeTmqcDACq3XKMJzpTfpG4QQ9OMZE/9H6rhdVmsiP9tO+uDf5Ih+xENhn+dNLUFBd4BBFMRjwZ62WpmUJ1v7mZQYqT9urWlGwAveN7jWCc8QRNbqY0uWdEJTMWSdjQp0gPr2d/f/gVamsQnl/w+t5M+mpEJ9BjOhnIeDwL2zAf1m58rxuj4Ol8mdPyU5G/3Iv0OPFHq3pyoI4RBcKzrMvszkdNoYzks/fOsKtY23j2+XG9RG1LKndPZnkErtpJkTr8+IIo29rWcx24Ur6hwB/mqpZ4Fy5D7zq1/AzucE771u7n0LGyFuBx4XQvi4Z51iNATv3IPV8NsZArXarvK1TWgRFpoMeyvfa5+ooc9+kpbcssAawADMaduz+QkJ6RrR5RvwDuAiYFbU9vt3KBpmULgQPlAAgQdtHwwQUetIm4b5J4gcaBNWjG9KHeXki0n2k6du5TD2xda8wDbWIU6uN4Q5rBWHIJAWCAvgdiKTx03KMahuPLmJuzhTsCh7Cx5febkupUaEiNJIe+xOeBno46b/3+NaC+jd4H81WpSuQgTWggEJEs6eifTE5OdlUQfpZ+RqP9qGIaixSkCltfoddUbmGpwiiU5tFuoAdaLwLKHywvmCx8kuMfhtpsOa+KX5OlhxuKPO6TnCLUinTVtOzXlD7/R44p2UjEM67EGV+pjpRcGUxkwzjdxCjoqECstAfEx8rgs6RyIOa4aGmGrWU775WLvqdB4dIag7INwfevItMSJ2g/ZkvpSn6zTzzYL1P8lwqgl9gXiy5FTj5+u9uzQU9ip7jLn14/PmDTndHkZba3tK55JRzyDkPoD5SlCUVDJ6CwlbLjk/sLuGHdSGZC6KRq8q+z6Ul3Z3Y6RlXEX17obxGKXEGnmOkCaznPyPWFBqmus3IGxnl+M6SJgwId9jYIBC2wE43rxJuptsgIImTTx/5lkKWQuFoO59zMLG7S2ElennGDe7h5XrmuLeUvulwuzAPRx0JxshvXGxqNdR2WZbulmghiv5sj4Q4TUKQhT7gPFLJ6LUB+uDXca/uzT1S9sK9bxOpBvVls3m8dj8QuZ84K+SCSXdLbmLNivxGe9Lb+2DuePXk4Vifg55uK7i+/cjGaIUvO8zP7g2MF5f0PaRdHoMEDmH1sg9G7BxkAViJG1D2NpF6Zi482K2teQ/iuxe6eR35xkOnS6rqM2wwGzmowQNS0OY5y1vzTDVE9LK21xXBb58BDUIdVe3Qqnd/U0obQWH+oIUiZPAmGQDc+3hpfRAvwAOoDkBVeu9rJQ2fcVgApXJ3QZdoeqMAWquyaflX4FRTy9tbp7WGyK9cQ2uPVR/uD3V2XRP/Ua7hXAJZ2ogVGqvIXC+Ka7NCegX0ChABOSyn2HoB7HWscceJsZFSPFSRtA310ttfnYcvBauQLUzXzNzDF+BNJ2Scq29YP86Ol1UopsbFJ9Tduze+bP0cNBu0L6t6MSQPT13XAV/SccwzmmqMAu4F4W1MhFM0DF2X8JttKbfzdM8JalxAfN0J0+sYNsKiiqdKLZoTV6CZor08u/3vUbSZA+DYcZY74kfGAn+Y3s62Z/ef1X/nVgdkiCsSZnFtGlScwnAcm0d+FHxFwDZ8Vs42G+OuWy0MR7UC06jM1ZI8e5u4kl+5zONJwbD53j3W07tAwAlrk0owBaYsZda6LxcjPnr3W9TDI8RddL3dmxrmAZeMwaPUwsK2IEcq3AXijjHEPZR5ZcGIPWFAapwUiUjGoozMGsvZdSSz8ppwRVgyRJFKEr40Xb2ykiLiyiNfMPcXaYxnrCecFp4cVw1BTux2zJ+w9ySTIHLkMFvmbYmL4APOsVgsr9RzTNFLHXJVOUoCWjNxXlWXN9rRr9lCALkzZR87UI4gxPhxojbpzbj3ff2Wg0bu3aep4FxxirqMYE5oXhvYBE7K3rQ5MC0m6YaTSsrGQX/WWFncNIByh2ZMQz4AiEpOEIVnzawXbH8MNZVOsjL1FpuduJpTP7SaP5Z4drxeHnyqROTia67NofFdpDukS4AhLhAGtfSGjCDwuQCdKMAaG0q/VasjJe3fo5YB5vkCbK1n7BsPsYhFzsk7nqwm0ORQ8vb8pKkEs5odQ9Kmjb3/Wd1EcsVGRmJJUjQYKmBmmg4+8uD2e0cnMPfLOxv56f9R5dBWOQvCJuZ4ItGg8NsAi8WIplFhDjELsHde8M9hRpzf/oAwev0kvcnRsTRX9bOR0qrqUUlmQ2cbfbv1egeu+qFuabJ7ScODfnCmaJxwieoxYGePK9TjkbqKg15LmRItPTgtG4j4YmCTDMt2o4TjG/L2mv9pQ7syLmySDQ8lqKbqwcVsJKJ5YJfHh8PCEM63TTrG+MzOefvSQ5+nolp1TxYXveApuB+Nk/0AYjulsNQpCUzQSQEKGJvB+TUwPsW0st7jD/vu3hqMs2ufGp2k33ySeW2zKyrWctWpO7YEHxQeEG5cULnjnJlZorC0tfM1Ox3UZvXqo42boT27aFjbwFmEQY65xb6gDZeaW2VruOBOBCchZY65j7aj7WNf/R0gu4x8yT2Q2OEH7vWhZCW+uDomz7CHalfQrzlg8EBfyDQzSMD9uYlQVKW5tPUXeeKv2sXk8K3VD+4NZkQDgRXuOpioJiio/UgTFZKCee/Q/oV+CO6AtOsDKY43JtWQz04yUZuU2KVRRF6IdsFRV6ddcvik594+0fcRikr/MbvBnb1yPd7e+pcHPoetBBk4NJKen0T5NuuNH1lKFbI+qRxYkP391l4310yIlm2bp24pHailcqEJ+t20+c2GZShkE9OKaoz/KhNkLi83W1Rb5b2KfJeOhYjVFD+nZq1IlxoPbQYMRcSsQrO53Wn5zkrdiudmIdZuFKSjJXJ4wMtrBKvu9OYELNh/s9r9lp3VUiGanBKNuCOIXCzbAS4j3jbDxjaj4nO6U0W4llNJH+zXx5afNpKE9gaFIeUj5px326KuizSWUFctOi2tS8T+JBzFAPNFOoOblVqZ8icn5LvtGWmoAp02yeCGcqk9U5LCdiiYDSCufTjpN0LWt7L0YHe/98L8rW6cnkXYgHn68m7EJc/byIrw3vVZk/JbMrLLrgfYnoMZPaHuNLD3l/ienhzXN0Kj1Vrw4w2JSJvtUxRttx8chV3MMeHV+Gf2ORdN3+wK8jAU+UILNLxug6YxgWjMfTCV8xOtOKiihkWQ3qAw0Uqvv1ji9rr+WF5tKQ6gpMAvwS46yoG8zDvbIQXjpUvWePw+1p7LYdk4FBA2LIwnc1mTTt+Jrr6te7lW0U4v5zn0xV0crIr7aU+LwFJqaIPHhumPwhL9Opp0tdpQPyvy4/hRc61OxsWCOPV7Nh9/1sDKwb9DDtqUEhPfOhrUt04SEdHnPJcjtwzPgrNjxmrEe6PGQA6gD+1QudvEHMyfQTNLqc5OHXvGu2meDilmg+rhEVJtkdVwavWYK3IHCnprHcom9Jzem6zNTpSHXYKiL93eeyRzZ4w3N9NMKxUOtO20KqsOseSDN/U/dnDm121EW2BIs28jEZh98pRP3WQEJzJQp0EV+A1dngfbKkJKnTseU3ZLfL8O3oyeRi8aBcM3LQ2rZr5RaevuiMIl4cqvZYrI9An6hOyGX/FD3B76k0aPDJP2mFC0yI5LKSEuldIKaVdb25+LPdd7sfUDqPEzUAg5NHArqiOouh2j2fB9DtJQj9zQvvsz4NyYkiX+LD13pnCmqB5bWgusyGmuJWt8kBfvvMN0Zz68iH0AiqjA70rffmsrMqwBrfVE/klOJkSNUPy4XwbYsvNdfpP7mOUsMp2QFC2vl9knX9MKk7LXWgjTUlpOG7m+4GFFzAJE0NNTKoJrAxcdEXZMDHcGkT9OZyJZFuSQpdt+81v1wjRauBXpxZ+XC6g5HeASwgTHxQBnqgONBxE9W99XsTc6117h23VbcY6C83A123ba0yX7IctzZ0hGIDqt5gWnXaw1FfDGVbn6LXXMlraUTREeWf/VF0sg6FLCZcbo8DJlSFRLfHFpTYlvE9W8jo0oVre0z5EtnwwfaQc/K6cJHSoowrpn6TgrbeqH255dbRPwmH9umFf8oNmK5dIU65iOQSOrIJfym71X1ulxSRavawUGHb+69GgGvbXGkGbk6yVoXD1HWefStHTsS69DhZWev2Ntk49Soa7mnwhyZl03DvZU635e6FbicZqNX2bE2xHSiOHV9wImtPk+2Y/QNivXpxRP0Y4qktIq/U5vXntiZ6i0zA+PrvKKebPpX3596Uz8ztbEXxd2jGloHpN4BJKvMvKPI2Ayr816LtETzo78oNdWk+wxNBHbAlkY+68auZg70ZOp7Bb6AXB0oQRwv8IWvziOmFtoJ4R1IJ0hYlEg4SO2pOuuAe271ZvHCznI2fFjbqbo0xabX1P/UZcoPFTFIboEnVHL0wlUABPP+zNTBH55ls8sYl/mOhhQA/fpSsa8QTEHj+3IhY+K2uCHX0BCpYih3Neo6ROobg9rP+RG+zTNRSKNlWZMdi+SPdSeq1leLa7x8CneHiQabuy+Lma8ZuFsq6lqOblsne9LT3fSYnXYj3E010JBGXZ2PxtsPoG7YGAB9us11rQckiWXV5LJ92e8iLedRJi+1umGnCnkVYcNz/F7+L+7+hrJN3LkTtG8gGYfWh/HUNGYqAUTTdXs3tU66D2RO/wbxuQpkoS+dWzi0U9EzQor859XZz5YTsjdpNcFT1QW+aNwqjgjlrIuGDSs84sZDfjziLH8Yj2u2msTnVRTyKsdYqSdZZEUoWRfcVZe8OJTZS1Zqtz/3s+h0N31ieU1IW6SZQZUYEfrw2ZMPxGrAXrTSM9CyACcsnqwWejINyHAHJd2alhwQ9uZpVXrOQedRKjqzEcC0piZAB2wkQ7Cyalu/cHGfytwHZsbCNdV9URuGN3jv3XK/n4leYuY9Nq0ZmSIJKwyVYFcoAee3TeGVfqNJiVJCCuCgIoADSSa+2UAKqbaP0o2ff08RPQK3SP3WTjBER6Xx3xaNYbv8kqsy3uGxlOmhAQmpBsnIYII+5nIWRN08j6Ed/q26nPichdd/S8JiADzcQ4LJ8lffeR5SFBeHznp3T9pa/nwMFsin1ruoNTo7k49pNZup3g91+L5ea+QYJEo3E2CTbiwNzaauhj5e68DtS06z8JkSbB1zqdwhS/DEsJpw/ZTMOyzjsUK5OJTuaJ7+kfLgyD125W1UyaPjLJtJJf9yhXiTgH/NMUdutE+5+6wECwEKatIBNFuEo0XjzE75kfxTi+cZJkJnlb73E2ca6PLrVLZKbbMau4iV3595JFUqnW94Dr5zBa1MarYVqWyPluPo/ZwmUOGpEdSoIguwb1lmCQYx2an3OEqpljIgSUvlOl1p63QQycRXfVTsG3xQG2qikUTSf0XL36+wxxFIfWg0t9RWrL8aSKE93ePsIyT+3P/FVEOi6AVS+xvw0A9F4RwXZVNm+dNPBu7h6qjIqK/RLCmagI/Cj2yb3FxuYiJ+5JhHpRVuiivsSUs1yZepmsqTJh/IMObGfghqz7XWY3UT19XUeUTo84sNvv7uNhsqPW65CBnuKLb+ruX+nbizqF8lPdA5zai71mTl1zpAUQWhFL25suLwGewrsZw7mBa4G/lY1iXh1BfgXEbQbA6NDL/Ruwl/D4lM4umUKIRr9QtgqIhDpcZl8ucQaq0AtQqsTg/HNAwACRhd5GEv8LYgFdYtbMibII8DpmhFbwX1PtOY7mzL8d3ApTTOP2Qi2RZ43Q3PHJyVn2EErbC6grIYwm4wFx1wz1ZP41G4uUX2cmooE5YMp4N7qrzUR1tPaO8EkcHDuavL4kuXTfjpYi+vJ6UrEog5QbEyIuucCapNeqek7AqZUzKleX8g6HIRNqDrCeejLgkF9IRbKvMFgtLLlsqikIkHlVEgnjk4PlqWEtkGoLCQlKbbQbR13mKEGWClsRXumwK47rDsCFiWsbK5AMuejfXt1DkP8y0+XDzluSZF7P9RNPQX7KF+nriFJTIHRMnYrjanPfRQBkMs3I90tBXhtby/bqrovJWheZ7eJLoOjwfV8ZX4cZAQG/I0AsiaYBk222k9O9h2VwjpMozGgqslWVMh/J3L7cK6awzsmARW+C/8ee+y5/xln2l1G2EWndcfn3ISdrMbXIKy7WErtoybORV6za77dgZ5lsVF6UZ2mZ+Erkb5d+9ixtcoWZkzYS6H/wnybs9m1fvHscNBYu4+ERzIn4zXKmd68dgOXQwgqUoS/hzTPvWomxpu0sL9dRGXSbYe8aaGxnpCPVMpYTvAoG774hJ318YK39Ub5v2fTUYUhcv7bTnh4NgWKRJOPhjbRGY9Be8qmi/ANbjQbfxt0LgGlQLn/LZIzHBj78ne8OJ3z+ONNM7JPZh67/vkiJtVnSIigLXmD0rj2aLE0z6VARFPd2PyzoR2TYINVTtssolVeZ/ON2/Uh2P83RbnhNwA66ztcdh8cRBsZ5dAwWEzhUbvDzUT3R4LH+oEFvkF00KjV45JnoWY2rMO7xaNS8egNGOf6F51CvmXXsv8iL3o7tgwY8I0NLFftLYhId+UQ1v3ar0rHdWQ5DMbRrzeVusl6HwfKOq+jsXvQ3Vy3CMQBmXTDqtVUlt3gYHT++Jf3b8nZo3SGlt/KqAEHGh25/TFiwJh/poRuG+K0aD95fmR9kO+RLutncPsOMWKDmYf1anSWBWv3LtrpTv3lWkwMsKnCWiNof37NpmPAPJUzcu71HQXNTfTDYANCgaJEzYZLsRKVeSmxxIYuWuugPGcI/8OtsxLKJN1+VPMo1YLsuUQDssNtnAKRfgFbKe+ynvn9olhx4CpOG10Sz8FXZpvj88ndBhM0DLv4Y9M5FG7bu65NtO2sM0UvpZo7QbWPOczorI6uf8panVuVfyc1w9s4kfjHijAuKyxfRd/teKFlK7U2JxniUeuP4OU8NBdhdnjKsZXWOhEPAuE0Ma90dh8oQvCv/Ms4KuJhTX3O06NVtUjFJNRbXHTG7l/8Do4qUZXztqWYAlaQ+tUOAIvD0Uh9kzjX1XuNXH4rg+jk0F8ebrCMzRdU6NDHoGLwQ7t1uN6i1HBT6TAErEUIqjTZJW5tD4fNJvx+uqToRCcteHvfGIEvdxQWL/VEjyahpjoKqu2g/uu6edFKUnLUn+dn8PEO6Eht3KLu7+p0EVYMZ44IS++kaqX+QZHTeH1QkA0ODUGcJm40XyL/rBHol6pxHFVIPnqGTLIoW7/oeti3L+OZI516lFzXyy3oHS/YHV6H2ksvD01HPPJiq/FjOl6m7qBIfl/aVtutItFaCAtGlBVdT36VCTztG15MOg6BHYIWTH20Dt/rD1pmi8nbwGeXS10zGlygyjr9l9MQdooYYavrUFmW65M63Lt6YBGTyyGPPyxlhJvJ0eDxijmD5m2Dey2gkiJEVSrr7RMtJP9W06dYbJdCn9sZ9hmJP5A6KymnHQlCNSuR6DmyISlT74glSges+go+daKtlMZEjxs43afj3RhJ2iPVrqWcX1gJuIe2mKJLHheCUPEfy6VZ209BwDjwqF9vB1czoJcei53Dugzuc8+bGS75ONB+iwp+h3omZjwM2B/lqgAim6EsiFHGp+MzECBPrzzkq++t32oE/InKReldE0sx2dJl3NeRmjJMZO4ijQJTy7EuplWeOkVgokaNh8x9dO6rf+N2fMoGEbaZHOJKUGHahQ3TJGjGQnOswuszi1DI2+djkzdFL3YMVVtQo4iYfsFDPDZA62K7tjVhx8na0nhq+vLx/9J3FmGRKFs4lZdZsPFoS2l0vU3eYBID7IiXqWApxoIChsTYguSfxLEShfnN2AZgpXCDxMJsEbVBo9vAsiIciVzEA6zQOe/BsvR
`pragma protect end_data_block
`pragma protect digest_block
1fcd11284493ff252de049c4f211616139bc6d62d0ab650d79f019fe6c00119a
`pragma protect end_digest_block
`pragma protect end_protected
