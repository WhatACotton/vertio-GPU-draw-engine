`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
WHlkEqH26WZq45fgVVRZ+r6kxsTkBqCYArTv8KISqOOWS8tFTuX9VoM1VCAsfUcE5CZ8l9qnV1ebwEWC8HmazT+BPf67NHJ86E7+DtH/IaLvn8zO4zNGBpPRg4dIWFFIMTzfvjNkQLAoSn2WRBSUnfujcSr+ghb2Xn5J6T6zeaGhfVMlUQDcVpW1caFpRZuiHkEmQoew8vTyUZG5Yh7I6y5IXpbCcieq0BOQT0ARo+obvjTzGf7vyWbwrUHV1r68Z13LMujFgr1cUv394LXVkyWcLJ8FWT26qiZP+CgJxFO/1qFVkSDwaF0byjLlX9SKh9dAf5oKRA30ugh041QhVp+YF+agP4kGbC1vp/94GOQFJuv+y/KaF6WQ7luPEZj5xXMoktL5kIzY7NZT4t5e3qHtDTsvsxZ6himxpAKR6vZb38os3PMBIh7rp72uaMG5lPMriV/FmXoImrY0DIYYoiPe58lCehO2fMdU8vHVNsajmwCrZdXeVu3/I+mKTn5YLHgP9He5KmE4wK8EdFDaosYO1zLNgpROlR5NBVoVMvzKLw3Pmd5wG3IgN2Hon3jUeykXjFz8ud6Yk7qgEJlWxwS/tT+Mn8+PsOUUUoONKShH/PBohz2ieqMB8fJ7GA1Vm0nGhiTyHt17ve1vldxg7SH3Tj9jIfsrrzO7UvpyKRKjTpfiCaTJRTNfkn/T2JBEA1zYwQ+DZl+CTkuuS5lLzmWVnEi6PKQJe1bba8W6NH8wqa15q7Q/24Sr4Abr4vy0XWbRqxQs7QqRxV7RMfjnf053KghX/lBECLpMpx9yBf6LEf1RqQRodfWrNb1ccSDGYWFudc9ec957C5yj7fLhe54HCg+o8e3lqy12dka54t6d3YdXNh2Ugk2f1+njuMrE9MBpDbwelipa5zPRXO8QdaRYu+/wO0Ax45EuRNKTtdXPVnqzoxchDuL5wHfNFArkXTcWJQt7HWC0pLPlwWjpCxC0y/sdFHw+hdN0qVFLKvnu1LVr14hLyJY2IHpSYR0RIF+oqtZESCNh0yoIIPIDY8Gq06stgLrt/beKkodFsCso6sKveb08IawDxDEqmWU+PfwpwICAX05qUmC70kbhJhCcdQESImH2sd+1aOnr6Jbcp56nQo4Hq5xTP2bsvwTkMSm+5GGSTn9tHrVIH7K+kGNAvCvXaDU+OBkDicCTPprufnCQ2HFItu/77xRokAM6T7PIMFFqP9K+2rC4NeStXGeZfMUTZu4LzoGeZrXUlEMdXBbJhYtmLhPLNsbmMwVJO2jR5Zg9Crm5qFS6xXLGFSlaTFK4bibmIxT9tVf/EmM4Zr8DXHH+FLz5v712WtCRgAqcsbeguwq8EWFwR1eEEG76gjXIDP0EbVtkm9V1gMU/+6FUyuypi9VUp3QGLedta+Cpt6guEk6aaN6iSaBpsBla3hxubHVsHkCOL8IQHHQ3nEVmNnUsSknJdmxTPPonVjdgqw+yFTCq4WDAaav81F+cy+fdIMRhIpsRn4TAtMeCL2KLP8nhHuXrJiGge7tPQCvqmc506pTtAYHEA8PMukjHWP8y9CqmjdepS5/FIYXGUty99Uu+s94CW8d+k1pqoK7lBrih8BXXH6w1xrbIdmDDPgA9tuH4N4l+dxiK3bZZ6toEYCoolYUeGxqQBni8Kps+9RFFUQv3z9izdOcXu/y5aKAAOPYFSLBu7DzOAVYJreWGSqPSEPxyYIu5eeT8a+vlpiGcY2eqHIYm0KICihWY35zclboBhRFPb65X56Z6/7bHfBXb7o/2JVpbBwEKlOZkl5BlrGD1XUNJcRqFuC1C6wvheBjdPVwhVD3OHf8oMvjhaswZ0ZvpCiR31ldd3B0ZVez3T9ebPloeQMkzpROydKHthDkFBN4FcsiAykc/4y5oJlMuacNSI46tYU/pvJW4W3oigb1rZ3H9dhRaPEQk+wApQ2JPIuU4f/8filHEI3ueL1FgMoMXJWgWwmsEaQLRRWbZwt1PsY+P/zbtWlX4SPBRnqQRZDrpRxo2UrxMbAqfpykUf8294+geekh1qNwduxFY8g86Y5sODS0BaKaCYqk0alHZ1sLDfCNQEjiwrXIVG0jz6RAvHp+Es4/++FCOEDYdOatzdDQo0wF2o8tJBpEQe2GA7Q/IuCZOcj2fG9ESej7xoGWHiWIOdmpaVVeUSIQgmDDxvPwjU9X7EWd2WpHymdMR48SjeP1e2FXRjFdyt3Vh/TcUWXTqTR3v5KyUvshbudkT0z2Hng1HFjOY5HvwPgqngKVbyUD3Zn+UQra79jygJHygqQ3Yb2zNqU13fv88odunYa+kiYnGRI8M4LnsZV+Z6GnnD22VKcxt1RogjGjjs7SX4FlPcyAaz4x1qfNzsew/RZgLFeg0vIhHRAH8McYDBec1F5k5zDF8uPhC9ED7uxricvru8exKNUUnGvcbP8CNjYFFIq2FqdIvQa5ywAw2sQDc22UA98jZoAGSxGclgD47DyzqU2unu+0TG1GjNnvM0L7Z4k9OTA2B7e4OW0TQ5Ss80i+C209Ve6VkbdFcTGibb78WW+twkB5eklbHi6r/7sjs3mf4uexPIPXfdnPFqWs9/Brxeb4o4ZcGdWwgiL1hr2AHqS8iQDrQ52KZe+hkLhDipZcje/f10833t8S+U5IwUlVaHsefKj9kzIE9OqFqoEyavaIp6UMsfoAIeJ/bMo2expqm2y5SUKOIu+wLkmIXncs9M3cF040oWHOCwlWNjgXbwMc6b6dLPeEvmx8jsyp3M2D769deErItFgAkA+SQq4gD7D6qf5x6h1gvKtc/GvAERfNDcDXdkG5q7gKnqBGYxCjTYiMaG2Y5oC2v1LM4Zh9on88UPwtZN+otrjqQSTD7kVlpyaJpzluzMeQyz/Mb0yvjPKif9ArHu8AYYtwBHhir3jG4NEPekbZJMB+5N0Gww0/B00nEbU6HZh4O6lVCPu3U76Qswj8EaxK9o7gR0v452L6CKHGPaATmqzQQxKGM9O/GvvtCx88AeuS3qRk0KgOi6hP3PouhvGRgIXJ2E+rfUwdoXCEEud/qN05LRnySrFJ36TK2W1mmuXoc4k1AiTIpry1dFfeUxtt0qfM7B3WxsxCZr+pVkgn5Xe/H8rQVKFNZhyOHOULssm6MyhbjF8JmP9TRBVCn53+BccC/s5o9XaTsW/h6Cz3zKvKjj8wJEpuciCVOL7luAc0UDNJdNKfP6VwYQQkQRwQnkau9m8qfDD0JTkidF84J2GxclQNA4XluZG3nhkOk3SHCBcQZM29twWi7a7j14XLyQBu4YNjEFVRZ3oQ56vtN21Ryhge6c6OXNjt9K5WArT+Hm65fNhiyHUVzq8QG6/9TKAN7NqwZ2+U8qA2twHV069ei41S9sfyuXg5M4flUoAPrfC10eXZJJK2xKeMR5NPuaAI8M2ycJm7EqoS763i2TL0GorHUyCtQ2U8n5krthIx7956GxSCHIl9q2WqyDQt0+H6/cKuU+du72wxn/Yltc3Ds91hCQJ52Y18EBGrgNJCZIgmRp1T20ECDm2NJwgUKY+bxxNcrkZlznmPyISimpC1PdYbWsOa/670GMQU17ioO0PXvcnqCHrDau+NldWr5GfGopuqBqHaFZ53j8EIzlN/roQ8ztAriKNY8Yd594x5R0e5OKOh0Yf+4xVQfrmSV04WMHv7oWlAraH9BDlzVRe5pPzvSQ/MAig6Ok2uu5ztipTW0YGJP7F9/EuOV38wCL4Fs447FBcnAovcMXQEABKaOz1b4VDLuIeP1yuO/YdkMd4PTIooK5kXDnmrrxHBFcDFRPIe3u/fm6wc2RiPikvMSe2pIP6IzN759zUMz+NgxU/C7ltUJYOF91Y4fbpk/8cGVbcaahto9ZWkjQxf84Mpjy9Ch4xIZyckyga2/3p7jj/oWok6p5RiL1f0zegl1UgksGDeg24wkABtGDWH9jRS2faJA8ruAQ3scjcOhOobKz3F3WVBFkJ1ilXXYh/l5WrWruZ+cF7p48qroPjvnE8oLap8J6awSOaw+DDjB527WFBN4qIF7VqEfXQn+9YyEqJ96UEXgRqGi4KEToZ888yTpg/XV/Oa2CGNKMF4cng+dOaw8DI42Me00eGfISdaWA0/5yJE+GIQ2dVavRfdvuP7LrzKnrs0OG6Yp6S0IPUqHxZYd+Uwc/inNpn6Vat3fWFkIBwrsVNQH4t5H9Wr1qOkhFcA5vLQbhxUgSjMfPfQQSIGLuv8H/sMNxxCOZg/yeQvheZam9TBbLUvZVzo1v59cu+SD0X2tvxm2r0SmOgfDpKZnghAfhzAzP8t55u39O84/mEKngQkSxp42BQNChlqidRJoHbOWBmArChpmmx2lk4b91YYzYUlpm/5e6qkwFBrXc5P/dXyJ0bzZcAe4ex4xWJNnVX1rePYT2MM4WKwPwm025qKNHoIN87IyI/8TWYm2K9Yg8a2R2eaIbkN1hqX1R+G8NsxmVFqQEsnvfu/IN8FjEeGju9U1wrg5tQoTQBitD3upr79W1xNoItFHGvKIf8dT/hW6RDpDARQFo4esve8IH/LhWfgNdruf4fSRJ06qhNwWJcaxz4voWd3h8/CHg9ZmbH+9WPeJsF1BZP1609pHs56VPAJlwWg0hBU6Z+oRBRap0JAOxPQnkAE8ocUjHXzK0BkTaIInMH6ehs/uYXO7m9Ce37LlnAyEZ8iGVs0p8Gw98Sz74+LKT2+QDKyy4ULS2teL+l9LF+SnFs5f4BS6hsi79nWwVIObyeWXy7YB9TJCS1AGLg6K4lxbKYdDhGvE2SHziCD2qXBmLoRhgnPKY7ni+JJE10VTs39D/+Bw11AcJYq1g/zbpktDACHrI9jTt+niQ+rg9yvRiKsGB1v4hPg0AHo2fA8LQBcO51atCRJ+deh/GyJJBSuHP8MlFaERrg0UCmLh7ROPS4GFk83bo6t9Qj1acV8Qx6OjuoiH6VnKz7+62zTzXZhMqBhU6XJkInhZnU/dWKjuM+XuQBGnTA1sODOMZBmITsghs8/WGPro6b3g/+0UUu4WiLEQQqC5Gb3voxQ/vo8NfXSiSGQr0vOInso+qOAuBBZrDkfu/OuMOfhFywCSgXfl38T2oIpgdu8MB4Xm4cYFW7Cpftya2OE5fVAyQcqCUa5DzxkmlYY8IbhKzFtfJCEZ/QhQxFxttBvRlvKDq/1s3wUi5GFre93HslV3cwcRXkCv84ZzpFm3x9HU0+R+tz+PNj0bM51X+Bh9Guxiift6D7VhtMxaATXZ42UZ53cfTScn0seOP0LBnzSLIKtioG77ISvxRMZctPWiOHA8sx9V/vAbrUhpWMS+dlOJhAMKARud1gYvo81pY71FtHjooBoYUoDn9vNVzMqQA7U7ZNB/tUWtovS6gAS7/7Gir4+MtLdDNJlNQK21iDTqZ6kN+vYmufbPGj+lpUr4+SE7ghVy/4j/0iQSnsjEQoSsMORpHTa4M2aieG3yI67cqbS6VqdBhI86ofdtiSeHjBzHn5G1+tKZ9bvpnJyXenOIyRffxPkSe0zPwxakdL3JT2XWpOuvbUNDQyaKl+Baq2JdtldOZ2IwyVvAJ0QND0/PIKHW4JccYrm+7SGiciHxQg22Uh6cINLbfdfvVS/Vxc1koEOczSFTkwwDff3BPTG+M2ED/dRkL2qL2p6L3BbwLPtjHI0z5ZDkaDrMSSRqqeN768UPztWxThJL0C507cyj+SJMK/2IZMEy56+3pHlEa6bQbtH/ApsKolR/dhhTq/HKsPnW1FLx6wBOIZogZ20/iOfmMeXEKx1+e7+ZSo0FST9FR68/hN06JkTDN7KgV+zyo+7wPZWOpr72Dl6aW9xZKFot1i9G+/BdxUiH8VC+8HaR0Yc3NXY+JnPPcy5/z1Na/YnA6HmleqAaJTjY0nu/ySJsNSrs/RjBAbzMofAlYnSnZJ2dIx7jVanQIOGnskPLGcsMcmT2vaXEn2Nz/dwGY8aLsyR+FJ6loVbjhbJE2eezMQDhpiOUxZCasJhh7wZXoRBptZ1HKItRgEER5U+eqC7t/UfjAlyTs/wncIY7wgIm1pwTEAKBo86syn35nqA2tY/LskZbK97acb2clkTh1bAPBbQeZ1ZD00tQd7lGjIeHw7VSHYvQaaWXcmBzyErrQB16u77wOzfcJ42qwRSmmhiUxGlKlDhDoQI9QZGVUra6N0OICtsE3ZiCbeWvj2pTL6CYDU3+MFFKCg24I2n13Q22hJxsXrkMMtaU11AW/a7BAxTiGfw/MTLNytxpBDYEtts7D/qUEli28OhOr9XsotWnFq293Rdtrtl+z895izM/uJRM6ifqnaI4VauuJHleeKLAjja2qa0LuBJcdzi1eT32jJZgvz86JRQU6q0llxQc0hwOycVFtGNRU94I2IIZTs2cQVSQy/NnP2QDXmbGi0YC6ZdvrGSl0SjK3X2yKC52+Hm8cyvYj+pmqRH6kGnIcnxcieliZQrRcBsv/5Fp/+zUyT1MSoURope0rsTI35xV1yV/eJWZPMctv8Cm1phkkcJAWeDV1p/PRG5ZY9rlO1s1TqEm8LAZBPtcwm3w0eaJ9MHltEoPS5o42VS9bC0MNxoK+1QMAeY43gXwAyegDwVgr2KMc/lgCQOXCBWe+5MFuQ34QiKfp2EgFJGG72FMYttO/XubNb7S+9pDHelGxMpnh0GSVyY0c84ojCF+dwSjRr7TqBH+rgbKqMvlyKZxOVER4M8kAIx0pRMwKveGPXQtZ3FrEmW9F9VcOsomq0WvDg8C1PsLSWWRIVOr4I6IFA9RPKFssZsb8B6UO8Rs6/bWR7NT6L/U03ehPgFIcHJ28ZtCvAG2OwPwn3P1t/BlbPcgOuDFXvsPxlJH6NyUUvgia3NArdWKkpKI7eDHQ0CoPGl8qA3R98VVqnBXnVDsbu3co7WTOser6Qp836DVFJDbVt7+azm1yxQ4t1zMzRi2csYmRrcrmPNviwWNVnvXRn4s/1xGmDcmNwD3EROc1qMpeTUKlcvo5F/V/eCyRbxRFTXQik06wWjMJ8aVjIjSlLOfBwHF4WC+kWvjg5PjJwmKQYCPrMZuCJAJIGq4EkNVyNq54lHQifEAEAMolFoUMtayEVqqYfm9gPw1ZIBV32VvA6YvNGjsLXHZkU2c7jKrnetY7uqywkBIF0pwA2qLScP5Nfd3zTOR+4WhAfTYBbtWQ+r+BwWyX0T74CrXOw5tYkqhQOgxNk17zhrMxgeWzKS8CQp2I+bytpOOwuIO5SfLwl5S9sHX2ynbDdtuqd63gMFZSQSOnE8dGamEFTOfzyLLqbXlCiOfNrztiO9gkCooRKhbBUWB0CazPMw49RRDgxDlcjnZLiEca08rssNlNDzTOJVXFRCNqv91xARX3BYtwY4bF+SCi2qBL98rp4x9mRZwIxE9K2ECAtWhwygNOIniZ5XRfwY72tga9q38W55zUSoLJqKWuX435L41zgK/LCGhRJrrZS1Z2cBqRCD6bZhuuH2KFgqrSacltVvXFgWFEiYQswMu4ua97GfbpEUnXbjoCHWRPzQ+AnYHaL7e9d5FUFsppHGg0dJfe5bVSK1ah1gUVh7jYOIoz5ZymeKb4Qm+7DuKPPMQtGE0dO9DvmmF8JwMi0UBakiTGT3EiCJJ3nEq9Z1RiHLhYNHGMOXWKvucDM2hvx7F4A0UMCK1s6Mot97cthFtcJZg/XRaXyr5wOS5wW4Y5mvmHC7xprXOYWArHz+9f/ONLVlJSi7frSXbcJGW6f1bOsTFTinY9G4suyNLrOeMX9PZpS4dwgBKVEN+iWO0eN5xBoVIMNKDy1EzyvA5NRIoHCDkVGTj2fZ9d03t42wLQgs7v7H7dNVmHhTkJioZ+vp/sA3VRYO1YGMV7PYwf0/ahch0DXvnNTC6k0MW9S6PP6sZn1sfFrKPSzz8xITT8y+H3QQ7Kl6LbxIwRpJesPP18XvjGEJfQTG4DrVQfuI2y1wIePFVkbx4Nna9O7yA4h3oF29vHff9HANalMzGGyEt8kMuoepH3KjW6qXd5qFhr43SCEzvYk1cRF1GgMXTF8hX1OvrmHWke00tefb5Urbcv3YjCHPHppeHpYAOXOQ4TYMqQ6QIiu9cgLfObxrQYesMWFXFqSD+xuqOiS9SzZz7VIVDH4M4s9BvirmssnmqzbPzk4t+nUzDC377jNfXHDuAygSKsyxfd4yK/t/RXmR4f2QE2QhEKoFCpFHRI3hXCaqU6n4hl0TIQYcVwhFsjB8f/tWXxzhQ+EHG6scUHYWBNBnY2PDeorfuqIi65iF85uvy0CY1VRQgyjJuJsAgfyoQApdinbCoiSwl9Tv48CAXG2Z/77RZWD8Okee1xPibeQYTrVmWV5rgttTjnt9bZCl/NRgT8hqNlr38NYNnEfEDptwsKlOID6KjaWj2hIc0DzwfNjSYus6sUxmsageFaYMlerEzBkleaAc+E3P0eWWtjboy01gU/cFd+hfQW1ISanoBqFu4KqusvDZ8dYnNQiOiJ9nKNYWwD4dyNbc/SigI0xJ3+kZ2/AyQwIGvKpsCvsd+kxtdZZ5MjGQeJRPQ9un+pB5ThdtO0RDAwxDJOxEmkZTLMlub+DDvnc6d6ICycT7Cx5EaXjurvHyXrPFgay8mVhY7d8K0pGsambqLd2XaQO4ifjUqwKA8BlfCmdi5c4y1KfnNojVcbNgbJm3oybIkrvxrUmHeYwIvbCidcynNiBCgnrJtz6iT9UAPKMj++YjGFfyT8uOQ4vOO2n4CRWkrOssG2+/Pm89lH32v5rccgV/wmjndegrVqOVJYOHwrx1NJAmbpTNH1C+FIpeHb0ySDey71A4vjC+RktIK/pFCM6gg9w4lzSWfQngJW0Cu9Avzyp96MBaIsLx6GI+w8hDH+RZyN58S6oN6BC3pNN3dCdvudoc+sW9/3a2eqKH5wqBZAmCY9VAtlTyxQ2LwmzQXKNKpZU7xlovMhF3CSwSMEwUNrBKP7rtLHAjab4+ctq6tLzHWzNMjSOfG/JCdyT9qI4dWjZpSy7egD6svG9Y8GDnEgO//CIUDP8Xux+4o/BocKuDXaP/pI262a8KJ7cgIhEt6WfCzhcjCFoguDmGbFSYg14hB0SipSEy7jiv0IBSAu91uXmobgqQRC1LpBE9aXNoJ8bmKG76h4ItatpjPduz/SEtIhRym9K8dr0DNC2RzkwBAX+GIzy+y6GNf31Wv6YUyvMMKLSwOZrxgG3YpJfQJADfapr0Z3ZgNYXIF3PZpJCPspQJKD0o+MnSi8pbP1rrC59WePBf+edmMnACJ4KO3jq0lZUaZAaNysXgMYA4bhxpM0gP0WkwKPhwetBAPX3/jbiBqrf48p/HlPtmMhnc95hoDwoLVDsIalmoxw31pfNNIFzmf4rNHx2ENvRf8n22nPkFhWQjsDl+QiaPNXaeWq9/yoolkIJV66CLEyjVl6uvy2a22RRP4XNY+3fHPuA7QrjGyIUdqKkE4uFfDDN2QkjVv/2+rYEe6yzbRT6n6SebXA4+Q/vJA8q5vEXXqTRAWJUnPwHtd5pmYl6ljvqkaC0GZzKrM9EwvAyo4MMyQXnFg6GXtmK0nOiiGDq/nmJsBZENdNiAoT5ExQlLUUcE6LdBTKdyAtvQjcmMWTMFDcZVD9omZId4WJ86LGk4hH54/hGGVz5iIPJXI1rX/6VLz3a+aWh8wuFIjoo9USR0t7mymrrQTx1qulmwIoBvr6SLAUlCCO9gyL+vBF3aAs/cxGSIcha/AcZ/P2JtPq+/v9y8n2nVJKUvzO5BFHbddkFharVxpygPmWLpSkxQ57ZOwB6ALt7YMvpX8DD/k+POivpslXFE1L1FsP2z/JHWLFztPxrCZj1KrT794pxdoaSLNZ24wfsVup0nYe/SFU0DWMo1TFoxwO7fU+FYXBYDn6J1SZ3qLA3RLbOJX3HoDUXsF0MIiaKKvh+TMQS5Ao8K+0gY=
`pragma protect end_data_block
`pragma protect digest_block
88b005d0acea7d9233c9404a9253324be9aef7a9377e40d32d965ef08b136309
`pragma protect end_digest_block
`pragma protect end_protected
