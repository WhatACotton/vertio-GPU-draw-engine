`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
f1Cd6Uoi/owqnuPaX4V91C42Bs93FnJZR6zAC4vAIDn6Q2W60Q9YUHuDvclhDFiCLC3kw7YAWKxl2YfqYV/lyu9l+Oy6HeWapQgcVVCEPRGLIznqm4AHsTcAKFWu0hdbCkbFq7w3c43NO8ecLQDk9nfqKBkfA0CJEZDaMI6ndHAhAk4F6o7Dxi2jEzfJHpssDYCCIlYnAyX/E0V7JpPB9Q0EQj9P+gfr8Z/ys4PSupyxfXSPgjIRzwOHE+mFCJYWBggywYLrjkY/JFAUV8BQtlm9ASROIjH2gn9DNQYTInKrNmBYG/pFE6N4PcS0rCVXa9nVrZMb9wP7DZwrdFoniMwG+pXECd79PV45/RZk4pNEpICiD6Ntc8O6R9tI2gn15EXZKyGDajL52jzq2p0C7AqINF0AXbcgTr4Y8k49t7/j3YFkNx5rlXTvceBNa5C1ejtRHAQfOLMaobr01Wewv+kk13lzSG8aulr+KnF9TVsrS3DWOlevNsVXSyx+NM2l2qJh7UMUXWgcS3hMyBit2HuCdBsYuSK7nB8iOUEUGsD5Ei6KG4wfm5sKOMo2p577Cz88jDrV3OA6Bg/v4k5baq1GayMVU2R2iovhNZogmxGv3qFlY42LOlHXpHGl/BvLDgPrVDwy73zG/NBFZlE+3NkOn1Bwde9kVVbIyK3GKcH2sJPZhGjdi9NOae7wm03FmRW/sKvNCwCdYlLucrsoQF6vLIs6U0QGaPcHytWUTC0TsG56mYP0Ej/jf0skwW4e6AOKYenhdCKeR5K3SmRwgROE/fAHuwVe4ckyBQqcW6mF+J+XaGEdj2a1T4edxb4LM1V1EHY2KzfiN3NBESxvWCe/gpW6roecHmg5r6MNyhc/wippRZy3/8zCokEyywXyLhuS8KAx4+P1VyrWiX+1/sFAckbrkPgHkRCSZHEBp+WLVyTfpQYAg8LlJp7ttFt+bhoKRGzvhLKWsXb0l6QL4Ns4FF69Trsvcp0eZzJQZYzaL/r+EGXyY4MYC2s5EEofTMRNqbjh1/Qi8Ml1PwSyHLw8axxhwlzo78agoRv5FtjTwbuAxrB30U6saNRtPIhTLHpSEUegcDYurq9Xj5Se6d2aa7LKMJPELi//cD5IJbeKSibh1Pyb6JwhNX4HYiQo2b8OQZ28HWFLcbbi2O/RgMZ2KAeU2CD6csdbCwEpnyazrOsdZ/0tOhH7pIEpTTSsZNNTtpXlnBbRU4iX2AijmVU6mujlPryZTmLQeUBOPzuzKLSwkbiuhW8gozB+3Xg3DF3PfG5dd3CDB2/c0J019DeiEb1Y9MkF5RW1w7mmAT/pGm4H2dUf/drUkyX6RmdFjf+y3bVUtvPyg3nwGrNNuT117iZVda11UuqAbT4vPQLBLO8g18CHK4MWMetCET2OTnAd7jGefFI7a8954OTzyPVc7jqBL7HhpDZFL43uua8GtTw2Dnb1CoeTUBs/M1xPAIPaJuMPszZlxJ6ZXjqOHqjQn9zLqYDZFuZZJIl1vYnFjt5/7EMQmR/TO6MqXwDZ9m+XlRbHADu+r1eLoeeAC2w6aG42B8xG4Lp/8RjVGsIcJdrxNofZopap9w4HmpqSFVex7wneXwFDakI1Kf/pArI2ABHvsWnaqF2rREsTndpXTAOXyGdm/MZhDABB7s3bIxOTxScjC62cJWbwoNgRVBTzwrHwgdGhG6ej6nOigw4hAIo+jpwQE2SmIIUB+g2IFH4YDef/pADdEdHJ5mE2bdQ54L2Zgj4oM3Z4ZM5q3CUBirMWdW4q3bDOAq7d7dc+3T/tIo88e+KjH8ZjU4hizlz/+tCEhMlbh8Wr/JFphEIrS2aBMCxjMG6FUjTXNF0smNr0rbhk/CGvBR8rI3ehILggdcFiBSBLJH9qJ03Fl7Q1B5mgu4hZYsvDCZxLmbRtGgc3/Cw8yqMehIgY2/juBrlOGLSdTKMrLD9Pl2vQUVTz4vv5HPr6KrQQ2OdPA5f53I6jwT9DZix+t7mLAks0VjNO8sYOdxUP+Limn/crRLOGtohdfbc4uzF6abOB6uL0B9V5FW1XS6NUdA7MNAsW0XqG3fpThR1BHRdQzuYBZHBUyIMV8lgGSV16k8MvrfryBIQD3VM828qVmD2xHMDE0W187sZOmyoVvqHDLOFwd6cjDUyB32QuH3bslVfKe9sG/lCk1OZ84NglzpC1ZL6r0yO8Ru06a+b/ysj/+c3iIbv72cEiwc5OEq/yyIvKwKsWHbiVNMxB/NZKMiVKkoby4oW5iCYEQDW2mGfl/8hEVAWocCZZH7apdiLI9bO/FTrko80pMeil9CH1LofQ8uk+1Lb+7S5hg4GvJ8CrD28oHZ/voNIHgenpl8gnToRMILzNdInT29GKzfrrthJBAYMP321wOdl4WEjydzDMVN8ryrKRlJaGfME0RvViGKqFIJRCfNViuiLVuvaN/HHCZrk5XvrRkI9UgXw+dtTFE0KixHTdNqdwInSWiLzD9Gn6oKkn+NFWlkQIITYLs35SGifdVQ6H3xH+p666XwrPIdlkSLe38c53eu6jYN6GHlXr5LlSJLStz8q5M7fGHU7j1A/upLQZgAw4NPVSbOjUlug/YS6qIZnSXHyK30rlz1zhjLAg5sqmBl4EaYBfaktdDR6H2TNwnK/WT8w/P6aQyX/CsjVpUcJ+szEKy2RoL3v7NDXVOPVIP5OFY5O6B5FQ5MgvmnBHNZTw5oSRFzBTkMuLT5Wx1hDRjhhrE1NV/NXWYawxB7Fza0A7LlRPhsOhc6XDKRjAEZdOOurKHwuGYeE3VBO1KXJByrPGaIiDdGyePCXzcr1tG/jX8ZD/6Zgt1C/WnM5XEhnCq7hHio/vP0tGc72svaMM2e46T5KQZ14iSCPwgdMNGPm7h2DJpCIomlqVbZmzcnFqTYDof41pvFy9V+XsouizHKZqJViFMmTJSweKgRREGJl/pAzxqZMgSDzfDewVMPPCUrC3KH4Vuzaf8AzKjkrv4gqjhsM48K6a7vHtEbNcOiLjfS9JRpVXLwVSnLJaV/QGHu9gVE1njDesqR1eXlHaq8cePCUjciWaqrxr4UgSzUuNB3HVmjwxKj0dpJtz9Qvk78+oRWM89b/ZqPq7hdkqKs4GlxYpKJQ9ofEyxEAz1ZXV1pldfVkE1wYoDXHLcwk/NDp+LIX+xytpO4p6QfvHOjSJWDn4+YZDHrSiNdulN7i6JGQL3N2B9biUXhsYV2vr3aj9gIRx8N+FeW/Ek00PCEIc7poNGLGuosXWYT1kHKS6hHwfJhIiKHIMRG2MheNFPcxUIVaCKmj259+jNO+vEUwCwCC1Ojg8YNqIZB8kxtAzw2dRheauTeFEEyIse+yXk4vwtZpYp2HwFo8Dw64aIOYyllVMCZDBB5Xij479w+9/cJlbpIIp+t9qt+v4xGX+NlTq426KOCH3pa8Rq+tm4OJzbmdu61vSv9Kigjz29k5GfC4bKdKrw/2pXP6/e5ayNlRcLEHtbW2HZRTxDN+RTuksKrO1r/kkXgC24srDEmAxORG7M1aEkapVGKe9MwC5n5M2eDww3oGbORjp7CdXCCAMAm6q5+cRmC1MabYpTFh5/v1vQpo78Pp+BILVOOq/WqTmX/p1pxa9Jgl095aWyQzkKiMoXFWReGCjyAvnjgJzw5stb6tKbk2PMTnyCZe/NekUxt8YDYujhUB9tFly9gQyvDGH0OWSxCgovSmFJxHtUH5F0PK6ZaigeBeQnHaqytoL3bcOm6XAgp3a0GO/yyyvAwcyUEwNSV6h3Ouf+UoSbR8UkzxEEC6VX7qMdzqrkkT34Bu/ZgGlAYe6tKq3BEnBaryumZ71vx5XmuUU5QW9wYA3sAxHNaSIcpLY/2LdXE1GBfxdwuz4F86dxr8RWsiP3M894K23tU+87qFUStvfSzqxlHEzPc9SCfGbH4xiTXvp4gp0d+EDam8xM72VLffk5vdJbq1LaIvSbnGCbbgwvu4X4nMT60pP6GqG1YZtaZdsEdaT8aweDwJembpzz1+2UbaPU5JnZYxYB2TD7Vl11Ei6aDpmeutAJ7kNJFn6sLnGdA90WEfrqoyhEk0W8rMW0mg0jI32V/9hgw+GNDQ9TmJpcibJkny/4hMDSAIGkbeqboJjiVo7y8Z8z64+tJXYxGsRSkiFwnVh3BQVJ1/WpoMt8nTIIcs6ITYQZtruxdRJ/ZfRpf6CQ3K7WszGHxuFa/VeOJR7t+aULqcVDt/bkhPCYH2iGknJoWRzIbCvWNDkvhd9iMUMAANnMSCG1wK4m1iYogIsDbrnvE7PjSGjGoBYg8DXZbK9qCmxlKLZONUI4R5H6uogMnVDox3O5T/+yli048NCxXxmU+hJnPeIUBt12WexO61MKz3haQ4GfVGNo8PDt7CNSj1nuMphWCfjp540nItTtJv6Nucxguglt1Ab8+O/Vn6wi+ZkJBT/OZgrm/MeHkXW4vZlkRhOC7JgkjkvKJ+qB5M0JSKmNj5BMnaLeI+8fXqs4FGnNXGxzSG+3ma3LOWJJOCMyl40b9oqjC3DAduE+IaIUXqNjlXvEjyyCPNhKD6LrcWfJlTerhHb+16cp1NTH1kOaMGG2wFmlOaZ4z3MO0fOctrjAuVg5w4+USK0smn+FUxPAdhp84mi0SvI//qCFUb0wdX8E4JKR+8DpEIaPgPmJE0UfiTiuEWTUUrc+ODhWN2mSVu4Q7MQ7/cckb6DggkXLJVoSjJxGzBEgo2wXObTjlzdJbzUnHQCgbSyzinjzOPBFLWbHhgpC3ddEkpD51OsPir8AQARwkyTLsicaMIpUiSSXHv+uKCmfXV478i8hBByS5aKhZ7UHdxZAxZKuCxry27zqMTl6W7geW6xM+AG35BKDQZ26gSrx6gml/Csfeqv5bR6o4nZd3drPvHq07MrZftM2ODXQwHLu5FakuWhpNGZCfHM0QizQ31gVBqzHuZmgqxaUKBFeU6DU7EfjU8wHceEwIG8UpSLtYNzldYgnRCpAtbO9TgOKgdSrBnBFInI+bQ6xS23q+tleEUsK5QqOTOPKzKwpdMRWiSrZnHXHGVfh37Fd03GN3E42s2iZP7P7z5N0bYCw2Lef95xDhy6HPJepwGl7Jsox7OR4+/YqmDAMmzKZFgpbGujFSGAQy+g8oRyKFAoQ15JfwFz1l041ROJtVqeR4tIuVS2VZifR4l0Tx+BHUtzsu5+boKJStK43GBW0nenMcEWqHVg7jBtr5QO6aUdHUfeOC8uyrUDe6U62LyIc2ZakJ9LOZ5wcE7jFWQTYsnl5x6bEzr/f0cNOVpoJvvMiKzUP5+asxa9h+Axd6155JFOZuuX4MD5HySPHNe4De4sGRfBcAAEhWmAc2AaAWv6UuzVYuDZsnnccaFtypNVCVmLLwCk1s66W3bTIidWxHMTAKUF4UnsFMgg8cp6lE2ridRLz6+Q5POowsoNI3VFkeJOVWEQQ9uHJAnBlBjSbmgmGKwkY9YsS+cSfX+T8wJ3RfEoJxg3kNEyHf3DfNCK1OmAx0bUP64hC+y3CBS7UQcDDRa8QMm1/HyHlY/kA7DmRxJHahVxR5AQKCLwJP74UQiAJQlUAniMaDdPAsUxriAocK3d3/FqoAulCoc4/sUgyBtVWBzPigHtpfAuyncDfOQ7x6vSsJ254zJIaj4kgPBP5E/mMEDi2S60bKNymEFwm10iRz3S4NWEfxrd03eDxTQPR9+51fg6phXLyZydYdmXuuawXEluJKtCbytB+z82aqeBnA8guqZJ2vp9DbWPbwue4xVtqTn5mObKTPrpTySuWLw8KDRCWC1GdKZy3v3cfCWR3QzWW+QcoI1ydlAKmY0UHHKW+7zJXOBHFqc0RSvL9CB1V7mZiTkYXGS5bFc99FzBC1grO3GWKVPUMJ54HjZu9rcKsaI1L3SNtSc6nTiT/A2KBsM8edCM0Cs4+aZ37yWgRpsv3Ph26cx3gOxHZaYtAm4KKDttTCI/PU7uggRd4DfhBjkQ121LjElIyuodPHbnt5wC7Z4OoiPVAYf0jfmAsxJWME/rCEqHr9xw4h4l8C9menh80iFLEJqRU6NmGxcpfsxmBnvgL/dC+nh0bfgUZKA7BTqTeKybD9rCr25JkMDVW7bHUHEk+50f3Y+YCUtp+PESGPDJpQ5kQ2qbtMYXM9n567bn7u+bvU7qm38QwVcRTEBrCDRjddexsWur5j5zxjKvY6h9AkZLQ4xrWsqRt6YF8vqoFtWi32vAIZM08bS5wqM6EKf2hmxSldr9jFeLKHBjw0mkvUqubl2mA5awY7bGlmjKJLQ4ppIqZFiUp/TIsWI4Pws170OEdB403sug6e6Oy1Lf5TQ2WaDdrSgOregDwi9zfkaANYKJBuQNCTXVWtJI00WY4TK4MT9re7z07btsomgQMcaioL/p8IoVP6yrVoLSvhIRVjFxJBaQS9u2RIOVzHFP0porqQLKhUkqKnugy6NIr/BDX8iDYHSry+MlJqBaKOtu4vUtzZ7e8Y+GcbGrzzpUBkzc9kcBAeX82TMUCJI3nPRyUMDCuNebuI9CHMiDHZ/45TZIH/RJy0+sePRh1HCBXjpgYEJw76isZ5kBudSWsML2++Fr1KGQAzZYdAPFEz8SR+2h7Bu1TMCMdcdR0wqmcX/GnLIZ2vRWkQSfoyb8LsCymVl6bgUMjpKItglfo+qHnl21Dg77BR17eeUBZkqf4xPjBhLP5ZGk312PGvG4PYSuF4fTPeMNCDby778GkFwoRIDY/uy8sfl4HD7Iv8oUxCVOqOBTP7YdFpnQQNWF4dIgegHKxPEIrx2doDuElosHW6x82onT21kped5IRaqk5Z+ZCLl0mxUGTkAwCDYjcvulAZEFuk2sH4yqWpgXbvWlhFMaDpBlO+zuMPKytLl3gi/ppycM1vrZXrLz+/xt6PWG56jxGIrCFeCAFaC5SjY+Z/q7fWDxqWKpNPK3uR4g7blxCp7trAFsOYxhaF7JvSUC/CLPyY5v5c90hW4skMDggdC9LkR6zDIj17APxdbgAgvXHVWRMcYPPN6CzyMUVcwu5yOCaw5lybskgt7AVFch9CxUaypBu35j2NBFBviW+y+qxjZIHx/IFMzn7nGbOEGXwtfwBraHbC6TabDeEYTzTlPR+ygNy4UGh0ha8tILua+KpFa1oROq/C8CHnUl4AyhGct4fRtovcwxu7pS9IDHhW6yWjfmhVp94DFuboQELZRUq0mB7cG2tPndQ8w4itXZHlo8rgTVFeFSY91NbPQNI7VItY2p30qmMegHpV4Z4PYexFLlrepz3vKfsn3y5vZb+hpVKWvvNzFcDzwgjujx0Ls+vHlWZQ/xQoXl/AZPSzfjo0KElUD7B+X/nw45qFOHfnLBoYy9kDkq+CNmcGdvD3W0wRE7WlAN73yjPKOgEo9mb0jlk6FU+t/Q2Zb5V9oaJgnCnLKcOlvonW8o4aGjnX2jNI19K+VIQyNnpmfLsTprkWXDryrwxmsGiGYYKIAkIFh2L4ZJXd+4OAHzUCcurIBwapEe+hgmO2lAwseOzmHSI7u4OPmbcmltBMc0wTKOedAFwEmt/sLMqEhumbF0ff43MGhYki8yVHCeBAMx0eEKPCuvMrPjOnaRAuiKXMLvtrTBQ0p7IpBH9KuWecw7uZ9CWt4X4UsGm9gwWkZUtkMnk+s5nbEbooyggUJd7UZssWIHeVfygbYlBHRSAfpRlt6SNtHQjhrsZYiLQaaC8fXGZu3iPlb5NQC5ePAnd+RH8RGWejj5XEsCNYRk08gfpcSfz/QBDvhOMSSlCvYK89oDGytpx8pWWEfWvK6Ach8lL/xdc3OlIXju6/gIKgv2IrYQj7qraXLXs3beE/iBFCB7RgjQe9v6DoK4d2no1o1cUJlulWh6MkTIAupRBBrz2+EUUHNslAUkGwTaUbxkO6lfdlmCYsu8q48BuPjtzE+9BMHUWP6RjB9M9W/OsMiWNHsX8zQi92OPZRUa0E1uPy49X8Dm6JiDNBK+g8cWgh3cJg5TJ/kAzIXq+0NNyiPFOtTM0jQAxgDhVdlrlcNA3O9bjLXtP1d5m9gECXUzEYYUqQqCT0nsZi0B+vFXA2lIt7LqrHF973L1N1G1XV7f7miShhyXhmx9REqAKZwiGUYyHxVelot0obpSREk+vYwuprSg7Fp/7YXsTS2BY474el55vmlu0RvGLe8JpPqunfstxMw00rP8K1rz6hGsOT3GTPgbUyw3t105N7qTbeg50Y/tQ8L7exY/4vEh1Rlu/I7MDju7P+xfW93BoYCVeYtfjAQtt2aVdsxag3qX9uaDMzGcKqgxw/jFUxc1E5+A9r2KI54JyByGFLSjbObSxQJOxT3+/BLsJcWOdUKRLMZH68zabRIVnctDDk5Scy6Oh3fRcH1TxjI5eDtxSLx1Qcau5JP4QOrSYPTJ+quT6a9r8NfWpR3LkuqDls6fU8qPZ5Pw5/rHShYjcqlE9mMjf+rIaykESROe3z7TJp5OFYLTmFqQQqqBDyr3uAMvMxuV2k9DVNh3FGdohlD+IgKfdwVoVIY9KugK+VWOimOSGwJlH5dp1dsMt9/FM5GRv8ol4gjvIeBKUmr7gAmezy0+E8nA78sTMQzHlp+g8o+ytGUFuAUCZ+hiRrBTSSKtrpwAmk85xtup2JAaj2tsZKJccEeb+/PwlC4sW0rTErclar5IJ57vFaMD/6LcjUXAlFffFCDYtW6telYkwbdAgfL6HljrcTMFOx7lWVcfhJUBlGD/fqMTK42rHkpP4WTf9n7GkprBAD356ceUwTm1JdwODNXpdhX6Tt2Wby5L+ti9mdeRujC3fJAvM0kOwOPdcKpz5s6BBqmriOCQP1Mu5qQ8MsHigCQOyBtbru0golH9MHvvsfmujM0si26BGYrEN93SnNlD9l3heE3Ap88wfSqrlSAir7IdYoSwduQpoQTsD8LGbxUupuNebMypqgT7sY0onNx3WKyqzFGivVRmLLdmK8s9NOvqmL5gY0z35Hz0lQ7bUxIop22HJTAPutCZA80XrNmuN8rS8q7QO25fs8gZAFzcnyB3mIM3/lSJlglGySN8urd+QjbGnJwNpwnFWIM1A3yTGJC69IYOnmz6uorA7/fOFH8AdGdXlmN8617pp2LPzY1WuZn4Cp9pqMyDvNx4NHkrZ9wrtmnNMmE14E2w5ajka4ZPyZf4VX+yg75wJLzhVoyPfvuGw0clBGsSeEtPx86CUMwOhWdqLtWSfLM/moY/Qoa5F1jXcLp59KTDPilb0mpYRRTOib4xenOQWPkH8yy9uA61JwekeBqbJ8TQZN2Gm3tbgmyomREoOnQ7tbGKFpGM4qj/ibF27fJi9Pj1wJqATQcZ8OBKcPNeG1IDjygZNK4BGXwR75Eop9DrCCYuM0X1ipwCWpd3XcCiItNK9XHfQoRqCShZ064Y9/MRsoLt2cVadpIPN5gH0MFKQYp4hM3zQtXPtZGl5aioJ69e6d2HlIlxl88nFfdBtIlaHJJQVm593McKCKUjadj9ANNcIftLFKgL+M/rlYuE2ygv/uDHc6bkX9y2wmFrD//+ufAY190rjFZr4XUIM9kaZVwuSec1ZKV3ujpLJQnRqXxK0+yM8ivUmgzUcQ43Z9kRVxMKCYA9nJSrPasIC9KRahLESEtzi6i7aPkeimr/8aYFSf+bY0ZeeiQlY/F0EHETdK6YuTNMGr0+vjGBAzkRWQsEFJiCy44/6AvZrvm4fdL6ic0wYcKgdZitdGlDW1n2NjBZM+JTts52/dht4eJxt9TcznpMfdLeNBkN9cbB5Zf955XMne0YzfKmcpIL0EqXkEdMWFzttzePbyTfVZ8r4bVlfPdYFSfK2ms9WHosqVq/anfCppq1h+mbpqtRV62EhZ97uFNYpELSmewzhOkXb/YZ85RVEfdZ2tOMA8qw3fyPLGIdfYoHhqNjm8k40sxN+4c+aYAEy1DhBHDJfF5mlxcv+uMiU7knCojzAYfxqhVBUE8X4KsNnzOLCBgnhrxUIMSZy70jRZhv9r65osEW+fsOvY5Tp5UOexhevgiwxKmM5zAMb52yS8gNGHWG8m2naFx1LroM/rXDNkNpUA/WjEzzqzr0PRFzfqsGRs3LO3XPmhCE7dwL+rYRpphh5iuzTdZckWDtQVX6eStxnSSCBN6bTVi5diu1/YK2U53dcXL0o6z4Uf7QrV34Ga2I6vabJ15EPEhx0AzQGDjus8I28JeYyCg2VGxTkOYbWPxJ0aOVusugiUchuCLA/H/8cZpET5W4JAKY8nvfSjg90+k0Mj4BIEqXc56RlMr6s0HGT3UFF43iM9ZhKDomkUNBhCSeVFy7AAEledeRjqpzkAR9mZ2ZPhCtZwWVVhibjEprq2XbRFlIqafW12TFOIE0GVcjdZeaEoyelRILgzsmGBx4Jr7+fjLNvi+SR9yMSCWuYltMQHO4+6EAu40NXMPW+Ldr6J1T+yLzKPqIQhwBLtogSQhrPrJTbxFW8L9ImCscfNh6bbsqqnCGYwdZrMMg98PTgAWPqQOsdWxsKExJzAfZW+UpPz+OOe/rWO7AVTFftOhWCrOJssqPplCf2N/D45JGOt40+/rKHN8N0KDAPu9Z7HqEIaXopU2isFEmPM0jr28/UP6Uf6EIIZfBeYGf+Bbt4Km0Cv1F9a5VUEKUMkoREejB92zg/1yhb4i1IwvVWJZis+D8GmaBy3tEPabRQtRoYYY9LuQ1sdeyLWwAKMKx0JRTjz8CdEl/tjAtL7mtgvVcO6m8AIN1BHjjJ65DZYfjFT7WspOnpl44wA5rER3A6km/6u+jPad7la+esQTDBwl1jFQxCHI3mOC4SMAQbs4uTm/iF5JUm4/qNXx1G9Al4BJ7pZCf4eQLF5ibOEGhE357YWGWfuVVung4p4ZCiPzmecy1+OAJdderMo61b0S3Yd673nBGnH1CW17Vb/ZB2Dwk/JyLUbxHkCtSV1G9ha/dKmnCxBrveaaG/svAlDbwk/OgPzWiUajtm1uIwKzP20s3qnpN7zEPqGY8VC8SWjlq10rgSDVnfARR5LECVa3BEMoTFEHpoiTrDtYeMoWl6sOYTJx+DTcZ1WEsLskSDNcw4SnL+W7TD4dlyau0GkB12JEFWKEyau/NdcyiPfbVdYf93djzeHZBYRciqKi1gqr7QrY3Oayi/i6qWmEjDcqSgSWeIThI6MhPVX3yDNY4XSm7lGcojrUEsiLFUKftcPc/qAaFviXzTguzf5b5Ou6eqAzVxQrmP6GKUcY/N4LC0FiNFaT75IRTZ2qqVJt6i+MRtkLPKc4yDeId289Klw3+6IGCuA9G7KOW4R3SaTc9NmbPQ6taGicknroB6NmjBV5ZjCUcuAy0bYoZZIXn5BMMgLp8EDPVX4wsLP3SGylMGa9fRg7w+uz/NuaFvatqyDMeUVDy5BY+s0Ehb8LnN6qwXscszMrMOOPaX4euS/FLOUic3BxZCYI2vowdSTgHoy7IQsRqBpMU3BkkLqSOV1AWh+WuzAfAibMfeK3wSvj5HIPlmrCfmjafQz/5nWK4vFbXn+FdtTCUnmPG0Y3V2qaGvf8DNvq7FcBVIj2orz+mM6xT2pBjJuY8h9/t0On/CPOd7J7QCdymKefaGy1tNEMJnA9Nadx8DXzdXEoCukenBnXQWop4YO13+DgpdomLDRk5IZ3IFZxbJnvzbNdUJahKb3jj1CS1SX/Y20thxf9FZoUcqpNMMo/gBn8nZgfVtWAxjUlPhkVgB45OOnV+NCu97MyNUQcuc6j6GIp8ByGW8SwuA95JDaageM+tM/lbJCJ26QLMvpdvztTqOGN3EvIFUMZswCYytLnk+THUTQGbgRdvmmLIYdlgzvc7FuwGA8WCvD6mD7s0pOG/33Hp269kJ1Dmq1eVb0KL1o/BSGhJ3W/DBeH/tms018anSgEYnH0NwPwjm1eRt71RHzEsgHCxV3qmvrxslXYDhmGBNIY8nX1QbAHpdwVaPdYjb3Mih3YL2pm+giINvH8RRCPXH61N46XzJs3ppTj7hfiXic11aeTYOaWWeg2M0DbJGClald2hMhkjONQqcTU4IzZCDyAghJ2CkpPhG8HPCRRVtHOgn0SuVgjWGRPQItKMZFylzQ7RrkxUwU1u3h9Fhz7ADDZXefztYi3jfHzfafm87qqTm7GrblW8ILVBjz+Hy/iiqBFVJ2AZSgNg4umLmhTxiL1f+70pQ7UdtDxgvCTeH6op/jtcTHcW+zzuncROvyZL/grS3Q4/W9EftMVx9g+st2k/QDMVanXHvYZyaj6xTXXQxNaa3hhXRKptKRQRnQfS2GulCUb38gZDZHPwhnIBAYn/aFSZyOtCyP/tdeWDoTRhSSLiFwUEKXSTmbar3V92utnY5bLSDyUQM+ZyrN4O5P7VIqxAABIts5/2DQwO+hGZZWIqReG6BtyhKciCPnZHEmrtXcY9U6k2JBwcyy4wsb1sQ/s2nzx/OWF1oiw5dqVClI7QjzhcWg2IkltfkcQmtVOD1ZFa8b5XTFbTfxSv7KXvXeRl1VSvO3Z4pz7lQ9PTP/4M3ApYvxPpKC7g5Pl9hNNy5MDsElavGptm1CdBsZDuv69XcLS378DdjNLZYxyzx/kOdeubdX5TCBDFc3VjhdD2wrtnxGPg5gfgLQSJkRoucvfiKgctLyDL09YCUzJFTHQvlqYuN2fCzqZZxU5zhFbR4zkebB+dVx5R/5noFv0EjreOE9+64PwMMeeFgYzoOxy8l9pobO2H5Ud3BRFu2QK919OhaoHj5ZA03lOmlbYY1Clh2eot7smubDJIZgLc3kBLa58CGRGisH+sLLEhe9gMoJqO9Xz1VeRpve/b+G6UhCu8rux95RSNVH23hA4OwEJcvSNPw6w580T85PF6XKlNzPMyGSPBAMxdMb0y2Shz+7PYUaznrURk9pvnx1f1F8Ngv/Ee6EPq2ebSaFgmRTSU3M1orbkPuECf7ToztWD+su9S+SVjsMtc940yS0nsvexY8p8maVUxz1qB+xzp9sCzmj5l7M32bglsgpwQ8rPdR5J/W62mObbd5kLpmPulIKxGD2GOkhjtvXDRrveFxNDJAd8ObbCTyrWdHv/GROAI/3xKADYiX5HDLTkX5L8cF+LIn6dGzbhbzfeqisM2b4UFSkCybdr/3vyJ7f4ve8Wjz1+RWhRYO/PMP7ZUcewNb+1qdZyfe/nWcziZdrLL1AsR6cU3OU753NjRF9IS1ZSfD8+Ryb29y5iKZUtqFu4Qjm1yQoLZyxsKuPSePArm5IRGQSp3muaZqfcQtJLaa1Vn7sw6Aj9bMhi/3fNo+z+TBYM2+7DPL6iwjZ4bgQ0dI35u/lPoaR/okl4Cmz2T+iKOtf5FnBhWqfWrPy2oT3Lwz4VV6mp3LEGT7FAMMf3tALwg1hQDNoIY4+U/PaycXp0je95ciJkDELo8zg2jX1YI9VjbnE3s3AGasI4VRxFfAY80YGSwlXPu7EeQMnr1sbn181x8EeDghEiJBQVyydMLEDFoZ3ITkFNrD4Ifi4QLk9bLMhUeABZ04VI22cAz1RD+CB4KIQY89y8P9gfWDTk1v25ZwWcJh2nyoC9GxhUMo6H53dkUyE2vTxmRaSWInBYG1siuWQtV1lVWqKDx6KP5E7RpMZ7otfAyGhye/+8fsEy58Q1g+Ny7zK5NSTqPpSW31BHUpyxovyKRgInagKVX9VghPgcq6zeX/XMTlXUwl3nREzYd8mPUtUIK2z6zt0gDKR5dUdjkFv15DcVqspzwOAQeAHbWD9av2DmFWA7JlkAVVouDwLTgXAl01/HtVu14FFzGGdppWKZuh/RQjRiCRcrj8mHmycJLsCGZPbXDgwbOefU2hI2dNQSqTgWhilonv4NUXRyOCpIGHJ1Jnlw97WwNczDG9G3zGOwrMFnPr9e8xZ4TtLKkeo/GivzgrfDB2tj1ko2fgExgYmJek7+du1BXInD3Vp3YkBog6wa2NPOJADF41gDdc3ei6vG2IUDS7AqI+ckaNhCvqp2toYXMZJRPWNpBy68pzkYRsngzazcLmDdodSKJGW1TyZBPo2bDTbyv2q7eHl7Hl7MU521W0N6hhFdEViGcb23zmokIdh1WmU43bDj1OSMn+JINHt6PlyNmo6NjXPyK+WZ7fC/ydU1aRBuXULTAdFprpUqyI6X3GmU14iZLiCYapiDubc8T8+X17Y83gCK9MVhTNFaBgLR1NjcnOIxeI6emViIXa21RWuZLPLYd75MgJP/t8UChqkFRMSsslbXgsTI0vWOrcZlsTomlOO6O+cC8qehfkzh/zgc3q4/Y3Pzfer+JsXl3J87P+7MDVe1Mthf7a3tblI0rgx0a+Vdly6xWu9RCZvUwMrDWzdg63///1zxu3AOXj8HvW/irtjwbuYP/FUB55GnlZMTnTbceEC4bRhKoO6ZBcpEliQPb9an9SA/I2MU4e8Ku7nWvdQcxhR64lcaWJcyMxPo1+Mju/nYYVFxHSC9Glr7SvbEviDZJR5SWx3jn+LPWIk5sfVQAMcZm49fAVGTEBHn7KG8LpEWRVkYltohOz8KakDOqho9vH/OXzOIZVISwveJ8+GamKFKImlFM3h1C6P6ZBNJ2e/lPbOEz8O7kfrpsWaeDzRpBhGaGNNm22Cgh/ZDK32Vb/OUpDtd9d2FG3t5lYN+M3jLDSyD/FlWGZh2f5s8bl+fJaWZ2ESCdqs1ZGV/5gmDvp6fqIxVpD/z1FEuNhNaFljT4Fh/DghXMi4G9mdx65aXUVwPjKrJZrRwuPtLuNTMnaErcIXQMIX0kgxi4/TzlAimCVvZOPOieQhIan7MHWzmUdwsGK7PxSQu9LFDrL9bfedIz6IdrJU9kFLw+Ol2j4TB1Vdz2/rIqgx8RkI+QzyWwfamkB/3raKnl7oEDObqX1Y6zZs46QY03qI7WzqTJO+U7NvONCSPNYr2NLkoRdA+N1NEbF+vr5IwdC648VVEjxGS3soUCGyE040ctX7HYGRyZIWSL5v2jyRWPPjoE4wBdflkcKYhec1G9fhEF5ROGZKyOs49zmAhieKq2kc5lKcDmYmYGNdaFncf1S+6/diFu6bflCLswx41jJJfch2wlsFBd7zO12I7GKwAV/+BG/n8ZECVDAU7rLfAjZP15mAWF+oNOThmog0QwTbYtn51IFbJFBF4Dlsg/opk2GKNXHReL9W7QnngDfZ/3lma8VxsR79rhZgxUr64lWGfghtgjsQMNl3EaGl+ZyDk3QTzte6Sw5NNYHZpurRqRge4SEsbPVPYgMnxej4ao2OlIfJLwLqQ4XF89OqvRyuKvBi0iSUAfgvadgNJoJeIc8D/hBo1Ozmsjydshbq7kMnEd4NPr+IfH2KKrnkC17BZWYnGn8koAuaYhjtw/PxyfKGOOy6/9QxHELGwBlzBmBF2PM7yRLhhV9hbl0TE5dnBEN9VDLHcVvsz9Juh3x1PshnaVGitUfR4Nj7TX5qhbgtRFa06o2lF7y1y6fW0ZDSFDT0mqNiieRCCGbEaT5zUYXtn03c5idIqrvRGoHK11HJ/BbVYKovOwAUzJEMxSQfdox0Fztai5i28wwzdyAvyg9JW0rfbyHLhu0VRLy6hU3ukBSfu4AdKIb2+sQHAuzELwjiNQPXSrd7aiGIXr+7LrY93lcmjf7ktM9gnpVS5G0C5Z5UhyXLg1sl+iA3XLglLyL+zLvgGymMpSx13H94VWlk3F2isEzXivWGU2JXDLhg4nDJnHQINFDmTMY9csSRE3s8IjivmV60YlLXU8MTWCnIJpM4JV+PB+yKLVWrxfGHFLzmXNShq24zog8TMJIsSgTLX+8h701S1usFsg3BSyOiHzqI+l/yxulH1LfjThUixN0ulsbRDbhHCfPqBxl0FB8RH2AYYB2h2TsTaWhItBQpkDI8Jb6WhqZj58PIvkFVdE+4Td1EYJb+siq+q25zW8cXQX+SDZ4U3K0p5TDr1V0r9btgB1YuqStPDQeSB+mTtMacbEzJWwAExBkNOixZOU6BwhPj3yLsBtJa9lK/6suQ4r5VJezrvQlr/HPCj18fIhgH8GMz7sE9DjSz1G8JdOXdXBWKEINgnhk8gl4pZhSOX1BVaF2xzq+xi6k03cxP5K4jcC4HQprMDSz05W02VyUj7hI65i65G1mhiYnHxht7MlA3lUcP88VivxyR/85JbpENjd30xg5VnplZ3yTIojhDBrBVHa1a2vhf3cbsT4UgTbcE/nuyfDGcHmpf7p88pw/wBikieh5GzICz6QB5Kyh1jp6bficRMmnx9ltwOaNPQW7T/sYlK5wnMLD0YFSe1jnyXmK6dy6wH4h3A50COfJKRh4/3NFQJE3/GY9tjrvXf4t/RvPcCQ63lBBzDke1BPlqXP+2Bd7aAxvJ6jeSGMY06iakRIobJGnvN0EAJDSrSsVEaicPsyuJTIQo0iQ6pW9gq2FF2vHC3mtC0LjW44x6qPKjo8MbyyHKqkiqahjrHjzrWazfWQuTnqWM037gBLl20f6rFKiV8sCu+veT7RfjrEOBILuKOhqnBeBcxyLhXYoZ2dz5SIU8MCGGvVQCIG+6/QG6ClTjZ3hoP3onTmodsiFYBvkb9YEwgcHhO66NRVeeI8tSd/VAX8/asBMRuYIzcXe2tC50YAVDM1YQrh0WxLdgBw95IVf5HMqLow+/n2NEyOL3bUqIqXoTmJ14Pfxq5lFUEj34NRci3ng5N2SQ4DCsdwwjlRoZCCn9Ht9wijChLASqVVK2ctrUuK1HeN3FPxLyeGd6eVBmGhw9xCbbKgrjBr8BEM1zQ5n9jn/8ws39/8VqPGw+a+fiopUW1DPI5/KYnwh2Vi8bFCsWUc/vT/iQsnAiVdRfIBNZ5sjtEM67wz0bEMBNgTXt8hAZ9ED/1YyavLCtcwAllSB+ndKdwkBQq/e03J7ug8LAliRp1ji20fastgSlpVw2H80LtNqu2LAwXbx6JnzpK3Kwz0cMvhsQ8kmsCrLhd3jfmd3kOg/54X/1xM9V0zYp4qEwvr3dHlagg6yKMJU0sPzlm98oXBHfZv+UJqprGIaqLy8T90DbtEPeW9T6dpH7qAT5V+Z0ioHeETmGqhKv1v48ZD1em9h4tnIsf8bA56gKzhx0+3Oax0bmtp8w2ejnnn4zTqdHUjiAzvBT4hWJX5sAYpJt9Hu14VT7wh/8s/0GQp4xBIwR0lVW5YdDNZsE1xRSWPZONTxB4rjCOyIaSZ5Q8WkyIx70mMW9Ie4faH6ITNmlC4jdH9fVInLgvdylcRI6fOdYbj1WFC3YaUmKVg7nJYU5BttSDnX+6UHDg3N0xNc+EWgkB4SyqgtKed+u56waoCQMu/sKVP3iVSVLyhR0odzCB4aS8pPdZup4n0jp/07UDcPNG1FMTdQC5mtXnrzuOfqB4fVwf3zcjKmXNVu5KTcgoCSMcaeByBA1rxmjm6hhwuRpkePDPLX085naFtHcvtV3b/mcbamCdh8Vhj0mty7OjJulp++94d81eR1dXSdIOK5utlgBekToVM3zo+1RAcQrRMEOkrAC8nxnK7Jh/6sSqGrSe2XPfsnsWZnkbW3GLrk/IWjoLC/zUJSjSRSQ3oDcw9pUAYuo5blfpCwAPPeeATUm4PUhZXhho79c9j8bvBgKMgGSh/oN0J9AExJl/Y8JOF4AvpoJajWLLWveIlTPXna12+YKYatRbxA/HLgyZsurPkeAkNWuOnj4pf3l+5dkGSEzFLw1lxpyyFcIwCjpxoweYzRrpBryPtqvgy0AW85Py8OWUucpMXQ49leAIbRxwIxjtkvvg64nzQNVTILxAY7fIn6y75TOU4qfWn5DgP2ewo75KPfjcssO4pDSlSmKR4ovNZvOENBtsqdrRSNCDkqySsTpnfMvXYFGuhkUljGc6IhqJJ8RLUz0XCReTFMEQgGJF9E3kUk7sx0lTjO9wpPXCOYiR507bofegVKn0w0Fcrl8+hojulCentkt0EiNqo5l2lERjMH+tbFIcDzNSrDd8z5cGoU9WqOfETxB3FpPVqhwNBs3xkaRHNGsLe6wUlb6XbHkUB9XTfkirRH+zocJ2Z4/r1zDXLwL21FOL1tkKS4b0dr8/RLC5YK/tV+7IocuhGBPSK8/1XQMjHWT8M+eIWeINxlJuC5F44d+bIjoXIOkR9+b6HOvqI9qEj8vfZDgyJUIZ9xfVc0+yn0dNilh2e6ir8xtjYQB/Kb6WmECPB8eF2o3Erixe/osd/ViGCFbIiMrtNI5wTyP6FUGn53qXM7KwoHdj4MUHP3tV6MYIkMCPvSVM/WdNJyQeNvNQa8dc2CmK7JE+14tuegcHejgchYq4UAkwPULpcPAVsACHn46P3K5UdH2P9/Z9xg0nhOfVVsCX3OK1HYLqoKWmFrV0lI4If5gbuDQEM2ebo1wknHJ5t53xnw/VPkFi/RBgd9SgxqjifdoZbbAffs0ABUUIGTXnNydcs+sBRLCgATm+Y2BtDtmdBTpKytt0yhkVipm/919wFxZLPLu174NIKsacQnlt84LfjN1UOyUCjQEVdinJ7j/oxOpIDBV3tAlR8XXvQhBY/aCA+LR8q2aUkuczHd8ybJeWxphJusTQbfUkFZCW21w3MV4pMjtV/k7gvvzHt2Nd33i7lCR7vzZpBqOY2Imxi4pc40PKugsJezrb4Mjoi4ehrDli0BkgS2LcCLWpJYmARid79jbc21EeRA9ljwnJjk+KhTlPPM1OWcI4clSWQwCuZnfqc6ClRbJe/q3YlKaFZV3Umbob8jRRmRbbTMeEw/SW8F57SLF1RPEvDaEj9ozPXEyY1z93HnXxoxMOQXmBN8uaXwO2QwRXV1dIxGNdp87NSELWG+n5wiaH55gMcr0+WXDt+NcPg75qYEbeuYTKCXevF+3atfgQimUM9de9LMaA7fZDXoTm/zW2edYOyikiy39UIjeqTU+lL/bbji2tax9kK7LSdk4CeG/3L7qliH4yyOlcqk1xV86g8fPbTxve5a6vdGv90pDNio4ni/2dJNj8poS6SA0pWMrnbWftlVNXEvwtjtF07VD6JJ6STTfPXPVUmPQfiKET1WfjS+V679ubdVLxNcWXh7ePWigsCUJZBrSG38YOYQVC9n9iXW0LFAFt90+NioE05K4aTny2ym1O0rB9T87T7rJV+eQPKZZbnIRZxtlLk76orQd48RwX+CIqmk/qvcZcUeopBcbcTJrYIuBxPDC/jZDXYB2+ZK2srbS5IrwyhMVVp4ONvZidtT6neHtNQ/eMiICAzykuuUFvrl7pO8WJ0ZIxjcxc7pju455zmoulYLmzZJ7v9Qbr73NivJIBRk6exYj50pVh5huBf+LU5DfJ5QazMKyJBIchXgdYls/5J283GCzAI+xCCkxOv2YdwsYV1W0SlB20Sor2MRDm1IjEUkX4xJxoVvld9XYHz/rrVo0Es8S0aTdsnAK3hQeJ8YTk4JCXXzghcxsYRrvKBrFLrZRvllBpSc+nDWBcPggOJ+tIoDNx7v++UkV1r2/eJftRutcj7AKEs1JxkWOSNUdBcBgJLVlhb1R7VptPPzbQ3K1vnZxvEZ2hSSQs9dw0vC0PQpZ3umXNLl/rWWsFHSbkghRwZq4yhB+9pSAK9UPiHWdgmS6TVjVFgRVEwriJhzSyXn3lbSE6+WtNfMu95+x7rLzRGF0wBtz8a0rhxR++KNj7y3tU+yZGKJBeMUVLuIzPwgYQQSMxN4I1eM0gdBjmphv8wRYTH9Tus4AN3fAdHzqUVPWmRDmdF7LSz5a1A0ntT3/kKTxb8dcJP8LEQS6C/HZjBet9qVNXv9Kdb8x0cqth7AuQOhkFoDOdvaRwMlm7lj4var5D2wvYKd0fzq23jVhr4D01Hpu+uCANvkE3IPkhK0NQ02dk6CaqJjcrNiApmVDqMQV4vvv89TICB+9Jm8YfOVX3T8wwU8k/88id3EHiJhG30MN6coP2iWclytDQ1b7dy1VP5cYZFqxqLkG5mGykn/TR2AHVZi8+eyUXqiV9ikJVfkQpeQ+ihAPHt7536hGHZ3HCC16b4Uqr9ueXp/j1DwSTnzhZevF7Vga/ydvI5eJr5Kh6pg43NgtVgmEfPkV7OuVKmmxQQvk8VdRItp1poFwQWVXlgxTqP4mjAPNacmNTL79wYbhwEGl59R3/0VXhDIsD1NGOWq0bXvQjeJDlsViLx3PNwzj3s/S+aCkeFpb6J8gYMTKqLcE2wg/nao97d4wqjxotNxoKYNj0osHno+IjZVrZaumuibVEVJZG688mWZhrGk7+tS1mIMTxviVwzyWMUWKHXUrBnKH/o7Zn7LiKGGDBXWNs2URae8Amxqeifm2zKbHSayktF+xvPwYOiSanQwR3EvSFNdqMhEBK8YZOM8+6vQ0Ud2zwk51JLvOkuQWtBVSIQwLRiwNxv7WqjyEe9Dcrpjjubndxfp40rJqqH/OTMYdgcMQDhJn3pkEGTsoq+m1gj8t3EJas9LUgiSM0J4myaq0WgsSV0X0/qEclxJmh17CLVJwjknb1rBww0iyJ9/N1DThqdqIC2ayolnktN3aJ2pNipXk9X/Jgs+SkjVLa2GTRM2LCu0xqkPSy0tOSgmqRGIQEjk5cCnM2Z1wkTWFSzBawY1drTguRZD+rD1IAGudbf99px3GcaAhTJe+a2+pJloJ1u3N9iP+o8T6vlEdL7BzDFnVfutOn3GZ6l+BWVZhp8HMy3Fdo93I0Q0rHlQkrCzOr7D96NCAOhZdOqbPbQbQIKsgTrrloCuSl6oqX57GsUwo3wMN1iht9fjIe3kd3WDKUyIzdvIITswyvrfuD9pD1Rh1UPsz15sghUqlXcM3OyPluyZVUU/9LElEFBOyWiR1dD6PikHslt8w7/fD//TtDCwLVoTKVkrRCf4DliUqVqVhejMIvVDCboXU5/Amf5R6tEMGs0CKB0ZuLISZzm1RcHVPyv4IhjTtxI5ldwTA/vR95IOtRketyh3nXQIal84TxqrvPFbd/uoltSEygHjcQ6q/9zQHCNjD8T0cQWoT8Tdxv6h19ZGwd8GChC41dF6csfmlWs/iq4w+cH/1L90BRxkB3opMY0QBvFETrQMkEFilq50mKB+997qJvDSnQKiVBpkmgn9A/2w22VbKFV1Pa1r5ko8IoudJWju0dhXxLnpHtgXg1irx/7BslBVhIBH3vjox7/gdj76Vj5irrEHsDJLQojHcF0XWyWdJBSeEeDdizPwmip4l2c7cqiLtKw6vsYvhMvg5bAdqIwz7rzv26ZVoF9J9QGagqINoFyLKdUahY9kzfhf36NNhdvVt1QLeWti78zi7FlznnLVoSKyvBbPxOL+QpOjhkzZOOfYmMKI5VH7BXqQ5FJWf41snVJ4g32GNnTeSrZ+IXSw35furW+kuY5jeQ9OknR/5gkuh7w/XH+GlIKYyOIqIxk/6eciD+Ka5kww5EVn6D58NqLwRaqJil9rRGf+mnh9/zjod+eUqZlIIw1bHJnpsUz501exHV7AUEVLf5qAGowlW+pbA6+my9zUFf9ZDPfwunFQEB1E7w9JTuNsNCsULEkcQR7nkqMm0ZLzWFbBovahDbGKsU/P9O5SjFmI+z7Jvf8c7ul+KKIrEzcXEj8SCckp0/f14zXLeepFR4bZMb3IspxNPgrVKC9kr1QSfCaoTk+pAgpuQ8CU+rJKZGp/W0683WgrhPVnOgV2iPYIhJy14+ikHEiifsQ0yBoXspfqtYIvaYnTdCheur7IJ80crY/lfvBZFcG0swsFE8n5GVyZqo4QmgPbQoDT5ymaVRogFXyIrfCO07B9kCIdC3gGjENHQ9DoyQOZQwNkxtMCQR4fstBN/Q89vjaea+sDFgVkkgk9dBZN5Mg2OaTIoY7pK9x26wZb74x5rBYIJuop85PXaQT3TnaEPX7eeMCuTCICAmJLpmPycWy1kR/HygKMVj0eLPnFyXg/fMsgiwlRo9c+nc0ykbw6lsIVxMQ1pnfI1TQGHuCWhbh4+4xDFIoNwOVK0xdQOzW5RF50Xdz64jGFMH1pEpyJsiOx2Ih6qGGSlP27SMawokKj2U8j8CIz8DoDrJAFQB9PeDQ9eTZyn5vHQ6S/MUQGey46xaXQCdH6Erg2Bw+kw0y5hA9KVecTg4Xyb8i2+oWIxU7mulpJ2cLXtTnav2Abkpcz8CWMhjg6/Es2ak8YOIRrgwKCXxVYL1SY4WHbt3FcpEm6jkjZpJNqMuQ44+MMU1RHaqYUJJZED0fK/4Zl5uGWpzcBtgVnV+FP+r7+GL/7m8Sk1M5hJqi0z3QHJaOQyom8uU6nzYc1Qexdx/+rwLezEcVkcD/iW+BcLCd/e07JPL4G0GVYWQ16mgPZmwpTaem5GZFQamHTUPWTC17s+2iVEBNPc5/hHALTBqg70qr5QyJJFP69CjsTF1y+XZDtr8JCZOZsIWxd3jBYMJxqSjjRhkNx8sPow3trTUtj6EGsrbdPibBhpwyhZrte+TOb8WPRS1WuvYYEwJCuBXxx8tcL8mXpVqs5HtXgmtspT3YmSwEVrkRPv1D333jR+4avAM9HqgxmXCRUG9oQK42RKpd2zPbCAQmSusoodORcVsMZqTPJHXPb64JtwyGXxjWALv+U4zebwhggPyxy8l9OIzDpHQ8SD9fwlcbh4KozXm1ZsAy0J9d/Winj0SOLVly7S989aM0QNXfBhgjtRZ82T5pP7oYKOglLdbOLerrwHMMbOVDUJ24+68UXVKNIn4M06hdTdTD/B1W0riTjkvV8wuHDN2HsCnsdU+IrS9XoAYAzcsL2sRh53j33TO1BufWB/goBU7cRhPvfNuDOPgbrIWwZtx45czHtrpngTQGcnLkYnwNsvIBZK9RRtBB69QZN5/TiZzZZhMKwKORXBRNBnBKIZmRTOq5+HmgfvkgP8frkNB4AVIsR5Bx+IJVxh9y+jaeufvnDCIzkkwHtcoUSzaRiMVN4nSElaC746ddztt+F5OnC/WnwCKgycKYBDz3rdXKJBA8Pfi5j/DkIsNuJZgIZajm2iWfiXO+lWq1KeBTivY38lhkoDhFGsk/JI5a2tbmUs1SyNvdicDD8hAZMLIBvBF/DE15MZhDFJAMoAx3HcCGvSLuNDA815eZA9zY2f90bVu4j7TQRimJXP3sszTe4FrT5xTxfAeE49bE7IRZ9enlpUkecr1FDiPQsvrvSfZvuU79MDzyBhPumx4o9p06+bjikR3zJozfB1tGpuQGmqG+vqCeIJAQF8DAS8hC8rRxnBRaTtLj+ccvJd5QnaPSxUDa1inNIX41gq1y1HbKeXWX7QrrGpdjJpOsHfcCQZ71JEjxfnoFIofeXAMCCso9YLqKAIrwCg70QvbdK/8qWekhYEPbOdDhONdqjyZzUMsQ2ILKtG6UjMYQ5C7Q4SjKQyt/2/R3/G0gqko2b/zBDkkrKM2zabu8cG+yh+cQ0Mfrwd6gJtsJlrvFTTmXxPEYLLbUT1buQyRuOmLSmWOd/V0B+PsxIcsIJRqH9w//TevQRY4Qtw45YxpToWpWsKUVg5YnF4ScGm58pJNCfO64MvagdNF8P51865gvaN29hmckBgWPSEqD9+RWB8u+xJsac5l8Fo7qxHcsVrNlJ3hCysZUaGXOsMA6VhWJCXtI/MUqGDxBA9iFvazfnBDeFESmLf/7SS1oiIzs2KO1gNJ8N7zFJRGdCM23VX72/uGx4p+AuPopWON4l5V+i0rYrMAbKblGIdIsubL1Ktg0voDnUWaKt2dCM4ygjGlPVqfCaTIjaq7RAmBifrvcmIPtfXdaukqfM6FzwQc38ssZYg4yYNht7m0HZKy+5D1zZimBG1TnEM1gRHIcjyOyzegbTvvZGZbiRxBkRXHUnp1XtQtSgqnfrPfa0Z1/2UBfW4hEDDMg7I/KhQ/yM6QhFiUiKiJP/NifH9UaHVz49cm57edUQXlZCFIIwqn3hF/jq6vUC8xstP0p5I/wEfm68J1HAgC/x5qn4ObgtQVqcXFfWy96k8PrNZ6Oa85YlPmENOSuvDYIY0sL8cDhyZrLDRyC8SvQ0R9vZOjcyyJUIh5cx7GRd9DkudmOOFP/VjjEAaPfiok5NwiCo6v7+wZbUyV3Pfc76TwJ1j5VC0iAXCmx2dDkvNnZBzuTPw1DoJQCrk2V26IBW58m3Z0NOazuCFIuqS+QhV7NZ1c7B3Uhfa3jdLACigz6XJawkCAUJgwXzoEo637iawEzlFwKJsbJjD2mpCJZVIQAG/my1evxNlm/bgRHW+r9nJ3vT4QrOsPWn0VTJgPA4rI6z8QUlXfFkilLpGvY6D+uzhgcnoy0DjZHs0kW0je+LrTt90V9HwZ0ZLyk8/0X/AXQN92k4EaJFbZYY13U4+PJKDmVxnKaFbzxLh/k9KysElA8/bX3L+uvUA+oBxsWH/dG7frqNGW8T7BQdNzcIToAzcXQq7KrzD3PQzVRObbhj2bfYT9WkOrPqvdYgKU8LSCm4eoXw0MRWKgD5220ow3Z24gn9X0EHNRjzby5EyS5vwGqmljCFi5lrfwvcwnT4cXqdsI9QrHA+OJhWaOw41oLlMOJ6vqHYxXnD/jgxcRpqt+H/u7wDIXpCch/tubXuQ/BWse0ISI0a8xoE7Jn2wqQBx00XiTwoRhpbHV8Rj8FCbN4IO+lhGfd8Irgp9d7nJzO6bBFgZqw5TwLy2Jo9oAaun/ktg6yvvZloxwW1NjYdj9NdiaHjtH6Wybbmz3Qf637XIpa3zKgovo3DmbuSS5M/xGPE6Zd9qQWIu/9P8GbC5X8L+Y2+mVINKk9LfqALeVRzxs/9JdlMktiv4TG4PqBVhXe6BfF8epA0TjiF2C4nK1aG8mpGbyDFVVESphl0XFZZ0CrESsxthnIopmJ+eUXQGUS2mA1Nljb7X3joLxEr1O85FQyL+AK0kSrdatHg30cLwoRMS9SehYFwv9AsrLFHkzeVyr4PPBbetSa7RpECK4X66Yx248SLR6FdOCzywd6mwwPzTNPI/dw21z/vRZh3fJWLSgmcs19TC929DzPzX0wwpwRbSKxMSbBUJxxv14znzf0i5sIZ/KiaLmu1U6I/SSLOkl/l6pBYTDRW7NPhlAj1ObRcpAQYyQFnT9TkAB18zZc+o20rYvhavDYxPeyU34PBq0+O1uczHyj8r5IaqgcwpOCiwaay8+TkgdpD2sU6poNhIQDqmDWkQpS0zRCVDnOtIdcmC+mM867IN9l+RbvCSCfxx4fgOXHg+1+E3k8CNBcuilcbbCyLlo0qwuKrPd82y9WGGJ/M//4hLSMjtB51Vzw9j+U20DLwBLi+JqP9LhaRqrUNyFd6A32gfD4S4YN5voQIme7fREP43cOQ+MsLvJuVj3rSqsS585Z2XHP66gKnbJ6SQk6bV/XVDeNguBVzh+UF3u2dug75BG/9vum3KZqyR59+Hl5eszt7sO9H7/e2mvwTrh8Sr1UoYHN08mvVR/cLKQFbLuBiaXRSct1flYK0yQgnUqqPsNAF4SL4/c5CQKLfbGtDHehZAfNnRlG/dkF1tV+b9ycvgjHgQ/6v5tfhnCcmSzdsNkeckEUDwyhqSD+rvnQ0cK7rROCc/ygB9XB3ZMlgizLxmUoj8ZYx22eqsCsaKHWIOtjWtNNz7RrdDQKvboS2FqIHDvzzkCTzcy0wMYVk6Gsqh8k0mV1lmiHGZoMjfQPRARrn1dCh+qrQdZKvS4rxPXg74xj77ZJUO5KXsasxrGSBl2/2tC8jteP9dz8In63EK6EwBYTCkntJ/8tj4HknGNyaSCRei+UHAc6egYmxQwmAvbCbyBfO1ctbyGq7SH2WbTVN1cOvKBgr4mKFhVI7dKCfNLl2E77NjMq+unEkTPReStTFfmdaZJ4ORpQNHz7bj8qLi02kk/lCOTq0fBGBucy7UxMXjxFQrwkPIdAE5Ku7Fdgoftx3R74EiQrq8wtmS8rTv1hkpK4uteZmtB/Zcy6VebAlCAMts8tToOdLKbomp8mGRSnMRvkp9XPM/7dXYa8WZ6rk2zrNW1P0BgUB444g5pP8PaJ9RQ8DN3fuxPV7hcMrwnKcmbnRa5mJ+C5i47BJpkuX7XXImXUQrsoxnafM8z6MeSS3Fi6PXwxMdFN+5IilQa7g6QVWrTPsX5tFFq4g7QoR8VyqHF1VrBHTtGBuDn2hB2DBl2h9QQ7/C+3Hp2l3ZpUYuSSW/eLSzESYbAZ9s6OYXqdGmaXpk6a1gqNRG00VdCYQFTV9Z2YsNb/F2pfFD5IBD8dGbAck3GrIwPWHAUmhq76vhogzu2cxn9X1gOuoZp+HKxnOWs6dNtyIOiAnAIveFpgI7tFdHkg7QGELVe02t2kjJ5r7Ctoe4r7wW+KfwhZWDpv3/H8VPulN3K/8jGll93RVR/BTkm7KPFJ/DzgqVr+q5KVxl2A2KvqbZMdEzNeyGyOjs1sQl+5oBCxNc+SFy6yhWwC+ZobYbGjcvq70ajntzCVwKm2ZK+/eZS7X9rk/6z9wkK1vHmSJ9rtJ5GVzLgyF+RQxOHM69N8HSjWScTOn3EB0M7J8RxfDUUm7VPeMQ6OSYx1VtN7JbZBuDYR5aZ17JvOc/4Oq/2r1jYPFvT3XrMSeu73GE8PfBAZKeku8N6NS9qXhX1hMbc4sJcuOlqZ+6qhk11ltQSFJZKY5peAb1J3iYm1PFoOpazMk6LGjvhbNQyHvBFC4MDBUzhrm/UM/HeJqoG3kaKcfUUl4/JUx/20kJ6YUGzMNjIYpQEGKGnJP/bMTGuZqUpRjD8p9kwLM2f0BfcBQIfUepZ6Gak3z4FDnAxT+CeogMU7208aqTIc213slqVBCu3aS4RrjH5F5ChuWGbdmjoBv9ivROKpGo4LhFUaVK9T5exFgXlJonmjfkseOeipGDW85vDZech11nnxdtFWJCpQtj57iyUC+bfICKyVprmzt0vAbPEhDMTnte+FFkAcNATA58oHCwcenkeK5XGMfvQIApLriTOaGB/g/07fOlBeQDK4tysivL2wcqzGVKdn68R5XkeHTC0CBdZBo+cZ2ALi+alc8PZt4lTVZgba1joN7F6FY3Kvpt4bfrLETgoTzYRh6qw6GqDxX2xrO3EFxoK95+7mfhMT0KdRKDxusbZMsdXchAo8MQWekyI8r+O7pKQbwMZozlw+GY6YLTyAiD/n1AKf67aQIhintAN37WRQXi7dUbXLf4qTFinXP0fgfyl+d4TyLHfqhbWTzQXHhX12sJACN/LJsQDUOwceWHkS3iRfuvd5DG7dhAuv1QCme07PvcDJ4oMFU+i42HdWRuf1o9Z1XBozfsanqvWiXl+MeRqkYfLgqBsz7dZLnbpegsciLLNn0LQpa8/odCHlvqzHgnVR9AZ+EVur6bhHH7x6kgHztekHpiOVqTveQbGhXJuJiVTcJSIjMUbvcyph+DeQR4MuGryFNLNDW9AfqzyolIRi51CmULQTAnF9XjAWCEk6WDbvHMql6KjBAu1Y4Svro1uMSlVKNtn7zgfUCiOheK3w75g1lC0ZETQcmX3eIywGtDKBWN6IKKbKfbo43LbM8tFZsC7aPjNY65izeV9aq83YGBAhhR2eTwwqYg1ve1pmqieHWy/NgZsUx3IwfB2OqdpiyljJmjJhi2thuTLgg+yQxb4HidNjI/kFUExCP3fwMvKM8zHRNUbRykPwDHARiDqQOMgY6k9KgUn5fMbVGibJkBHQYTX4pMd3HHHQL4cUFzWwf4YKpM+xYUcSqJCdsbYBKmQAAM0c5HTcws3xMCA5EHBqI6ag31M0S/OcQ2Aes32V3WjvNvrxwjwsy0xJTMp8ahFh93Ia3qq6/bLJDdHAe0y63s+WI6GN6NRNFZjUGsNdtgCuwbb6FFcW5tu60GhwUMCTWp7068YJCK/NnCWymSWWAXYjUC8ERKPDir/1Xdi1iEf8B0ZjicdEy7+l046aBden0CpimzP8PklTIeFoCXJXyAMER9JXc+oee03LF14tJ5Tpngaw6IKTPfnsk0EZt1owLaRdEn+WA+gTFpGftMuFrFV9g6JC9pmqYKepa18cdT7pbYSPva/AJ0pYMGYtDuOHXSrTbM67ydoW2ww9qwzbBfFFz3nGrxp0cn/vdTGzccM6Il3UfQo0OiUbDqPhgiY3vHwVguRqvK5vOP4qzhUSbWSCxGJBVN2l1xXgZ6VNYQXHaQrZyT0bfKFNiv04uOjZ4N6c5kgc/yv/Up7FWzpaPTF+ZO+czYzmEpJs+kiC2DUdg1pDLCXUApUmmOLEgV3hox1uZeROg8DykRP8ce2S1lfRfpPNPfKwSpFsJviTnZ+AqW16dsQck0JYmQVLNrv5zHFDQin0+Dor3cfX2VRiIcNIo0B82JzjBfRB1D4R789/qscYhivBlGctWRXiH3QKZKyuoNn2XD13QupQgJUnd+/XSG8tyVihxxcLv40b4bSst4qJrIEX0qCDZnA+AxQcSo7eGEiVGXzWThWtRcpu+QxUWsug+bBnbwArJRF6zzz7g07tOxyic0xe38YYmYx0FshD2ZvlJw+tDs5xtPuprb62Gz9rMfjHNi5xkdjDA6vqgKrDfYpIoXJCr8C7JlxmHNEV5Xcvke3gJHyu8Kjmxb+xQdSjyJ99Hto3blcnuCH+hts7ANmPBORNZroKLt7sNaHdIU8brFVVHhgNbApP2MNQyj0HVaIxVj+4/Zeh4LltI2syNrP63A0s9U5mEg00+gMBcXY69fg7gB9wMMWwKoTcMIdUN42g3c4v9XYuwDxTPCtXCJZ+TIVp92HenlB2UjA8BIC43O/MhPQsYkdwCRjF/Ku/P3Pso2nPNllbqX6EHO8lnmopp1bSXoSoinBBdr4YimTidnO0N27YQW0jSKZGDN9qn0gG4gZ8rHgOOLNvg5jX8g3LzrU8+7mSNlzlf6DAMkoivl0peiwNCmMJeeCy91CxCVOA24cOB2gHqgpjLE8AaViRhWhK0UqBSWhfh35eP23qflROT6QuoK2S1lRx1r0wujMtfM/auRcy+OU+bO/lEdo1kNhWCKnusH9HUEDIl5x/gDxxtL9TeDzXVYCyTCvz959wpB7cCpc7aQa2cYvfIvpWUQwtUBZwjZ6aEkDEi1oKXXIums5D2ylgn7oAaQIs/ZD6aLVqJokiMYRmE/mvnIG1S5yDGkm6kSiSZJh6oOwwewaWvg/QOoQj+61OVGOX4UZbrJupFnz9uBs5odlsmisV1J9v1qJTUHsSdZohHdo//EsVdTD/IJBR9eHrV/1W+3c2n2rLRwbg3E1mpx0ZtLT6EhjbauoRgiANcVcOR4LgR6iQMoR9dMxb4LcRDHoLaxVDJBbbdCWllHLjzFHJ2qjStX3JninskhMvM5TXwRfE8EwB+BWPHip/r+W4wAQPnbSPou4yTb3HIRbKLSAOEivpMgt62FVEwuYCKviWsWC/NGOLPVg6pnNFNjWcFfpsRUHJDPin2ODar+OeDlDjfZC7zTWP01RdWGCaQPjQZG3333vUVcv7hEeag5GJ8nkW+FUrHPUSQe57cqMofNL4fHiJebE74jnnwZylzdkLu6iDdLjEO7woVXOdAUWt+ANfrTxwFhlZYF8wYrR6MV3VXRJLMwA9KEAJC0S8PdgWboqmk5gaSgfGgPMn8pSWM7d1X9/QW59ndYhseKfaMz7Prg42UfmXhVtLtzd6EMa3MXbdYZwu+KSobdcdMF/K/vM6ZHPX/4L6+HeHtvgbxiiXIMc4+wsSpT2HLxE1WPrFr5d6LKG0lEfxY77mqnWIyOEUuWQMwGxshMVHH/sJ4kWtwndCMRKWQ4j1/87opbARpsJ8HY0y2LmVqLOiYuubRQ1lnDcqvHbBHDNF65AqjWYnKwT2JEp+voQFc4FVhF8fsoZzaxHVcmraCQ0ei/vekNXmfDfuQCCrhhYMyLxoK9Rl83R3HpLg3YBsX/jlc9G+K+rRWd7tloQ/0Okl5b34pxJVXNr0OLYoCXA01E1YOoeViOBk0RI4NdxlOGi+b294m6lanD7jVxqLxv81SUtTH0cVAM7+gA13a40OkMaP1f6lp1P9RsQg0tSIzl0uYnuSoPDLHexiSo17oHPyE7/wkn7J7wBnfCsJboS3bnEPjqfejlCgWcDBeX1rMti3yIqVPGoHnzs4QU9vXueaEokCDZE0CbXyy2Xya6/IfqYAtLuscYPo0i5XPMxOihCanJVrkLxQDOZGBaTO7RlIFb5tUXuhcgNgFG2nFVw8jFIYjN9VPGuzaud4T2m5vTdCpzoT4htifFi8fhlq4nMrIevScqUWk4wKPA62LztHCZjD1ddWX0uuniOfeYt1WoKqkb1buNJLvROIeFg6A6uDMU/2uDB1cQsOc0v3mfL5OAAeRrRD3syUJ7ClTkdtV1W3hMayGigAs/A34UwtznDVE1xseWtadLUq51VJ7L0hkrEAMHv0FtvjYP58kNMFbR7AhSxxIY9/BenthiNSZVE2EfR/wiGmyOoIzPU0lsMvcCeIzIdFDPp2WiQ32fAC7Ar1+Xc6ZSIfLl6nYT7d1O2vVJFhU4VrWCwx7tT43Gokc38fzDn8PCuTe46n9GdOqDfrOVMGJ8RJe2WHfkttWm45jAyy+dIGe1tXC22ek4xmjb4snw2Vm7Y//b+ke8c7beObjuR3sg988sPTpg3Mg7oPbspAPuMwN4AXzLlv1bU2AnZDz6h+HkwVyurrsYS+/ufRaoL3H7OOGnTUYeK0C9Lby/fMiSUMUqmpexV7MkwwGnWwkGJnhTDewJQoA8IXrEMG8UQdK5OKYlWW3ks3/ubgUIrLydqZf1UiaPR9LCD9VcLAsGH37uIrCj/B1cXsHOwsezMA70ZAREvRKJeQmC7a//O4ViC/5w9ig8rc8/laXVbYAkV575OSD1DfzrRts1nfQ3FUODxKosPrOOP5c7uV53zE0TzBLFqavINuwbgGNx7gDFYDXVNsnlVSOzx4enDBgbD3vQjVMkKdZj7YXIIdJDM7uAYLGhkDrN8vpzUfBEtzZiCUiYb9CfApBK2OLe2fn77S0yvYBrnEm16hKLHGCm+eXflswcqTNrJLwQ78IQtkv4Qmz2cqeRV0O+01hSNrP7YCc1A6xQbXQSwkVt9eu3rXs6qnMg6jcT892cU6utD3lYc+TqzZshpCSOToSKtUqOXdjqckK0xg8gFbXS5YB/f7URKfDhyQ4hOymGAYbuforPmdUF4fM0n6MlF05a315PFxl6iZ3+s7yS32AZScuVzBkHvRICEYxOeBjZeWzlfYi1YcmCtjbZYK5Hip/m6Oc9o2lHH2e+u4f4cvOYkYucuousjXFi0Fovqnhab10kN1f22SbQMkw19L439RYHdQWESyRxSWurAp4y6s/wYSANZKqymKNhQBs6B6J6ueUn8GL3ROCBt1+RzaScuaZvGxZDUvE0zc0eYHAVXcEu8HQGkFrEK9fsmKr0wsPMPeNGOB6wywrxmXaFwyPbaqMDDNQKqo4cN8SCp9mcaFDMK4PRZjtuRMRR5BaOJzMmiXw/sLS7wC8K57v/xgE0iJHnXv/qvEXbEB52Yr8ytcL9oS0dgoHzDfD9Z+63a2W9ZBI0m1JjtQKlld3AXRzWmx2tDOb61Y4rUtTO+IOJxcFvyI2SSR0ifqOrCJu9xeWbyXF8B6c8jSslufkuCcK27wWffYdpvv4mgw91kTQVVXQ766svMXw3twgdixqz19uDbbOnPX9u/TLcbvYQqBlVYPa/dcd0GKnnplf4v+j+9c8i10EQhL2/a8hBoErFQzKwfiMguvY0HZ5ojI0RvIQlQvNPgX+lmerO1hRlttYwtN6TptpszdvKI1H0oEd5WeM4ZEytQHwTGwi5xBaV+IWfQARKHlszGsG4/VNRPp521dV8R6rSOT35r7im8+8F11RQBed7CRfIdIO+HCaSmoqj+FQZPd66CgZM9N9VBiA8Td0S8jqWQI+347ofLUrKsogbBsy58E397aOtuK6oMetFSVJJL2Wcs2JMPcyLHUKasO32Ypgu0omcoa8Sknd8dJu3J5UfiIDmwwsvoLKGFF6SM4cFOoGmWjm1+SN4lwVqd3b4ALYgyZD/eo2N+PKGdc9Pvg0jSvA51/kYohbEt+K8gHyrXMKlhTR/Kaf/LYse7vDILXmWoGohocoELiEYyQCQYBrHwggkPWdks9w4BYMlYOLNWVL3LYEa/4tQFfxUlkb3PCDSVYivzZ9RejPbQujPlUviEcXU6L9xnEDLJ56H6UTkNEnlNtlGDUmUKsDBbBIqBUKvoolzFRlmE7ADFg8ByYQBeivsC1Jw9nTPv+LPLC4Brh9dYJ4UL4U8hlRsAiwb7miEQYkWPrEmhHA5PA7NAyqg4J36BviNiq1Ut82ALQ5iDZRIkXECs6NNuhmLlJKxCJJ1mgrWgllh31LdWRXzHY4gIhstC7ptZE88KV7x46JvCWVaVAcLze+Z2ElUl5y17JhgxNJf3E2Zrwe+KHcuc3jwXRabnqciwl6a/GW+wujYcD5jy2GemTH5padJXQzpP93E6RPxE2wuCbBSpxGtZMFK5PIChI6YKOu1T3hqwehgTTc+aw7O1+ctYuVAJS/NSjNT13YZ6YyMOno0hRu2gWFn/FLAOs5umD5wtETFrBGfryEb+QNZWMGU4FVX00x8megGX9xjX2guljUJGcZjgt7r/LdcrpIHonOa8wyonDHB3Us9GvnGpHyh7W0uxrjTp+H3G8rW1/In8eexlaC/qAuuseYB25uFRm/xPytrgdNdz/MqC0EirxaIDpKP19T4rNEufoO0kPmBvsC7CB0GfmZpdV+0hjhNlgNPds60pLLbS++IUUIoqLquQEXcRuOW8K+vSYgiBOwV5FNKExR7lD3j9LhElidG8HpbV3WKeB5VHKc6Kreb2hlZnxYxSZ2J6oFDx9G/ahFv13WsddVRIBAnzkZES+KCl7lab44T9PclrwKoJ76VhruKSe0LHAvcB6X2JHF+EkTEpfGFxHFhtTHzdzlDeUZw03RzRkiqoLnul2BPU98pcbLRX/kNGOlzMbgTlAHuZXsVLB/zbUUV7n5uiJwj7QStqy5Tx/h2rqZ9+SBB9ulwknBnuJahKDvwEitoR3+IMDgFFJ46AgPqwGpqdomZMmv8ccjyD+D3F+cF1aDqgIzPK8fFWAj6865cn1rtCyTQZBFvTHHoq7lPZDAOKH6MrfqJXK9OMUTjjSwDXHlWIM7j+o3vlm0BV9oKstuNv2dVSupEyO24m0RXAnsEKdWgv8njkioKo2Y5FyO7NUmnsfd24s8BpgwHY6tcpVd6NfJ/Gch4qs9M5JB8MPasC7wD/Zz7bA2lpbVZHGGF/LZEEzH8RGNaRqWAuLOx7FzAWs8NjxTOAX5kdxxnFyhAIYZd0iraNZ22ulTeO5XC0gz/Li1QByIjReyvkrAtJp5we0s/OR/V5CSupL4nwmK+1SsVe9hYKzpJ6K1xpyyOEWIGJkAD2NbxQ2snhKLgD+nQYnt0aqMnvN//PZ3pdJWQTxacNj9LybzyAyGykduYnJTbIZlxwSvFk3Qi0bvPShJ44zOxBJP/bOxRkR57JP6WsasIRRMOx21N8AbO0tu7ufQos5gK2DCqYc/AfCL53NAfWvniE6Ob9rCkGASQnkwi3xlCFFBaH/b9HgnOaqNfmPIzJirV2YmLhI58OuJFt43bDztEEHQ2HxXU46k7mznf5wPoUjAFoNhRaAyEfhyhiMq7jsKmLM+a6hz1R5GcIPx7mu1QKT+jwGWadCG86JYG4lAG49tAty6qqY5MVpBmI85Xd5mUtDRTWZj9yVVEtjuSFJFf1MDEOcceiWhcvMnqTTrhrb/ZTzILqH+Rjx7ZNkthl6oBAvn0QpGP6piHoGZPdBEDRsrZ73Mixbbq//pwDsk+y1+Rexz8qXLyAM8JQTRF3OC95Z9WalUNZCPVGs7RcPxaqVAuU0xzDtpZ0N2bNeQEbavoGhD/vBBeE+LJz1LKN3a4XKPkCONXIjBJ3SQjB25u316EJ3dAEhnT1uoJqtmMkLAZmf+maqi8h54LMjK25W75is83pwQzqJb8Ft3ymgzjpMPZODlnookqIKv9GpmVsr7uWyNDB/gRuH2uDsjNNukaZJd9Qo4odf7t4rZRp2h1IXdrGEyvgNgf5WJMFY/MMlETf31aKPy+yrGWrV3ev+8M66I1/BXdp5V9O1Ji/m0Lq9uYJt/u3nshmAex49No8vmYQ3SRfupCl399qOstanE4hU0XwVd6NPvbSEsGN6X4vTtAlNrR4GQeXXn92carotv+4QOOlnxe3C/2tcVRqe+MilhdVpUuBGVxIritw/j/bNt2wQBhbPLea0/i11hV0D92TOLeS7VUqPunYrbH0pQ1sIUrCsNYJRO9o6+4PvB81ueQAgm8WP2zzPPjNWmDV+sg3r79T9IGxAIUwVXDlbYOgGDN4BWcnG3wRD9oYZTg3rQ8Qe+e+lTa5MybAdhVyJQC6p62bx7CiL1Q/8iRmcVxCc6xflW1eG26ZM3+nbX9UKL/AI1xSTxP4u/G5XCV2ufSd05eID1re5U1zwa7Yr0t9GaUwIdv0iCrLzLUgsrYd51LqRMM5GA7RVrCUdLDGySiQA6wubDBzXzMXCSDRbrJi8Hb1DsiYZpktb/dE8N85ukCQdOYaoCi5Uezzl4exfBVNJpv+pUnd0Aq5HFOEorgxvk7Jkk02npCKPVuxRDraeUU9tXDZookk5vItA9ZFTCEdCo4bNWqUgl/H9wUFQTKZv37Fmiwp23EV0oSlKwgjn/7UqI/YleMmyrJUnp8WaSoY+AvayAKA9jGCOcKL3nzmnu+qEwY2BDPUqbT1ZEeqZsqRDZSeiQRwGY4HbzQop9XDafcBgftlLkbOXpQzjZDe8nnZQffWoAPjx99ucIUrzJdV8xpBNMaSUJJq9QbnfTrx4fxtcr8NSzEj6uZV6S1BJ2GswjnyraRF1Pcv4h1TBEBo7FqAnSgBggoEDYInTaEP6taFmnvIii0kdVlCYr9eQBtrxczz4aPlrPWO9TGR25+3y63YdusFbWOQEoHBaC5LJb4z2cQ67OpEhg0fhDP5SiJGHwAYbnaE7IZzP8+0OZmb5tCanCs1Bo2/DrmoBGjwnpl2ANJ41ss9sfcCTyk3TpMpohR+okZJ6RKc6Lgvt+fCctQzFeGH0ts9trLdf/OwRsZYU0fcFKbrLZOcN08jL01hDBmc8F3KuRMiTKml6aAZopRA3Npcd9QVQbBjEo5Pnh1RZeevH1+VUsGo3buSLJdswzO6FXkNOTzfXJj6TFvQq29LTtJL5a8SzY+vV0IMhOUPg2SCkJW+7yZepWFcaRaBCImCNgyLrp+pop15Qg1TzLgEGYmrsT3vSlodIcYpYk0fIJpsYnC8juGpkPk6DA7ZDjDdsnnj65fESABduiOidXXgXaYbDOVRF42bvco7Xel2GEGjXMWUpPAh8T6jN2sA6X1/oNVpOTYSfuSyyCP7QIuJsYNgWmqqG/IYH/+4fO1yW1Ey7kl+9DVrnTHnEeMXlc27YoaZh6P5qaRMv0vFrJTXmC0nlrlMyaPczPxP2OalSlKSavoIcy5ZmdO0u9lWgie32Es96Rxv82JgdWSb7lFLmSc+mVXTftsDppT1tz/U8a3Svmu7czD4oemoituMFBMIQzhb9mU8DJnRURtJBMInaza5tA4AiBOtDjq/hJ8cPmfys8JD1Jhw1a+3/cuERC70Oi/ghmo+H20tlObhOvard0hz6oBj6kiK0oL4F3IQrC8Pqo0COWvbRqYnFS9VMGHonbXJf5uW5PyShqUxOWHYzrm5v42Z3dmUUMJ1pWoNFBi2G7YUcAKE688ieyF4GAyRwiMxUi9j4lcOOI4fxzakefY1omxc5QIBwkwjxcMlCfW8Vpwt01HypDIhhuZSg94eces/xr0aLLaz1PQsyA1rQeqN6I/+8u086D6bSLXcIKWY5Xua30/TBlKJ7KYGLxMKQ9vCdBv9dDUrJwxxKfOawTginyGPRQ/OHU0/TBE1q/yaKsxj5j/lrzSQOm9VqcP/ct1v2h5SYyyv4V4RlwVDDP1a+FspnfWSkR/B4hBdu9DG5Kk9mYuItCKGsZxYHQlIq50ZEOcLnftSkN7oyiUtODHahdVprB+G4chFXOFPY2kjVPRTuen89soU6N+rdZ7ARlGuZfsRx95fnukOQsGKZweK0Wu2UCqZk/vqBeCs3RYZtuvzXdRCFReSvFFdVs/FoUpHumdBPbNjmq7RsBwqawBMyymREw+Pdb7CCsVPloGyBc1wO5+iAIaD88XKzfTgAl9jyCaEPSb31s3Hpvxt+WJs87+SGpecb5NgiKcg5gdxfXCYG/YnYJJX/9ak35B25W/RBrnQsXfHGo37DmpYbFb4CcIpScq94ZFSwHWWodH7JsrsOB17BV/ihMHnviK/hYvp8UeoufHJjD+WbKk7Cfp9l/Alvwz4Q7VzRw2qDdEQglE2+OuLoT0zYmujw71BqB4f2nF7Efa9283mIsjG1KlenF0UWJ2bvbtsR4ai2Ec7y1fqeVvXGRXyGmtnirl4I2MBW6uX7j9AvBefoUXJFTLiCke3yeGSQNaurMY0V7hSakMr+PknhULqXWjsXaxFRfEjr0rAPWJytClN7usyTLZ+iCJO3xGzoT6p0+tauTwKsiD49lUBGjC7zrXuHEMXtOLwatqBNl+DHocPiMrNQTt5MxQr/K0KcVju8NQA4PS538SP2N05HbTatHmS0K400umXuNN7AXu5dx2+MFOaFc1xoFMTBrjBSZ2ZQ7BptL+DIHO5iVWRKvWCAsIW4WZnBIoB6q+to2Y0loZOFF99g759mmvOs7Gt6Vfp0GLVhIp6pj9rk6On6fq7pqr9iV2ursFmk4Z1/laGC705kcUg6naPc/8eJCwTmi5ixVZckLp+ninHMNoIsnzrA/SHyEpWO+EpQhBPNCL79vXxVYYHzoUNhFNibmuxQbOY+lv2Hud4Eq1DGKeG36I6eMv0XX7Fcn9hevGxvfLW6rcIhOF/ORYIcPrScrN65/Ek9l6QHoCT53Ttl/D8EQ61Y1Ys6f9Ld7aBf2k6HuCEWE7z3R/9agZL+L/Q+QmjWDw4ORBaJsd45a9UZv5rjiEw1TKT4+rLzhEKeX3HZhycY5QAF5mMix8t+VmQJ8SN+vNPgM4+8nq2BckAL26FZDljTfVvGXAiDySyBPlJPcLFWJX1fc0JKG6vAS1klLT88OsAquy1ZbTm72qVrWQtJYSz53ycGpmzBVCEJhGg9i1IYZNEJGqt84c03zCdpOwnMuq4Gin9hXdX8DiH4W8Ma6vww7WX1N/jzkjVUdDRFFgcJEJt7WWbe37IJdq243kx6pUYF/m0QTXi717PcTt5BLQvOyCEHEOZfp82bAoUMdELOSPVf6uaihlXcDGNNRkVo8VubMSbk6HLNdlq0PWIzoPGokAmZtDrK4AeiYRSv2QLxWbyqV63tUMNZvEVDIiybUDQ+jqSFzJVlg495dbkpEr0yyAYsLsQndRHz9wa73fvSrye7f2oxkRgYYWW/6bjhOj3aJvFNRWK3PL9zFM0OCR45DMVxCqGD+SGrXYzkk2hJ4xv50zNcyn2jxod/e/+1FUixXdWnZEzgf2iZO2u1jgkxwezdCBvw5QXnZc7ooA6V2VSjPxpGS1Jk6z8tQdtX8fg1dqHrgpb1kL/9qcdbooDQQ6jh2Fxvc574NanDaBoutSMTf1XzoSoQ0hLuAL8gM6PR0FIp5nIQzYMtAxN1yfhSVRgYq8588qzQ3eHjXEmF1hC8bKc4BVxVdR40e3Unr/yf+dE269oFsmfdA6Ttd2Qx3N6XvKNEwdqN6J29lWmiia8W6fqZC9wdTjkpTRnz5lUhZSzuoqMAgi4H8BBkzvLFQalsPDcrxf/23pK1f1sD3GmSy4uqADUTNb8WWzubFDWeYhk4xwT4MpnmMxTV5k0K4YUDbg4AZKbMpePnBZC1S+pXKblKhG3JaAk7RtauRTaaAiqdCgf2l3g2QrCO9iADHbchIGw95QvzVEbcCXPoGjPlYrx4it342E0purIXaKvu5141mjA8sUmBoPQZpNvn4T0x8XVsAgZdrdmmcW1o4DCpOZ0MR164cXlVm7FhNlK6qDp7MA4XXseoPWSU+qwjdyxcXiB3+0wDwhZFu+6YGTt9jsWGfkeFVhU5Px6wngne/TZEC16jSVkkf6CxNn0aG4C/OihVH1pAe4fdgyXf9szFp5RpCzKTOEkvxNGexPbv3pQLx+7JmDSduRKYTcGDe7BrnGJgRY6JRki4e80f/0H6UggmBg7lixMBV0oeqfvFFhmFB543eLOtDtmhHHFeviJVXV5QIn7LTvxVOF0XLL3dIEtkbE9ONbSwMU+US/bxIR/B4/amWagQWzAqyLU2a391EzdMEsmrwgzfNXN1WtpiS6b5wV0BrCLhqulKO6VU+UzgfPLktP+hIlvASCRmp7sKMLK97OWxpX52eZWP/NRPk+Y434t28Yp/5oExVWTYbEGzVqprIOvcAJBPQplwv4J0NxRcDgiBPg+vGsBxL9xNUlL2q3n9bKlFf1IrunJ8ein1ZSN8v1relucmV/dwQB+0zvFFnar6jD2gpLPeheIU3k89IVP/7VL/DBTnyz8MMM/nooHk/GbZvraeQKUA04o6oONNHp1d7Rd1xLYdx1JlNMopxaSwWt2kPuFHdNYFHSWyE046kFusZMfs6yMdQ8MHs90bgLrWOfAMAplc2TWi2IqMQtyheeY7TLwfMApgNB1PcbiGeCZf3MUCp2h8fkbuDUtjjtTBNQkLTWBwumw9face9rDYkrTU4cZb6Sb1K5KLKh20YescM/R0Fl4wYoVdSVUBUH9M7RwS7QRhSH1921PLlxqizCBR7SvNGBbRRFhhIOvRy/vtVx/zPFL4kLcYk8o/SnFQn6bYrQ1agkLPGiN+NIHYDLSCVdm4QGOHcaK+NUe6LThQjxxczDEZMHo1C1qB8WWx45EADzpUqBtf0h/Pie2YunHnODqirYduBiCKlHTYSF483HRy+wNCU1ku+XogCdgglxC555N6VlDJasrWSeSuHypPpmxM1yoHrADd2J6jWf8wW4GfxsCZbSM4ORN7lvcdSm3QeovQ01ypgPdWvVSLSEjwKn3RlTHrJV+qoHQ83CLnRDJ1llkhAhaNhFJEnS1uD3pDKoT2oVKxjNwJsQcyf6MlNpcFoT4SeMmXiRreqDUu52AkuZcrxMnA8/BKlr5PiuNQa31FbTDlqXKea//AvVO0tljcGBt+4Zrv27/3+OPzCzXdF1M6mfEHA1/elOqnhhGwR9qwz8AczxY+uHC0feL7lTGVlMjR3qUO1BmLKl1vH75F3NnF1FZyD/zyeP7ul18xksTdC7hjAPPbEEWzgQASi2wtKYXdp3caboX7REkd9R0CAgTHYHuSZ2TxkHXNCDeNqyuyP7swwFRI1F/MvqAwfDoHq/OKwHK++E4zWDP/yER3Uz0+uHo37H9i9sX+YRr9qwDiZVCernlLNjOnoZEe6YjCs9dmtgweKKJz06JmS70l+/FkpTFyliUu9FCebzE0nRBoMEsSEVrT/Vim8rsjgInZHCxAmTGzTrQCydya+8mGN8Q5zp8N5hgHk6G+FeVsIqHHC3qkGZgwFx6VbkrNhgXnM9Tj0Qdg10uHh2BJe3UX4lc64qH1vOEgGpslbAH+X0i7QaPOS7TmkjQYIvCGpJSOKC1SiP3QF1bm43bCmws8ySyhp3q1ppHOzk4tFNEhnFxx7XVFngOj8Kiz54y+U2vLvpm7fFhojewWrOwgZ2Cuhkwbbi976UJk0degkN4vZ3bosZLjMFENvVw+qRSyHBraAx0lE82dQTpf5mqIDDaf1JuHzfKUSjYGfumFCyy1MxC5+3BSTizHlGqlaLn5TQtWlnOaobs54bulDYqp8joIHMup1sEYuf0o7PkSq+Zg22kka0+umsZs0gilSj6xr1gOPzToX6+mIIkKwbtnMiwuzm2396rO0c3ZEdes2zJDR4ifTCSnNBTl7zGhPFUR0ovwpUI4fGlbhc0fsMgtliNsORyP43TaeeBSq38BZfelAYGAk56m3KEBmGPGSIUQzgcG7zYde1qHgzNmDeVDNZgO4/ATmgjP0AKI1g1Egh0MsXhwpeZt1bOI/DyYTGfCljiwRHyudIA9BRgiG0hbKCOUtR+jUhEe0AKIKckpb+eW20aMWQnC7yUTn+y/UAmncSPqrXWJituHHNvcmXfHTnnpTt17E4uFxiXc71ADtI7q3IZwnHyXNAsMpEGZ1Novkc90vKVq1NNRTKA016ZpbV5OTzTWmFfBdCbKyHOSoP6pXdy++ZWvA4KPtQK/obMbMBHtKbeuVHYqHrc22zdFNM+nyBhFpFwZUbMDIsZO5kNf8wudM7brwfXWBwYPEYY3LD8AbC8DS3p4KfzX+LAD7mL0bIQGjM0Za86zeturN7yT889GK5LEla+NpaIw/AcRLKOA2jp2S5zI5dyNgXgoSN+6xEHKe0fmeS/QaOx9FkMWI88kRHtdsqVH79DlHhnaKFYjuaXy6CRYN8yBCK3H4RjjEeYYrJIRd94Nh3/yQTA59z5b3MQA5av7WPw8pbV4jcq+j0cLF6nNNfzEDfrX6b4M3YHB0bUYtS3KhB6pSWIEEjcc7+gwmR8j1YEwQe/6WxRzpDSjCo6EUnWzYdDF9xgoX2gPTiAsqgy8Y9IiqdhIOD4=
`pragma protect end_data_block
`pragma protect digest_block
c02e6342cf2c16fc9e9b6fbfff53ce1f7a18a30f2cb56fa5345633c5a4096463
`pragma protect end_digest_block
`pragma protect end_protected
