`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
/546Xt1i1Iq2YUk60dp0Ck5+jT+XOIUJNoBzFf61Nxxj6jHcFk31DYv3QunDm4gxRl5SGsGLSAogReN8wZJtoe5iNgU4YoLzElaG3NeIgGlMsPJLre655+fiO9m8cNDM2jVx6oZowUN3Suo8NGK4nKKT96ekCLkl8rbldzSA4IaF0yIVY58TM69ZmsY2m8+GpVDejgFfyFffQ9az6XUEz6uToCqRZwcfNmIaKlik3dgX9ZWHtVr4yri+YdSPKNrz9sCWv4xpIz7jsb7tGUvRDOOWW7Q+V2Nb2y0iNkIAPHBcfYLUmi9wW7FFkGRmCV3k/si/N/4f2dIAJfHhqeGR+4qNabdLP9MvnTwGTMPgx7aigclptC2yVG5Kw/CIzTnFPSsm+zncfOkFQyzjRFmx8q8NIcMqqCwEq5nC7JwcncfyAVZIZQC3R0JLM4yKhHeg+iWb2Mm1upLZiFMf561nsq06nAHL4rEFpIRJTEF5J9f1ZKmank3ddn6DUMR94oYScr4tQkpw4N5tCGrB5UGUws8aTn/vIY078AbXV++NVMID41ol8/7o1MzeM7G2ATobgyFqsDoj4GhNCxgU6p81GQkTl0+lqGKmpZGJt9yMJ0Nz4NZcl+rQdCSSmIt5LHntKJnRPs2z6E8/txJIBFnEnlFbUEaebX9ohE4O0oKUDVSB99FzLIAyaHd/EdQcvSQk/BAZtrV4oTbh9poulzb5Bx92XN8ciXJFb9EzdYpnnKXRnUz7LhVkd2fPP+1UfcRl9QvuKTqOl2V3Z487jcFMrya5JYf331gfjfYY9D3g9rBaiYmAzjsnPA7CYFOiY18RmGS2TyQqc0nNn2d3u+kU8h0octnfXDuMB3JieWuEQ2moQqxfW+sbCmjpm6/VHgNn5dVoahIOLZtY8LtZHD+PHGesAqYr2EDrbFsgNZNVaFmSg4qq6cWbSXAy9llCvCInLqUw0nB/tEFJnAwerAVDYlf4ZJgV/WClUD8VqGjIYt0Lrd00z4RNjsrIDSo+81LqIA9sUUIlEEACMr0Rbm/Bo1hUxV4bgJP/MIvJ7iWTACuYLYZtsL0vQHzyUwhi/gN5X7sE9j/Ffu1iE0WSBuzGB3zs7RLpItSV4iZZvSE/a+P3BMu/Y9obHmjk/ouufIKujSI/LhClGkSMa2yo4X7mVCyJd8weyD0jxps93E185ra30mJSn4Jq8BVptuAQMSwgzFR1kS3hRZP9lIcCKe8kYJUKeo5bEVdl2WP0JvCaoZpAIlUxAe+eqED4Q7OGaS1LESjKNnvhXRWHXoB9s2Es1w64qApNklvGqLAJ0vCC6uq2xUXjjBCDO+Aq5A8gRV3+lPts1iQraNnjNxP+mVAkPeWrwEjclCyK6rzBYpr9URzZUvhDvRW/7/cB4f+rVJAk8oIZl5ngCh56XYRKCl5JB6ewzQSDfICp5dkMrd/jDB/P1cNkRh89aXA64/aM7K48xP1OVGE79Fa4OEMgyf4jiuGfIvxQ1Zhx00B5b1CbncAqT7ITPUt3/p6HnqTHRYKM1Iv2ECicxup9fqU/vl9kPLexqFyf5zriv5O1yZ3/al1qkqXrSDZDjzDFzb1pwS7k6VUsAy5BlcCSjFgQDYGeCYuYVl4xwwLu7+VCN0D28t9T8rfYDxlWv3yrdz6ZhbVf5ApCsOuswvg3NOBTI7IBcWglnn9i1q7LMZcvVdlc7iAaJTHCCy+TdwvadJZC3ASKAUBthifqmpZbzqVex9mwnPL51hEzUtl9ZIW0b0HuOAvvFKDLToszOfhl5CaC5xtmN/uXfnX3kTaxIdbTUsFbJyyl1L3SqxY/IdMGb+NEXJEVXmBptH7XpeAWLeVzRmySHRf5162LuPY8hzZQ1GCrp494UrcgiCFi4A/6HdP1WEX3FzdQk8RDN5VYg3Cs0LKJ7eZLenEzx9J13d+i/dFFt+kRgvBmc2Sd75bq2ZWa4Euq1n0qECL5DS+udl7fpcm6F77C995hoHyNNvs0Vjq4tfp6jbxV7bSL3LEIhWB+ZP+7TkFaVVB6kojccHbnUXtZDycaZXNAwBgPuSEIi4VyezqYnTmT5kp9Os/kQ6FKFSocMGp8eZUsw1SxCQML8Lu1GuN4PVCt66xY6eciBDtPrRlbAukkpCAxmE9VF7Y7eI1kQ0M0HlXZeM3R+oQtQ9lvhTj01PMXGVnbCeY8IFMbCp5szx70O5SBfYn6zB7Ar7Rw1vbIzFIiEqr+QOMF75vFR3idxGuWGpSAQhRNfIdsWBFhp+YKn46DFn4B95LDjkV6To6SNuNnTAQhy5xC27LK5iSa1h/ej+hUbNjAGlXSwWCpFTU6E+d62Rrx/l6/c0UksUNYNh5B9GmIf+DAUEPZwm2vWdYcOvhOhAumZJdJH92IjA6LEDu2xHQmibZSSQsCXzZVdk1bXV4HVDf4xWhXVG4Plg8wHLIF26V9YwhAdUfPMgKkgfM+hjaxo01EK+hT4GBaOunstSlcEAyppHnvJoFVXcQUN5cqcJVHnamcbYrTFcypJjX4iw+Rsrve/WbVV+Y3brYps4waGwrUcJv6ZSTppsnYYLEvM1weNim+tB26XUvd63awkmn/Ygd8RRZ9zX+di0H+pv26X8cmnimjMq9ExPOgonAuJ2Z8TkN7RowXZ6/64HUICfli3FcE2x9MfUPh/I1HId4wr1Y6k2LIBIvWCkPEpXQq2wHQdPmerDZrkyXkIY4BAftsiKsmr1J+690Vtku6/fVPrsk1fwum4Uo0FqjX5c4m/FMYnzLk9UTgbcZZvG2c4SI4nhWFVCfaw/7EXWgCZ9KbQa0JeKKE4lOsEt4h4Bbe/TJ9NboKk2glBP1zkt5zauGU7z32tqkY/e02ekVJpSY4BjVFlVQRJMkM4vOjOu8nscM3mtVlVsO1X921Pf6WGQcxJjtnhlgV3Rid38BHSfKdqHCZyuNerE8ODUDry8lHMoemJOdZ1ZGHbuBTaLEtxdBLgpbAeAzAd4il1LUuMFbC8HxceSTXSPXK8UqsqEansrDbv037bQY806OYbPzvKH25utX3/RPPrHmlz9YEqCtdzGS/yQp8wcWJaktZzvsmE7DwEYD4yTAW5E0O4cn7zJbZcCtgxr6V5rx3BJy7HrP9/rcG5ErJLhmreuM4lB8TJMH1YJ8DXFf6yxYPQf1H5TV1vPgW5peeRDk0gwxn51ZG5uoyMjpm6A8FUjDbwj7SDRONCEb8YoO8YgfxMSfKz16WivviiTVbrLLceNYpTJYXLv1VP4zloThrTjGHOZ/7QjcN9cXIbt6dmo3mm7lE853j2WVMGcVU+m6SBn5+kJsm1I0XfAGX+jKuKQPj9WkicnxwDhQ9wOk7SyR7PXC4w9m2p1pob0CTUY8RyXoXIjubyA6DG6DMSiGJbdDP3lBCpr/1EWhEVQR8XocIlNFTUIfu02OxyLFLmiHNu6qp2d+6wx3rujk1xjOXSr7SYssFJ+oTPVNShxrlrnSOJmnENGUEd94wtCs0Vzv0iVJZc7UYWBOs/pXbycqUZKy2GyrUA63PdkJOtufEjdpBszJVE4GLy1RlC1OBZLH5J+rYrnkBw9v/2vUVi6lU5VkiQYThM73Fcc9kunWzJI84Nk0AR1EWYREbRREZrxV0vv88FV7LlOC2tFh6myJIjmZUnsMH1KBdMyBGbMIfiTomuoH8FQL3rINQwCikOpwg/w5ZwtbQeLhEdG4i0IfYwrPN86cHL4mlBlhiBEwyIQFig2Bq2LGtwXab7aE1V35JCmK3WQhJofbP69fOrtBmvfRKmGN/yrmgCOjrfNARLjaMMOWLLhpCEcJNoPnwWIIyrhdyOR3kZACYlGbwa8SkSX0AEpGl0D+zmXBdISU2GcSCYslX0o6gCvTTUQ/d65ZYCuJ09gqC9+OS2T0vKH6ZWUwwio0Iy0oYm2c52RpTKjN6++uhCgGX4Kl2bNF0wAbA0gRoUUOEJuP1CMQUiYUd6dCt06FZxuGvEMoXUVQUkptJ2C2PmyS6s7ajrSwp88zINeMQi6gs0rQAacns7CugWpFUVqgx0GCI2BseGEgKEY8ap8AWPNULpgN2c0a8fTc+3ES1ZQ8AJYLeqwQk9+ZZByNH94PbpjKgHql1DZVDuWFGkjOR3CuzWy2jiv8Y3+tKtuTJqzGYL2klkY3xmgxPe5PKZGihW/rbGdpGcrOsXKJPVw4Pnxgcdjhyo/TzgDAT5EYyBHEfEqMLbwlPmJglpA4nHMfszPk9K/UmfRhxtuEcwPUZfCFvCWv1wCKmx7+DZ5oumgo5+fR8jClAWt6DPkuyq0GamRn0KaGqGT6kwdpVrM96z7nrBJFSDESqp0W6ghVjm23pamA6K2GSA17ZgwuYxMSemytlPhntgopdj4iYikXfmmGx8B788/DKTm+EI65fG0/YmUNv8iPnkcj736RNgDnuq42/Zs11dSUyy2zyRgOwTO0fuNSl/RvHug1Q2j8xoT6UAryOk1dCaA67iIk7IIV6rxwprZH9bUcbaV1QBQNNezkrRy1LX0W/37JQXsBZcJqBts4ATdalTIgPS9xMJwtn7LJ7OVN/KYjkaNAyFnehCpLfd/a33Mjvb4YjFInIFBrFgh7P3FZ4mCIPNAIAC4kIjbTZvz+pfhgrXFrwQl+I11peoqisfFga/OJ5HUmfuPDXvr1mD490+OpJu/OM2AOxaNzUMY7A3HQnAlk4AXvnBBqb72bx9UGXftuXxsl2p3LMrmvnFUy/YiWcBOfkExm6zlPKvcDMBbkFtS+24sPTVtGLAL25gVr8ajozwAK/P5wCmFDHBwEMTiV5QEfkaWivNL5PwMs6O02pdhKWjxTjDsfxmKZWAR6XAS84IY5jaW5bvh6DLYzqH22RRkKzGuQxN4erb3QHmIaBYWR1k3zLF81IdVWo1ZF3gvjAw5WIoeGZR+nA8QQc25LTEJn7c7Hn+IRkLHuV4ZQcn8juaJUVIy91sQ2aQ2sgIzvqM08Qb58NRRCDWfZe5iLcPsp6GuvcT0Vd7aMmhDVv4ItNMWAS3lFVrxSnQro+cyONXrT7j3lwaKORo7BU1Cp6Gj/cs9ETQKhAxGlDcJsAL87ZMLe/EJyiYQCiACpfjT+B06fKH3YvkG+fjHc+8LQQVLAG5sr/67nPglhF3VXJx/uqP1deYKCfJC94XcWaYNMslHUqGBckuNWxA8XCWwexayyWeVQMtjwL5fYy7pdeK8zlVl2+UdJBbQcfCZQsJSYv2swbHU9RJIYizRH0QUQ4RiC5O1V62tCk0mBQFPG9eEoY63oV03wSDtin3SFe9d2h6q84d7wmpl47PSsvU/BAEJq5Ozie15gCBUX9vNwc1/qDA2oYbUrOMdTzuqBCVyFPSRWjo8ncmhFcliOPm8RVPq9TtZoymZ2OuDyWARlSDVTI7RZy2rqe6vcCxgY4f1KG+CiNuLDT+ym5Ci0c8bEuahWGmdYgyn2Z1PUGnKuht+7LSfJXdtoT1SXq7PSdQGAnGBL54e+k1bX5v0ekKxzstuvPVuRYO7UxOhz63JJexYnymxnablkAGrBIpwh7YY9XN87M+jKuiU0KqFGAaNZ3RfMBfYj2xhTgsDYY+6sKViW+v6PcziY/OrpYfRlhqzT5jHDjtklmSuONQeZvFt03S3DMzGFDIGCC5DfJRv4qvzS3Xw92Ztxcehu6+qVoj7jBFxhdcPQoI89PZqRx2rmRp3WumOabcrLeMOHiHfFchX+QJuizi4kkfYMO6xrtt++aFuaigrF6XM21hvS/0VLGt1W6EomLShcwDuKBERHLBaefjltOvLc8yLcVKLcWzeKo/+cYUvkP6TSHw2fFNO3uGXYgNqDQw+NYHv296JWqjcZiOJUru4NS7hNK/Or3WrF3te8gTKJ3dgkGn5E8twMxt5GR4vxh0FOGtU2WhTE+dWEK7K3e6kZfpdiV7QB0zGE9g7wExf+56zazRIlbx5VRzW3LpdWfT7/2yprjskYa9u8tKS6cpXSSq5ujNdAK7+LtAfnkVytGPaFNcvSkLRr/fqHJSHVemKq6zguE5Dm9u7wqtWb+9R6e4hYgNVfT8M/lRNmJGzR3IXFeb8nq3sUGQcygpibDeXUtwNSwzjfc0MD4qikN5idvW9PcUtJI9cnF9bFgLFoyIJ/0SGJqMKIwfSXqI2sYvdRA6/HU4KpoNt/kd0EyLF5//ji6AGZP68dNp+L1VvVMo+B2E3/T9mjGJErmm23Z5Dam4JsQl+PNdLFHvkTMaMHFoJZo/dbbRBQbdOhzpf0xAhHV3fvDz+EVt1QWTSUPiLspjfnBBKNIwXcpj2+8aDSu/EPaE/mLmjWH+7POeXhduIFPy7hFA2lWYzMZ2ByHk7uKxUj3SlkY4jFVPKXsrVbsQXS4o3FvrckHmg7GvH8e+Zm+pTaaUYKucxDJIi9Z+oFO90PCFl2ODmUgkf03Aoh8kV9llERUjOw2qN+zHLcjgNG+BnJANVfyRQW0+McZq3zlLkXH1HX5Z0oAfdb7pw8zLSrR2kKBT2fnnDJ6BvTj30OD2mqeWDe0dymKMciwsJ2ZaHvrFS6wKPTufgKFi7tK8LyiSxIzKWk/LtbCqvQACTuW0+jspm4+zzXwa9iLZHiE2OY6neTYqyTpO8CNld/c0fmaoGtt8wKSSfHIjLK/JNK9quXWdppFRKvG2M2J6d6vkQmhEHyEA4FUW6ZZ5xbHpmXp2+H3/90oYcjC6CC1XbYkJYvCwXIYPwMQcj3YgBlDPbYNXJZiComvDUn9Ufy6eSdexXrEIzDg1yeDx8N4vmKMslZhgpQY/xgqy9w6xgI+MZT5+UWoKuBuAEJ47IXZVy1x45x/o7ADqjMQw07+NYRdCLexwefK2G4VpcRTooUyIFW2uxop5JvwbNOo5fahG4yFpCUXpgqCU7oQaVahN8j7vOz5anmHFpghAiASDtRWL/wE7KtblKxQlzN9dKwIt3R3dwouc0u5BG0PRAJt9HMH9kVKKNo/bXrN7kCx3iIjq2fX7/B1ihMRHOW+EtfGjS8DFMuJAe7qxWr4qXW7PxIaNfV12mY9kPn7OwJCvd3uAB9QUZl9mcj4D/bsghVrRXTa/eTDtmoexXexLlu4QeeGdbGi9FFEUw/052HbB/4XHrZB9zGxlaxZrkkRlyszxiiL/iqdbPH28e0kynYKqRWHUqg8nIYEkq7cd+LmgWJ98s6th7e3kLYyTSFPumvvfUTDDrM+cse7Zwy9AgiCnrR0vq6JVN4yEkNWtt+9NwoVIkW08Ny3O4USj37XTIIvLzM2ca84DTsBIbKfrO0yBQlVTUvpfPBzKLeNFpCtFaTnvs59xUSmFc9IK7dk/aC9BX4iiq6oVxyPbMw5ARR7PGfp9ip+H7JpcZRqutgG8DCQoP/jSNAKO4W2T+eh3S5fGmecA5N+bZ3zNINK85ZMWhDXaMHpxUfyw3AMA2X4nsQF5vsctKqjYqpCGnwIWh9aMRHTu9cIkXuyhBqZwjTHv0WqclFlZLdzXY8VVeVK3Rm4hkn3rv59jzvnh95h9oKXUlB2tRi4MdTeFEPDZarCG6goygVDnB/x1OUp3rl04KwmxYXhLJIl3KSnHXf3cx6rGNLTw7qhylfsgY+nqPvESqZS2GeL6OzLPGhB4yJzSaFEuXEF6SBOYcgkW5W1kvvt+x9HGGkabvEiZ/YZTH3lv6sZvFTa7Zl/sxiCahB4UsTK0RcLqawFXzQHiTAdh8irsAXPJCksSTkTZSNqrHZS7gDC18BqVWKGA+sALAa8c8p5bB0bYIY5A6WfviP74oFy1zeztodG8xHCSfHUGPc5Ckc9Wzqf5iwybXif3sJ2ty+knJ8o3H2QZq7k0LpnQw7h3GMB5ka0hPgevQcFHQDp+i4I5KkdxBbCbij0uxHcOFiWMXh0jC+lh7p+DSDaV3BIiQIaxjm7lNzqUXVXUDABjfFLoX8gp6oLkwce/Beg2woi3H2gorSsb5YqB6eFl6btP1Nrai2uACshSrB37/UfH+qgze4SBds+ynchC1oGhVh/6jXWXrYbTDkm+lubdP6nOohDYLxY1iB7C/r1HeusCHB5CCf79hgiDAtsZ1pow4lO2t+1QeQZD1ISPSI0R4dh/DkZ7wPrtjeSm6jbslIaI2Uf5aQcLlEthK2v0z3j1af5jlu0YikNE+mG0GwaO3n4B8L4nUZTaa4tx6M4iOerLLpGupUSap5LiN+L4ezx1cRMJBwsULnOlZAXLTGZl9Ht8qIREfl/oNu31iq7zHxsa7sbvxRfOuIDR6kNOKJWqhqRzuFP9VZF/hTWv2QZWBWGrjzlJW08P1WKHQXLg0FTFZZpkm4tJNBLFLdtiaWV4+GARDlVw0Bf/ESY4u87ckEHdDgrNb897ZMmidioRPWvaMOnsAEZEI4QYYuOtLlOio1xOf84ZjKcyEgmZovHfgV1/iT8CKF7PiaYdsg6kdPpgkWjl/TWoi/ErDyq6VWRuay2mnDlT0JmutCvLJA4n8HKojHIG1fu7XWQnKBbdBQ+snQhiKWvv3fH1aGEo3XJE3Z5dpp24E5zLJMiF9KpPXRblJE/B9+ajxUyXhXTK3IjM1UAuP1MSUL3bHlj6PaSOejYikCsaOD7uPa/POIYj2GD+Shsy94XWdXfadwLd19TSwnGXB4OR2haPZlNttcQZaBECTKg2m7ViIVgVTqW/L2SNlg8JxiyJp2A1iqqnKpbAIAtKt2IHHyGEkAYNVsWqvtSeXPo+dE79iL9y51wBQoFD3NSfbZhURmkuI5z6Mzd0FGYCaJWw3Sul10oYUFKKtYePQhjV483O5b9hv2xfiXEAC48pd2VmfeprSpijl2P1btDkCO6drid7u/BpafzJs2hNcrUpcHEF+Tuh82aBycUkHYkHD8U7YnqE4Wl237+Ue8CAFy4dFTuKJRWebNe467/7+F64HIX2pa47a26jcX2Vk75Km7Y7jcMNyzt6Xk+hRcau7BwgOhITJwUEUxmqNBPpN79HD+wKo3ECdZRE0PcRnWuQkCETAa8qrJZJftPEO8Qz50gneeUg34TNbCQkXHmSPcFv0tpJJ5bVd1nYyMYJunfvgBPHBoJaOPIVUqTaz5tLruYywi2N3jKrd/1mLNH/coB1m+SC+6HIeoPdpFK2xnMZACtiWC8TjwYVVxKENmVIUefROxEdtKkWGPmw0l4QHxzCBZlqIhKbSnkCaq+t6hbF/dp0sMGeDIUwbB3iAfrVyms05vFLj85uKd+jbjtiDkU2ihOTVFudphXAnyDKLS+CXxtztFTstLHQKuDa0GHJOWnM7CqCRvih3B4uDa+qsK8z59wWP0qsFh2t/GPWkh2wZqYUG2mZ3LwOLQbAqCZNYIGNx9POJ9Rc+0scEY2IgIi1eXBE7wre/f93v593nDNCj83BbxT13eTwO/gYqzIDltt5unmqRQ+pIMMijeFLTKZdySYlAvDZzWQcDhnksS2Q4YjQhoNERZoTGdKrdVNZxgrN+peYOteLSgagVTyE8ng2hVt1TLzRMywFZtRBhJpyvhnCqTpHp1cESRmjJuOGxppF/2vLsHIeGzOvwKUfRJy9aqBvvxpn/APJbcZktC0UZrWApwFmluTzDe0oxCV158s3StY7lhTpP6lNb/yLQpGGcW4lyg74Fn90yenmCFomZ/HoIg1RpadtFFqP3YgTk5JVGGJBK/CJUkM4E7YsOSOmtwesmYCdr5OhbD5u3h3r7OoK8kQiS/cdjXUHs4MUGdI8Lh/zJmI0IvmkHScYYq5b1nDOKcO5yNReFmQlq0KBQSDdWp2yL+1XqczBMyt/c0IVSo0hhBJ8gUGLyCa40oLJp703dxQ9pP8c9oy7R/ArHDUyiXtHFqlxTMVntwpCDqwx/bLLh/HNEWQYaHxEJscv9IetYIVgWXBf7fTmmMAip7aK3ffxVPBxtfpIpfqtviufeNWTQHjpAkLDBIH27RpaNm1JstaCGgxJJ599Ng36X4=
`pragma protect end_data_block
`pragma protect digest_block
40b6b9bf2888f8656b20d338ce7ab65303320700c1795e1c8817defacd867333
`pragma protect end_digest_block
`pragma protect end_protected
