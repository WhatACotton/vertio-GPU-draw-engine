`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
Lp5jOJWZNr4MH5CsQaeKQlYOUYROUjxObM873qOIG808xmnJJZc5J2gacioWQvMQNdq9QzGxKo6i2itoMl+5WR1tTaY2nopcHuwgzIkEUvIDsPE1VHlF7EfEN+jr0dOeagysmjwtKvK4Gn0A4CevNQZcIJ8bULZitepFJFHnhRH57vyLm2Ku2JajY0ORpZD7Xdw3nBksfm3gyPblAn7xcXJqrKSAmBfYT6HKMLTunKS654msxDMsSbKnr6oRZUwnecNJ9guqBBnMZcw6jP2nw7ksBCP47PkvrYI5SZP5LvudT7L9/7polhLbBfODOrVzHfWApSCRKpIyxiPauxkyVfbGptRuMPxFBlmWxmOmwvcrvRqWytq10fH4cYWxV1f9MYuLPv3bpv6YVRo273BRO+q34FoZNiSY882l+XuQpkkcBP03RLKyE8VLvdptHdZ27lEzkOOVJe3FNH/GU+wxil/dIofUDJuxsB5+N6oFf5o0IBqMLAeBq7wnH/7fzIIrxYx5ldTuhnzbNSaymxe0gPengeOq+eoEW2rRhfq2OAeZAFkhEsIwW4YKjPayz7hav48xl+Cddux8Y2GbRnIQ8GHc4ljp7pYaHvsYUqr1FpP+Kug9KrIXAnrST59zvf0o0fspGtUkdySqxKGMK+8se5pTa36cJCMGbnp4y/VYOvtkRR1zCEktRtnClwBVJTVs6GEmsr3FV2AQ+WjMPu/n3uEq4557AHe0IqfUtFSLMr3MQwNkTGEdBTz5cnoztNv2vIvhL8irGF194jpu/LaO7ZDcJ8nSVHdkrKNUGHk1/h6LE01ombc85WrtQbBZLBW1rOK6JTwxGBDsYRqfhGqSYfAqWz0VjUVTmFlXRo9szVIRizeYjVTICdNro1HXvrn0hPUBMnTB6ocpLTfeYiCIPTfmDNsHvM7wgTC9SkniLGHuo0vaHaCdl0tQdjx/Fhyy0Q8WJJ7JWaocygfXJUe25YkoLzr6Tn0OL9vtzPFA/iIBF5sJnNn78qeM4bWWs7V2U6PHs3a5r3ey8GxdrkdDz/BE/pSoMygIQWu5M2/+JeEM+X4kIXHq3ruAKM8YyBb67Bxc86lnbTam9uITMJ8cchZzPo4+1cJDi0PBqVa+RrAIQHl4Kfxn1kj1QWXnZb2hDphJgTzzrut6aB8pB8vcdSpNLx0cAkhlVn6oCffLSvGiTFPhPUocqwLfdFvVQ76oirVR8m4CKPM6PLUJV5hXL1QnDHD8Gnsmu7V5QpNlJnj8PtmIHdzCm1TT9dOWTXJcQPFZTpVjCy0GwoDX8rRXv+CBJd9qVZdxo4bQV2qsYIZgY6qS3ms8Y4Ls+JEScPFT0JJe2McIFDaum6FrgDoQtTZlMn2pbmRzfJIaiua+CK2y5wPRo3n1M+1Oe9arMpuS4WxaKaHq66YBMhDnZz2JTNJRAlHkYIGNT7ENN9mJIa8BkYZpqwfK620XVKhwWUKdJ/SE+x2YI2+QYIo1Fvb6RxFf2c4qm3S8FCa5Pfzg5olg3SuXDtULknAMl6VeFvH/Wj9wl7SLlKqgE+57s5RutbOizOEy31DJT63yd86K9+0nPwbEj1rmDeiHwRUZXGzKwOkIbbTZ09HQ1V7iPOUqTYohbEqt6rgZzEk0UvQlfykWzOMUNPuMw3BLR+sHYljaVLpqzF43mkHdIPM1Lq3yHiyJ4ooE1HCjTUWeMDltMtozqP30/j9dBeO4d0ntHPicRjpWlESFQ66/PruKQb78a/A3MM6r2sqqKA4S/u5VxnXDseOIUPvuSjJUVHK75p5U1OBWz+RqxKIU9eDaJxrv6KBjtY3ULt5bWZKMzD1sQUVoFh+9qBUodP4Z5YYTG2dopajs6cZ8tr0GMlLN2QxK8+nkiyCxegMLpCgwJdsjj58t1THYFoedlqAJq10iehioIX4HfYhhoRWTgJgk4OigTYOc7+M9LU1BG9+6bjefONH7HxMZunK66KaI9qewAXAiP7/AxzY+0t3dtB7/D8yLdfNcd4OhSduSKYjx8b7T+lSxN8lqTZhWN+gX5ThEBUCQJmu/o1r8lqkSgWlGN0KFVWHMb0cuqBadSht0G7biVTdEjB9Y3oa0nsA5wEhZqEF9rjyrknoXzOJ9MZQkRvAfeWHrq50GllHew9rB6cQAmcoYERL6BUCqN/iMEUxDJj4Q9NoLAcBkenTSYgoTjVsFd7mdpisuts4CZG87kphak0MhfEzA6lHy5daDqAPlLkYxSfappMOaYGPcEU8qaY83WQZ+wIi9miQ/Dde87yK/rl9HyI0//3qK/k6WijWYUPgkSttpRlsixLjoNahfk/mzXgmov3HN7sqEsPcKpkvgH9/G4MJqFfIRZnzicVHY/pLA3e7PboBHOx03ZPQzlQoVQBHIxsEvockL5yEXAKdCumuG1ekRfQgeLGwoDKW1Ej0BDhlyXDMy0DXuWr2tQwrSO8kj1D7s73edTe1ttAszIn4HnB3x7sN6DG06QZ8P9T42EPVF3xvvU1YiAWx19oEAgQbxB0ZIVdQg/ExnFdXxq4/6/0iTZ9pbfjNnAR7uMnOuwttyLwwrfDVMBDs7EYQA7nO9qdSWBSIH73wFNLqSTEEHJUAGrSlJvtZEa9HlwhTRJeuJJxKwLmOvT0rEwP30OLRn2uCvbQkXDMczl0Cw+AsImXUyRw/5h+3DPR8txP93jbQimiNuzKfuCBOiomCEpkp1bFVUH8Kkj0FJHs5+uQuw3+zXPKsZ4qqF0DhKif0e0kd6vcuJ22POTNxUJrWZrSYKy1gByZUVxnZ+oRfSTJwpXat411FwunIkp6eVA2W3FONachyUwPMWuPzOAPHsddOzdKHE6ff8oeh+RfrcJ8b3KefuoJ1jMmYhxqCc7G0uz5KFC6Oa96fT1YG43mTbBe5OeUfPQXCfauguitJJKU4XsSDBaPZfiZDtKxGnbaYCvg5U+W7xDZBzx8N/sMrnvZiuO9JVOKxTnJPA4u8YfRNzGtkAqfTBGD2NeI3AKkLS5v4jXwUQBpiy1fBBHr1S/+zq8ggCk7vPBHf9FY6GHF2icmRfso2qzWCJm68jLp9VQ5BZvJYpzjvFnoCXoUX81uYp+cWB3NuSnx8XJtroDNgb41LLzsi4P5ITDcfu+vOuCoLY9IVIwrAXAoKlZ8+8/RdWPQIebrKNPZyCPnLgmpTc0cYN8LdcPdCJcw34oE4UNFjL7KV4vOXpaRtDMpmCnt60UOvKpeb2sWU0z0wJnX0tce8ECpm4vVI6wj9FOYlOUVHTCioeNczwWFlJYNKrXNgnq9eBK9huGXLjF0S7shM4FLINUy52ZnPeK6y6h5y61aVRJC9E16kKkFtu2GimR+x7hDY/pEL7N/ZKhRHh6XoAPNXAiGBj8qNaK61WwAFai0BCapJpwVWTyUC7Mzgnl6os+zwZVmx2c81psWSk7r1tZEFoqfimObJb7+uHI32oQif1IQVY679I6u1meI3z48xHr/1qdnoXGQ9gwp20sMJltBBVfyJuomC90zUCDYVJiyKm8bY6laYVIMvUHLwhi60Ttu+FeAWRt4P04Hr4abLC1xJpIobZhUDzZfCE6qsMguI4pIPuA+Zci59U4Ff0ndLSzhOK/bHTtk31jnFaPJ5+G4+J5iv3ddjVePVAjj+1zrcoFTpicUiFLdt/cddXSZP5DuVlHzW6Oe2TOai0ZgQiwHVBgfAtAw/YZnMidKvZMkUjiAEjCqQJ/lFoHdGoCZSUtIY8hSQ4M4dBqzOnnjTY2lZFNDPe33k0KjDniUdibeb3qnvKaQ+Jw9/kAR7C0KIinA0ejcd2T7KFycePqN0buPxdHBiwHT6TMHlenFFsYU/vAxq1oyT3h0kJeIR8LoiiEvBV9xVo5EB9p2ya4ommuqMm/1ESbUFUHlbS+6+VvUr3HG7fEnWg9N/oVSUiMaurpNYKbz+oJmbLasTgvlZjw3c9/4vcAb1DAS4bACJZiuM0FaIX6Yzc6JDcSXSgy/S72/SdTQbvU7rSma+icPaB0POpSIM6IsR0d+tYLSo6cDfZ/Eotis/TSRAyT12zDUcX+RaY4qsWr7h3iiLojGiOWhtDIaYUCHKgPuFkT4EgvRQAqYjwgUdaIVEWOMPvQ8VCIFiGgWsDveWcWjK5+wiUtpAeo4YrpEfRvVjChNTaiVitysiPC01iLQLFA9Grv+is5jTwrhNGvfToft2gJjFrOjifTn7QPMKT33GvJHqnRq0Q5Hb+P5bqOzRzdO9kFOBioEktpY1fud5lVFjgDLzU322vAjFRhgsDSNpJAvy3Ink+y4l48VPk49CFrqLOz1PqsPsP722yjui0AWaW2F4/JKRvBg89XWrHIH7l+wqAWzQrWw5Ni/Noy2/Zk3A0+lzayTIZ6JBjOvAZULS5ZPyg9hMxWw145PfqvHCG4zKaLaqoBzgAwBF0GfH2jMhBDg+rMRGTgI0v8cO2SOr8XGfQMRDN9AgPgJ959pBbB5plLBAATgDBid6Pvgi/6ru3V5ZjqAvNbt74eZHa9MzfA3nJPgZ0iH+xwRn3wJ5ml7QxVZ7s5OoVLZTCbFyTA2VOjBQRsCqzbsrTegYGSxe4Au135/ieknIfn5PJPykIi0Et7h/u3Yf0kKuKBvks03ObkAKz5l6b2WhaTckXz/tK5vkCCvEIGCxAN6NKRSQS5G5OJm6DTm9tjz9jfDe1y0hOcbaJ0nyzBhP/m66NxHXg28sTFv4RsDoZzsA1Z2mKVy0NAeNmT+y0huyxc568aVtToVvXKiPhaq5Kd9bXJQcvbbWtIzafUQAM88rHM0GfOe2RnZxpqFGuVPP/WjWchWYJQEXwcaQtDXCvrHtNk9bNytxZw4I/KT3qU5voM04WMByWOieoSW/L3g5ngT2zXiIdevXhpenBrsOv3GYEMtypDcEfS3KhpFF0OPPOk/bIacD97P380WcyGvjj7Dk7MXZioGQDtt0r7IAccTHxrobmezSrLk9PkSKKL1GQLn+9KlTEN8XBB0umEsg9/HsHjWFxlHIrvM/IRYGIEjGMBDTNzboKLcd/3DrAgkWj1haWzjFmHGhgtOTwGhK+fL4Asd2TKiCrETCwq5rsrFks1DU5z1CdAXYfwyhF2YugYsQwM3R3Gs933Yp4n/77cse+VC5J4RDcMXKeSRq5DkAFjTF77eI33THPJihJ+KDQVO2vf8hdDnfpZJ1ozucyoB4l0MP0TNyVdBgJ8TQXhvpEkRbDQlUz7mfYzkqW4m4do/GvY8EKcCcho9gOV7xR0N23fudR5hivKE/EeP09hJCAxf4lHLLt1lKIF8DVKqloIA19IHP7033e4PQK/Lh31B2b1jCJRSwcze6k9Y02Tj1JLruG5mu0XyGTNH2ZyD2BYQW1gAvrYwIyYQOsoc0d2jZkE6Tu/lpl3bZ/9Z+lwr5hr/WW560V9PmS5O7PvAcT0zj+1FnjcGofCFLzeqeYaulxgSPyYFmB0xuqnWGXHr5/pPX3/v+weUwiRly8/ufzRqvrz62t0nq1G8UBzQQimS/vVLwK/QyiHjL3Tv5Cl4qbLn5Djab7xus5wwDomDvhQUKBI1xfwj2KSSgZSHoPb7RElaxDnWZoQWJYk9aAiTsXacf5adBRtdgZyRh+pA0djl9hpocnkVihQz5/4t7yJfSGMN1CMnh9MMScp3BFuri42anv+qt1yu0g1zKsksrqeFuG338aBY/hxKmV9I9gBvwcxIEyzu1RDMXya7btby0o4a6ZyZt3yWPZIIS+eLI0/1vHnaNWBzxbUIlKCyPCfe+JslTF70aPzrGWPj5k+W6nzn/eRuTQ5EZrZwA3MaPNZdMlKfEqTSgMQSvPYn4k14jl1ttXVNUNljqFusPog86lydAHBkHZd3hpxdChJF5+IEf7M9NsoGXl3UmSSB09eqOC1MB82QitMeEanMLMtXmdalcVh6LGai1H/5CXb3yPrmCcSU6/4mNJ8OBnIbXah9o8vpNQ8G6roBzNrFe9dEO7NFwPtiLkDQhwChfuC6SQZ8qExVKKQTcYcGA7HShwiC9MZOqEP36Q9AX2MPAxXTvNJKH4CqbIGTcAquwr6HMk650P8FjYS8NFWDh7GKC0Wmb0ZGJkSfZbG3J3Z3E2h681/hzneUxRAVVNdbGPeqWqDG5IVYjwDoj+85va21gKmjtxzjcZgC23iXmfQU4N1TLW3jgRDkVlKo/DJ6H/U+eGgPwbtTPoHFq2EVhqhEDAq2QA3PSHZEkuacnjuwRhZL3JMz2nBc4r5eKQvCK9fD0Pycyd/kbYHVL/mD7+VNCLabRPnIopykPsI/Ff6YIAHw30jP/dKpmJtKHIah6jw+1R3DnqUfVBRgz/FdYWxe4oTmj8yNeAR8zxJE3UnLKiu9oL1dU32B4KCDQ50MzSP2aCKdRkqUd+guzlbFye/H85aW6Vm8aF2kDW3w4m2VjBm/M4gGKrmIG8vC9UdYlqU1mVtjhxBIHowWUlKvLCOhril4cATX36or08mZhzVSyMrtbpp7Xm6baleBUP1m3m1pOp3nC0f0u0lpyO+3CK6F9veXqV3l6redxX9Ln0LPIT5OHi6qjxwvVXbr/EkkGhyALFM/WCd+jPFwIXjWqCSB9GT7CxY+mI/mIdZPxhYIRVGqXztYdsP+NPq9AXwZKFAl9mC2JY7dzTaXp4GesgPxrg1fkwK2pTTTPKGIATzay7bi7unlA6TbkUfkGA0dj0VwxHgRx+sOjTdBtBZe0GZUCkNhQn3AgfjLTSTdCVvSO7Nroa1igoaGF8uho+x24pbhhT5Zaf5r3b4v+he18VbbLoh3krTgHd+j0rEblDwQDuS9fLPXIUIvs4TtYxNEzAT92W9Z9wE66v3V4cyXRQStiJl83YX3BYNNso9yRubLz2Z513nPQJdkTVOm5Mk2Y/0YNJ6BozO5w8a+knldIB885wBeHnDKRhku7pypo9kmJN0G/mBqPCmaur3zBKAty35tkokz3IONJAA4Txrb5Ti1bIba4P40wJMLg5Fokz3U2SbfWo2NkeIOldP0WyDI1Gd/LGW84VTpOY/J+nDAv6SujLJ+AJX9B4xxTTPA2kQ1pgsUn1Sjeo4Xw8UNuKuOFioXo0FY12B9CWyyo9LWNpK7wHuj0X1P0vBg6klPUTKPfZqvvG/gZfTstshgZo6QIt3Fs+g67PYaJWv2HwkIKWZ50+cjSEpSY5p4ggRaWtZ9SN4NCGf13TVeX/aS50TfEfCW7inVLCfNvf3N2juierPESXil2fhdZgBapf4YZBApdIAZ4NpDgCyumrQFGsahHhfEGHtD2avZeK1YT/eDo+u1kHYBChiTNKaH/Cu4lcP1x3hYp0H6Kxf5uCmz3L8XANhVGfFFV9p7k1M1kuctcy+JebyV/rVHMBrLf3S3WUm8n0XLFTakkeYoVwASCScVkOHPmFsEvgvEgyYZAFUT4EcgmAxc25OFOl72VRWiFqCVZaQGDdumQFjFZZFiMQaFEDlkWm1hXmQ6QtgrLask1tBj1EyLKpKjVTHkA2LAX+4uxPUjPQBtzaOuCpy38I+Zgc6L3mYeQ5/ExU2JyiW6btP64UAUIoItPAr64Tg+cPt1HLYuu29ypw54x+zEdHseOiL85FP5l5x6GmqGf85zIfKr44btTKn5cCmlbKh1FFg52Z4qnQP/4tI0kxSdoo6mHpepjGwK1yphYV/S7clBqAAR3SNTVwoBnYwTLPIW3VMC0/Hpk7nuXbiib1p9KO2naRwonEiYMMpnE3a/MpwTWkPZASU+dzuwMqJN1oLoEhe9vToWv2oKCsNQy+0msFViHMYXWwKgWUZzObwTxtyO3S6qto/x3UlsE0ev6unzbS7Lf2LGpW/b5dU0OqSzykAEl5ehh29Khbf1HpJaYZRS5U+m701HeEzO7FR2A0S6A+YBaJmWLDQiE4iXpTKp5Y/Cye54BleKpPUe1THuioFS/ol+iheX0hwCumy7/sU2NRhBIczUzZo72/cqPb03ywYGVAMMhL2VCie9jnFKnJK1lu4aCLhO1Gl774IwzCnC3E+tDqGFl9ljwYIA4l3QvEvOhUAntntjF9kdtuF219mbM8jjoqiyhM7UI6ORZsriqIxxK1py6DU0+uIVxFniA5GRdfQ7A9iK/VDRgv8RHthAXf03Ut9vt4qVwNh7bBrMgESqQgm5eM44lBdyAKIUxZwALM+vtjs1taSX7Zx21DSlVI9bDTvi1q7gO37NVtlgtbFcT7qb/CmGtXVZW81fcvXViz170Joj9fvqUKs4wR24YNDR71+ykz/RjJI7DACJ6W+tMT+LsDtocLEE3HaAN1A5O206F+sjyEMrj5r44tXwCuMwU7a4FDaYm6pz8Uf5fsMIvfcuTVIlmYNXEWPyRUug4v8+U91q1/CtdRnfChb42BI/czkzqdeUHWI3wN/vJ5HdaPYeaQzKjZhR0nB7FSCDT5eass+IAlsxY8ZV7D5rLuUGHkSThA/M0Pd4pAzfmOgS5ZYUzuCD9ZY6ot2E63u8RHv3h325jLyca5z59W0WTobOjZmpRst4PNbng3N+3IlqZF5WkAPkZ5V8DqYmWpxWSVZWintDZguK9FMiub4aU+DlYjpymI7ArFYIpPlJcMCYHrxntoYdrNL6Sx7G/bGRi4DE59J0P/yIzhMgDitBkY2ahojSgLI4wsGI7AWep3Z0NE678ATNf8c1u5eo0x0PN7F3b4AeJhFSJ4np8y/w8fEXhQmlt9beFZC7AGO2gYss/0GSHax3JqnacMwhZL1+ENndFQKQLlfDhxnOC2WQR4ScAHedBIpy3eCQpUtSW1KbEaqJ8bzEbug+ZDXtaS6mPbeJSscOQvtlaFJNoDVyBY/ZHHQLjFG9cY3x8YXk4+tfezoxhzL5GNP30F6+DFqkuNz2JErvMbfIl9huFZPJhlqGunSdJEFqJ5Dd1WMfvZuo24PpJAs8OGX6l8VIhbmTjVPBYvzksk9dPRJ+l3pQZhEmTwAxcbbEisNNmdqTgDLhMiOR/e3RV8lBE8Y80Pj0DDp7TgH0ZesLr/cNLJyIOCruk93DjtKUJbrUWm98ckRv42BWCMemhNX9m9D3SvW1J/JUCKxfabp8c+V0CvMkqDVY1UkD7TfYey9OhSdWVk8AjdB2usePlBDk52SvAxsQ01piIHAHRTl24R39QjbWSfaXJ370D4SyGydaX+Nu54EpuFLmh4iQ9Ks3bkr4ig580yvZA4LUT10V9pOKy8E2/LLW8i6iYoxwMYMP/xcCE5fUttlaqjthwuKKdEocjt2y8PyKrdYRqtSowRLsDOrzmaFqzeEtFoztAyhrkJkr9KW7lQBDMwqSMm38h+YeGyijV7HqLsajNs1ePrhY9U4Hn+nfGI3hUX4Bq7jzzLdblFMzrIGA3DcDOb890bQRhtd6ssOhL1fXUVTZGXsPrCng57W+hpvsa52HY4C0IbOpHUwfSpMjhjodYvHOjmhlXIjgCYxUUSyJrRjTibF0V6ztaiddJPkzmAbz9J+GJy5xhpLukXfxc/P+TABqdl/iYi+It1ocyJ2zlsQs2/wH+YeoAsx9Bueg7JUDRrvy/29+8Bmi/0Y94WD2HuOekKdsAl7VwJD+i1CFXgpoHjxnJrN7uQmQ0Iujs0QZLZsHsonJpCu+cw1IVeGJe7IZsgefyveu1Jg4P21fRXgyM+19gTAbiEgz1dL+iK+jIE+I0gOW7qfw7MHkoTpAVSgWE9UWXPfpt5BPV3CUwbn0t2DbjdP+1R/i2wYWD4ias13uIhCDUie4/thSb3ezufwTBcWFgJD9V9WanPPA23IRbK2geChYiVniHH3yFMhUp0CSn07errssRvgxTipOKwBuLPAhc3cQeZXhk0N+ndz7ZgzJ7P2PFS5J/fJl3CXOXfIGTGrVTiNjgZ2l1yoXty+Tzfqjc/g1Uy6XIsWBfGtCFnRXYQH0mhOQTBRAyhu0OkKox+ZSqSH8cOqvHcLAzvuZUX/u16JSulzUC10YXPEotinFCpQqkdjJl2rEmZzTEN7pNCS4ZN9rfUOnhwZgOGdNpkPOeAKUlEw1ZeS1IK29bdRPEVxoXzTEwDvGPaVONUvBBrBUzn2VSi03qi1Jk6aG+N3sxz7bbW9uA9zp2xwNhfn/CePTLZA/ggaaY6cPeFIUjSXzySaQ+Kqe0PQIs9CKTnoBjAafOy1ICwm4ocpQMtoO2hdZfC/nhIuk3Ei4HchPka0l3+T3HUimDsS3IRBLIZpGd6X7VjTQ/1IXB3kPtj9BLmDNJNFxBlfprTFeLm9lDKPHMTLl2bgRcP+lgyN/L1/A7Ko2YbPvWkvsglXsfRxASBvdhFiq2bkrt+HEeZaoSAz5xuVgM7zujIeN1OGiTJYLfeSkcEsZRs4Ol5/d0wHfeZVJxmvRJhfVj9HnrZg8jGoLVo6nKvDW+T98P8hmL95JyMN1pHvW3E63T1Q0aWeyeXaiBVhXETgmkRd8aLX3TcaGgizkV7QzZDyj6bfJiSf/BaXEpFs8uuupK7Jf0p/WSXsINSs7GR2+yrhBuVcr7mJcEJjBX3el1L66RB6/l49RZ+i9/pUueTYyFE1ds+OvWmc51OZmAK5AxT0wgIl8xdsw6GCR1ixhlh8GpDpTDJOtCkB6dOGpwLMOJ+Kf/61DuyZdtE6dK9eXxu7VQh0E6VoS/+LAjhWo2GNSThno5eiPRrprt80G4oJxbxRqFnhRB9ZsjAxiuBG+KM/ue26o3S1oLTeYQrWmXJUKHhtZZxg/QVWPuOTBaFnDMIHgRbL2Zs5012H9+kubi4ISebVf8j6xs6pDJjuKVpaU0PKrG6duDF2kGaj3HJpc6/B1cf0HNvLq73wzBGHLmUapXUJSKCDsHLYl2PW3Pz0+8MEzhy1SOdRXML9DENU8JEutTUlESQAXMwd9VouqqLgDKk2P60uxTNpNIImh0UUAVl9Zn9a8R8oasXyCRmYT/eWD2tFoJe2NZkqZaBv8A2WIbCf34/jsH5ODOJfJPyQbDYWAhcynSsf9NAwQGEY8L4NYXa1qE9cV0avW+clnydwhtkpvQU18OErmklEnRCSMLgcScrfSkOADyAxegsLtZsFhWrK1EQYM1cZhh+4w2lwlIjm3J9CyQNmZo+ruIh4gv+BzL9fOz5Lnob+jgaTDpH1hAR9g+HiAiIRAfmp5LLfIKgw0LW26M9KdQ7pytM4uuGvFp0eU5SrF0DAvzEZLMSxIgguGodoSMFwLOoTLVg1u7m/eMXbPvjOPdMAaGptl9ZyVl9wsijiN+0CuzlQW0cUnB1cBAKYR4TLsVkuIIy1fw8NOg2WB3cGeEJDZWF+8LCJAdtcI2qtvq5RXb1LvSd89GW+0xDcRA+wuKMJPtVr2TKqLbn82nEkaxDEJcgLHeoFiGQmBU1UFSJRWr+QIOPNNBCy/y2OCfWBvzPzBqm39/YhHHpyWnblp89+p7aoR9mXJMFftaCfusuF0CLANJa73rAhfEDCXE4+6fOPQKOd8n90HdFTywamKDjxQdo5z4LCGKZnmRkZE2VdqnNHw3b8CC/asbUa0cQlYjrxDfYcHqlaXHOjUmzIclXkf/S5wY1V7iyjk3gKMKE32gl5QNyRdZSTEVRnX5AlMghAjSwqHi0a5ah3PpkemSgQ40/ji4zQHDQD33c3T+qOljK5mjr/a17gmivHOdzwreYnN96wIh1qyPvmvCJ8MJvSZn88nF5m54lOzeGBA2XUHTieXT3MyOmrSKyATfS0pBY640JgntpfLZwz6xZOYQfx2X66t4ElIaAgZFPZEOLdrrHVS4dLSZnFWf/j3bkzxFgr7CwohD1n+11vJ5BxAulVJkgHXGooF3RYXOMPyWo7CAkLrf2rYY0on7WKzV/1KoN+E5iz5GkFJRZAzRbL7OG5jnygLpPBkHBqIRRkHweEbXGYkCEDFSrr7qltEPapsnRETgY1Iaa3zaZNmWhafEfzVPdIxa06xX7qaGVbSNnrwicz8KSQm6I0MZQ+AY5gMrfC8n+doH7+Kf7Xe93UxXvPc9NpQjhSHaKYGwEU7G3q6OV6brHBe7gv3udSfBQnRS+khz3BpD3wQ0Pnby2qb2iZNSdr6zI8Kg9pILARoy3cYyUhKAxTIVDnybA1bof++N8jYKSY5dQEJdkRXEVIykG5LaoDUEOmZ+zhtd4uj+BNvH3aM5ZBb3qHUcWwFY0Fjeylw7xVySOrHAXNXP8mOtKHsmLvuI7WXU3xEFUZecPwfCUM+epysAgGy5n8mrsnmdjVbgQjLqmc/hinSxuD4xK/T8JJLplZSB5jzPlblnb2f7tvsfhuAYDFl3KUClwaIdEU0LqVkUHS00womPV1DAavH/KWGJ8iWwf2S7YdZkfDTHylGkv0Uts3ZQ+Njf3h0fQ0/EWDMU0RjiX6XgRN/j2q6GMl2MH6kqmV6c/Co92enpDojrT5ftkLaihtVZl6qjQ1R9RgWMsjMi3WxCvAbeFdzRwSuzv5pkUsOf8coUJC5UXtyAszOWj2e07amyvSNCDZoiulttZvOLTWjZhWovjU6CTjGECld+chVJGB61lIeFscNxP/oqwDVSFgwAQhukXiHDgbLzNI4HCuFEIuogiaNDg+1BzSwX02FMbTxOP9clfbJAUQjBLM/+GV9Zub74u7fKsjWGjHwBfusKCyN6htWsuPdaQ4JIAZlEvzSLe6sfrsmPS3gqtFVPetN2oVocgwq/T/wgbjLcODvOvtgF9SgJkEF/0ZJb/4Hj9IokCkjuUjNne0aHiUBLiZ18kcD5tejOiBy/PKU6cFquYOhSOJwZOb4/UUaC6v9EFZNtnh6HnPzu2cR//F7Uhddh40h73lGhjy3iXnxYAa7o8KVNzLK3QdyoOHJd6qgPkDlcRI909svEF7NqXhK4dkWIkAyzhWNqHBwfeErYhN1MI7s51br4ZwtD0HBq27eSsgbZlEzae602TznSqoWmW7HZKUr5A6H2JGm6UhzIx6K5PpAxQzvTAyRMKz8QsLeC1uuijMUpHvVzldma78IsTyEPHMCTgnzmHNv0StRF8KcxLSts7BzPiSEGUauHqVEu3IEgNFVCXHxfb+uA641hzQJkV0Y2BbFi6e2ggVE6k9LphhkdfCnIR2kLXRDBbHntPe/UwvriQFF/Lj21SmXsRMtgmjJEkmY7RyOTEPVBePxi/vvE4lbzjOIvCG1uVcTm2s6HHeVeXNLos5ijuNY03svNYdAZmdXBUpPxWYuh525kQd9syf1AswpX4mKSaUdpEU5fzOXmwLO64OWpV+V1iaAFqXynST1MbUozbuygP0sMADDO5VagRAUSgBCD4GBgEAJe6gWenyk3YJ9+L6ANSsV47fIm/mmZTId36naWYbn+F5iNRjSVyxvyzOyy49veWy+KEF4k7Zw96K7xeZCJ+cX6/kuQFcmCJTB4Sv5+IP1djcOqfX2008Xe0cTL+ZhZWsz/MqepeS4CALUG8innxuz7D+Sl1bj3HMsSgGJ3vlJGcsIEN4/w2AxklL+m1E2fF1+XW9gdOekgWgvnC7GQ+hHWfM0tjzJhRaScxSKj+IFMbdqsMt1hk9Obt1Ej90DipdvjdD2p5SBMn57GW/oZb62gejyH3GTkFeulQgVB9G9Ru03rN4lHhVhQFpIfMlDAszMPh9OVDTQqR5c0ldPa8AIqZHHJiex+GAyzj+iw6mP6VJkmMIhj1c93dXi/Qx8wrucpDVoVKjMu32Er/j4J+e+a2HAQUSnEcrjmIidQSQcgzUPmuXFGuZKJCqUy1W2ia1ApB9IA5a3Jb+tgsPLoCVuRtxTjl81TdtL36o2W86M1V3jBNantXxVK4wBrZuY/wuqDz2BNBcN5PINlCiLE0ty2RIliN6GmqSxuUttsxfjEL3Fu6kXrXLacOa7lN/J1w9dog4ib//cjT58vtaB4utm3hdfRMAtjHB5exnu7VBnlzjD1+qx40gdUpYq6TAnMwoE2Pvx8n1KsJaDGxucFNDxSV87LdWyWltA21/syPBecb0s72y9pp9hztbLwq1Q+qM4AET1fizKw1s/3ds7PfEo66N28p4IFK/PI1bUZSQXmy4wbvRUgQxSzSoSMn4OcPzDZpvXf66qIbSG2vJkNhkh8iT5dxw+qoHVX+6q3koLZ61oAm4M077SL4GhCg3wRdwt+TOrCevra08fT/WiwesWbTPmLy/SjsLCW3ZEh/oRmY3ujr3gScTgL4G+ev0kenfv7+KJnhnGkgo9ypreTqoymzIvREXqLw3DtEdTCafZtceIupIghrMbkCje1p/w/h5AcVBtcpWp7ZQutXsaM5sn8ukZdXquInWkuHDbzuk8mq7axALJHQ6BluAB4dOZLShHoVFKjQjU/V97+0l/E091qEkIYeAejiUMKFwr3i6jwUbfbJO0C9u2mn+2lOiIMOm+DrfDv8oD474Tap7EJ/pCAsRq0BL2/ROI8M3uJp62Ou/KcAK3W8TzMRPOQ/RQqjVzpajnJOfyaKfu/a4l/uICnHvRh+3AGKzq+o+OzCdbDLu9LOGtQWnOlSdqdETCxnITIURLE53BGVVZY+sssmZXC3mcNMuhLFquNdROP2PkKnlhkYoMxcY0a42zCIrk8Sdtjv3c8ivQmTVc/fAgQXRcpp+OL7sSkXxKWQlKy77TvXGwCwcloYfXXQZTcEXwqJ6JRCqUcRnC7pGMsuSmnQp2sY0lpxUpNmRZAX7raotod1s8Pkx7UH3+9qpMBSB4+IOU6Jgpw/BFoX6xlTaGOAwdxT3Ng6J0Cy5E9QTuDC5CJFafg8UlQKo3Kt1oXvwCg2c+QsxUPA8Yz2+qppV8U8fdQasOjIITc6H7rClEtc3hnQkcqwEwoyBFh+U06jwyp8Kp6HstZBJNA9FqmQDEhSE9lFUQE27neXPy0UFnsD8iWVrDKSFpuYTIbkmzsIxryEfBxX0pUqKiV4T0AMEfWNJi+Mnl9yLvUuOVPTDa5eWSzHvNuiY1A3uJ4oWP9ypuxP17jnBuPDLD8Z9iM0RbPyp3wC+K2un27Z98R9IwnSDV+izgjpEHtcCxhkNFRYo/mYeLXNRivKEUgD6fKf9kphGbvoyaf41qJj3Ak09o+Xu5f1MINWhMQ5x9Kp/qcJd3OrFTMzX+Vai0LX4h48nZIgTymECn8G4TrM+fo/DWYcmqwB8N5ZoHErgND/mb7BtSKppiwMNe6kmnVDGn9hJW8vn+uZ39WfDxDvYdxTFqS6dniVM3tp37MFROkXtHHDAC2jQuYUFVQXw/nsIFLpLIu98yUw5fhfpS1uP81qFRMP3AZ80uTghb0/mEIwLbc2wxCg0X9oLqnkNLbM4FzyOsgajeAxVmThySw+qgswtbu1RtzmoLirjO9aXpNebLjoZDmD3fNiGcK6kSao+UcTekC4qUIYU8oTDdbewz9XKKBboeaP/4v9smikaNxfFTyXXXDI74hkmbKH7qRRwlU2AHBxKwQN6ufV/ZYMTYqzuxGc7cOmdXnNiVDyqL4en56jSlh03dHP7k9SxQURZMNLyMi8h+v8jCqwKwJUmMgel3ULfwJASjPlmac9RUGMny4DX8N4aV8CA0BsPiMeqy+hJLvBIdnBX6p0e6SIgFQ9WqBc0h8tF9d8MWEvhVsm9Ka4nTw4T0+qQciSBgQmLbqtVaYuhpJE8CjlieCpit7pKAXfp+eE8lCO1R07vNlIaYQi8oJaJERzXiMZPaUbb4NRcp31+67kabtQNRu29vooeXhX3U5XTgnMnibPOWq1B70eERGuDF0lfvgAc2TqJ/ZePF7siFarOAegTJHApJVBYGUdOSZs7j7wOak05MIXUi/KbLIUHgVGdMa34p8N/BzdD58x5muyBBmVbFZmxl+zkxZoH/hNWMEnwZW7nMBbdgZell8LGMXoj8ppTo5584TVwTV0apGqC4fK5IFwC8R++dBHOCGTbf47s++FC/QsUjnsBJFi8r34OatpSNVkbMvRc12x5X/Z0BcTnvaXn0POi8bKPwuSMPGuS95ywAW9812aIHrIi8Jqje8HcbmzZdEO5C5havcezy1s2I9e8UVxVh1RZUj43BGczwio3pKv7Mvky+YIWcZhwXy2zlCPUVtn2Zo3KPjcYXsUrvzHxf/qDbrYImTnMPdNUeL0SuOoBORHXiwcQMCG7+lFoJQnmPB6HzyJx1T1XWF6vDICA4ULSYRHsjLw/QuRcWw6aH7n+cKc3knU7w6Ao7By9wYmsAUQOfGpz/d1tnZq7LG/UDL4Pi6nSdILHFvFUvI1E3rmY8FpQD8pFA7vCpF0zCCAfSM7F2fAbn/AeEh5/6DkaZeQ8owIiMLHda7Exru4AVthZEAAv4BYYKdr/hos6zsddlgLTHiHjfDsXgD5IKFYUw5464A9CJTPeHIvD4wzlec1bgKxLye/3AwuEEobva4y0IABjlYU3O7/XdEzL6l/o+Xu9MoWUO9+Y1cn5AFJCxTNrjaC+X0mumwolk85N5QVNU9fW0d2O23HGy9DC2db6EWi8xfwzz69FETuZJTdM/b7SC5gb6nuzBaZe/5PzZWXc5LrfO00dqSAiqoIW8/ziD3yVbCZnuUVmT/j8cQlzVv7V0ttoOBG2aRm9w056FrBMBE80w09YzDzo7JCh3IK2YYNpBqrjThAJDoF4SSEp1AzQrT+wbkE9Q2oFL6jVMooO7cXBClKaCyYt9Z+if76BewcUzOzaPPON9bS01v7e4Vt3jGguOrKObptZNl1nj0te+FJMrRBDCffL7hyZ6iUSuussCNkJPiTwiz+Fd6VQD64rfmkmHHCBY4t7me77OVXFD6kJ2V2Qkw/V08ojEh0nksZXLfC1YBV4s7iBzal8B6H9Ja+5DUz0QJIE110z0ESGIp8EKZOs33X66kGJs/ogc28hvt99JejuNQCm+mcX+l8UiQB2DJ378mwGkRmF5ZUEI+BcDw5BG185Y83vloqhe6vRB06DCtSnDmMXG6WADzCYmmyfUJwKux/1tvWx6tsVQBprHIgs9GyX4fdFfKfySAnK+XaMwSHRzNpX++2iARHcGrPjBxnPaWPAqkVEfRWNlxlzxIfosBaK/PT/2nQuyvEHppUt5B9IozvU++XTuG7fl8d9Piv6kKx40MJWhw0roRArh1SxlWCWgi0fF58kaOg9r/oau+fvpWyWCQZGBPLSAjU4e6Hj6CRuD5A9XR0mivXmhf6XiFwS2dN/6ldLRDa/d4g8/YKC478zZEceksg9CXLJLX5fEeW6QzOfbjOm/IOF/P1sMROUEVm7DTpTwInsmL7jqN+x/KnpdX8I/V09AqTQCd82PejjqoESU0fwRjRlxivsLccG1+foBcDuhVBHwY/Ek+p5/R7GJ47+68JjrtL9M/nY4F9+G+Vi5gnwZq+ZDj3sBLzFMudxiftZKEXsKKU29cKUsdM8GIoc/EXeC5L8FoMtpejC5ybmHTO14y8kgz1N3SFCiQaw84F7ja/ZjusgMOcStWlA+NE+MCh6AGsqT0czFwOZJW7TWP1H/+SbQEj00OSerbTzzvH48J+tHOkyJeN4OJVKip0NFNFu+KBHu87JFeASQ6iDHq8BSxCo8tGfr9zRk69e6rpMdFEtdcEwxsaifEGBj66cp/GySn9bVSXLx1tM4g8zTXH6JNauFcK3cTCzGR7oATePQ1vXWJb7F6JJp4VAmQVTTgW8aXpmoB+zK8p8t0hVn8Y+i0gAlV7EGOwEcpHrGSmLTeW92YvdEZgDZiopsk69f3KBIJmvjQHfXoug68CUCuXAGk5/c809kU9unAxQPcb3JELDq/FNZFFOG3rehoU5qW1zWnc1SJmVl3jZG++2jRacDBNggTVmhLNdoA6t2TLIglSNbacI9s88ELm7JIAVXpU7joKCh6hLT+kYXxWM1zYdHZlY7KZdbKhKl9X49FiwMryU10zOZWmlTx42Mafp1ZtGQ5zUtFqsVZ6JrBruJEe0rFFrBSHMLF9sX8b5WhvvTVXjXONm5SEOi8s8ZSwDnQO4eFxO4amSVIJWL80jcO+sCmxGfujLkiHAi6PiV8VOAjbjDtxTZvNG8zZ7bZIsr42fV+ZsZ5/tXCD9XBvTe8bAlMEtUisiZ05E6eZHiCu0DEqT+ouvPiRq3TowKt09ypFytajYow/sEisVCByyVVEb6iFDemLcL9yAl7qHmoj25XjS7A20LWiOpOfkKXV1OUlgL2cXPkL1cgfTGrxnlNYJPm+6RX5cxOF+9tk8ywuDOMBYzRdbLzhcbrF2jAL4Jqyfaa48hhLd+SGHI9GXT1DDISJZzmm9Jt0V7xKl+wq7HGk1pEczEtCkn1hSvitD7FBaW9Sf3njvgoxRvDMSyHpeS3Lwkr23eRwSUQ5Am6/vOy/VlWgZxjH+r1rtAPZazQTgiLOlLmajLdllPuydq5yju9BwSFtUmAtgf3dCV10VNXYZnTO2WNYi7vhTNP+W5JlSaBhMdy0v+KuTiADk8paB05rhFLDNkODBrjI+z8tynlaaTXOLV8hNPHdmQNuojKB81zzn0ohDkNfh0NVGJ5kzQTxKPffhHQP49w2SBmHYaI+GtskAK6NOU3n8d2EzOXDmN1wnOfPxF4+XLTVmghGGOUOCHFh26BeI9DdHp521OzVEsjbsP8HQPSyZbPIQZqjXjBGomIKRHpPqdqx8ndhrTQONdujO++bp+lJU/LcXXns0tNRuJqiIhQFdwRExxmoqXx/eDyNpoE28FqX6llEifFxP7d/lZm1LYliYqiaCAkoE9OeUng22Zvzmj49wbztsl8vpzN/VCBE5A5hQmZA/hlIohFUnsQyGsj7rJVU++/K3v2V7RMIyx1Whw9hguaKhz1o+CHJ1k1rWyDSdUq77tECcNYc0iBs/F+a8c02rf8oxnWQQwL7SUVkLkvH/TEBg0gfTsh691PYMBCOmBkNgY0WeuQSK4jyMvSNIH4AAv/P8QLvpWuejAJSTnYcfwsDiveP6KexzN3eI76Suawo9xZgmgjjyfnDfgv6i3oaCOHY88EzC01Pt0O+hIH/u9Ch+4cq5Rw0uA5ch0PB3U9tS14+HzIy9nzhOeY9BIbE8r6HjXgvIa/hsc4UNb6GSeOazqbGhQ5Wy9qhaXL5jgqGDVi0STcT/RrQG62xLgx9q/CSSS/7h5CKS3N2uwg1NYVQfSZzyz3+X5kbCqv5cRz56thAIZ171wBX1Py9fi44iIKVscwEB4YcHaM+0tisFc2za/MsNqIoJgjkK5sSZeBBxh+AyivslFyPHrDvcDvSQ4w8COe4xGZ0/XE9AJXOgTM/9FuLegEf/NYkejn0nrhXPd34+UQgJ0TBB9rr1zYf+hJA+iSlWa0SfRJ11os44UUc/XoR5nXlu0Ypj9e3PNJzEqug3qwAxTQvslGJv1jQVbBwt5UXbu/DKWt64qFqvfVjWq/SGMbxroLdVxBE2FSTFJhG7cg1uFahLimiJzPchx2j6/0zWcgyyIY9gy6bfSlpX17TtPHLD/I6k/sT/puS3176dUO0YGTRRYZBoQ6BNT0GKXg1hwatAez/daKI/A6AtTypp4xqKoCC69LCuF0W+HcmCh7EywNqMQXHPBkUDvchGWwlUlIDbttkeukF4Ny868SP5XyCSBx7/g/CIdIyow7/PxyAxeUTONc40A0YBAsZrRtXCXsoqkSo9fJd5O71eXP9hgxK3a7OK+oLoPZZ8Lf1e/y08BOXcYnUcdY9NSZbNuTzRvGTTeDjipqGOSzkVN95qbeLqjnMkNCRhHyTMBl78b/rAoWtsdOZhhlVgm7wjAuy2UJEy3dQvaxNShZET/pibzB04/6rehVOX1vwWvfWbNRnXOZ71XUzTEDxx8LKwNyqfsqwfja9CT+lLQsMDj2DPbDyh0/t2yjs4ghMlltjMyqGVNHXs75euYCjPjt03PLZtu9mI90kPc2OFNSsgPf98ltcRNSOr6UyyghB6HSOZz2RqBthRwfq916gEDKA9Vra7Rzb4PZPnnSewDlmAPKEYuvi7p/42GlqZy15L//oYBYrZguCH9qm50x1ZQiAChCFGfTWliG105z/I6oYe9muQZsqFYPacumxju8GW4N0TZ9wDRnRqE/LFUj1lp09x5BXRtF+BbpPU28yZkwIviOaJ3zkEZJF3iklGH45JOK+GVQ7F0WoOiLD9Lfw5w4z7qQMjJLM8TFyqtE+e0raAJgPgb97V7KJLDr7oOuYIC2UJ8sP3IOn8XXzAdrHZLVr20V9AmCP5qbZWbsAF+jwMpjN0iDrvMU55XfSmQ+kscswP2/Q0PE19Q+UoOq6q4xSZbfuGiWgIlaFfFomfs73tkzsOCj5y5MxLRdo4zuBxJU3oicZ6Q/h5lo+hcLTJXbJuzd1OHlB5EnYjHtle0yoN2zW/MPpGdcbzYGNL02Yx4TI3imaCKih7I6ss2XRuYwXpRevbgSlHRlVb1JAlAcf7xym+F5CD9n6g1pgcPziD6+Vnn46N0qo0UQ41BS4hZXlNZs0hKpWEQgDS3jnWx5Upsj33zNFovJwski4I8w0UsRcu+TKXDR+iyfpL0eFCiGNloyueorxTeJHBeHPg5YKJqPrHcAkmGak9vqDKOrxx9J7IoCGk+nBMYLLxZxT/VHJIz1dlnhrJzwuYW4DQybRyeOcKLIlfODTUdG8pBgb8yzNqc+exJTJntaiz85AjIr/x6rSL5kVCGbRe8slCgygh5+eCGafgjK002CKYZIg5oN0UXtaKPOOnqUHe2cfCITBAJExNeTlI8nRV4KPlv5jS8U/GNh0WJ1lwm5zubv1u/yw4lwWJWzBCTVBh2ljMOVvt/Vo5744ToN+pxUsIxuIH7YoKrGh8qpON7AM1fA2AN29PFHID2Qo73rJ//K10P+M4yms4Rhm2oHw1iAXglnoHx9irVBSPMyl4Wdm7C+3SqnflJ38AQtmytBQs1TwPnYJlpjZaWOF6nBZ1lZhOlYTe6xufRL1sHDiLmJOzbQJ8vt/wcVBA89Q/eDfQcN9bHIUg7dRW6eFreGfQYJhHb4v18K0+Ils6DhePnvfD3tFM+MIYfrGe7tryj6OihQOKhEpowJoMij3ribmJvhuh9NIfE0yvbx0JBap6YMsw3tPAQxXq8f0h9+SEsipfhYsGZ0vwPX3GECSdSY2HF6S4yxew0sIUD8NxKsiokGI2eolA17MQ50qUutk5BNCPV+QRX1c8dVcti6I47fPBWnPXvLQVAaQC+EcqoClSMARQ0DnKxTEE+n/KX6gPn5+iCALALNdNI5AFxvTzoPZj7xrWxXcIIIWesUcyG0FIyYN6J6nyQoxvf2c/7D7zj1nyhT/6mJGMjxZDBI+t18HABn6ElawNM6yVTQFWL/n3lvngGd8imm7BIuDqzZuyh6KAAH/iiC9Lae5/0/VG4ocKYNJ/4Vr2nY+8MWtHdmvmUhDM/2Q8mo+k76WLdCUywPTHlXIOdEGKSOU+Q4Q6U9Z6qmYVJF/JBR2HwMnQwTURHhiLSAZvEdp/vfB7zZNlsOWUm6j+0W9xn9zi+XcyGTdl0MVPgHHgnXzpGCYITRlCPIaFt6meznZMUhIEg+WsQUhIcCB72iSV/7eFId13FgTjFDd3GV7jvQFPRjyuKZ2h8XK7Rdxzdvcx8a9FT0l2hBwwEpErcszKvA1iJ4h7wPwz02p379EJnAolQEeuCs1mtMSN4KvetKfHhhIyOn6NvAOeTxARsycHkBIfSVpa5q3BmfrFnPOjWUsrfyO75LWyrWmZlKjowicGfA802Bfw4JquEZklOY+xwQZI+KvUtyi27ihKSdWbGczNpyhj0oLHBHpTqljPQDOVW1JJvBooQgD77JOEWOx5js1WFOeblXQdDrxmDAV1m5C7dFwQbsnfnzD42gSWATGEOzyYUzIY8oloSiq2/IH75s797a/tguvBwlLGpzx0/tWl5CDcRosxiPXCaz3xkP51BTDtnNBmoebFLpKvzqYKFTw2O+dvxfcIvZZkkO/7zuY62dgwlcz/vS7mMXOi2oqz1ePmEDGHlJYNUQdaOEbeZOkad+jcei493vyKPgyfGhI8rVou16pHbota3H33bdZ8cbfU/jleJmOg61ELDiJzHc7GR0cy4hj/8LXHoyXapqc1sKRM5y5NoUaJ5qR8dsbJtSHHatY3Vu9dy5k0/lCvZt7vcZXU5N4WM5nyZUMOG9dkWQLMYypL9vI6lcD++tmLVM/JeofTKQ0FRLzG0k2gMAYdaSiq/mB1/GDROubRFFMKauuJ1Jxj/vEG2lPcZOCpK61GKbSC49wefMXA1qxHnpTah2/fhV1QC7Ac/BQOGo9Z4BssqW5bl/ooHMe+99sTsiODs486hf3oWdelazYdFI/NFWJ/UhpNwEOwM2Gxoy6WXKMI/tAi97HAaHKOyYBy+yRAGYXNo1y93gwhAp8H5Qys1A9YXsymHPQkg9j+rP3zjtOXtwrtmCbr3nWoboJniPv1U9UTO/6WrhuvwoEb2Zd4AseQw/A4Sl3rRewJyOehdTWsRNvo7tvkp+X7VwOesMs8BDi7BHtXyi10rqlPn5LsRtJO0q+cMOE9WhlhFVzYFEvAuycZqUmfMzsID6/3z5sWf10i4CRnXJErtFpTUlffcve/8hvn3OFVfRIe8RijkpJqzbL66DK5sE7HN/Th5nC5BaVXQXLNnjwUXiEfZsFn5JvT+oHm0l5I0STXRWOT+atg0uzfrKRKwffc6OQC8wkonutZJjH8Isx93/2h5HfMNuVlh1HY5viFAwqklx5vrVtK5LUcddRMnQTSTFKuAeU+K/mxvyzaMV/kDmIfUlpvoLPtJUbwnMvOo9FQQHvqL2u/ntC3idMOCKi5j89eoR+0ACJBLLEtz93jjDh6LhDhCsvLxLk8mUVvjurA5jE62dzMTKWTRee8nY+i4cxhiMr0snnWvycJnqU4Ov8Q07R1E2bQMPFM/zfNgJZR0VYWKhxw5/crNP0sHJys9T+kSbbA9p0Po91b4tk1KR8I87+M852AOhPvrUlP3kSaWwSny7eM0r+s+JnTkuEx2/tX1N1OgC/fUs/3YgeJIQjITLQhtEoU1S07nowPN6N0ARWeXfIHRebYRreXU7WCzgYed4NWkhFC/TJShjJjZEqxjoxBOtS0+u13ldx2c/SW+5lorGsVO1Kk/zmvP1qtUYydBoh30awUdSLzJ5FB7MyNVNQ1lyEgsv08mYmiPsvkSEWjvtAA9RRTk9EscI5KaxaDX2KeH/z8uxnfXGfk2i2bnZn/C+5wV/zC6642BvchenqPjEulL0lk4tyhILbmlI6yF4FIAleojIFEIdFiGkC5WMjNU3Nm+cy0TyC2PXpv65QTW8axiNQ2HrJB25X8OrFWPehhThVxCkdqPQp1XoTXgR7uft0hgrLX0EavH4QuWoSpvohYxHesoZH3/qDPTrGqOK9hN0qfqIga3D8iJGd2tY32LQS2dVgsOr4RyheTvhGwFxEXBdr0OBU5pxKo4Pn5r3QGijYmZXVvR+OAKtkVjhdH9T3iL6RMv9ebCpUD8EHqX/cgqn/vrvgT2qzM7tlzqAQLAfsdokXF+2MYfYZQVAoaloMteiYUEoZSolhP6T8N16RSWFGpcfMw7lfshWoSqAjQ6bxfKKFc/8rCUUUtyENlujYOdAueGxSXctcQigCuJsDhWww4TxwJbLV6/D4r++3XXB5vtBP9q/My/hrIetPVMHRKrVRkrnkRS3LCnM7Ilhdo5wunC9+tjHnFQYacRNBgCiI0zzhafY5LUHzwcRGRanynNNHQCLnq4Yo0upVrFm/s6rvDmQv1zO14TnvSNoBbgq7crKDbIMjxunmD8ife0gCmCs0GadJaeT03BMbMxkqYTvDAqtYMYwVWnfaX+FZPvNxwNp3wvmUkp9TrsJ/zhy1lwKbsWGnKY3qMtEs4XyhPYV5SD7LtXM68IDcMveZIvOJPDQPsyoMiadI4Tf/xHZA8AFErTg67TNhAAWYnzyOE85ImJsHXqIf1QjhhvVsbn+5a67NthDG0fxODq22mxkuUAJdhWsFNJ4APOoGKrqaI3XSjLI+10V3R3kMLhTYr5enBxTzwhKOV/cvc28B//BOALRH19BuzuqZmW/sLRyikFk/oBtCq3eqVJrb/jzxJEjLu+Oh7WuBQTvyh5GipRdLrOCi/4oYqSdbcqdY9uCrZu4y7L4LAr98OnYhEOSV9RRlIyZFjYTz2RG0OFnae8REBYnv/16gVF/GrCKRlfq7vJu6mARZV0XI9+mbiyR+SierlEZuaDsmZVKQwIXuq6PCbnvjT1iBFEl5REMLSsj6kiJSqAhG1LxNZwd8WxHg+sdnnmdP8stJiFm4HN58aw0Sppo69G9AhXxWzpzytZ187fdfiDfCV41jskbozOcLuWM3zZrqy65At1N9us3DgssG8+X1i64Qq3jQ/d825EVayLHMp8auCsNI3LrgZtqWkiOMKM8IQAH+5W/SyVQJ9gVvz4aAoSvOHhUpO4vQO+4/CXYKtlk7woyUtlnhEhuRWrdgn6r8+DLMNH+UOqSfkP6b8c8z/ro28KSnbezHpdqtprs3oqw/kD+L6ZdrdIT8Am/iFzyT3FcB7RU3nB85Yw+ysEwiAvq97ofx0ufYrMfAja2O1/xIppVT5R6UMNPpoa8jANBaM05SWXt/Y5oZCut4fJzXQlJbf4IIbZcuC8pHlnfFrDnVrkch4m/TYgv/XNkjdizOWTlSb2Yba9qoaKW0ckqm3lSRRJ3ERJqFPPetm6uUAefBVKLB3JueukanTucV4vc+wnjekRQwFX3vDHqVc7oF9Z4h/Fo71835iIKuCDKtwOyGSaJ9DndYOsCv0E68nKCiqCiRirIiu1MYCylV6Od4mWy+NaLCPi+6x/OzR4fcm7QYw7dkmAzwXPoJWg3hNHt+MqK6bRq9xIQN9MKfg4Re2Q73GeDwLp4DevHjnZ9QD012YIb/LBsVSvj3wF5dHUl5OnJyTzCm32+XL8XtasG+8fypDJGlpWRq0k+3+t4G0Ac4DGNlZE9gqHeUcYQyK68JhpMuQ4fwg1PUUmy7EuK4K7E5YFeogotZwScqIeQaYhg1fTu3YB64/ZQOVS6BPBpBk3NxhTghRnGD1BkGBvExNpxTHY7qt3L1qPfJ4m6mNULV+AqTfGvQNGidIVElmUyxB2/r+S3btdBTn34qjz5GuyIl77jSK627/Io+Z2wmHo+iuCARLQhrY9oOAxaloUtfNkk2wJEytURtv1dfOgJ19ZakV5NfAYgKNaCUiOF5KQ3izP1jwE3Js77Qghnr0qXoRIU2AThSkOrbIKt2IMqiCeF4HUE+9xvPmFBweH7uCWMLMc2tMd7dwxxhDr8gWh8jexMRbR5T1ETeiJOPYWfFGsAddCO92VeQcnP+uopbkOmWcIpZDuUbElb90yTh/LlGUZgQ10F7aZWmRGZu/9cEX80x1FsEMb+Mzn8yzgerPcYCjAHSXdc3eTfDuURhNElwCYDryTtvJ77yfJG4o8JhD89fkOZAmzDkC3MyLCrsckGCKCdYIqwmVACGYWgKSwjpLvmUW06FFtfwbacI/mOX7diNyt68HESXQWYaSuXwoNShALrmHX9x00PZ3EVdEFs0LlNugJRiEprCifz3CEBRRZhkk0m2L+LnlRVFZ25HzaQolZqWcxQcX/kqMmpe5LlkpoypU97SGb6vF28AOVWsJlV7vyT109lUGX2UBUN3ch+sgIAccVjtuHeN9fyOrg/ymOr4Um74ZwyAGOhqGhAX9+2usdOMDVK5DY/yRv2x2gWcNhJAj2DEdnIwFdVdfqQ/P9wjOSAM33uR5pvt7P2oEghmkBpg1fwHz0LEKHuOLZlDT1wLqJx6Q4uJ05fr3bHamGjqNGROUKvDVWBJO/3ddUV1x6bC27EQ5Tq3oSeeYaXm3hmoIRy+UjE5t+YSiAJKXcEydKN00Aljpxaf0b3vaIVSEAuVJfoaS1l9waJoW/8VKY4/r+DhQpxRr/lj+TLcTtdYu7RtQ/14y3VoPAVMjEzMnDlgr6oZA9iLWARoKVikPdNcBn7SVtDDG5gRWElIPzI0jymmD33y2vvRIAge2Is3V9l3LABlPxdMf8aHWEud7cZH8qjuB/aH2+PAglHiPzcsiwwLgW3/JiDFmYZRt5ga0JMYhPaPdXvra2W4CdqY5uLJXr8GhLCNyPYK3aOXbeleE3cRyJrLZePZ7lmyquIakEFhIvcwpZXFgf45MRwbe0ivqzFOEVAti5o+/storRuufbvtcLn6IxWJ8e0aafnrEONoCzbkAb/kw+pCo9H9nbWXTr+3oQiGJBwezqYXNxbNiacq5EAkFMwhYznTjpMnZRw/FoSiLFpY5wOpvkenUaX2ljXgv1lTPecpoOVTH+3XZhtBGRcHDr/AHJUISZSo5hbAn/7VwwWgOYy2QCGzN7Ems0psZCLy0X/CeQKO4fj3dn8O6zMAbDyBKxHtCQQFXnBe4yZwB2KlQm6H5t2obvpaEqrsfXAjIMtcR5TPc3RwaBsM0vbAWtZ60OayP0Ac5CKyrjqhQlC/YHvE3CFxq7iLOh7x/l2dJEjB2ijbOhlfJAyCr3CmO3cOAbIbas+JLwfv4S1NY0G5P5pby9CHo0EGI6qK01Mu49ymKQzeQZSzl1zyVRIcOFQSMOSrCuh4C+grCDfarj6Af4HzZYh1TI1O+hWPrIfbl4v1MhGr+fpahu5b/KCjzOStV9Br8Koc5a2MrW/Yk03Rpd5BxuPtjvsfA7AzAe4WjVsMQbiYUcBIucMD0x71YnYj56+A96WFy3IGKxTbiZNXtOZ/e8oP9wvbFUdCSe1j29WlqR2U5O1vEuGFK3mzRWxZZulGJNFu5fE8bwhqThQypcKsTF8jbBOQ1vt/F6NVTG6moaRPsXsCuktf/xBuCxSXyTN0PcwC3jDJpkCWt9UTudvTARiKAq89XaOBuQmUaurrV2afan2Zg+KihaHeWw6uSvsyY0LNZI+r7TV89ed8d6xwCz4ErftlMlIfCqXxZP5cfGBMSoAUkUPgS1AeiXiux5NiICh2yZZixG0dSoLTR2e1bHjBt3yRVshKoIEQV7EoLm2vLNMQhsM7X1SnV5TyjmxzmiIzgJE8hzI8sTLDnKAmvynfd1J5jT5MFHub5IOz5hsZ0TpWICxI9lMBNjGQdN15qGmyUW2mHhuCpZYvqOidrZmluXvVqW/Et07bLKI2dRYpSiVTUty47EHuvH13xJisX5Bj9senZ+infv/0ghJV76Ro5vKOGj4+SEcw0uOuPmbofnLx4BUyJCQTRn0LkK27Xc5Ib4oP5OqGUOHDYfMyiR3U6etWU+u/Nrgxm1EzV/T3FWR/NfPEF12api81I8jNAMDeGO0gToRUWTnKn6ZUiOMJ40FHmYdXrGyZ1blnvAgfLa3jeEGVrtaBk+5TjnkzdiG1Yw8O8rbnh5xukg+JcWTd5b2y5Dy1YVvar5B3wfMUm1prHB2sAlYrhi1SlRxtZ5kN5hTLovjacZR23USLk9BCgB/H587PbB/gBiHqD4keP0vyoGfnqFwIdAJCCY+8LYcC0nMigORLkKOn5GatJoHfzprfAy+Y224u7JrQWW/vijzBA7yHiNxwDcs/2ztxUxtwpHJI+AC2BIzFsb5VgHrqnoTGKcQpM1W4sJrJI0ZohuXJJ5m/OBrY8S0UJaz23fS16ysLpFvnTiRqI+etrGpqQDKU+2o3dY7hodYDyb6B1JWFuzCMWSTBYAjk6DcHJmrKhv+osbmlQF+DoIz3+5k/5eh4sE5jZmy96YpPDInpH347qAlPMT22rBnIzGm+SNhyk8RhniS67ExsrmPwubLRb5Z7Ft3xcNBaFWbUiP2dBtt8XJU647Sc06CrKMFkLVnz85lNpgob8ZO+kL/cAx/J5/kIbXQj7TfTWCIZXY61UoeoiDaVCXB2V3SmDhV4ECV+mwevCAMheXjHAaeOvt/gDa7Bi7Pcqe+eii/hIdX+W0n/ieWtgI/xPIQ4AmeLTzJJzYerPMl3cFD1moh2MBenEeQLh81pF7u+gxV42/W8y4gQ163AoBN/EA32KcORoLWy+rvWH8FYGhepYxjQ/hrvy2t3i0wVVvvZtv4f18r8txW33jx4mpN6S7P8TIzMcrIFycf/RoCN6BWPnK5QvBhzGbmRf+RR+A3hu8hI6ZRTanaDj4euLcrJDPcq8PpF5zgAfjVhgPYDgAb4Qp3ZmZEzUCnLtsVNn1C/9wt+BBah0slXgbcmEtNBzJpDTGa3vhfWIncAW6uhNSfU1nmKUFEna37fueq9IOizD9+GSlg4H6UoBVlZdrtT6aIC6VrsfNrg8e3tPa1I1zhwKQogDps+65Q6V5MgnjAiKwEnNR+PaMlu2fU26I+FnNvGksUTeLd+LF6WSNPOG8PpPhERnmTPVOpLgAg0vZK8hN1RLlbdbgbavB89XbiiH5OKYNbqUm+NM4102st+NR1I/xmUzOkhcdYsAw923ofDELFrpGDznO0s7BN534mTk1K3oBNou8umJuPxQIFPdak6498FvgIih+dqGPHIHxMVm3qaroi6Db3pxgW9hFfNFBR3khMW4nPjYzUdEStGUY0/3RaWrGqcD7q69BuAmLRiKq3eNWqvBudUFzzxFGpD8NMfzs+wsY1C5aUTqRcwh4ea/eJSyt6Amsgt70wjZO5JjW78whMI4GwVe4vUhgarcHg2lHgE/VuVlCpqJIqTHzfpqWHz/QqwKbCHZsbIOhanL0pQdgKmBQTvnAJAAPWShokClco4Z4rgzzqzgAQwMPAtbnlIrOLKXnS/eoPgIBXipUdoWLBUpf56SBe8IeMtpW/VI6pQYVEAdnbB+yEk9j76Bxzm2/ZjI5xyYKcxzGi4cmhCt3I6PnFks5xbbno2h6iaeO9rDLkqjL9KgZ2MXZQRNaTwgMp2k6aIPITssh4rTSsYLczSdmpsQEKyIipAJq5HJwt9+kASQijl67IFVrkaNJ4MFZDJ0QRdhmk/uY3bbbEmdt9wge9AfKYAJfHO+bDtw2PrjPVaduUkA6l17z9CdYbLOOoWk5h+CmotVePMUSKhRAURE/i71Gmphz5XWqtGoSBKgLiBw7CFShlil930Syd51XgRPmY03IZp0yHCFKEZWuX1JBLwbnXCGTEcpKTAAxqGRnHE5Vyd8vIh8JCZRgHq/KebE0/4jnpPlI9G7i0mDi2OYkOjsJekkQSmJkm6TFV2/G989xyfnD8EGBugeS60lMARv3AWm/2CfdGC8FbZY6vY9riTftsUfN8EHI8NY9JDWGGnGWHcR2PXT1c5UzbuZWa7ywl6aG6aBKgof3Pl92R+mDa8hHlvs8izwVbc2RwBsuqceb5MJEwiylEF19uOeR3dJ8QmAcDVx+Wx1lvBIhNebz3ZM2XW1MD+/ErfY3QIrpHOT6q+aextYsT5aLcC52Tdu7vVXxX+vUDw5MoVj1btj32TEoSsfUpXQs5XrhSzzuLcnqMQGhbrjI7zy0LIVB7VpQ/TNWMVe3FxROb7hsOsnm4p/g6blmD/OgTR5g5+A6Lby3kvchrB15slOTlayQaFqMvA1KRRxSVm7TPEomfcaT1AdP1KFPJxMtN5Kgg6Cxo9sEgA3jsA0XUpPWGBciWyaa7S8kcffMnEt3c5yyV5Kwwi9+i68Wf7hCoZx3TCb+yEpmgEkmxbGlM3M87/UGXGwO3M1He9JcNPwnCRbW2DnfCJQ9PMm2zgRcziy1mUvhBjLP1y644VKzR/TaoW7IU6rdCMPjndKFb5Jhxa3pJphw66Ii7xNP/TnEjAQQZgadoZ2PktKFyeiRREGp+8chDRSzWFQK398Rf+xTUJ4DQO+Mt3es8C2nHUyJ81skyzQNzNh2auTKNzqb6yW3YsF3e1ywhWmZlEmBfhWDBWd6kX1Ezmt9f7zKshv9xInTCpTBGrKPabAMNcPttvUEpaRGKtd6ZFVHV7Xl/ge4nrDjs0jynnpemxRibf6+UoZv0aM+5Uhr8K3Yfu85qBdjpeEnN2So1/R3r9fXS9kZCUea2x9wGnnwER8wk9qod0H1YhGOJdn3ymDatkZcaZQimpSKicSN52efP+lDZyv/FaHxhauIeMhP66cVjmkSddUXhWtxbuJnz2yVxunQeV7PbqM4cbweqGeYdYJ9TPRa4uPQeTFxgJMQx7ywxX6Mx5ECPJVWSc2ajmGTNaIhtcmnILCjHNZKbZZpfLJJD176emHHdu+o9Z59XmjIfIvwUaYV483xrhr/ocN1Ywx0BVsxR8RINN/WUIqfX0mpewHv2qyB5/j26dh/yOuifb2k2zwyOIQKmKbR6iaQekKiku+v21h51wlvLujxJTd85ALgrXgUO3XFzVfojxKAL5n+ozvor/UVBBtcY7oaPZeAfafvfLOoNX4aEKLzILSGBfxFR65cZOQnFFLIFi21S2kYk+UqecVaqjRZ0TiU//PF6HLS72GaL8p1pZDu9IOypINmyfol2JuzWiiz2F0wgGKH1y6tVddSxwnj2wSiP7QtAbcnhigHTUKNLWXpnXKO8G2eUACLJT3eQBalMKx8o8fDijlXG5bOGm1SgNXKEiuj8qXzOto6Zge7PPsjAU9+yB+8Xgoq/a77+c9ozFLWHbqOe5pEhShZuML8AnMEqWFLlHriZw2S7hZlKGp/A5eu4YJyJx2A9vdjEi72flo6Ka64S0yexViCZKa7wHjtHSGuYWTTu+vQZftEffeDl3tlb0h5D6mbA0xKVBuVxI2U7oa2nOJHdChoNREppja0PZE8su6dhzDerQ4AEot48+SseXcB5mXvqeDDU/r8vd2lVQYR/gYDXHZwdu2n68KPQsBLDPCc+1vDHsNJYN8XAX689Qa7fjJwuyCThTdhrNZq9kNXz45FV+um+YRECt0XBMwqVu2wxntEXpej7RT+tFS+LvRZQJyw19c37znrg0u7SC73kTnv6YEFs0GTxPrAYHN4eTln3Ri26P5+bD2WZopm8G42sjX54QuljpUHa0rrqrpMCWfrM3jmFJNfoMOv9Oc0WunJQWZA7fJUbaIRiDuz8Fj7c3CoIoX/VMSnfb5lrdJ4+2wm2wxQ3SSdjcVTHVU+u9n12J9RrwIo4u1nlLRymeKFP9V+iEmpS9qvyaJuiITspNW/Di1hKW3zc4uWwBLkNthO4VAkGPUzMehOi1r8ow0Jd5lSvORs9BTcmyXqmUdYWWwC8DQQO3m6hMMFPgv3wGunrd9HqQRiVOlGB/qorJXcFgfR/b+iqlHQkp2ylKF6xbXb/xfWqXNJGzj667s8t3kpPg8h6m9jjzYi29UsAjiyNBkyBqVK4x+xDsni3Ev/mYC9S3va/GKojthQ5xfjKVjA/dwSdV1ZIBEVRNrioviWUZb1pIlcYEvO1kDXzcDLYpA3JhvWeGEAP7YH1/c1zeGYtpXG5V3f2aVq2BRoAD1GzTokOSqoI5IFWUHo5kPn5UNMU6FnAzHeMpGSBhJwjYSeYwnOdkrlO+Uh1Fd/p6namn/f3g4TOYs7psud4kMXzedOIq+jgvn+lJwhfkWFSxcdDP5NnxK1BeUPsDYrdqAKMP6XUOemtJa0/OYgNeQxhOmqSeWoCZgoaNpcZWmdLdlXd4Y4RrISq7bNHHbAYFrN9Q+2FlzeVKCwIHJgmAIBw6RZepvhK12jkQW7ailsuI1eRK9A4+HyENRYQwGGhul7nVpEh5GOYQcYDvZNfExa02VJHHfd7epGmKDKj8gGWYPuLfGoM+3UVtBs+1hcBGuwfjJJ/aTXZOHkhhd8TT3cjJ9ME7HfoYAlFkXqSL9+h5dixyfIe0JfYvyLIVWnWeDBsjE/oeMAXCDtkmpOJSri3rI7LveVZ80mODZOE2F8Bf1Bo2X5GScAGgsYviVjtlGyR3qZraT4Uzc9JYBG9Mw5b6N//cfJlrCME+fO8e7PGe4Rc3KTabAaVLtjNyxNUF4O1YUFYn2ywv848cee/En5hebiy3vMHd3Pyb+nOXnjzE3cac5v2QtPyNosL8JLEEIHeFpN1EJ/QjIwRPf8qM91Km2HMF5pDmJBaF3a+oCdrlzOlVsQHm/Qn2Bw3Zeou5yjRhSR+xo1hUa8eylIcVzWby58U1yzTKr+mWW2I8XeLru38RD2YwA3ADee6fCiBO/vY84eehOaeThJMj62UEajMVsGOma98Nn1i1W9bSjaOZ7DEXCuN5PvorU11mxeoDAVrAbk5NUXt+SbEXYHWKbNjig2oc0q5GFLGotP+PUIh8amAe0qCYAbzrNaqVEmi3mkmah8qhbEXHXsRKQMCFr2u0mGZI0w0NE0AF0uYApe8QXxkA68jVC6Caf+qHGfdlZO0DsoBNbblBudxEn4jiCye054L2fWTA+MMD5uG9CSJWTo6JKpuHajQxPo5Ir1eilOtLbL9EEEX+7utgeOyajdvl+1qWekUGfgNIlpgpbauRC/GUSnkcU9qx/S2jEJwsVLMS9x3bgFESKcvgE+QrQo3QvIh7bB1MoJ2EX5wRz1I9ATS6t7ts6MeIItewjiJl1w3ioQmElFFmMr41/ILasyO7HWSYGZalsobbbF0G85TDIf8b6xVLKBbEIbesUp9KY3UuKpvYWCPWv2VcvpeQLiinLhF6gbqE95o4r8x9tEb7oFkFEgnpzuh9svyHJvQECmxSOs9hTyniyVJq+KuGh/mYxY8KSh61tTPkWDvHk+ONKdyz+Mfxl8j93OGqvBqdC0L9uL2mY5pnmSt+YN7kbZIeJ7do2W8k4OUostJ9SkvqVdrxnI2bqhLOb7LZhsay5Trqzr3HwNBSHCyUhMesStexhgL6rKJnS0n/X8hCGavzt9nJlai02kO7ZseSlF9uvqw99nx2Rj2AX+1LgMSSnFpRQcqokkXgZL7VUCpYYIfsAQGoXCMgztwEByf2WFjZy+lpczpmdCRNaG2Zh4mtyohNtp/WdZu+gHxlDVPHWxtRa6uNEGd8ORBCPTGD+VwRuvbbXtbKaEYGhkbXZ7icuQnlISyLNb9nEgeK5ohnmE8lQVj7hH0G1K4OXlz5H0ItJ35Tj1NysxvyP7zX23l2FXlzu1pUuBhEv7UfOcz5xM9Grb1xMoTyu1nH9nEKYbMfiQXRuphK/6S8b4mtlW2oPELf182ontsSLAItDtbHfPBc90cJ1Hy8mrWWETOpmlymbBGsps/ktUyGQ4RJYNW25gS5T4GapKaXLGPfh+UxHktFuryNaXbYF+lx1JZkmCbT9rAXGWz2TeV0Yoc0HYbNQZkMaCbI3QcTJ3GhNzL0X/WlCuESwHbmZhfC5rstdH7WSdHWmSNrcuplW8vBB2RDs6WtmNxqiyi8m+xI4EPqy6nGHFzVh9/Gpf/EgdSQwEn33R33lLjB2kipZib+vSIYc57jbgw52bUBnNbHdX5hjQcr6li8WbvCKoZ8WWsY0h5hmMVJeeSpNziUeoBy417sguGxfOWmUkesf3qh0k1QCsistGXWFAUH1tywG0HFib9z10R7+zn+nwyU1uC327B+PG11ayfHPR6fjbjbTTFiDiucD3f0YABxPAc5jE6yiuk44mIO35LM0meyicWueorPfcNX/ftbPHPEDizUPyJ94IwX+iRW5JVCklAH5yBCR8KAJtUe7hoNOn2qnL2a87jezM3E7JY1aztILvDDFP383/s0GBjB04wKbruZCDMSZCfFevhpk7talyfGvfZZTQLN7m3Y4w2FyV53OSZhyqKG9Q81KhyCbYoeWKUqRhyQYb1UAd5JjWHWn1ZTvZ4MnVCUZPM0hQOao+9K36noBxzkUVqFCNCaT8UfwIVM9ktMYeV1C8OKFaPNSZdqPaSYrk8ASw9N6zadfBxvgXVqaYinF4+DBwtvjJ8BB8odxqmzO6bwc0ld0Wga8OiVuha2RZzrog2oYRlqM0CiTV963E0wB7SQsHxocF+t+F0/OjLYXFA4ESEOszicsfUR9cloptqoPKduFiqWdCq9bTCBqf46+08aV5uqF5T2umuYwa4bhEzEJDhXIgfLzAXZeqkHa2zXFYloXlLkK1Yji3ne9ih3jwHMjhcN7JxKyjPYmEFkt37NrbXbWmq+vCHnLhw+avNBE7nSTD3wOmzRWiciZiCO3LCcFoEk4huXc9tIt67MhUR87xXnYsLrC72SvfG7om36O6Ini/wvLGxrzwBCj1cZT0hjL/DaWy3OTT7turY/QR+D+itAgUXxhvI1jKu0jV3geqYx+IPjNxAlzG0udiQZs07ctfWd7oGMuGVbn20sZJdBkLwJrubcTRjsCb+NuX2lG4IKoBcN7cW5cPpwPrctPrYj8GxjbPpMmiQn5d9DOeDQ1KHjWob8tkyh+rqunddwDp8MZGsOWXkH6Z/z1NsWmKCFbX0kQlvmk38DOpF/HeeHuXE8InkWjmxEguIRA3i8//rFWtsoDwMlpg82zsQ/2+0Z8L4I85QF+0lbw4Cf8OfKqc6WA1QCelNmdBide8QBn41xVuu1VaNhbCWdmRTh/ScB8doacR8urWACVuw7+0OtCF3DMBe+nd+/YFhjAdagtW4tZnQo0ZnJP6QrN86trffw9oSu5VK/YnweA1GSirSkJd+ymJLZ9IpM0RnhHMvMeGunaBKQwVnq9ldN87GamSNnzUsH3Fqf5DYP0UWbeWZGLA/IzolKH8zIRz3KqQgglnidCoNWZv29FOUuBkNsNtTMEn470BItgaUmz50n0TB4H2voMEsc4maNTLHxVsK7LjKmVsXn0CNkL6L7oeR/GqFIBEh9LEz9EzWIdlEm2n+QEW3cIwgQ0ucgYfiD1qfRPMjSpWuUmJdlOiz3kaXOVpcQaVR96hzCDh6g+P0ZCTXJyua5EIZEiY6cwxBHg51svUkP/i7Qu3GH2qRpUcc4XAQ1KDl1fkqUIyFGTxfH9CA0uNWbZdJkGe2Ae22W8maZzbDJuBlXK963Pgg4wYtzeQRaF3FU5PLFwI6mkIiLCJ7lGBV7hFYFufHIjEWx45d/m32xN7s4Q8XSnr5WQczFPjhuBRbRFM7bPDSBOKcQDh4/dUVDTXc9kx743aL1zrgc2HlyTfQvnKgfic/U3sJHvdAEKUo12zQVGRFdjR8/BF9KvgcQAhAMjNgC8H0LD5H2aGw01w6VvVfyODCO6qO1eofm2wI4YU13QCjuPuzJ1aBtkOZsFWQZBuIoUiK4qUJGIuRTpr98xMGm5HWZt45TSuy02D7v1LO1lg3kw13ImxvJWUUcFjdwKtRT3cmAYb/WlhwnzrjWYjdLUOX7U3GhbgNm70l8LKdVnFqKFD2QzIpY1/me0DlIs/uXUqcjVtm8/2DmOhyQiXwwZGt6rH9KoUeRPVQbJZXRZvbM0UgIlRYzMDmYbM4qV1lVFiFBH7YvYtnordyXo9KY+rk7H53qeMVmfwoDucrWSYdZWnFG9K8xGUG8/HYWTX/KTBUCHLUSGuX/HsAHZksiIQ+lyBDtBW7VL6NPDFErlRViSVBo6SVQr2IuHtUvf+vZXu65uxRqZHiMF3nSaDbOt97U0UbNuThz8oL3BndT78DL2NBqvXSW4gujRyrtK/VBahqc8zNIzVhjgp8I7NsaxJ47pt40Y4D3FPi4gWmI0U2ve7R6WYnWGNLyrHjuM7jWSSI+wpiMDNHY9d5OXEDXR+1xDzCIVyA6IpZUuOXQLFXYN1N1zzs+ELMg+IR4iyjBIlYN5z1SCoMrjKyBcVL6iP0CQuBN6K/IoDenLbBLXq/iBSEMuNwx1B7U6u3gt+Qagzeb5HKzGjGaj2I3jnA5ZGLhsGl1HettMkdo6+lH1Zu+bhjgD2rDQz2wlnQ5JJgoy4AH4EOyfTkbJujuoa83knsxCFlrZvxEZmJFKmWRUgJ8BT49ARaHF0UYSWcqMN3zCIEKrZXVTLTAEinArXtseFUSXjgau1bKhvJatI3NdTNeeSMVlQnEneOPf8/FXlH7nSI5inzQnGDpy1aDkN3A2WqNxjNMKz+SxFZzahA8mMdQPv51vzxWDH7k07VX5C3CY1e0LqvKVgsB0fFPdy9aGlI2FQq4m/Nc30m2HHfiv2iEah/2krYAOBt9YjQr0JXihdpka//zBaOItp9epwJmdPOHt9+e+2rYxylI23Iid/1IyFu3GSZJqUn0vbhvoR1EbYP8Y5l+0ZIBrVfBt8Geh8y1zit+zY666tJZs7jHlvDzSHfU2MghLgbZKC3nLZ4JtetwglJ7xoGyD/kvZLfMu6sk/RgwlIBRK2hTeoUicu9ftCggrCPoc6WePVWufcKT212ADySHnPwz+DKHilAqJTBegnEVm5tFyTDiEL5MqqvDg3le2sbLIY5MpLR2vIe2oYlzQX/nuKz3vAgeIpU+By5NRD+5F6RPod3fUg6bMV3RgpraGXef4dSqr9PnA5NSuFIcxM69Ajogxy6m+Vlv6OobtcpL+h7hxKfBnWSYSx8hk2Lmt2+PD3Vf0tL4DHPp59ncgsEa+vkG1dypCESrTPoEHl1yO4xW7kUbKUxF6GqxlUhOt+JFXDMHZvdoxUur9zkS3iR0qZy5Ivc18i+dSDrrim+qQG4JplR1Cd7OdKB47QUri0nkDETn9KWCfeQlqvwiaQXaVyXN2wQSRbxmGG/tso0jQ1asTNT6nrVe139V6d8/FBO8Qe1EJzA8C8JGNUVCmRYrvqwMEfZN/4SKYHFM3Rg15YO4P+xWJxaFq+aUkh8+ovVI67laTzZWu2nq4iorBNGwKSa6m8eW35gBT9SI/Vw2hz2qATMK4KCPAOjJMfzac7JNR01V9+xTL4iZR9dK9hFuNtmzS3c46F6NoGr3i7CqWnIbBxTpbWST5tRJigHGowoHcIibgfD5hUqFL/zWglHHrLlTA2aWsqZZmXGakhZq4/go7fQLuyRwjM1pwUofxuqpegMXm3NhOyE2k4aG2dR4hpGEuvHTunWS5vhI1ORV+aPnJg03t1JIbXOlITHZsKF21J7Me4uhxc1q1fzjj5xvqcF1ERlM2Cj1yBgRHBqWWDgcQfc/c8WlBhJ4Z+yx8L6jiiLkBs6Qi8/ywpV2OOUsdcVVymG+IH5za1dRMBtsMV92s9F6Wu6XxTTwUCCwmYMhRziEo3OF9DYsMoRf2xNkDXk0ZNh1YCf+PZl/OnMe0Ts5IdUBeN1rzToX9O1LOgcUVh5xLPtogelx8JJbueAch9FAx5GWVjwyVbGBhO1BK4q2gsplzVYUWQ2CvH6CvZcOxQWPGkm2UnimYp52ealQWoJVsp0fujNvGQMILztF8Vopzc/GD1KnmVoWAK2dh5lTsb628FzHlZqNA8nTkVg169eFXTf68cVJ4oU3WxmQmkvCFJqz41MPXNyW1UK+mPJCysCJBqdrQ+n6tw349sMNdbgufsjk3i5u+ukBxuV6t7ynVIVK8muRYRni/RDs5RvJqULXAVWZmtkb+2ErgGBCxiKXHboPVfUS8Pql9CXb5O+j+kDe3OKbkvgV/3E5kzV7esx/gRYByoKY/LU1iIuTCxJ+lGA4PQL/27vhncyBJoVZm4/dSsGr8SHsdBV1K5o6TDRdJ0ezAAe2MT/Q3SYRn/U5Z+XcrHYyWTX2Lq+DgTktlIspwOQZdb6GpnE2tRRqsi0oM8Ul9AbHelUtBFVcQqtSSZ77/AXmbiWM8LkBPzIQrwPhoApXo6a8JBcqL76Hz82ECDZ29LgrEVtcHMcqsRGP2Qkjt8rbX8bf/1Iz48BtJa8tMiit1L5BaeNfdFk7QAUEFaIbNJn8LeNdTjU3+sEmLwHa+2j6daO8oGQZpiAAFbSMMEwFazvfZfZcnbh57tHtrygDcI5q7yVHh2mS/ceTivdavqRpYnGBNIMDya906d9kre2FRhlYJpxNdmplgQ/dL2Su2sVnAL7w24cgeEgIa46nnOVUHlBmngmqfPGbFFfzWeR17G4sx0q+vg1oOj8yotG2Jmjtg58e0SOd9V22O3XEfuRbOMDGvIRPcTlsYC7tr+SwIGmzfpILn+AP8B0dbEdpgNnNllS2l+Pb6l+mLg2DgM5oWSF0i0h+yPHtSXOLmiVpPa9Yc772TmYRA/LC1vufo0qxgMbrp9wYZeVJaOEWkckTgdupC7NeEX1x0qGQFoT4QyjU/k4BlTFcFM0HhqZlmmSGrLOIYW3xjqNc09X4mRcYPXVigovBQ6nnKMdGz70uQA7DAzfhr+jEuhhGQ/pumNw9RSqJ0o/OSa5hx+kAwJsJdYRybFxMlU8OBZ78jBhdfuqOw4n5Ru7v2ZvTneBzPzzMOgAXzu7ZdOHNwl87bpBXKiSYGqcFD9GYIyowv2y2bVlgktT5qqyMbTKKdSimaj1WZVYxnOhD3CNjkQyLSPQH2w9z4wkjqHN/jQfsRsJ0dGEE0ETD9Yc4rRx7VpEaHg/mUdX1tsWnncR+DEarYxqHcT3+DxxwcZrdu7fumhaKpZ+kfuERcXI5Kt7NuaK3P4rkGZv+nNUDzlCi7RgnECZX+Ydp+FSHpPIzSplpVV/55V628xM66zNZ/kEUajU/JS+IHOcQf8qtRtYckoLLL9D/75+BUQDlSs2kAq4kOOOiBvzb/ZK8kZ5yssBERJIFZVNkODZHNQ6w+2rHO+lBFF+GWuKck0HgUjPoRKqVFJzWGdTsuw/Vu90cq66YXHdO7mFFcgIYnr9n7pRpvk/Np/YI6r9Gryld98jpCFAPxX9QvxfbqfYZUmMe0x/SPjy5+v9nJHCnmdDESEO8+VUNuDezzsYI5lt3vy+zZJeOcKz5QKkXA+Dt+72qWcnbAd1bHNM3k3mC0m3NlK+62KbhaY+dmBNdzOZycKZGrGq6ewILjyBjesEn46DxrO4fdekg90SqtgcJuUhdvloDAAkmg2Np71EikQW8x+Xdl9l5rOl2CUKsI0OT93vLnqjsRhSMbqU7lhJ1OCxbPQBgImjBzkWIcZh9utFnkpit+dBQ+fWZNy66KudzWD56VC4dxAh4dLG0+VKAA65Y/DANjMmDFTWSFfwwm+sbpg3sINol6+vC5X+f+aQsPK7rD7ZQfJ1tg5e0stjdQuQe+lUyLW/8MZFqGksq8gS+JQezPJGM1persAnXyGFxxqpBaGv6PX/lZ9iMIN5VrgNwzlPhTquY9W8A3TLtUI/SFdKvSAFmRBeLlA7V3vm2aRMut+m/FD8O/8o1gnJo+dYKd3L1negOD4SejY9hnkg4h5Mo6rKu9krG6+Drw+B1njVY0Twzo9bHKwiKaV/U/cagf2EYIWSxlES0ptZs1sBcKyFD4SePJKK3PBttH7DtdCJvQ2EsWc8AsKW2Hm7AAW6Sg6s92/Tu3ery5nQ3vWVdZf8X9PGWlyDDZ2uBqEKuzaxIKS5mAivyZRun5iZGKql2wPuQpuQ11JZieOxw5r88C6dQfzJWH5Zdfzh2pwve0a+FWYDRRqb69a0kqFizDvEvOILLok5VXJGIzbZWPyLWgmap1yLxHrvz8e7WIWR/viIJ8EeaRCelYxQ/tkvI4t2Z/nB3BS249ePizjU2oYLN1Bb7pjy2/E+LA+aW8zHo3pDIXAF+nv6eNUmARObfLz+m9dQHa7PP019lihUIAzRj6e9+4SW2N+XvC+eg6wIVTDjxStufDxPzcYPDUVEoWITFZVMe1VoTj7TKIBnXOJZvvNWP1BtR2+adBFDgZ+oU6juC3NufyUH3+Isfi3YaPU/F1/njU2wJa4IKyEOTGeiLDAszeoYn7W0NaDz++NDXcF/nxjtHtsUDulkXsP604N3nMWrChVyvot9ZX5c61xyf51AtdE0axr2+iUlRD3V+VoBfqUM45oquhZT8VXYELXkd2r/fq5p2juXYis2qR09pGnQdXeJ4qFlmiUJNIPskU01fW25jkYkvQCpcsUm80962XXi51fzMy9ZGgJAOQl03axMO2KTqNoWrg4tIpE+YMbKlyYp/7Gy+xyPC4xIQLeIg8s6oHOSIqp9sTTPXncJ3IxtufILiJYS9vnil5eaVt6qeOxiGs5F0ufuk73vKZXhzjpmMGnN6jinmSmcu1Av5a/QWC/V4JYladqg6iRIWfXp5Xg2SK/xXU+kjjFP7o+nEnKxBUhlWlwDlQg84TnwQ5YCmfAdd29YLhI0zy8o/mkeA4EkWIH7DnhmLtBBPJoxMomh0wWJ+L/XnOAlJMMcQj2h2khKX1uWpNVFEExkjWXPSkl6LYvi2PWbyIabNiAhlUuv6N1a1w7dm95I+j8L3SkMByUd0IeCJwXpUWRFebqBo+MWnj3BC948wWq+LtMgHbIlsnbZyfBf/+x4YnKsh+ObvaS+XOiiVTdHl9GvVHM/1bydTNb+wOl1XFexVf72tYYWuqUL71RbH/4/JrtUs0annrzrUhnsImdtnX5q48Nzg/pdkPzFIqolcDJHHNQvrxeth9Eh0H1H9y64t53GYUH30v0LOfgETW+o7lEVEx8JfxChb/DSo4ozBTGbTe7vF3dLxzM9FxaT5egzROTNm/wmAkRY5BncLzy2z9JFekY9CBuZ+Nva35MUzI2g/YZjbFGta9k7LeSI+BauZgsT92Vczr1hlob0W0fORemqL/3fXhe135rXhvukXL+wDDZPY4rNmPEWlYb9zsz04UPu5EXzVET1rsmkaTOjx8GyBigNTD/PhhXELU0Q90ertysNXGqpdrlpAjLDXpHH9aqSeKyFzOdgzewyvI8yYitzi/11tTMEHUxMaChoa4chaVMro5kOEetEXf7q49X4KbfWEz5n0DRsXKxH6oWHy2gR5Um6uZ4HNPRjl0p51JhpCDvT+TDdZ+8THYcyQmOH2sNw=
`pragma protect end_data_block
`pragma protect digest_block
34b860514a15a207d6a4cc62747615c1fe2a9e9616920c9fcaac73df1e05ea4a
`pragma protect end_digest_block
`pragma protect end_protected
