`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
1C28PaN71D3tCffwXfLlKXt4xJFmJmn99RuOkWAjN1JXqIZrTgzTykoMf+Es6knoI7eHd9jzKQtcBMzFedgARDxmts0F8mM/0djNpFxp2WZuKldi5l4y151cH3OhFayWfKesTzYiERNqkqI2eXCI62OjH4kkqEzb/6p4pY7EXZVGtFNqS080bEVdYjOfL4NKOPJ3z4WqL/0++hQ9fzd4Y9RSM8bug1uTck52PSfs0rmD1zrDx28xvYipwPXggmfng7uixR16wHUz24Tz1IqTTXvZLpT43P8CBgG77pQSXwTe+5dC4fL9EHG//oOH7hok4P1LgQupnfk5n8c4QldmwCyo3wl4vnuWWQBhVoww6OPwJm/nh5+CUSHO1JpTT8O7CT8ZzwLVt8YDPl/qmLw88omUkGpJn+IRZZnSIT63rEi7SCuWvBrc6+nUAdv3f07HGRRH1cA/ERdsY1YFGj/knYHu+l8wcoiXfti1vdV91fb7fxwDW6xUrCaKDBKm1eRDStT+lJmhcBCEocEDkV1hz2DIB0+XXGcC1w3LUuPCwP4BS2vQdC6jBqz+9UuikJd9vgWMFswkqVSHBIjQ6vcZbVdAjuQwP9nuINyXqEQcpkoL30VKyWI5zyvWJlWPft6C3NvygDJ668CY2cUUGTZ7z/r4cTXOuEHyY5fzwArb/TZvfbGk9HbYK99k6BJX6rDPD4XexxUJnAkenxZVrTXCMmx9HUuxQSZC/U6EBze3YXDsH8O2tZIQS5894DHXbZktTnVVy7EQCY9Xj2op6to2CHv24POnI7iW53dDKbnbWwID2B71tYsqfg/nTQz8FYrt7ruKMZY5XXKkvM5dAMWJu2h7FLkcmO94EITb1GwbigK5SXw4JwBOFRzcJHWJ0n5qLPvy0oQVf1Vo0uihilCjOE2yqHLPDCz7qi5IwhDrqhsd8m17ucOwibUAg1u52z0Gmzk1myF8HdpVAd1WFp4ZECXKToJWoY5H+KDQaML4IZ+SSoExqsM+gt6rgTp9shvO3aPhSHN/tZ+efQIWweOTORdQG41LvQ9nzoAHSo91QmuFmeZYTYC1o5S8l1LR3aaaMmuvS2mMvwVSTR7RrmOgLljVCXTrx5ajJlBwF9URemufidOvtY/ZFkslco/N3Evkn3wSNclJ9rWgxkhyUqILSPYU1HTiC7pbgKe86jd/6OdAYWWjOugNR0kWl+dVEw9+q0Zehll+UsNjQ2ngyySI6liPQ5MqNPCSq3cskET0GfvqFfr8BRQSjju26T9ha7OFpm0mMWU1/e39fSk4Arhp9q4xuD0ze4bcDDq8VlziURtKtlSWKtQQEBgO3furoANB0XUtxPtWbyyIM7/inE3Qk78H0bX3vku3ZGowzzuRt7awbbqFeJ/sTcgPGEK/CQMi/vlTuE/Ipi3+mLuNpxH9YjwQepcCUqvrCpd5bETiyIxohNn12JasB1cwjSlOSh1HvSQ/yM3wDBgswbT4Ke91eMEAQ3kWNO/sbP3lsN9FzT6wVCHmkK58fbHaQwqqQN0ZOxGAQN+IbA1ybHWM2Je8iM8UECB5UQhWAdsMrNNOUKlwuaxAUM73LzVIRYKydFVgBeCNMMuIF8lTJvLILkRZpVKxhmiZ7iNc3hf1Xgz7xog0o5yn06GMJU6pNfgBfEOJSUpgjShtFgoOzsuNFjEOeAFPCbOaGNL47sIdcJX2EWtXevRdaxToDAfnNwwlMZSCiap/OS1hOmuyQq215ee1IL9S5MXA/yxhJnozYbGqUVL3Gigal/OJjndmGfp2ZRs425MY4p/dJ0VP6FUbMYJ5gj+0KWDtxHqQtHEnBH4Z+x8EjJWZ1UCbsXDpkPM5ZKXd2yaKs1p/Zks/Mud5gzhCvMMLILugdwPVFutZav0P/xYz3cg1XI5QmXWOBGlcg1dfjviH0VAQZby0TiRJzibcSgrIaYVPxlowFgWQ5e5J4AIMC22ZixucAxDumjNN83er72/ySvnn6YeFOHJlaXF0hG9o3ldNR4FY5jFCuCDhNQ0d4RewX3U9iZWDKOry2OLZ/WU6eYUUbIglA+Q4HA58MwTK6HPHiYiTh4lkWUYSPJkV/8xjJ49ouIwvd1aP9dtqK99KNQki/PlYbGqlO/oZ8QKXax4wb/KdSc8XjWbjm1d3G7zmwoKfNdKGByV8zP0C4J2FonuJ1q3BAySBLLHMK02S1Hu4HKihwm2pvTkUwUJmubktXvsrG3Eo764LeTtF3JIIcifusyO4TiDh2YDxisIhCuaSDzGQ6XNgFWFXt7Y7iafwg7rW/cGO5sOTeOHYazgNJYnXDo69Mk0FeuMJZ0jHTTmjP0NL7Phc2YvcMVXtnEO+NCBC6nmHQHzlMvaNALrkFAXvF7D/gHM93mJI/JcicsKImp/ob0rjUykC8/h7ZVCT0QsDZ8wQi9JDmLULjj+csEd3eKO4z171q3mEE+Kh4J3jJ3ofWqGCV5aKQRl5138Vvi2QEuoFKX35phm5S9V0CEGmSlNciaLy25TegW83/anDX8vjAzG1bwVHmaKr3KVJ3sE4OdYQhpe9q1mc5bGEOijJpxr8vYCyQ58iGi5SrZUer9dIf6CxgjoQAMr2YpdOVSy+K0FU1Ib3Rm3T40YTcB2tdf/0J4R1BXo1pGyH0L50g/CRZYvla5dvPhWDLhPPDjxwCwb3/xElT7o7T2L+oL6+Cp3L31IaBoqp/B/WF38hZLI2ReMsjOlyd/Y5ZbftmwZPPGsv4koiMyFivFJWMD4UxBw7fkP1HlJIPitLMwYcrIMoAjN87oFLGu4WV/1iXL+iI/2Fd/f/fLlar0qSYcXuunc2HT6xSZspuXrMFQcWRZPjcNUGabYi5lfA4PI2xuYAwR2/KrAFXDOlEK7jzhsjj0B4vnCCiQ+stJXr2F3W7RbmZ55HFKROKrByqI8ECUeLfKtDa6S+qWSCdsrm4E3ueqqqqanabz/Ed5/opN/sRFbzRO8cPyO2T9gagQVuN6Qz2/BvdNSF1QpDWI3vIwyE3VkQ7Pxi9o/QxsoqKfVVTJ9wLinbUfljQo4nogJ2LTVL+An8speaKStwvegcrqZqHYxRVDQ/2rAHaH21xf78mtf1jvJqO+HD9jycqFt3HP4BHGh6BXALv2QKcmoi8WiO4yGS/B0XKKzEBgz9T4BwutoAe/x64UvT/9Y9EALTQOFVDCabeOLBnhSaXrHmL1aIcPY7bPlsKxPHfTiUsYLGxxQme7cSmvlRXQ/PcZ1MBQ7YV1KypO4mJtbbn/Yp4sOXOtwHZUH2RJWZN0J5EwRCz/94mrIw5qtOEUE9ZbjTc8pYTfljKo7E3cCd6Q1zd8Z8w/NEbsoLRKkxu1CQTItu2UlrX3JPkQS7t37/rD9DwLqutMzhpHuOZbYqqDiaXpkAVY3WEydoj52zRqf2MMAF6hCltZoIjBlZL1Dw2wj6dAP+yGIlHYQgRxTHFFC2hWqzuDNfajYiCVfhkBFEhVGnuK0dlTgwsp1rFFJ69rx2a2zPjDZBQMaALEA+oQXQH/spLnMeaNYiqb/SIQsQ6cur+mK+efUe8Mt8E8pSgfL6CLuoBcfJsqDEtms2zdBgGE5KxNvzivd3y32//bYitMaWDY8M7xPlNZyL2QpbI3ErXt28evCQ5oMhBgmHYjZleQXaIWZ22M9uG2z4TMRNETM4cS/c6FHB5COM9IBdDwRUVRUUQfEEY/w3FVzsdkZPMORGj6Ju4u2oWFIP/Bj8JZOgKCWXU95jKyywC8SFplm5Z9XOe65aDYWXNwnv/IiAvl6X+MloftHuAV2og6S83gpo9ZSsVcpxgYknQLTa0e7Wwgh12+5O6ylukRB8LOTKQN29we3QCuIqUE99KHZfV39+n3pP8XncLejRy7kn4EeQlaxPO5FZJ9tmVYAKJ5zgU6ifu4P42DXlRdAGGp4VGPslpiXzVscUGl7EyrQMl5FMToHR2TlRUZQ8VmcM1QfduqKV0kaJISE7qZLhYBVg6SXRE7gNOYmL2i6edzfUJcALDGgAGYHIJjsxd9T/j76gdAbD3gTt+CFpOkyZn+EQSJVsdq5M4I312AX6rtRKqnhc9BN/0aSiE4XnHmTqxATwg/Rwtk6J89UEug15MrBYBDPGOCTnFa0MoKBS5wICFR2yQpx1QHIkYJAXMgRpqTJj6ktRLwoC/b0+IK8RsI96vaLsPG++hYnhB11PGAzLWXIWoW2vHaLuybRM2W0gyf/W5t7Z9J+RE3cg/XyC51PdXJGDjTrKcOYCQ9tczTC6kJlxOE8dl5VsgK96Ea0ajFEsUOVAMbgYcXLNTO2ZAf6ULKXXTUgqQIBKAHaGei7ZTZxLj6LWcAC7Oi+UQFLSb7CkHlYgqD42yEgOVZa3PNxNmLW2qQ995Wotuv3emyMI3fmFXb48tXiGHltm2SLVOXip/LGfnW87Dtt4OJkEOZiVKJM33J8IIqv8LzWqpsmz6FcogPIkabWg0CHkIKF7nTzOrYJnBeXfR+12rxLaeIWZy45dQKp9NrnzzuVcNG5pcEcmCozbZb8eKDqmNNUYWs66VOMThC69WzDq2tUJfTJS/TRNkvntmY9Ti6aDLAmIKAoInUODPrHIkX0kKu1O+AOcdPcluT3//HugLxPnIaVCFSMK6PsUlYQN80wfe6gy5CFcgXdner3stCet/3HlWV65abw7gsQPK0lPSycYUSD5cSe9vn1EFAwHB7dEMAnOcKGMeOd45CVyvG8H86O7T9tiX7paTE8EaORD3fnz3RW+nD17QYEargAOSjBjjY2WatizPFO1AZdVVEf/pjRHr6x2g1Oz8/e+EmF4hNxRvJIYv7kj8VBR1OvyqSBZRDm16UTLaAmLCtQrR871he0LtrgiWBNCtE8R1MuP+3zHpS2AlUeki0iwkY+7Ml5m8S3CRMufCdhUTXD9bYuBPsLvOfwISCe50JnoF4/QTFezx7q63aC1oqq07NjNIIJzNZF/K6+vHtEMiKV4h2JE1x8c4avSOq2WVBf0VrQcqoSCpUNuffEHqdWYmrPN6gLGJoC+xlLyHDvBPCOPbjtTrDid8xrsR3D7u711gHWSeSTPtnflTDx62dUtySVTPG31tcX+hmcP7edHQ7X2jABcV+5rK07kWMmn5jHFIBieY1qyElRhEZiFkzFNQbrvei4bg/KrXPZZr05vGmHgjWnwGgXkaBjCTSoypbZr+uaT5bTRnHfc0UdE34kUg4Res7L//muQx45yhMGzPvS1g3NjHwE0wosv1cf31jHWSLLx3gNKnpOylDISheLm05y7LcdrdeYx0++IpaQriU1K4ngruZmrnLxRycmj05hLg1L1T1CGHiHEGU/ikiAi9UU0giEhK6dt3dG9pb5/LOH5yFnwPTniIdZGjKud/LZwjRPxs36Pq8lvh06unmtipUW5cPYkC8tlAcDImGhTiJssO04CGuCVKGAlOsuoinKZNDZIj1u/6Ky6ah00pqJ8ZS3UJzjdUMXAw77X/6DauxKU96P8yXTYAE5NIAsmkfL0cbeEQdar819kfLHEqFiRBLX9+HIeH17b6iGaHXAH3xQioU5LtNPpiq4apFfifbRS2Ml++Byz0z9Y7n4UVrOkapirt10HrmxehuAe/9ExECB2V05Krrn/8jEB9PQMqG32qVCapq6LDDJMYTkBnIZHxL/GeHuWm+megAgEBV1dnzUCrH5EhVi5w/BXA8fOPkdJ0YyOLHkh8YVMqqhyopLeRR9ussZ3b/1uTyMRW4EPPN7qtaJqVE6SuPlnCZkL6+rhrYf3WdViai6dD982sUIeRYPc1P1/R9AXKFsbAfUtiRexFyTTiaR7jfN8y0sE2+FJGzZQtP+Y2CKWZ9zuZ160M23Rd6ZzUVTBfS9znk6XWJQ7u2Ww5rlu3lru87a6Miy92ECzqlA5zIGsGPjBIg9sYMpJhsq1y/0sNxeQ05p71dRxZ1Hwjk3xhCZIyGbzj/8FO32l6ktAWseYZl5leY/yvGOB9ccyOlBwQtXp6hZbBJg4/yBIGspxgmXi/OqgnScfvJu73AmdqzF0RhnlLKPsnlNV81ROJDNZ3QVvIdV/kkUov8hFpTJShAs7OFkv+C3ePlkqbU8IU/nuA9i6E0hRd6AHJwYL9A6LVhR8N0xwCSNv5JSzT5JT2mbZJB5OP0xUaNsKOqjX7Jyhraf16pGoaLZwHABi6I/xEUy6J8xhxXr0XCtVo+4rCtvkR5oymb5Pts5vUxXDIY+jFnlYH8HKLHLpTE10IojiwGZXKzChj2++QmpNhvXQa2geJvw6fYhzwjmI0kfV7ztYoE2SUt10vmmjZjV2lQmhFY1KgFGnA/dabzlGicdpQf1KVoRxcfsZnRpI0L8Uy+0nLAjWUY4Bz33MXwU4yyKg/32zaRy0TBoK3H/5Kf3Lra80Mbu6iW/H1xqntCDKwkrDQfxixJKd32Cbizcm2ROkL9iJXeAgN4UMpskfo68sQqIXgXUebgELyB7j7cYdqLLIEDG9EmS4CZwIOQI2YVLI34Mb4U6FPDjd28e1qwIDI1zg56YhPLbinuOl8nFnihsAtuZs7LJQCez/9OjBGAw64LrChGOZPT/B/AGQISJAdtW4qZH8GvseDRoN8Km4OXb5+orPe3JHsmzOzwQ0k13NK7mWdncRuNsupzTn+r4aqF3jA8aOLkcoun6k9lZTIGSM36/Zoc2w99kYaS3cW3umJAtmJ94vkq4tZNOyCI7BMeSeq3/725LjWfJilQ7Q6C2rh+gfbJ4sVc6qUHeSwha/qfl35lV5xJofk29OQPh/ebjVSBBzjL9pEpqYRlPh1emtpX9IOfAH4QbOPzCgHL8LRfbmZrEAkit7c+9/YE/oe6ClorQy0l95AfcFXMALgwO0OZpPqBHUsR9BWga0DHLX3NBQlOVHX2Ya91n2WK8mFsTgiO0iQoJXBDmx3EOu+9EjYgCpOhXMwJBjHGhvuUXweXEBK+d7nq2U2EJ/xmAcIOq/Qw06vrNkuAhZ1LZUJgrAjIaSvsPMoX0vVojDTQBWbhQ+DMJJlveaVHg4sJ1kkRv1VZXMWrXQ4BgUWrZnfHeZ1CXfWkhWHsV1GisBMd/H7Ixux9Z0xjAF68D509CA5qbXJKaWvchiHzU1SgMlftOgVQDLPm1dQ3PQJpsLQKHa3W/45fgnKP3JJAP1fRy4JtVS7Th7gzji2jsJlMrvnZvxLPpa0/oXvCwwDY9zOizdfCyebwlQ6Ms7oG0481nbVNhmSavV2a6GdccC8og7nvTQ5jDLATitveFzMd9xr6pBy13n1/r9JiG62zaPP8ubLasGkSD1Kfb222eUSx9ggAT6mN17qtgQWAvS3Y9mVvlg4VyW6CCOHDwdolPtmFDzdZ0m82o/2LX2LXO8ucjGmEvGM7z5JDGqsDF8Q5k7kGC+2zrBvVHPZLVdr0EME+5MTijzSMJVZfncWUnFb2uABqOd/bTtGjH7aFSI7ZPYTD6pPr/mY6zRJxe1xPmnA/+oJ2hyg/XpL8xN0zhw3/XHF7Qihk+PW+yLScMIiV+7YGGnGUOTU6X23jArEMq/lV1Epl+T1tfpdziGWh01BDUhpLxcAA3BHRfa4bSecmDfhAkxHXCm5PVGOTrEEEYpe73nDF5p5LBOZPfJ+VMkNvrX6kKhoA+3ZoxrTiRHc/ocYWmp/LYdz4x/uTbxqBvt0ehI5nJK7H65W9KeQIib7mc9ZRpcdBg34drhi0c3umSxanLhvl2Z3RVrWgB7hL6qR4pfPsbE7dUfDH9zYkWbSWBQNqOy7QWYgP7XKDln9ERljwWGWUSdpUrIPlfimab03gRxF4NRrv7smFvfBm9JHuF/NEztvkDh2Kg9uBRhgJMjCd/2BNcMlXJs0MqDbTlIA3MEI5XjHyzpjWMsv0tvJ5o8XWP7DpK8uXTLoqQtQlrQleiBiE05uurcDD2l9VtU+dbRO0vOfY88xpNlRwX80cz1RdeXiD1bwaGTuUBzzHogH0lHZeOIwWoVfYxXo0QTDT+lIfUOmr06vOq7jY9FylnqkxsB/ee9dR8kahwMmz/pFIQ8jzBynMZO7RrP51zApQRWcysl85Ues7ng4hbwcU05elAfPy/hAHc9SqdNJQ9F5FV53LRYkU8VIns5vxx04oqjoyW7DkRssJ3JBSplAEqSgKvbdPPi5mjVfcimXhIaD9mR8OI1Skp+ElH8WDlN2sKiPhJQcHVf6LdR7sXyNLHqraRi7W9Zt11HkKoHdEV491Lv/QVKKDBmiBT+ppQnhviO3Qrl6z0ytwpdbm3RDBjm3Zqy2nNGmYUV9N1RvFf7jlfV4vnuzu/18a1EwdspclqXdXBy0Psl6e/B6bsBWw3iJzgMQqYIWJY5BtjEuDm3Y/o339tmMPpyZuT3H09karzq/CoFMHMh9PERrngJDdgpbznNrjS5FxDaWjQL3OLMqkUO2s346/K/a/POB92EAV160riUMbqNQCAHJDVrBRIV5nBgjCxA5bJt6Uw85FNJdlFSmlY6H02jmKlY+cRQssWbiT4XbycPEMYurkvq8a79hcOKVvJKBvQYdoZvdlK7BMSSe6gTOU9TOBudyDiAp7keByyZzrF8PaU3GpL5yOakHXhMtl/r9u9Q1Q9V1R5oKwPrEcRXOOe7ipgZ6moBIeqiM6dUvBjQ7LkcxvjQ6MyHXW363AptqUrlxKSB+CaF55QOl9CZlflVUy/2YsZjM4YnjhhWO6r90xhGILBU/2uSi27l5hRyjRwBj2bhk7Bs0XUl4w48+5mK3XRpKJUjF6W89bPYgGtZIYBHYacIVy/iX+Dg0/x3/2uRRsCqDWM0ElB+a+6Vyu/yVKEq2O0VD0OG9Qe5rw5OhZQDxha8Klgo2Luubq8uLQPaCiAYZTrq3TFHDLpTuwSUoLwwU8npPG7TCbjAGBC40KQiyGZH9cyuENK3ikY6mUfPefm2iSsixBg7En7Xx/GoKG32iIQDTXPpgMmndLyZQL9sWGtobl9yUbqbOO3zgHYXiLC0Fk5jrc1b4x04mMd9f/R3SE6vgh8AI0agZWadr+8BTGsSGTXQR1vDHja/Bd0UcMWL99x3O0Hy7b0tNOmqO6Pumv8NvCfTWsYlJI3Wh+HjTtFIgKR9RTXX4gFlh6GK0JPBYtSqWtRzuvQo0bKbd1TjUP1DsCTi1L+gJiCVByPHwClxikcFi6pyxHn9ZpmCvyIfUl9WQeXGvFyzBoQMPxM9rM5HfyPODMLZtgn7JZXMX7RhO8wriIN3TKXCWMaDSVpz4hdbyG6hgtMOXvJwDM2VHjsK7ERm45d2Ho2IP0PDQ5E0c8MsfcFwYmku9lv9FaqP2kWxH7WdEqq7eKk79FL7/q16CW0tFWaf+LasNzKbQkvF5BJplSvpFEIvdEEmOtYfKY6mI87oMW48h9QUkQ8i4SPUuRaZVlq9gUgc+JqAomK+UpW5C+mrMPISsMA5w9mlxC7a8Nd/nR+fWG7PkueOluINdr781f0Pxsa7ktqbCkx1olS82w9HZWr5r/7s8NoRrJFZZ5ejLfwYMTIldRaPj9dPTvFFM+KYwUWfeRB4enAikz1u7NV+r3jlBPiAE614o8FheQTG6SPrg8burraVeQgacTJxkX4X01zNy3Ljp3jfkd9qSumrQ7SqKISpo1IWzArQ8dekTmWEkYUyuGelcJYMyu345JNNYCEP+6Zp0oyprvqFQ2/pbieP7TWlNiOe1aX5e5f+kps7vE8fpqWvoK5PtXqXFVTK9BrOXTIZAHQCHwRJHsRaa++pQSKsdQF2ohvQ9z7CeVay++mrSi76KLz5eYCO/VYuiCuyZVzwOvB1YdiXP7kIJUj60m4NsBxQiSb3hWwqNqipHQrz7QYEc/PG+pKr8unOCxKyaGvhCamuaPMfEwMERu4x1tj8d6Pb/i18ZrFnIfxuTnr5zc7iqkXE+NtmaQKoMRQ4lG8qo8zxlSCKMCXxxDkec4B6p7BUytSVfF9zV30UaXfPzfTJzV6LCB73mKEAfF1EWgGmB0VlrksYGpDq/olB29UZApmnVqg+gdw03y+w/ywR6VQQPXl+5VCLcApF+WMYKCbanYqq3t2D+eJOsobNWCeVUshsq6cWDoaUzB4C+HhwHH26GuixZRbgYnh4vdi7oH0+wQgqt35eZMDe2cRVbfn+r9rZGcVL2/q+Ui9clyat70c2+q1bgQfIPjpBnK6xk+JsU/BsZe2a4cPsNVHHvVP6AiIsdD9AaYYh9tkdo0JLouKicwn2PPq6Gfx/uES9f1OseYgpfUc9T4S43p6ngJya9V4OeT736SPmjACnAuedZBylXZtFDwOU2MsjdTh4b6vb4/uiSFaYjCL3GZ4CowcG/kDLJQZhlCEwofr5P/0BrtgPSNsR1BNG/mu0SBP1lEp3F7nuo2aGralSUPMxd/k6etTV2Cnbn60EgC2L1rWY/6lNOCW8zD30aQQZh3HAT3WCcB+Zih0gCk+OUDiESBrlgd1MSjXHWUqOTD6iXHxXzGysj34j5c5NvNZew5e8givyWtBf7V9jK2wpqo1l/D/1SDRVk2iH6JvW9r/ww9fIGaIGddpejy72EDlGwxlD3CMcVSZZGJuWmOo3R0IbKe4qQW6PsS2YqMSFuFXmzoIQ/ky3gv5EtYDl+QiamTvVk0NcMZtuGkDXX3wlLZgHNVezSfitTGq7dX8XwZAJ1t8gPT6qkHi+uguwhtz1Ci1LrduU93uK8Y2lnvjAATwJdomxFHkwktBPCVnCc6LE37zODHpMKMSwihGDwYs6TBrlE7o4KfDvX/ji7DAMTmEY0X45BrGbZQWH9IQcRULGkht9oakHqzpi5dOcB5WqApeakmFGM+C3sPvxqu/w9QhYdf7dtfl37TzvjJ9PSmutO5+hOOnos4FmZf/opkS9Xakd2IvX9Kx2RiIWpMC+A4BeR//ZgOnROBrHRVudTZVZaUvkjGKvN0tT0BfuLlls8kuYuwhRtfUOTa4v2BnF8WCs+bq3w1h4PjBwuhXNwYI9ZGdUqAAu+W7qkM4ls+6yqIb16lgPKEiOI4zOWb7MQm4usef1nyX3ivDQRLKh9q+f+4sXz1V9Lu/1JAM02rivOamMd3BKxmL7d1izGWCsDAdwQkKguAl6HsYo84E2EQEmH6VqJHNAz8Xm1f+oor9HMD3dbW++OMKz1oLavAzjeYZ32Pd1Q9FwcDRWP3jHtz99lupIv8c/oov4c/TMD0KT4inZbDNm/AdgN4EfNHBRpenGvAWnCUeZpoK9vQ+LT1kcrqGsMco9G2CAyLYGJARJK4yWmsoLCljFUN6QwBNoy0biThQ81Rq/EyHMPkHMBu5N6LOxTVCVhkIfnZyXh7EY8xiet0ewTvciQORtJ25xzsRTkMjXw30+gh8FZ6bjyQLo1fCGNBYy5u8dJup77OqoXA+yoUBvtphb00/mwzSZ0V62xGgg074OYgCoWblg5I3/Q9IH8xJMURD/+lsICwAVTkD2j4OLktLCLowcpHezK1oHVGUqcMTQRnEfqydO3Y11xrYuvifhKyjcE3s6l1OJrkYphIZHW2YjNERERu330ZnUOYWja2nhvQ1CQeCbBHMbmXWg8PYRyYSO8nROSx8j5JYGMp2VRju6hymDXpx+4RUdn7Qx23D+y/3P4/Oyo2fSRcJglpgGVbuUwa4Sue2bmH42wvqs6MdTtWDq+wVL4A1H312f+GGFuzinSEfXrCPVJ74U48QaQZR3Gvo7AKrrQCNzEygA1LDKwWH04Vf15NIer7R2TRP9DOVMyhfb0Dw0tKNlr9gL8an3KP6iBjf73cW6eUES/2IBH13jWHLdPk72hXWwUQP+HBDzq8g545BmXHHav+npZwfWlb3gOvIKARvUDo7GB1smnEvydM6WwKJDbpoqvcEa/Bep6FaQFIhxsl6eg+AJZLSDm81xKIFTn0Ef5WsCTPYDgDpXFZSzmubOwn6Z06XYGFsKx/WAMp1YW9yIkoO+yJK1mIyvrQnVM7SGqfJUuh+vbt8II6aRQE5B1cs9jtOFKsf3OS7F/DeYQWnXoMct1Qj8fLRV9yNGmP+n56OwGyRu4f72CwbWy67snp5FLdus+wlKX34yWxt+vrYq3aNdq1cpoKgN/OYNWkf3qOFmJRMX9ar76mig9/GNVkDXmwvfJNlw6cTWYziCfEvdDRaSYpIZGn9IaDrSXR7COy9BSYdfPRKW8UTuIWZe/yffFG7qOwG6hMdMH0PvM2CBT0kr8a/+Z0qcd8QXePY70lXTzpPLWLmgCz3B/WNn2DPPwRfZ9Vn5wU5mZ6/Mzc0M12r79HCCnATj3mCq6auls29T1adlfEeeUGJCOZfPRjTMztr4WljiUjoWyI2ozFLfvIlbUXZerCD8T3uPuF+dEi9vI2SHMyRkMLevQxpTwvXNKQSV3D5AgWNNpRJdS01XtC4OwPn9Jhh4efWFSKFb4Hh76hiZkfu60Q3ZqxgJPYCxRSqaxong5Xir//JbZclYeRLv7PD2DXDFEmDB9WidORGpXLl086qLdt8gjegIvvVxRCrxinQco2684nrH8qpOPXCW+DXK1Gj9J0OXmmq9zjlE7NJgK6dsXqc0JX34Lc3w6cO+pXVrNnrKusIbs+rBqF7c676S/lmNdCOc1JhcMSdR7FRBRgdi7wdiaVLfuRQDiWPmAZMb2aBoF3oFwD5wW5CUbC1KE4v6mgIjPQDEg5reX8g21hNs6x1WLAvyn8UQv5CW7L7GqnOlq5FgFNklanT/qA+xDYpbOZ2Y5I6aT5JdY36e8tkVdK8J7undem0YXA4o6KFQMk/KpX5aU31XGn02y8YP/0CPNFNeUDo3VSXsYbGwW62TFXBGAS/0FDPQH1zYV4TNII4QyqyJNqug+q67tCgg0noJCdQsN+naVoO/tg5QsZF49Q20eviD7cb75EoOJwdjZsqx0q77sJOtBooqu/DBNShQ4XYUJ80PcG7mKhbjR/GdfW3peeHbPUHnKyzeoWazII5M9FaVYkzuDno5cqjRsS6lVBr3kh4pwS4J4TgVZqy7Cw5hhde7FHngU5nu8iYgXg4kNpAJSssDFq5zAUrZarLx8uldJQXfT+ENPNHiAymWjvTIcRbiM3F0h7U/encerkI7/xF9zOISnY+YxbmWwlnBVbJU/l6EPnvQ4NCg074SJRbWaZ4aRo6BdH5he4IV+7elIqeQHmYdHouP8NdclT5pgE/n4nlHgxjdsa3JyayYIMy4G4vBnEKMddhYeTuFrzOpP/uj3hdwjmgdwD5baW17RTvJzLuaRkogkAvub2KpTtDAeHbo6MF8GiWxnzqecxxjDi+Dh8TfHDjuxtlLZ/ObY8u3a1lM2leVZg8vJbfE+SuRnG+LFSZtjKmkVWPEem++v6ZyrVNBO8XSuvbiR01FF285IwRXZNj5AMxwd+pe9mEvWOt2uuczNr4FfYXWEUyFOgQ54BV766iACcOqGQoTsyomMPD8TA8EGaBPaKYjqsIHT0OTS2UgbWwH7AFTNREkyI5h5ilSDktXtoRvDKVeo94KDSLms+ENJ4RCQy/q0PIFfEfwgzXV5cHwwZU1Vt0ItqoBY1IClDKw1YqB7nUIGCKbIZSCRq6f+Ihkw5y8rEsxd+elqkSzJDDJvdRao0uDeYLRvJtxEOtxTs7iICqsuMo8IVt0BlxzgRuM8hPS9Ghmi/3IYQ/YZixkDit60AJhHAfyDF3UTswVdwvTLAhRghrsdF78owM7NLQ++ZwojMUlHDU7ZeF1NwhYppx2v5S0bhC9gGhevr2xiCuDKwHGa78loJ3yK79sVwHrRozJgupGC0cOsuIlkUVOY39odgjgWcWb/nVr4gvKxcq3/AyPD6evMwMhip1ITf8Aspq2DfCmHv6h2Zs7RSaKgU3WnI6LWhEldugc3sThwfzy9LKuS1wbQNIK6w6a1IpJ6U7N+lTfjCZ2jhkZaVr+fa+VrNm1kucj42eD+hFBhDDvUH2FpvMxHcCQjcGyZ1Gey3NbX25ztntntnvZH6DeUBVDgzsqYxVmWJUioGYMxyZhE0rpVeZtIMBT3qUYkp7w4DivaSdLEkHQl2PZpj06YoFTHBV3MKZQZhWnjlR6WmN6tOQsec08yQ4mfPqqT+0XOns1KTunUEOTdFJfS35RQUj3Sjxlh7TMg6xF9sxQkXEselTrUoKsDrcX2X/B6oPh5+cOL+AIa4Kt/BBTt3msA2bwAKWwxP5IWEUm0b6IPkvPZ10WFdicrwr9ES6QAo0pOxqWvlzIIcHlQ+RPgBPqExADPj/hJArMpLKbA8kt0e4o748xNTEW6WV6pqqlzyR7QpjB1ZJjRIPC69e+Cg2eLO1vHsRC5VMIILEO7lFmhyPQfUmSS1XcoQZKEe2zfxy9Ss9qAaQ2DFoWSb3Acm3knm9nLf3GnZ1Iw7Lh4sTzzCB/SaxvlfnIOr9lzKbmarg3YmfyYvZV/d+Ob2avn0KRd6+xldaEVlC8Na8wx1ABISH0IT9UYhupBNR7QVAWdhL3gMlld9C5oBG8T26Xx6NqU3ojNDFgXpQLxF5VacIpc7ud9TjZDrZz6YRTjKEfNf84Zkbblac3fVKcJsF0tMGuEVPyjf6k5FRnrzqvWxqpusKn3vBcTALb7YBehS4zPFoJn1il3B5YTECaHO/xCU6Ugr50CCdWWUl9D9vKARlGio4VImzEE1BFKxZKRtXWZdxGYWK7pbJG0KgrihD5mjak+lZuzq/B9fSs1YAifOo5ctg2RtVWd6/vjXEK20B4tf2WlVdSvzmQI+hpQESIkXlekIbvfhYhhKuXKhJrOFlfbGXH66rSZKn7P8WgvB1g4H0PLtyW7NjwmO7E7DAf5sJcLmVmLKKNMO9B1DsjHjpjAtoDDRs7H7+VwLZQsV/tBjBZO5G79e68UCa9qIVUqZUvP6nh1DDOGdbpXZR0qET6f9xaFlRYh2KlUMBoz5myjGwpKY0lqao/X0c2QAQngQDX39QLWlKozs9CRGtSJDNW1y2gHUEbUa2rsll+v+bnuyh65V4g2QN27t1AckGS4bSa0z/W79uJALDrHlc2HczzWVWe95qHFv8I234OSF5fh/q+fwwr2h0YYgy47wsWm6p+ZIzj5yjA5s9PxQ0TD4zQ31E0pZMtQ8GVvCHB0/6qT9khPnoh+glRtx6w7cUxsybyYXqHUps88f3hEB/StxAE0gBRYwPy73mpTAIOdCTYr1aVHEetworqNlnzWzGemaUkaJIxd9nW2+ytAnlxb/aPUFoCd5Tgq8BJ7ndkkrnevNinPwHDtJwgQmKl6ei+GYxSEwEQ0pUl8wUZgcY8jaBexPvE94wEcX+rDY2usDOUpY15bM8SytVlvk8RhgXUpYLRbP75ELTm4vCsed3Z3qag+C1jnd//k+K1zrX7sytbvmoh50SGMiv4jjyUnuHht1Bq9pQHVImm9m6sfZO+IaEnNMJlTRphyQzLQ0jivhJ+PHr/oGOBGEO5G+HeI9h9vA2WopN2+DpsthPymqyuVCe5gTX7gnqGM2Aw5C57vXgSaE+iugdu/n1fqAB+/KCNHeEMH47oXvRMLxC1jWffqlWxOakbggrxT2t8AhuZVjcqLdq8ocfS7ztTq1KV20RlMbIx/892A5fkpaKj9Cww2eXj/3osozdPeG/mEVRBUYNVoupcCxu+ZH0at2Js+b6r/cNqMf2IBus28zYwGtsyS+GCNIkuyMuiALSM3IX7GlbuiPc5iBda8YKeLNHT0OnTm8iCsBvwZj2IwQZ4kh54dpi4nMGKu2zjwHzbrguI0Xv7VEpQdcJeHR+53sq2vNIMtQ7ml9rHm3cqX9dArd15PWpz/gh91z2PVxmbOfwyCjZ65ECC9P53T0e512bTXyjULgYyfC73if1ZfSLu173bsG4BFTcmI0GHVJds47VWw4pYV2Ej1XEkMI3E0siUsvOGi9XSXYhXhwv/JrV/YrS4zMXAtJKZkbE6YlPyu55S/HTZLCu9mGMqjbMXMeEvEbKLtrzfLjtVj4fNR9V7KCsuQIVtwqZdZXEIfPrFg9ViP5WpkfjB6VGCkR0Gut7+f0M5wwBBHR1SGYPSQisCXOwu49JKj4GQ2XDDI/oxAdOCFvskBuuA/lJwARsn/ZRveB87Lh5cqC9um9kkLPaGIpq/vOfOpBMDaiHqm8VxeGKqRbt0jfJmvdjANcL0MuDbpFjQP8bOw9udb4gPbjAC4buILnAT01ufUcuaKhQPZgQvxaa/e8UYRuxZ2ZkHrw4Ki0nzEYM8Skt5iLdUY3Ppobmyo/s25i0U+Augren67pqdHE7oGexsdF5BnELI6s0AyR0xls+HCR1JtoOm17RNhxN1ErSOzvRkIy5qnEuMZS86GvI7hBx6VT1QuQrLNJouQRsInBlpP5TtLyIWWONCgBQA8SHaq5O8jn2HYGuM9LuoQKSlnmuBZqR/K9eli7HDRD2uBX07s2tP3CY/qbYkinQ8YRjc+TVNFXklwVn8piCkSHkhnQ3zXkLMqwUMAdT3G9iwfBA40HbEbzed8U7hML9IoFa3T7Ea6/x5uKg24C2HGsnI+v8mCcy1A7XuTkbT4auMeCzgUgycWHaCn/UvzEiJpCij6ljHA0tnm+E8mZB2Ap+HvCiBaMJoBxJI+9lArR5Nkns/v9h2yM0SZ5y5Ih+USXXel2rr3o2Gl26/xZiG3R8e0Oc9KGBOuq/LTtdgdpsObMLpOE3tB0gVEBIu8Whj8ICKTfwe+MLxkDIEO+Suy8UTr9Divn3um+mAiH0pFtPYrsnUjOZP194X6fvxsnzLYWF/H9ZkasoOY4ThGd/SR3cNT18g1uOMSeNVrt8KHo9sDZAxpzhp7zcwidtXpj62WkyGLQMwP6/C1voGjOE2yL1w+2BByR7VDo4/oFEI6NgymMgoB3m1ogFWzzWWTpSFh60cAprj6t0fv6aQ2a9z0ZTWMyUy4oDT+zyl4WB+k9zsWibbYl0IWNrYDDMcrVcpGfEgCX+cZuzL47e4C3/9m+Xdeh7zEP1eoXdnKIaDwWAA/b1Lznt2EnKviPJrLGfr4exTPJ+hoFCIKR//TEnJWLSode5Jx04z5Na1Mw/WwArSSBFMEg7i2+Y+d/4b2KttnwQdYt/FvXuFqIfN6nE9IeGM8blhZkAKPjMt+j8NMVrYY93Hx4lVfA80qvi3qx15ck4n0XH5LTOu5a+3czbL8yxlhB8weRWqL/KIccS0dND/ejsNaW5fLRUSbtg20tdcXcP9wdwCinmKneVXnXHEwqwpuNwKA+N5/EY/rFVYbnk9b+TaIZloKe4d2CdlmXk6zCiRuQwJEFn/Je15QMvkg4ZUZaU4IN1B2obFZ1AYhM+y7eoZmx0EnMWvcp47e5cE4dr1jDoxr+7QwyzoZ2KTvwWIt5SsUPe5gObt+3kkkVH3KbP3rAHs4Yz4U/GqZfCNA+JiXcH4IyxVuVScrOdR+ClTMnPjG+XUUiQCtHD+u//FhSg/tTd/CT0ky6Z/0cMygUib7k56njumMrdev+2sVZIVbT1SAxyZhFZo9VkkQgOd6mcMkR89Ej3OjpMKYGMOX7hY/62FkMkOd94Fiv8u3Gv0PMgHRUhQ6jDyLv4Qrwv1OyCaQP+t+RvddXEOdlR3pHcw85ErSYeKlhUf9vh3BphjbYnQyqdDRgKb6tAg6Zty6VggkQ2FzsBnAdutFwsRn1M3cyI4m8H4o2Kex/s8iy2kvfWM5YKsSIrRI5HPOCb/sVZ/PFXbBEWM5vidQ3gU8xQsu0pE6y+HOAqHf7eBlb6903aPpYFotgclXFxFo5JoKhEc/eLhSAbyEuv91b3GPL2bngfI2MCp7M3rbFUAoyik+q5FnPC5UZn4IkIRBiVDC4yQbVTWprAbGGF6biMCW195zF3NrS+JQROWkz/UmKWzOo1wiEs5G6Koh316BkZRpBN9TC9xys5SujG1kp7ifOZ5EM9iLczzkYloCp6eDNLFx7efwrImDdD23Dq/PHf9cNzMD/so4m+OAf/fwbq8I/Fbw1zdjg9spRcWfW1tqOaEo5/zevyb6sUWgnVkd0s6Gj5iGV1Ln7XwSKls578WKhub7OkBb5iUJrLSJQUuJL3Uothl1yjDibVuouQl6XuBE7pDzpfo6dQu67z9QXr903E8PCioBW2UHK/9GDz5jg1AcBdeBe7N0g1zBcCggs0G2Pn3L9PGyDkDlcpqvnliBaKG8def5YRIbtLQTuT8b7jOrpX/xE3dEJN07eNf7CQtJZ/tFje4elOPKK4ye7e0d6uwh/VFdtNK1NMzh8qI+zDLHc6ERVWyQ4ytIoP3Rfnml2eEYHSNYbe27n1PzN3/icx0fMifUSECjW9V3GtLkKano3LBQDhE/BQ13QjT6YUfzF58GBGqOeZDOnCDx1TkSPg90E+IWK5DE4jpD+GgIMrlqqnQYDAvAauT6t9Azy9QfDJSjvqmGZ25bufDYC6FF4Uq9Xq8YAKwuUwKUP5D2j0j9HhBaysCHkpuvFPGCX7oGXAGHokJ691dWHnC5a5/otnHoo6a7aYg7ggz3TefN7wgm9taLIlxTjJdyygZ9/126cBnRT0YjUlVimVztF3KQLs399LT/s4+zUyd2H8/LCDirg8s2ofhh2IAwInpLkMYW3bgQyGxELme2FNuGM9wA5G2b3seWC6wUsC4sza8PuQW1I3Rr81/I7Ho9r8t2S0cc0yUZkUFlojAjw/K3uyGnXXyo3Y07ASNt67obHe5hZqkge/cTjwktu+4pAdUW3ZvyxPsJc8BLCnLnDX5vyuWoMnKR1ayiD8/KYTLoCE6Ej1WCqxa7yh9wstq87m+qwLTqAk9byfPaCGZQ9llwjKT1OfnKvTuwcs8qbX/tmoM5UcLKPmLlAIYTp8hK6Oodze0oN4Te77/Hamu4QEiiRpeGjrD5YiIJGy7uvVxkDMa3hawuSF1Rz7V8dPwhtYYjSB43IWmQ4J/l/HTNHSCPOLaKZRe3rs2+itabkbFlDK6FtDzZ6fs7IFC5tOZryA5MjPL078a2CkyDceKntO4mCOiFh8kZkSN03wCcuDoItYkY37LlMa5ozN+/shnp492Jp28slIh20k7rw3DmrVhPVOeK8qm/gTYyKh7Jm713fGhvFXXobQBBtd+NUn5DzDRYx3x+N1FchUzWqsB6ojvfqcqSAZdRuvXnTpGCDFvmpg9d0hiNZsFYhIic9I8vqlfUmgJMCwiTlufZWFjts2yH5tNWxxloeELU4sqx96nT3wO8+UMn52apvBvJUcfCReKQ13jP31rW9kfOQQxC3Nii//NkgHf65kGhWB2kgmzT0ENg9XMY4B0eWjPxbdRqVTCwj4/7R9R4wFATjMPbLdvqgLORoVbsFk0riErI/kk2ACtel6IQH/z1yMUsEZ3LuCbtJCHv+Z5PQJmNuU36rHWlHQGpeNdKXkSsbumyJBLHvFZLbG9H1WWxZdbfo+cyIFUzC8UaY5GyMLGNIAHcB0BVi+JajGQLcHQqt0bg9BktR301fiDyX5DP5kTh/3AHSRm0O25WGKtwgCN2vmF7n8NGV1Towrt2lqWjK3icsoMucGY7qQvskL0lOgtIVEROo6xyAGy9/3psPPUCcruvOyIkBvMjB1aKUXepEWv0XGWev7LYeVzOabMIc+pJ8aoaTYzIhWHW7YTDlXJfibikL+0AOVtUojYDX2zCLHAzibHuJrnQfrbQ6CUaHNLrK7h+qhwtWoGVxfz+lR10cEtCfKoo0K5PqcFtKkfwogUo2R8lp3PI+HM8qGrlRL1gYx5uqqKghxjLUhwSmUoxGVtNOnAsohza6rYxH0WoOCPbZfK6ZegpBeFMlKhs4Fw7ZX5GYiOkOgeBMBihXmq5STkLYDxsvxr5zkPpPxPFgVahyeWVzyiZ8Npe7vzgk5nBnB6xm6UWhTyFDNNEsEznQrUQPvd55RDvZNnqH4eHpzImvM9eh/a7Y8RhGAVTxfSbJw5Hw4lhOmmWwxXmT3zxq2U0tvQcvpa2T9i7JBrLb9F8gp/u8nizPaWkxZhae1krvi0phXAIebtpR6CmQ39a+hed3uiF9sbaeLzFSALgTmPTpqajlb1ELg8KZTPr0WseBsbPPXfJ18as3eHBGKADBA9N6tBWkcwK2YvPklV9aCnUxd4QGNJIsqHUGjHYZ/fmsCS9vSqTw3fRAmeGVDfUtJOhZIa8BWjNBzZEOjrcVEb7j9123AsoSc6Fhr7pCF9HbtWMxEsON/I7E3gbFoa0EBf7chO1DBSdsp6ch+BzmTa6ZNfR8bGNrCHs6ozMUXN3wntIaSFN02O1nPZVg1tTofR/hRLtXeOG2Cn2tUDtGn9CDYgTcxsgQnjsJJKO7tWxoOepbeDE8m2TkjdByy6akEB7NUsXLgOam33UzP4hKIK8nc+l9sdOubpl0HSJ9xVdjip33UDzGfAvQKHHHLP9vyPyn4KGomCaZrF8opRX/kFyzBut+fQa7ZtP3u7TqYkodCsuke+dDsBVoqS4cYT6sZJkAv1cxT/vH0SBAHD67p4zoLt/aBIgwModsc7xfKm+zFu0sGTjjurfWtHRxFFvrAGqy0vi0IHPnPagBMJHCIPQj1Vfjs8SBjj2LTHT9Xee96KGLir7ja7q0WOlM1wqxkl5q5c2Haq0VYzxdBabhYcGR4Zb4/8tJiiGz4NziwcWOaZK/4rGkafQlS+p7RBgvmt+IuWK65wi49G6LmldbBjBAaV4EUjQvrL+FKQDq1HahKRI47JuNVDjIfILVv/Kpz8KzFkC73G59ptlXkWreioJi9yu1SbIYX2FNW9U42OvRsgnYkNZ5+NxWtfg6SriaJOxXtf/Uab25H2O5luTPVxLgNDI3/XTEWlLe04XtSI+dezhrMeHs0Ho7ZdytTShHntbLq8cJPNkQoJyFszhlZmHOWs5AwQmWE0JHFayMAAMcOCS3rIlgXtcOy8kLo8Tv5bYj5KTRc4ehXQfmLlr3LO4aJnXgQn+WmW1XGeo9jdiwrkcBYsflqN5j7GfcZBEnswyTG0+p/ATgi/Wysjmo9tHtngSRQBlAN4+GlvLJFBAysgpjFSrJgtI5vuBl3YZrCcyBV/YiMCN8fkMQGq6H4/4hd0jA/kPWkN/e8eOrirHTefFryrGLvMMaXGQGkbas+fdwOg5+snigwNVumh/Obva85XjE5p4tIP58WX4fvotqICfZWjtfSIFlQAOZr6NSB/qVYSBvj8/6hkUNTSnnJifSl20BuBSb/3afkJZCyr8/padBqcs/lQ/SkFzc40IbvsWU+Mtu+QlE9lQOtutInj7/Zr1gkHgaoCZ9CcVYyZQwOxA3HfAp0EQTIZB6w9hNam4gCtzEvCFXHh7kUQE2qS8uu2/hLhQu3ug0QnxwMHMrYRJdrLCKb7oUqLaG7GhRpfL1HZTGFeBevAGaAX4E6HgR0kqXx23YHS3mWxZ6hTa9lzEnszTHukuO7jeeRq5c2mL1dJ93p8DmawfeLVp6B3/jo39GMHZAkKmXom0tmtlSMlrMQEZFUXwVjZ8gs9Ypgkhxtln1cbf+3VlT300QhAuLAJo2ipxYNHpVXj7Xj+Z9KCkp8elsdDwvSE+3lx3tOj5PdLsVN2HGVHNCB2pO+C2wIsIfs6ex+YvF8KDMRL+F7oRsVq0JjYIpWS0CgXIIJL7HWCnSISG5/Z7820fk8Us3xAlGrOCMA9yTJuSJyChrCrzX2Uj4wdodJUOetwcDegVtKM8OdzAJpO2IRSfkaUuIXJakAfd+V+ONRJZHyKcdK7NBse9aq6V2tW8Aovqp42aKuwE69g7vhi3N3p0xqcGctkQVGlZqne269asUJ8pvlOJB4dc+rDXqaqrSbk6QM5gPMqLOuL/6zJiuY0VqAB9UY6oko1WExb9+JHzP+jy3HC3pEce0L4nwTN4lAuhJ6rU1hwsUkA9tSC1UvkmXHiZ29v8sLJEeZUGDZeTCQGJY33rKhth3qhTv4mXrB7Bf9PIHMbuMdr88j4GjgFFLh7Dgk0fdCGyVaesewuAb6toU+A8f1Ho/sIIAn4YjwpQ0flYFgwBun/cj39catgMhHb233l552JzY50WzlPaZgzyRDXLB7QY006H3R6O7I9iP5q2WhCtOzsVvklxJlEupYnAjD7A2n27d4VPlmslyvyKr2uLTx1XsrdHjsVi9ohHADSIOBDTzBk9rw/I+U2d3tAXRislIocvQ1sk+/iJ5PNb/6GbVwCur/AUiXk/j5mgUBaamW2XOod4NWZ9ufxAxxFUMvwSkqFWG+9GaZY361Bhm7hkmKI40g8qG5RM4IIhvbbFpxGLrNr6xHEopHoXIzMU8PO89WXwyFDkyizTyI7BmNGJ5Vg6GhoZ6c+PzRJhfOWNrO8Dbr0L0CVZyxp06+5GVUHadN4MnuY+i9Xe/xjPQBnSJzuG1oYkQKUapi8bwbz69V5qu2jNWveZU5aKZNm4Ph8beYSx0L2FVG9++LMSgg3TjrgrqOy6NBWe/wBQaDkpDbJsGDcApdX+7mgnIwS9D3q4cEsRiBtq89eWoWgmETM1BNWD7UG7DJLLdpJhbfjGkU7tG4iGNk0zZXrp6Hylg8ySbf7bsHh4fVgKgakGpsHyQEsDZrrTEsMtlwsxr4CigBOkQZizE6u5+1jpP3VxSrd0/WXH22DuteyS+ge6x2Ver/2AW86QI0K0i7Zx+vUZAYfDhJcvIWuf6oasqMC8HzEXryo5nZGgvErk+R0Oy5SNd3dFx/Z2b4xxIf439iF0s9hs2yOzrQ+f9jimX/hQ4es3V+ZELiDdOWkWWYmdqD1actCII9A5xLkddi+zHNmNDPzLWa/Lmgi46MWsiHUpt8k1W5ZwiCSDupCsHBt/JGAiApuNTsHC0PEZ8Ktth80Xv8QojxKwbTv2X6zxp34R20b0GD2/LRW+SQorwiOjArHMtGFYQkhfK5n415FTGOp2JmrZDVR3wxAEyvQQsVn5BZ7o1kSHJcPTfmkqrcAbnMi7fkoJwf5rOYYGlaUZk3zeVOParSFhsW3e0STB/HThpExOzKRsOW3L8Arn+IgMH/4ouHKy74V+8AHLityJct7VAoDSXINhEV33E3c1ZdJfdC/LNA0PfqtS2c3j71WWb+Qz6Xjk+ipDVXj0MMTWelzopAEs87u2t4SxSdlsvHlxk/0Q1xdAlKbiGSmg2/EC202df4OMXb5KjGxszxf0ZoZu4f08flO9YnK3y4SPmstCHtHLg3A2y59vU+FQ74wa9V6hO5NfNXmlyU4iKg13j2Z74E8UmGgxkEUQMyizwu1LAqpJmlDR2cJxkGi/dRIa+aRwTF9C9zxeBmNG1mCmeQ58fnjVwG3iUfpe+K97VGeJFYmgMZyXdU+n7G8DU/7GhtySDQ77DPl7owv7H6XALiKvNjhM2PF7X7ypxVZ2pSTJq8urL7ZzwT79ciun9IYDEfCnyyXq+gDTIoM96KY4KA4D9vXoMkoaomO722VAiXpF4bgV3DyT3bpcJ65mFprNYmp7HNALAr03HrM7RzN9ZPumKIOtIRHy0uuZCUX2Y077k9ddNUxEr8B35PTmY+UN7HM0Zxy/EXQeSyKRlx9x5mwoBCUlE0OrWDfPG6xUVPwHEe4V7xmn3Lto+7QP3UhKxdmsiz//l8ogbTSQctJdjOeoVKkPEGCS5UDB8hQkOROBdwunlldeut/GhNaHkO9RH2mzvgzOXT6u0yMoiNUm98r3W+QrXmifXWjYwgVjUPPB2cKri5LffNVghGfWZLx6+GgRoP9QrnDAl+YWL557L0dVO/QijohlhSAbJqHiJcMO34CLaUWOxU1+XazOJyC6CFUz1srGE/LQVWmtqvbEd8gUpAhcx4ubtUHv1EOVyd7PnDUfu34/PIG7dc1XST/rbsgTeq6dMcD0QiyzdZmAmKot11t07FXWb7NSqMSMGGvuflZ9bKgGO3Cqwdwn2nVKV/I4z/Q0ASdYt5r5Lwe5lM6cxGRGQr5QnofDd33iKKBvcH1XbBzSnRgmcy74dxIatIYEJNlVVf5Hq2Ul4NnMCAgp+eLKnX2mgbh39FjE8yOglGxBe1hU+yr0ttwn2N7kJ2+rMouJQkcTNr7AQhg4+Q06vagaKndfY8vC1WAmpGvrpdF6qY714bVkSjd/j96rnN5T0r4wIAIrqvtIG8Z+goKFY+E9le/xjRIhSQW5bJVbCwRsxYRDetg3ha8DmJ2oNRTqhQ5cvjcHKs1pN7qIiTbw2q+5vZAa/TqXDrYJ1FvPxcuMgAPdBwIT8FJ7Scjo+t1dZU/x8zQUeS4jjle5izf/1sSbYhyyWmCWgRsfevCcX1CQEGDZoH76Z2dc9LEqJmVJ+qgs9friQkuzdym8sgzgoh5J4/N6zz5gxBAAd9bnzMdcgA05HJhowP0ockb5CrwsfZdG36IajqoDXWVrLDV9pFF2Vp+t/MH+fWyPyGczvtzzKWHfJt/Z9FAh4b+ucGtW1yUYWmMGUG4EPRG5wqsslKWksns0LH6FejI0wC673Qjk2/PNI+rChNno2CcRrnBTswsPsq3yH2mnPRLaGFs1lfycfNf3saaVpumDgz/f1+X3o2mlpD8bbAnhzUG7Fb+j0mqA49hRVXLMB7hYdLP9zAXi0b/g+U/pQcE2t9K0z9N8ntzaw1UsL9oFreBfGfRocw+JT5NVIrkzVG9dUI27TjsyP62fSKTrU3Xrw0NxFjv4ZTRBoIAr2fxZrzopEbuGucLCLIy3DbcfxRW5Pb0FX7+62xTe5XqB3oN2dz6qLO53ogp0DKcpxs06hX3C+nU1b0sq5Ecpl13GfOmViI4bVJDXP36AaEKIR5i5KCf9970+jezhfGuJPpNIvzOMTGgOznpvurGN/+3X0gTzDY4cjcr8247HqqMka4S6fAwPwY5g7jd22RpC37uGzgxPw7Fx7W2zy4tm9lgWponzJj9hxKeVQH5U1iklrOsbmmG9nXFwOiVxjpctRKkBYd/pBk7sg/QdliXHnqirzVlRzGQQC1Qj3EWVfrrHcSaBaaZro2+yGqO7uxzHLoIragyzBW+W9ULYSjqFCeLbvL1FypZADaisCH5u3bOEmIA96B/0ZDWbzgkf7UAmq4q7ArbR7BxJtQmYLh5f1dEGQngNN5pVD7Q4RS0y1vec+ci8Pe52fTK4YP1coyHo2KmjkMvKSaSTfUch3Pt9PQLwrlCyCM9lsLp2ho9xjyE9aJMdKnxSqFjO4KfpXSHjFBvYdWOopBgXX1iuKcVpkG++9Qog25SqJKfwRgejDDoSGo4LnyNc6+ZnJoUXVwFEtA14pbE7XNvVDFCB9e0bVEssoEe5cma5WkjIIzi2191m1YGVeO1IhIXHJUgyRSg6F5D6mNX99F8xPCynHMfdjHnOwRKX2m3EQ6xb3B5oQ8CG3PtgDXvUf07HLy4XrvcGhh1P/AofN38G1TqD+Khl08lgLgxIkFt2x8o5rLOx2VZ66lby0U1zWMsvSEwL38hwWkyYxYmmx+iR3qc1yZYRRnCwgF/T7gHB/axfJyM1oLR0b3QGAw2VEbUog1jLz6cWGTPfbSLBV6L/5TRjFamNYJJ+UJP/yr7lE++YDznv8p8V0/O3Rs6OKIkpVWloyIu5z+UGHdC3zDq6HgyyNIkdasmd8uhy6I9GuC+/5/qp9Wvzo7F8lJ3rdsuJ5hrjVBCWIB8RccOkB8IXDBdxDGZBICZPJ0HsoMI032DVlK0rvkoYhDJqmeGJqrpsZqpFnXz0uHzp1v19zsdz/tFI13rQtKEfiGFmDd8hoaFtywgZXkRSYg+J4RTDVs49wBWim0mFDb+uItoBcGiwnAlN125qLtAKT/eccSGV5dqpPalhnSzgMTjmFVJMQgm5kMnHXS83ZIH3TW+8eoNMnPNyeie3HVDucOJ8Ea4CTGRc5bePWHX/Me0v8xV46U9hpwTUCL/GGZs8PNf1rPKTc2y2F3PizJD1iSo38FY8x6oPVsqjqSIVbzNu8tr9VJS4EA1e5TkMWAY6kEkiDia5lELp1rm6o6xETZ6rNUl1VScIOS7HlLr9atDvd01YNYKndUarITrl4A9wDtQSvHg2K+Bs2mRolBtablgHwgUGxsImYpVAvcP4yLjhcpeABaif92+5OU3caY7vzKqcCxwjSgPHNZIxMGS6pAdo1spDlJEn/VULVRdihoMXAsbKokvlVI+/txFtDObh+F9hujeX0OxEn2QNBLXlxeUXSyvBr1kdD1fPV/OB/Mu56alNtORT/w/Y8cX7qL1R+wdQf+PixlMxNKdH3dObjHs4LM9ySeJNyYNx0EuR8QBJIR8LNfq8m0leoih5WE7Er3cWKRLQvqUC9I8s+3YlZnZGEyY8GWy2RtR4CqJTXdM+AlrO5eTkI1ozc5HW46nSo6jsazFNYYommh5XcqrYLqPHQz4XlL9INWhcDiBWQQKgWYxa+6Ih7BB4NzLWzAENtADpbspYEvhroKBgk7dAEcqs2Ynbtdnew0PGvRi6Fki05IiECycxWuwEtObMr0u56JKCtZC8DyUJM1snUQDYIbmw2uFyAGPKiDJ4Cjzh1yCS4TDZsfdSRTvk+0ZZJfnU5jP5/omCpshtoZCmmeuejC7bCihn0YEgiUSvICghtF2d5QuM1XuhF7a1MBmjocoTUrmeqTGkoYEdszIaDjf5nzq513Yv13xN3P111afQotsZf5b3x5s8odj2QmAsA8sgIc6TPgIlUEULw0XL8sxilVj+KUPQDdLi6hoFLuiW9uHNN8DY0hmbz6fUSYdQNG//4K/hMtz6WlvOVQsrGIFk8tXh1UqQLyO80blgpr1/EtNNtGlJl8gvdSUA+Hhar466yDWajED0ISD6/DzmNtHpuzdV8wKcPam9vIGErJILG3yWrwEuMHvG9Fkh/HUqr+bPmoeD6UOB8ECoNtNE8cowZyKbT/4u37LGBF//JTaghuZphIRwdJ79HcPvhgvpwzlcKpQ1d7JIQqtrZbaNil71XBEO/e2qcDrVbM5YvY3pjR5Nc0hTzQVNWRPo1rcIFED8fbt2JE6eqRkJFCMHUWsOrdjqoiHa3IOzjwsKCCu9yhLosM1Jeo2NIriKCRpR61Y1qehn58aZqscpDiNWMBivqduKWM5AXeLjyaFf2GWbgIQybuIgIuznbvlFGk0eEPFQeEQI1GS9bvPh5B03RTTnkFFKQ/HJ/SKP4rG72sgUeumtIOVQ7BONOLTRVcgsvxFYC0dQeEbxiSD6vhbgJfUCzYQ1DXmJY+faIVpKCtHpv+n/vJ4+UrfYgLMV0NlnEjUuXGq1q6mj0jK2q+5FoMqv27C1AVkhH6xJFEXvWR48KniLuPm6mz0qD5YCHWXvhikitTSo8uxcQS1hlqvIb31JtYfm0Iq9Mdh/+Fbl9s+cie1Q29PVWam0kvceAqzT39FW5u/b4QCT6BbtEGYG47qPkDsKlDjQArtTPo+3u+Uy9VY6LeLAtAYb8GFlbmxvxg+45FcOZIQSzkzY2t1CcY91c89RM3Pzl+mrtjAItkjlpstWJ9xS9nWC+D1K8NTze2NXj1QJaY/XSJY4zbhu36ecuJJIlmkhpv/S3vjzShdQiiN0k45hxzPE2BRHyvcwIZ03B9w22zMASVR0OvCbdwD/XCUvGkfWYoXfg8IgXMaHEIkZxOQQPCi6OFrz0QicZrZGuHWDaiKKdIZ8U62nYhkj0Nw1Y4m3yizlGBqa27OAXU3bzr0S5P2ipPRN7YFcpJMP2xOC5/hbmPEZxqihJDVI8C8lTd4+IcVZmcZl4CdBB7OX86ZpHq6NbU6KaPVaU9qGZYu1IYRM6Cnq922p1PjTY36hs61HE+HfijgCF2GThZ5TGpWRkvrA2vPmx8kak1Hn0HMieHFOBodDLj5z1EB6IEEwEipDCxCiW8J6BCAyt9VyGQzdnJJA4dVdhwxbC6OB4ZRB729sG/xPdZf1sRqAXRmtTrcpmTITBPWLsXlXZCZCvePckj2llwuTOmqzxyqYgKqyCPs9yGFqI2VTTbBJtguPAxHBwWEPUAkSoNauYNa1Yw/xvKS0evYiW2vM6EGyT0wjpCnv4zHXtsA89XTE1y2ydbfRwyiRUggs/LochGVwuH4/z49QpVV7SdBVBh2eDG+iFasKU8hmkf0Po1XRoB/3Hq+RsXaG58PbeQCMv0B5PpdUVDVTEZgrRp98zNujByMtspVOA8Qkq9J0+zqF9ucQTcqqceToAnKbzMtyzmcxXitvw1y/VM8xkhBDLqLxVMQOr3L08IeG89XSuGpwsrP+na+zVHnMw5JH4zVvomOpaOTPAzNsp5WiWKSiY4T9/J5n2a7V3IS2wRIBQ3IbTvuqjescj19bXS7L2jWkUUJwiqysWzSQr2yszi/W2MC89QAh3VZDo7OnSvd8kNY6wdYnxwqkUfT6ZeBdmkCuOVO0/zAAeEPkLGzamnsdjrlrqONoEqnvyDcuJy2BYMhjfTQV/eXyPGbXW9Zm8nV3c9Nv01CZghTuWReWs/huZlAu6Rww5PLzAVi3GybxJDrj/8zhWCIP52ZvHSZ9eodh+12ppF9rVZz31N9E8PG68jpWp/rxLOZKwIjHWRVZCG1PkzIZiYXte5PRPP0kHV3a+foz9TgoXDMyPTwBQwClDleGHhdopY82qT0gYsemea8yScUoaUEtKLYYJP6fFS7jjvsI1FAc7EHceyI/riUD6Pf+inQhzLF2fOhTHKRSb04gE2f5sNwLXBFqk7KPiEBrJkYBXo5CQvH36F8zQs09LFLwQgVKRkhi9wWMGdB7te2khfLoIqVOInHOnmI5rkXpZCS5eDkOcDOnP3mSt//tyzT3qyPW6lP/TNAZTHRg6dqUb5y+bzO6O96Jf4BBUzHD5sOAmhBGEYtq1tfwiLPh07xCJSweCvjVule420BsrnhekqFsdm1FKRtjNQAvoyVgurKH1nNzIqhLhlO2FK/0DDrVLogtlQJouYFfn7bXDdnePzHIkAN2PPOXoGRvnv6QEjSAgSXPmDDR0/yGp9H0piZoxdkkksc+AcSvSL94WG8hIB6xTZo6Uz1lyc57yUltppoEWUIpzEDFtVYQLZQ4lZF7CFLbK9SIcHfb4AbXA1VXVEJq+27m1TSqFJTnuLOadG/5uU4vjsvc1yi3r+ppT+JKUTjMVlDAblwypkDam0b9wkwm4yu1BJfvygSsOGII7KwtX7677B+ypqjxsvBBLFrIqVFEBOEJ4+5OKueQUWE+JzAJ5vh987dvDnmpV1qHT3diM5G8j7GtrkTSFZvcdFgMReMRKw0tvx8+9pQhFXQcC+qwXUtvi649fzmx/7Iw3raGWW22hb4OdPSRV35/2zceOl0m/lUgyYBny6EJtETtA2ST1jE3gtjucy0Jt4SGPHJEaootpkI3mOmMTlQsbbxZzE23lGehfvUn+NQdMp4HHRo+BUsEieMOMPcy7DkfU6NVHpnRzN2m/NwqZ03/MoFJu2PIeeMo4bl85PyaobdesZ1+eUEFFrw86EZVm7+s/3ASWuu8u2GS0+yWdCB5L4KHTxSHqFEypSV+WzEAoX+zhU1t3rCagHIktPzS4/alOZRuEtMN9f25Dis2oddLyQKni8SH7AdGyGLungD45zyHKjFmNt59d7u7ey6gEZFN1SR051/SkPUbMvpw8pQwgkDWg/t18xhtpmFfWbNwD5CbIlG7/+UxI0N01jkJbKC1fyG8x1KOb2oHS895Uoy1DQ1tQWnuBVHDT8VqlWb8jGUMx8DTmeSvM4na6j7/1sRiJI7GOV0WIjEs/aY5v551H52LgdsBDak2bX99PxdAjoseQuAUUp4CTO4Qwq6wjyTAJkxG/EDU3sAZf7cAXGSxmFVgBCqal5HQVfheJUOhTsFGeXWNTYziVKM1xMl7AmJzsKyIfJcGF51HrLwxBaaSio8dD7HTTe+SGP6iOxvbgmq5xIWzFrdQn49QmKbni+dmwCiwDBXm4FjnWY1gQxPpZJOV5UIKEAtybk+DycHQDy9Tw10+cDsMcB5mBcPrCbcLwCob6AXrmHHqnuVTVAaZwlFXItKeZp5ybbz0ofbjiZK9Q9MiI+Y7qMgiGFWNtLUVSMlz5N48igRfd2uAwx16pdrh2YpWzj8mu8NufGtKGLkeg2RWOJI/hF9k8HSnoio7ty5yljrb+4IdXGuZxa5olSUkOW5V2bLZ/1FKqScQUs9RXpbIAQ/9AcHB+WDuKXbSZrnc3gC6JVJp2sQ+VY2X7hVJqGpNgU4eA2VVHpnILYwS45NTW2vA3b0CWK6vNElsE7wv87iE4qMTvmA0wsD5YsN6euNkWii71pRszC65CTYmAVXpoDrinZ/LTcl9qbxAMgj7L0GQ3IP9bJMjIPbBR7m+PDW/5CW4ZmN/LS+jx/L5fhAvBw2D0nXzY++7a+D+mZseemtCPkYJE3Fi/Sxc2saBHAQYoGHyqzWn0PeKUGRIT8CfI9j21WqBrRqbYYOcT3Dh4M3mYLOcIy/MfMcG0qgmmNiCh48vHO8gjYqfBZdJreHIgPS5YLrki7g5kfZXGikSwt6Po1lKFiBhO6AsMRagWIQU9pSQxblW0SccQJbufQ8WXCLQEjJRtw1m7gLKlVquWItmBT4mIRVF8pBGsL9/3mAzHym0467rQiYK0YA7kVxAyX4pBAPdawOWRnDV4A4q5QAletH6hlpcMIWW9UE+qIauoc2MBgwbOi+07eWEeoelg5Lru04UlDS9f7mNRsSfxZyG4gtPWm1O9OfyQ0P7VfyEf1EoyxZckoBd2+dlUC7+mFjWOBCgruV2wunBl/NpqLqn8S4jvz3fBBDSCvPUdRoRktKBN32P8+/UyFGGyQlSpzaA3gaLQY5DA2zK5HIXsxxjAdo1nazYrvgS85Opt1SXA9AdrQLP3B9AmgzVehsrwxpE2xF4O+RxNLQLCRc4/K8jN1XSNy9Ehq1ftzmEc+HoNbD6zxftFJPXxJqMtU2y+xiFbjvCix/mXUkNl5RtWlKod41d1zVevb16M2MH03DgnHehuIPY4Qxb8P6Qx50Rgyty5ihOaR5f/rdMF0pdf7I+0T3yE0sStaaVsbOiwk1YtX+rMkCJfSq2wahMTRQi/+LL4/s4uaxyFtRV+vx7XplVIpPOc19IXjzJP/dwhAxKga4biOrJzi+33fu5OpCQTHXxW/Ra+rsTi1TYly0TGn31NfNR2YzWWhnorCTMgb3dqdAwzToPt1ObuPsoMhAWQWkHEdMFF/ZU5xpbQMDFaSbqP+SxMN+tUpGwhwuACAb5zYKCxfv26YBoLpaXhgaYNbRqCojXJPvBbxnCLjlSSY2UCYQgPgXGaQrjE1JTKo+xDtU5eevjCkY3pAA5AIvoKc4lgHvnHcODszrcqMYOiZM2t0x60WnXTwWbNeVx40iXmSefLQCDp0SQdsioEL8hZK6J/NbLwpiGGX9k3ptqm7cQoHjzYRtGzRovSnUH15tPiVFlIi9AXQ4HGdjzxxkyqVMQ50d/rsxV87bHt9gqdJGOCgE7mJ9zlofvIvqcSOYbi7EvP28wMAMj3sl157tUMAkZUKD19G4TSI0J10EjyfYQ9wjuPF1kp2Ku+G+mdjYFeyQBcw2f2Pd6M4ysrjJnf68SffiRzmsxFeg1T+aonR0ugyh5dkkJ8XJSQcDNR8HwGfN3b0F0xNDX1N0yi13IjQqzKLVSwGglmrFUiMyUP8frNVLXGB2FlzgbsBkvYUq2LVnZ3PdLfHOM/+Dxn9uMhkHdV76SwoihW7n/cTEFS/BZtjhcUPKJGJw0QayM+W1xLSo14cuvWl6AIz5SVGNKcMVrXUd+C2yv+2EMabPiIwa3rc7nSwcOU6uMIfgiMAFwhnNoJqkZI1VZDFUB8eBTOLdwRPr0HIFy/NtH54vx6A37x8TO9npVX1tek1V8BJJvN3x4scfUj0rT536bl7c3VFtxv6bD/o8kNAjolUQcVrov7vExeCo7HYI54GfaFuUvy+8FbwlFSuH/BKogD1ReQU6QB6AQ5baZc4N9IjPCWEiwY1p7vWdbbCskXrNMbWd9zwIO4DJUaILT8ngYe/i3Bh001KmTbkdCQRbPaMIC9DmvTIbmVa9QLG0kcGpq3oASS3Pbcd2GxvLyofAGJNgYhvWHf//+uX1QZXNTNoK8lDkfCCrGDHWi1015VsRc/n481c8c8Z8LDKW+/7RCQ6pp4hQhtlZANPKv3wOBKBRdKRq2rxcl8uOXo38xGuVEbSPKEUBXFOpasl/AHSd/6P5HhQgDzzSctxKpEw8uj7NMHeOxBwYABEWhIAenpWSU/eNTkl6FSJnOzwTmWcKfWHsTH2FvT73d5gFKqb4st8K9t2B0nEihpEi0NQ5ZrTuqIXePgPDfKUcq2QcR8OOaqgccNFuSpcbvxtIRQERDKk6/Jal6hbPyLr/q5UBBFVTVYh6heiSAyl/lZtqWsQPjKrMg+lDbQUk2ZBiKff3YMfiH3xgEuyCd37JBDJms4OPUjksWlrcOcXYC6svr/uN3wWacrheY7RWpkKNZ0eNjEKznxmnbdNu75Vkut4TSD7zBrMIqasFObgo/L+zgzxv/ebFiT+bqZNwxrisxkpsS4UR7/tSePV5ur2qkc26mA868l4A5LfASVJUMXj4+prDnMyLHrzNTmMPb2IEIqdqRpN4VmrH3ziHUnxwzPlsDOOTWEYg0Nz9zPzLjeZF+o2Io4+K0tfhYxKC4/vHU2bXJTTDeu8s1IG5Npnm1D8mvmPsPrD0euGQeApnuzz/7wawL1AABJzSkmNKQt+3XeZYHhop6addHL1fTcKG7BPbm18lk3bYmU+rLBEHH7BO6GCrX12ctn9j5Zin+evWN+IPF9qwu5uyNaPDQpn+7pQ5BpCifhP3hwXepYl+b7SxpcG1vUzo+EqfL4NRB8vjemwP7l9NHZJ7L74tO3rmP2QZQ4ahv4qVMKrdxvIhvIUbbGTv2E6a21IZgVAc3K+oojLdyU6SHgoOuVkApX1Rlz9f16KYZB7ndMFnhf8U+qCxlofJn71P2g5wZChq3V1xI2wCIccY+fQt8A/J5Z2Z1pHvo7LlSmMWAkGzSdHoQL+HK4XkYgt4SOlFgSbCoExS3mKG7dzSD+CnzIbzEx/aITfKPefosWmGu6/ExRhyuwtF8cTI2SD+8+HUoAFgDTPGIMVi0b7OdWA2fpP/3/enaS9e6VmWEY0DdMc6LcD/1/ok9oqHNBDHc5WL2zC1coQ9H+SgBr4IK3bNtGBqUFHHNS7qNUxVZypQHy36sOafZLpAU6yVx/mbsDljcI3kN0p6S23OtIQmBQKKOrda9nyMFpBTzT6r6drNpfS/C5R/0J3UPqCElMbFP3zPdaKqxVJFyS8WCieIZ6say9e6tkgUbVR9q9lbDYz0WDLcKkGWCYs4G5+Qv/y6d1A1TxFgzh5gVT/B8v/CNfq8o9FM7xrFchnD22YMRIWONEa1j/bm/sELERyxqoVxShasiHzoemEPPJ39ZAKlgCBaTCqYSSkAxUSWg6WBa7kMCu3S3iCJSre1J+0cyBoc3UENVz6nxfZexi8z1O9gIXJHeULi/lAPFgOwsenHu9fUaXk7UhTRmiZRCw8EQZ3Zg8iAv7a0uH6iz50XZRxJomLK7ZpVR+GSJ5I5akLJaJW0kDDTa6xltKA9QSAJ6knoIG6DDAEWh/wstm/rQlwYHEgFEjXPAAL41P7zlp+ethcibHEWzLZxtAbQ742xvIt+kowguRo53CWFG/8vL0t7kRPtXUKmiqPbPVsFjF8Jp2jn1Az7OxRhwknJ+suFzHfCNPpkPeO69PIXoBHEcn4xz3N2/bYmuYW0b1r4XYjSbQEcFhGOXm8AB1RLwoivKuYClUnsuzrcSsCjFOhgKIrIk7udh4gMqpz7Vu1uN7uYZhZMsfSE1Dm0T/lyzNKZrMyep8Opr337cJMMEt64WPyCuk5/Hy18VP1jPPG1alIAzzkfFDmJ7GziKXAVWUNfgsDoFandMxiwZVSfR8yfouJo196QRPlBzf80mG5rEIPlV1Zzah9Fk0a0ZYU3CBIrxwSBivlq03XV9SgNJDTwFltykmGjfGpvArEQDhK7uHG4ZB0A5EJmjO6/dri01d312APe6mehj1MV22U2dwTyRXJUv28VzKQHDbLi8EQmiIvyOhvaKyXPHxHE7LQ/qPyjJileIQmdJdRemWq/Ci5Hr9YMFAQo7FnZQeoPjGsIXtMaHE2csDKri5X+b87eabRfiLTbDQHZZjT5NOeb1fxA/jPhm9b+u/9RiwV4Et+8VRAnsDpHrL+h/gHY28Kv1Kf/6LH+nXu3dx8RR+LIo/pFDgJY2LMudO4djBHbJ04BLqylMWV1/TouZJecTDt7e4IOSO5zuwVGnTDkXLj4hZfkm9vjw7OrlrQwILb3uEeAH4/md3jA/1HT9ksC7ApcMv7oHbdQkeMcBIygEWTqUL8lTyss5MjfskvMh7gK9fXD5Wr0QOHVtAbRoRsG9G/VlfL86HiHsH3FIx35T4n3qRN4r64gZ1XBNlMPsd8t//F3nQK/PadNOgyZ6ZZNXRHg5QoThBGzgB/24Q4UsxZAPFeKSC2f8pVbJfqH8chL+RPWkUdnH3AQiHd0Hwm1wBDIgHISsf0VfddhNNYrkepcIJM7lnsU2Baid5ZmlUizCa9fhErS+vTUvEB3nEe19jl+6HyJ/n/4N8PZQ3YiaZQuJQsHDr1+7N2IBl9gNA5UA4xcmlrHcXX2VQNcGXn80EUFDO7FYCsn29eCqr+abCWvmEaAoIxytS7ZzHYK5okQxp5u2JxkMumJDc/xyfzit71d8/0pGiDczUdRybEvLGsjg4E/vOSsu0hNOILtcN+0+ZuUwsfX+7R8YSZJZGdOCR5Q7+ZgzqJPnmKmEDepDDGX3dJC2di16P0IDIIX0mSSmpXLL7V5SvUzg3LKixMuI2Q1wAz2E6cvDinzWfLexbqYja0VhX8BE4pYb5u6d8tRQjuU5IrsNohuVofL0MN5K+zHDJFfHUTqrjj3QyymeB8m2oAFtnuNoJKIS7JwJHurywJ8GjzgJdzmi4d9b6rs16pePYNPpO60n6PRFAPG0BzclD2hyCzWR0vfpii8JDUv3IMZmIybpSr0sbOhcMhU2tyuKOTeTJDWzXwLJY6+mKTqqaosycTnJryJ0UkShyzkLF9JLa5yxkR6NgsE9ItcB+QEs/fgxqoUac9WTCx+AkcrFpG68SCFzy1Hscynvu87EuwuO2Si6v6R+OeeJXJWcZ8UrzqJ3WuuE+CKW8V/G2+VAsldZLlw+93jj7d3cxSY/8uKYF0JdxaHR8UE/JG2+sUmL6bPhLFiAi3eb8ZINa0g2VydDM84OHdfxwtFAAYIwu2mb6/jnFLFCkg4VIR1rRIB/IcxnOVdB8kX1btMasINMHU9M3MCdwEtQbN3b6Ja6In3cRbMuwCCAuqRTWFIFwNhJJk6fQMajxhhBfmSF1TT7sCFzGpi5XYDh6h8L3zz37x2K2huU2P8Q83Dx4+ne7sTfkKhmyIENttTqg9KqOJ57+YLbE7aR61PFdrVfAp6pD85nwQM61nCUWsZaBh155xS5sr0PCryKeU4E/5GdeOF59xYAW4EGaXIab1VDLcpeBN35q8+uFYFNVPjMGzV1BUYPjJb+9ODgihTL9gbCcFxBl/KfP6T7pKeUjEc4VYJAtLfw6Z3lOexPEccdUTuC1Zv8At+KtjtDOcw2Pp8Zrugl5REjFLpoQ5K0umkloZ1RSpJl5Z8jUrpML73DJ/Q5/Ur+SPNS+jmmNpyz6Z1uyWp7gOThIn8IDd2LilIiB8Z4dbh4nfToi7FGwNzQg8P2pOcuwfy/NP1Qb3TuirRgAl9Sm1MylkvmY59RltnfqOS7Ulicl98UI1MinlMo8UZ6KEQmpgyIeSHp9JQqt+LxrycFiHuMFHJzlUQIrty24h+Kw55NkDk9xVU+qub/eI0wEbwov/KurBoAsttEHhUS4FkHKtkNcqyOJ0/ynavmTpBltAtUiapokdNqUs3XHhKCfxZ2uJVODF1512W2tpi3Nx/71zIwXP+nTZMA6nKf22hcX/8WsNjcJwV1eti0oY0eaoL4pV0QL3ylhmaKWGksqxnkkhFfjAQWdhwY3wGWBRHdrLCOIeGyZde+TncGaEF+LKmMT4xz+surIcmSLgCZ9ODirk/sVPwUJjAcn+CyZM/aGwPpY3R7LBcAbHH0B3CZKHLqaX0qc6uFWm7sTW88Xp+4YOzDwJGXT7HOtGPZGaCAetc7LIOTRlKSvlyFaMIHo4rvYp0/amQ8akFFM01YFfjNoRGFrs/+TK/urFNTC0siMbAzKcTddGEz/t8QtBQkOR4eruEb47hB8tWz5KKYfBicy2IfJjIQeYaii3F60z1M33I5IGMLOMdNJyO9PBBDi21qagrJrhLjRgg+jhqJzKoomw7BwnQT54pe+7A1vxLvSdb5LR7SVouFgVjVapIdo8tgGf6mf9t0zqB1rSM9dF/bHoedgLZlgASlW0sTk4hGquE3f7bOScLvFVGy1FKujm9rxZDwu2sHi4BonzNiirfQpgKikLktCygQYrKEMlOHiJtcHjbaG8z1mvQ/ZHXRBVGYhAfAP+2OOHmaKlpVrsTCHMdBXyLZPEoYGu0sz11vHVi0r0hGHoku5TZTwTPyGUVlecQ6GxthLJ1YugY3IFbLOkqfFiodxWpOZzfH1O+ChzNwW+4I9NP33jov3/kDzbxNSImcXPkEml7bDFlGOXIwFkcMR3BiM1zQcAgjiTB24fGYxMSyRVNUZvx94NAZ9hX3VM9VyDP3ysbxSoOL12TTkkLMtkHM9tfMurOHPSORV7PNO8OaZhsKkf68tmM4sYb05efvKuELU6hdAaL6ZTds7ez5BPCfSxJynL++mKYc/cf6ACm1/JRGFiGfEG4b1AXnaTg1nWlkBUtSjTaa4xWNjvvR5ziwkVHSZirVEBxqtCcVPnwCzmOrenxkQ1Vf5nnJaadWctluyuVnxrdF2LfS3Ud+BTSxbGmCsayD9teO+adTEVTYGw8FDOxBV1DK5vDPWbg2CFtFMG5XCGo2CkfJaG5IHJTEGbY1pyyBXWdLPDBY3ApKk2OEOUg2tWohKo2xh+A7uB/8xeSiDfHEX6gdnGXOfXXsiHqyUQkWFHNqPRAA0W2LHiqFuvYSbh1flPq5qM14NKRoSjLfiYdFq+FM2nTs2fTIxZNUWHuSTKnRBeZnaCf0oSdVbflczOn9vivBtOJbAfe5W6wM3PUHl1CGbWTj2x3ZhPJyeDKjc9qY6RBoY9cJ8DetwP5MU7OgVOarVn9Ge1RDhW51i5By3hvHmCVHvx1qQy0RyHQWMOYQyUI+H2GQDnOTN6rjafJlpIcKH5L0xTzHJ2OkA3LxOw19RIKoslFHDd1coXtMROz/STKqhANyCPciDh9WHAIDOz1dch5kx4j8oxh5LtoKg1yYT4HYOISQIlg9DHTdzWg1kY+4zJXdeEJ1FWXOdIVv7J1z214sCFnedVAHe6IJUZX/qAMVolYomuxa+ZIoAdHmsevVlUjfLstkMXorhwlq1h01/ux+MEFeTuT5HiCgtGgAU32qmlwMM41iBxNXi2lO9X4LYmDweRTawE4eX2YmCJKhS8d2MyP+z5ExPVYkv+xA4EdzCbKbqQnez8FQLBGCahoJXdl7PZRZFpLFHAd8Owtprk+GBn17/DV+XHz4tf0RZlttrhVJxreRC6N+FBkezmLyFESqZtKe74v8zgV8NaCUmXUImun7Z6DR8l1i661W+zLs7SUk9M2HssOdFz1tlu+PPBe8PovsDyiDzyINQA84LsMd82uqbJ1xk8jhfdCvKsROAzGCcqX7FJCqyudKMsHghT/EDb9HMEYjVR4PGi5DmW8NyBWGkN/ESNJ68gOTnnWtfs+cqLYbYwLHX0a7SvaLVZKNcqWPGHvc3jIYUyps2g37BYqwFMMzZMM4eETMUQQTOFdJuiMXwqkToKzkZJXSETQSt8YsreAXcN72N+qo7/NqwHChU8FpAUBwvzF2jim6dZ3Mxwr9fKY2R4LtkHixJQX2v609FTy9nRti3AkX1/m3YdRM1UDUiVxMAU6fR91wkvHFpoXq+LNUa6bwKQcQF4qGoSQHQOWn/VWCJdWmco9kbGI/dTtJRDmtw2uAmXTDrNlXDJvJgqvU8kjJYAkoJFedMah6/pk91n0HUSCN+eyzHWNQM380UhAkTg/MSsld/OC4XtHEEBejX2cFEBXiOfsmrH+V8ZO4OISij0FPhzy0w+HcHPD6p/mqu1V9DIEoeLxoNQJ7dsmce9Oe78Lp9HLHyBz/SJm22YdZg6/0FlJp2RwHQl83DZ7U/HHqpjBuiTRhTlnzA+A86XwMGxEGv6qox/ELrdWohUb0koQB4vAby6M6UbQAaJQSWOXdfO8NS71EMh3e4cOKbkpeip0W83LF8Kioaxs6oyjOXGAuQZeaZwETCTsC1f5E+n09hOIuc1oOQZsrmLYCGp39M4Faq70rJQKOkQ4LAkVMbgU2dTORJddAZARS6mmYDrscg+PQvBtMm6Nmwu1iztusif/RWSWS6DbRvvNe1O9HZJ2w2kmCg2EEUZ6xuRXAaBsSEIdFob7/AL5DrZvKwQlhGUrofEA5G0Y9/dwA15xA7PDaTHrDSauZchig+3Kv8ejRma0pPtmh9lbwhKUzeepOzwLkkaKXnuO0H0hzPufJ+rAl3b0kYlPHQBns5IMfOghg65EM/TKC0HEbdHKXjPGqplBd2zZ4nlHn39hfpB9lwmbAUVN8b8QaxBmvzGlcst2gzK0UQxpzKyO1Qj/Zc5hcb71NYWY/ycLZEYtIf0A4Wzl30t7G1oiWZgMQEnE5llUBvPRS9i5QthvkRUuZVf/cqJ1DCgdF3x6PhBCwjBkLFp7rBCYi46YxWIELF8IGW/jHlIj0ta9O0RLu3fGzxPpElphlUPPuzw0i/mLPhymYhXi8i3QnIUItvQyizo9z/79mkXDJdR5TssU42l8tiKedfRBILtuXBTqqsGkgEOsXOTNnOOTalj1uOwDV/72wdGGIG2DkAO5Me8AJmYgAbRMfT6RLKtKKHbdwGNrmXRJEmUSQSuwIANnMxpNQkhlr1z+H1yytPbLLcNLuUG1IKVnf9mfCAfEB/ARVnDbtrf0SO9291ixzUP6Gsa2uOh9NJfHZRZfJfpAPBR++Tma0Movn1PV6NYgWHdqGHHPyvTV4Js9ZA+SNy/P0Bf9QNzZDzlKAaItCPm98JkWKARJTk8bM9p+LHFV44/jwWZb4Xc4cqV85N23FIlk511+0NC3eDX3qGxwsGp9TdmCeIVsNZk/E5nGG+4Absy8hU1KexmaC+IuxzxGYcpi8RcKGpKsKtlPD7VmdUAENSYcH9bHKeqsLS/UqWSKdQCobFmCX6vPXVlX9FSiNT7zN0W5mtQGUd8yOOz9vhe9MxNDww3yb4VQtBPBNqRRsOok9Tv8k3JPAo2hWUKQSvkrQ+I/mcScfssKFQs+so6FJ8kD/AFpnynISpQ7B8E1lsDG4PQleumEMqecIBtI4Ua0XQxCadbs43x2QhHLYS8PdtSfF24gkbHPYie3p2HnIDw5oMw0JAmzgKZdsmwyUpkS4fpfJSpG/7ri7kVMdNjRyEIktjued7ZmA1jDmjB8tWb25qY6zj4PKkA0tRKL3DvE3RwDJrUTar+UCwPTJCm2xk1vcAF8nqW7ZTVZm0ylSbvecVuD3NoVMgwZezmmquVlEWaGsUrj9+/7W4l1tTdzWOhGSe05TWRKg1gfJFVnnXAu6aJa+tchv9/TnSeQg10cUpQQY5eEQcyfz8+0HC35vzapcEn3nxaDkn/4vl4oo82GZNQUnpc/AKyNOvVsDosyDzhczx5VkOVmdW5Dq2afbhpAPSZ+n1c6QCuNnmZdrMbNLdJ9LTTIO3FNJibxX+4pYwPw13XjIwwOHI79XpnpuVe3WwsuhPwIGU12KIROqEon9xadSNBEmUDs3INoQkKVJp3/7b7gv0KYCKqpgDl8JTVu6HCWUDJchbH0WIovbrziKSED2YYTBI3xXER/jEYRnDe+WMnLLaiSdEVUhIzrZ0Vz4yk6cCn0aMf3cMpRRBEsbraeoYLWwpI6+GcYlTXJyB9ExPqz8c9r17gEOAaeQkqzojZ1w5LtqBbt+TfnKEqgVVid+rUKr1jST/R4qMMLw9RXyVBVUe+ZMn3+mFpAQAy93HPzGuPFn3mnaan0feY9wzSpV0ZXQXzKrTOlqha3TYWEZt6SrdZKjKuKQDavJADtDiY537GkNW4PBawwccwZz3eJSwXlZMdUE427iMN0+zbQjic0+lXNfOF8IZoE1jImyG9wdzImDUovFbjYV7ZOQ6agrmwh7MISrVt3j3/alfb2FTP7xN5WwgcRv66WaJClaCZ6XIi+LnY9ddP4o/Dd8deSFjASJcV2vWLHyuhZQ+aK7ttK79htyItdVbIKnsOwsjRjjLAITFOolIus/XzjvQI4fp2yWAG3f0Nxws7ybjUKDkqPlt8wqD/r4WxCLl17TgDdQGHl77TEDfj08hXI2Xk/JPk0r+wU48CzR5LVY9IhNb7m1ONlNAMU72BzopDvq6kU/U0bKRzzT6JQymhNdHw+vKwcGKkUNnnzhzPzr9VTnKQIrVwcdeb4Cvu9QoSsLOOttKFSLcQEN0JaonvmNamCGJxdpcZPWGMIxIi6ZYsQxy3p80VacqkHnHxUahRjgzXHFhnMUcm0nGvIWuv4KNrCB5nLLBd4psG0BzvZ6bTDw8CU7kXkYbjDmo8r5Guebce+A417Fa6aExm5GWs5arZ+XI4jAJFOU/t4metSrGogAk+DBZsq5dY2mF69ESsc+x4QqHdtZ4UKbpbf71npRMoe/oSx5/ooo7GSIcFIqUDG7e+P4hsLtQzYwZ1RGnzR5pOYrYjRR18TWtyX4jyx2ZIXraiP0SGnhJP6iWtG7NoFhpmWh+QhXMrfsNRIEp34PKUpM7nlpf8TVxB7iy7500wG/y9viUHT3bmhmXr8XjgSGYFMvXQUB5rwybSDAIACMVqM0RW7UHEuvXdECmYSweF/mFlRgwAR9VxfojpoKlsL0xWUOz5u7avHtFtizsoDR7miZx4sM3oI+vAoKMnXPXQjKkuZG1DAg/9FIimA3u+nZ58RTp7DIOp81U4rIcjSx4QRiKwEOehPTwvjWEgDY6mqPa4l8K8/tMhqwNkvARJeXCIbQ7r1bsmqFE/gg0rP9vwexzGKFDoqtRfR3bB2A6vrs20NBMeV4QPVIkSDHWjyC9bQbbWGKya6xgQBkPpsH1rFR9z2mxSU5TvE7zYFeRq+RJfY3I9SPsWbvUxVqg9iHsx8NcAhIkyy71W9DWak+zPGINsUZBtr1z3mzxRHsu1k3BR9nOaCplK9Z1lgXpY+ch7bD51kmDdeSEaltpWUqlYXc6dnTLSC3Bnk+BuX6+yE0RFuz1onDdd23+5JIpVDq8QJV8ZbQCYxmL8hbNyKuLEeElA51RKBaH7XpnmtbgaAyK/2lCc+qw82u09eGqIsjnwTS82SdfonEmux/j3N9sM9hsdpnmov5WEETre8d2c6jukNDO1FqcXJ9ABppeMPPzmkaUgfwTRHjBBzfZcp9YajHZkbjNGc9ZHHDOtXZWG6otQfkjluuMfr+HLDG7Kx+2Lvw5xjBre39MrvB2WXWsu87Klg3Uji7R84PDOmoH8+o7JTYqvRvp7jtEQoYaR1Q9rlc1RNYbWkrMp1Yebefnw8C3RVtAfmEhuHo2iQ3oNs3aCjFLuVR4StuUN/7aTvMEYcsZdgYb/v7Ch0Xgqwm2FudyDAiMVKrMNpFzqHnt3x0cZxKgB0nAcgjfNE58abg91BnoLoKrlOhPOLGp8sf4Y6C8+WXKyr1G85iFcaFDSrM8s/MbII983cAOF2ibLjhgyYtyo8hmXf6KBPSXJutYWwWb/SvISTbMcGVh/2LX+He4bBqb8V4/arwDyw/laL8JTeuEejb1oRvPomk6hinSCH9CQn/b11SnBagmXYWIOXOmbmzXUNQooF7L0Y4millOyi8CX+UT+AUPRb7K1JbpAy5iXzHbCz2AIiLD3dX3u3Ws1XaTFnxiJAJ4/cfBnhvie6OANxUqXVn9fWc/IErJ8+xWp238OQtdOwdpA19Ea33vGpBgCx5f8ZTogt9vRSktbB0ZKKQJW0UMa+F+El3eolb+673ePPG4bTPHyKEIq0HqmpY/uEo1EcDsdM4ad4zSSqoJVu7YJsm6YbCbpbUbpwNEheniV1iA7k+nWWBHzoxT3MCWGV0y3LeOI/X03gtg0yfHvpcjYveinoCrYuhaudTtHNIr4zWn4NlFvwm8z4+NXxnhYJfyiBJ25J0MHO4iIwlP1xNG0GJkRINEk6m0Gm0+FKJxhskam3d4ZlFANJLNsT3bGXw811vzJriaCg50JlUWkHPBsqaRTqBUVHsJjUh3TpCz/tFvOHbCodAOMwwXM5pxY0lrGrWnl37ar8theo7m61zNB7Ia+t3dFs/8doXEEtAjvQIFDulh4RalFzc5vy3niLN3BFWZu5FMpOG7MWoo8OHtrha5syL1hA2J15a4HTBYnsphM6Uj6EMm6tnViEF3RDhCYfrFUGTd0Mat1vJa3TppCJ4K7dzC+y1b5cdWvqz3AP5mkLQlAHL2FfNIPgVohk5D0xTzpP0X+IxaqmIjuh8ocyvBOXAGUgJqKpH1s5sHDQSPjUtbS5XPqf66TXYw0zbsvEM8HKNZOeCYAHZcRahoTg/V4ulXgoX2H7ukhapwKijUo6pkggpAioEQ2IWG4UgmXo3b0gFC1j7fDFS+9jqvUv2eHMWtGoKMW+Zh22z7vqgx/lNCDUnDHM8YnhG9SQOs0Cbe5U51ZhO9sSIR6WyG7zBgwgaCmRvmuoTQKR1BogHmOMc8aFIe3CS4QR7Lcy5W5NKL/x2NamHq2i41OkYsmL9IafBcH0R9BP1B5yINcM8QJYZpkFWNjBNdd35/Q4o5gb3cPF+uClYlnMxN5rosPVfQMwP9izkVGVJVwSVyC66wXMmCPUiZh6SaZqosTBrnaCXbTUYTlMy8jXujkwvcg9WSTNugILBq2bOLuS+XYQETsi/WeUvWmh59FRjcQwLImPsoIgDGFOnVRanfGXSLAqLGeCMTwrcHsE7ZzVIynN9BF4k2YMpX86v7jROC6ZApu9+H16RI+3RIVt3ve5NHkv/+M/mRUbsiHKndZqrU9R4EkpQV1E3Molqdzrq8IFw79WIa6z7WKMX21APMfvq/JmTOJcWKLrhQ+s+UQ4TemJJ1zdpG9HdPJKxbUSC4zPtEYfWQunXrprhYT3oHgNW2S746qsVYTDrBYKtsuhG/xp5JbBzhkMTG7/HbI5Up3NJHPyM03znYC5+huExnHRuv9qShx+ak6JvNZF0bAhNwFNfNDWp4D3tHbPP/FQEyCfP0lKA9E0+KkMYsLkp6WaG8PPoqAhYO4VijUusm7HZIAHqa836JEPcPKiHxoEyTZgLA+KJTKWa1AUr2bqQVIhlZmJrbsDtGWPmpGtFf+bUHSlnefS0u5SxxtTOdpFo4lnA+APRw/tEU41wHO3Y5be3+cAqbQW59WkQOj4s9Ftk7+OaFCUL0bHjGH6l1hvNXKO+THYfu71VKtPz1K54hpZtk4c0Buh7q/xdgc8xlMl0u9V5rleNty3n0p/tm6eUi9JLKMPksXkFjbIu7J9VQ2Ue5qDLUXQymyhWUgrrKuy92ZXYSoDIhmuztw1aFZB/XZAh8p9smIpR/sIfatLbgmgnog9+2GDL7oqtu04zIw5v/vWZRhg2OFnBiSN263572+aqYzGgj37lrsySsGO02QxDNsoURA6XhN7otBrtAlNaK9zke2P9SEM9kmfOlLUQEdeqWQsXyLALof6FV0GmUe4CJV6paHn6BoTRAiThb6nMmBcicL2l8l0CBHWvjD/XxY7KSloii5KaxCPXmCZ3qL4xrus+cQOx5nVgOxu7oeEMHnMb7N+3H3NdSteePXpm4ILpdpbjcQTYeXZAjMOhGQsJ7LK0xW3EdKWC5HAQ/rYr03CffmDJDh4dTEaR4FOXoWNQ6Dw6g7ZPXkrv8RkCnyOSqw/bGyTXiopHYSgR9b8xopiye7a+L4AEW+DpXvkfnpzZl2i4oihltr8jTJew0MW/CbAq4zvnR7QlIpNyWZ8nHkmGD/HblTxMGuEjgyvzl9i81apqeP76RkdH+O4PzjjJi0lBJekKg9ZIf6NXXM3C+s5hTuLm+5KBqugr8VU8A1VJtRqv/MwXIYxar6EYrVOgjzf92HK4NONSHuV9tcbu4e0XKNBep+jx1hL9Aql+eNthoyVsvXhm/pMMICJ84PIB3fnnkGjM+rS+ihIz0e14WKi+kT9IEWdJadK9lKS/Ctr/vqqpDelvhY0prTmPl4HWVbPuLvFL32UQwCKULXfmASBJabb+uxI+IxfOPclyVN/QLQmgQLZ0tiOuIOv0zxAgGBKra2cqfSS9PJQfdfQXF6dpU/xV+TtUV1KuG9WeocBJvt+aZ1n+6itYxjuYYu3wBwJq27t20NF6j9S8TvlnYHZbBVoRzLMx+bJDHkInnfZfa0LlIEnGe8ION3DxjftBN4ozZnI43FOxwRgu3Ipe9BZCdg+jK3Je0UcHj2EeGKHX8Aq14npbaGM3o7QzgHDKebWQ5tqUb2WxEkHlWp05Nhs7InSRgHPHl+mUn8CSKKlmE73DU3fhV0vPpfCGXZInBOepcGlBX8wOKDK0UaLu9R2f8pMM82RTPIcoDm7FIVZ9DBLp6IB05ihFDQzho2TaUhvUmtm4W0Q6A/qcoOk3W7SJ0kaYJMyVGFjFyRQOjNGLoY1KGq4LFhAQn8iksREvaEmy44uae/11hGL5mx4iDJtBzmm1BLvUkaCaPMTgSru8i3wZcKxBiiwRWXUj1LKzDpDADpAA8WrDd8huO0XFjv6KtfI+d9skPK9f9X0sc50FxDVUObd+qA89xGwq6dZsVEp4KMnahfh9wKfdsgn57BBj5tvSo6sY3J+ymOmh7cc07LgX2l6tomwOgA0raIE0zUtQVreDygryGdZpjPXZ4HE1hytiCC8aStD8F9Ff+jHtkTuhu1uyvFQfCPTObdINmSC+0POrjeRTRYt4h2Yv3qDWKJen4wScOByZsbHgMR3In3RCc/nQLESO13gvKD5bMUm64atHNMxMbt3Sm+vPpCTTN2ZgDWQK++oHE5BfqsYbOpKiqObpyKFXpXHMwj6GiA1QV9cfdc441EppmpEMT901Nqzw+borxyqBxpMJO38AUazzyfODTNRT5ry1NS0ORWUM3OqZBUABtD7lXkmkTVBjPySSvcOgsioJg788hsImxxCEX9D3MpIKbJbsDtQGsqwSJwNeTDCgCM/0A7A3mHD/Dg5dTp30xhp8MmAmqEXT7bGDy+6ARDJcjojYHk4cWmmV5D77onYZYoYj+4hanKmFT8Alvncg3k1reSz84ykL6Wg0FicRpV38rdZfzdWcl520r23qm+ByPBKas6c4myKrDHb5H/42AfLeN1wdOyHciQiCQEJwJgdudB2jWL7twFIgjRIe9/P+EIoAIzcLLnDadKDHmvbp+QXRsEuSq4/uTF5DW6xz64Jtq7eW4jqeTW0wlfWuyNiO6HEQ/7JZ0snolaLrbb9GvZsYNihkwsK2darbaX4ITrhWKn1jgo+UZGcXAeNPToc1NrrSWsWfmDF67oIN8T57vT7JSuc7bsmHSYf+Ie3UHmc3mg+sDFEdeqMC5i6CSpdMuoTyNH0Ns03uHW9BbI/HkXK32ze+6niRScYn7kWTfds55oRcrLizap4CqM8Tw+qhx5H6K5/ROb8pvvB1m3bz3hL2KpXosG0WllwtRUihg4GPD0HjILTUmfXbG3khC5NXNdu5jLDxxDRlatDRAsar/MUQu13Vbby3/3S7hU4AJkKYcRLrEe10bMARj5sGSzR68XzZa0PDgl401NadV+v7CoWa3zlMtC0/uRa+TIoalQNllZMuRbur5WPNa/cSc/YU8c1P7kuLhwHFJp1JNAbkwuANpQG71wBiLjMMZQS7TWclK9rxeW62R+GA2DZ64FOQ3qknPalJ/gkQb134gKnpR0aMVTE1Vfj4OLsW562OcNHlgRLV866HOszOaxnS5kRymxe9/wMd/dkMN5GGdno+tA0idoDrDYEy2dgd6DgrpgMTdnPLV8jS39MOqJVYWHJb5pKaNsvStzLuDM9oGLhdbuucFGoeoI9tIjQwmzjFdig3miTeRRqeLZpIxL738CKnekncJKx4IEwSA0Ira/WnahX0cl6UNSuOLexIkttqR//xxe/22t84y5FC26JyCMh1Ho1FCz6aulndbK9hsY/4APSHwK+uMN+HBVHBqp4G0IRwbY5074s719DJcRYvoiiDI9koQFnD9oopoqugp5/JHaVphFV0PsLXyntP2MHhXUconL8zWFRZ0v/CkZpDhGBlNkWext0dXEawpyI5YZB3SrqblJdCKGxdZERUSRHL2wtJLu9rAlCg2ozIxFJYd9nan5re0CzboBhTt0c0+SedMlRp9INDMGjEStNsaZ/fNJFcfLcptRymvkC2EkzuryBBVWoaMxDr1Qpo3FJjF2UUzZukxyuYOYBPvI8qoziKcj7YNaD5j+qzLGcWpQa21WFArAaSV9ClzzDzGvOxooVxiigZTfAn3SuN5BHGBJqlNaDsZW+zv6q7zflDLxqhMo19bKSn2gsfhj3Dps17s4IwMLn4X4bJ1ySWooKzOiJ1Zs/ZWYuG5RzTECTwGgk+euy5Mgeu6ffFOmsPj8qffuboiwPNeZfnqkzcXK27VdlLDz4v981Mtl73xWZzW4VgsQ4O3ISaeV44siXoSlfZLOrBPRPtLBSdN83ak6LWC16U7upc5Bu15gDGZjX7zHopKLEd8u6ni6O1ad53zMue0Do94u6s2BVWqTZFYp6H8rpMn3kf2zHS4HbNQyBWn6xDLwRS+f0iBM/YQ/ORh0KurcIMWk5t8pjlxipjaAIHwCxkfrO0WScH2DFB58x2LkXtwfpcGuwnnWlTCmHm1E/ajDkWj+yZC9HviijNLANgOl5n/t+pPa5pskZWQ8Mqx9Q4ImNXbOH9JQ4xL+FRLA5/+nxeIc6WXRqetDnkkq7MeEwNfHQxEY2fqR+jHw5hjCj+jfJSjXHNn+8MUnqaQ8amfhMre0vXSeYaNlYzMYGPrTKGfy2zAsISVRR+8l+PQHe6xy29+578KfQOW82R3db0vAmuvaR00pM51rTd3L2qqWZ+2PH1QHzmjqI6TaA7yRlXsw4ncjJ38q2/YdgtQe8QMQraz8gh7JfME7PxRO9oHZLNNTP0KQQ9jNzsMvHYWjscTVp4TwrEQ+lAATzglZnH4t/pn9mawLxH6+m3mEkWz4SyzCVT5ZaezAdDjptTZPH5yVSlRfLe0fwX1SBxxGDd52Xxj7JprwpfqSDwlxvu/2AYfXyit1s3oyMyvCvnw2yAipMmqfUU9aB4JHmgeFuaC73AIh7nfq/+dbIHIjoDNmuG9QjOYmdSe7ZC8WdbZuew1RkD8Vnt4+uO2919ZejtKDn+PXR/0SDOD6bCyiw4e1DHy2bn55iAqaMyK6ug5UxffAgJ7L1i22sQRHrcUBy5TjqIhpsK5brTa/rvda8UfIeZW1V9Xk80TtU7kPQsV9TF3eyc/wHQRE1fLlN4/B0Jh76DJ8Nn56sWiA2xZkXrUAFvt6+ILRkySGpnKgq/l7jQVj4/s5dqBfTZxuWNdx3ktzT+MjPK7zpQyqNPqEBX3z6vW3UBjL4sCUwUJkF23gZcYYzTNo2AtIc/V2dp27pWNt/PEHcuRzX410tOTqdRttV3/qD0e+faBUDSg1b1z7h0q67bd+wDvFIRLeic8WVS5jRqsOn/e73IzOlWu5UGEqWzQHXBp4tKAVQS+emJpgF0oEM2/OFh3Kq0FEAhQun1IluoAs5bg73fIeZ0ePj6F9EttAhbARdKFi7Rekg5uXc5lMKIy+lpFTmv+R2CNVRftJg2jadb2oACxNl0j+Cr6D5gkJ3uc1ppiH4vkbd11/Oj5FyG0w0P046Z1EvL7MqtkD1e+qtiVPo5boySVtzIIKchQjVD3HsnEtYTjjHZK99aJqdljnKXL8+7bp4cA9tYyvhFuuA4AWV9y06c22jkDVXdONNfYKyQrxG2+YfGdIbt5qzquohSTmNZxX+/797HQVfQhRnfS+mQ0SB7y9SDZZt3/NnZr58hLVaVZIhAt4H+8WRwtpg0pcUJ8zedRKeqMcm87prG+bfvIiVuu0UOHlWG5cCwhoh4rz6hMTu5HNXee0xte59wu3WgdnpoRd5TLIC8fumzQuMw6KiiJAvY0CmUYKz7wIJ0hdq4jfJJMqaaYj6nd/BRKm4r8KrDbwNpBA5DAs60lHc9pGqYhh4bNY7BogPd1T/45UiByp+3TA2hWTnKOpXdefM5qmVBmqgtiH4CtEoUzgTybPAsySxXjk4EoXdGlZe4eDjiPWb8pB9xyEhvPFMmb1A3jE3fWt1EK1HIYx3eVc4Lmr+pA8SNVxtWhxE729esLgy40wai8qbtTgxDqFtqlQvZZ3DTWyfrrKGQb+2xOIazwt6JXGpB6553mhT8lsfRq4YeizZkq4uYyezqq9LUza+ELAUlgq8bBL7NNEI5bqqNb7DUJqxkqHYR3okVsBbe5fVUKV64SNT67HkCzX51dp4gZgANTAnN0z18nFzZ2EAp9SOVWUXJKfA7s0YAIlWEltB/YOFVNwtQq70zRz4WjPuLqdA9JpHgEoMfDcWEBkEwlQSgvr9ZOOLKpCxkofPXmAoQZC7/KvMfGIsmUooUdgIZlAxfbJTuCozYv4qNWeYbHpyWreEklmGbEAzg6RjD2dQTqVGQ5cDGPviijIrbp8xdm+BEVim23eXC+iW+5QtD4M1DGZB7djNM8aEq3hAEDm4eAmGMKuZ/XZSSEdWT9/YaHE4UFrSzRc4m/rolWPW+uwzWB2CxiBZWL8WM5gVjWtiIQ8pLi8IjpmqtowLt5/kSwxRamBDxLG2oADSzwSwyGDAYLE8/n1Q4vfHkYIA7gQiOsxWNVQwPquxchVquFnyPPeLD3RY24JeY3rU1kte+bCTD6Pf2FegHAyn+Puc7vaVEXZe1Ec8ILZFwqvfxNE1XbTlUB9bRywkE4hdcxO8V2HzSGXmJyqRP7fucg616DgxZc2X7ZEvXT0TaP/UwoUeEPwMyqstDMN/huMbV+N+INi215prTBTVeJ0ZjTqM2LekQXaLs8ZCnzU/+DV6rBOAV5TT8Gly1OY3eyN7yLPPpOmT5deq8XEku0Hp0GRyPKWk70UtpdDfwZ3ON3Okw/rcmio3pufhfE1TCdrcF4MNhgmKqJBp5zqGYu52NP+GxdYq1y/1uQ+Cku90lrDojdiUM/0Wb/1xSWRsRaxswUxA47UyLyKXdM0Lt6XzVHm3UkhhOQNYeE6jQaTPYXcdPQ6LAPCIBj4ghsDPRJi6Ip7/s1aJdaOBL5ywcgw85Bb8vB0CNi/iMFTMzcV65Fc1IjCoTV8269vo+4fheS1K4RBXshhPp5+XFsoePuC9fDp0zv5BnPHc9SdD0GvcTZKJCN+DJDFQmgyH8wF/8JXJgtb5C/o7HRVaPE9hko2IqypY7LwJl52VbXNmSiB1s7puY3IRrPqCZVwX2+4NvDR2w2Y0dQcRgY7lR5pK3Xsxfr/LUa4YX9tFvss+eOFuS5gfkGjP69Sn+AC0gVwke30KHON4STrv/v4CfGaZkLYq8sbvUwWjh3yHLAZwbTDwtnRQTS3WmFgGU7wyjaVbVtywDR9CgBe3inRZTB60FDuZcrLpfDIvtprPnKcj39jCUeJF+TtqBVD1IKzhizPpeeSF3ADwRSRtjyDb/UFGb7/2bSf5mRUosmfTXRJc7SoDifmqYiLoiVjXugIgrxD3QwjH241ERmxLqAzZ0FmnxjGmn+rxHHwy+R7PDYPW+kdZaFpSqdUMhs0KKl6LARK/i4jRxDZX+rE+JUGQRKaAgJxClpMrJN9Zg1k76hCgu9snup1Lg45rSwK/S35AQncHZQ5E76iRj+2dAn4VgasiO6Oq/iOBh4cFHUi/E+bCsiL6MUVfAw6pAgvdkUVQ9b+0/g1LmeOhB7VVDQ2xGicAA+lKIdhWSeIpDlM4riS+sFY2NHYE2PzWgyhHKoTJ7HtN+g7FuFtxjIA5kefWiUJBGSDia5Lz3QZjtC8jY2lHRtRt7Ur9V+3hqDHq/se5Pw5TPReRoMkiQ/N6eVLDu16+g9Nu1IvoJG8WR1b2w9kBrn91W2r2sLPNbqhO26WCNMv4JfK2/+Lxh9mkHChQ5BJ2P3PHZtFfUsWHi9lQ2/tvgozjyoJAv2DYxxtUM3KNS2aFhD0agSn5hGkYoAFuAKIrOIOOQNCSx33kSncAoxFMKPWD0mUL2h/L9bV7rLRJlIKqM/xxx3VGZhwyxb7nR2fxAoB1ECFW981vMFpQv9+1DYVfoX47gKI3Qlmrcx6hLpuBLqG4hvl49nNTbao6ivcdSuYTYm9oNRxjJiqpXOctWupGwVMR39J/iWEv8DJCbQVkS/Nqww6UZeVN3MAmnOlPKhf8zBybFck29KoKB5AU90NPf0xU+RoViZoKkg7yoevcf6zEw4QgXg0GLgmU6LhfwuXqhhl3+FpqC+qYeim5T9qVCCAsktzQGSSCmVBuJ6YTOJmLsJoeKZL/YiVAHuGaNELqJxHAgMRauP9f8enq84fcSAkdRT3y49pQr55OVgDSIxFdxICXw7J9bP+V0Aqk0xCcb6yEZPWQqEjG+cTV/XCNXSmXVjImWZ/h4MWBdBlL4fQu2cKYcwhwY+T1WG0ON7CvFT0KjaSlPzZy9uietFdzdLT6GSq692leiftmHrwXWZb2S0P+yQ/QrLK7MMbKKNEccDU1FtFsIP0MAa3adSsEZYWFiuKsRhn9fqrQHTW3svI5kga+ajUVASg3mEMnaKJ9+GAvWfakW80GSqsZDg8RvwYFtgwFcvguVKSUimI2qmzovbxdxsPvtrLwSz9vnUYBjWKiQicC8bhK2qgx8AJ/KgPNNJ9y4P1o9Zs0AIBRSA5f3Xb4GtMmbA6nI+18pk7oJ0v7hJqsZVWr5OdYSZkGKGonUH6tf6KDT4E7sz+9QhII2+sjLCixJdU1TihLoSeNHppUNVFidIsLOG/He/XAtoY9+UTGZwZRwhApMlXDBYwn4PAbwv+O8NtN01yKPPtnaekCoNk8BZUCfVNO2gYnno257ootk3D83BxGzalz14TX2bB2fWUJLcvc5Hz3vh9EFGYlwWYfT+req+uzqBZxnd4PmoCLz6i5mp9ywmamVcmBvCBIqDmxWe5ttZ/JrlKrD9dw9ILR/8gXFFJfP4w1MbUMQG0rocWjZ26nBrTuZmQfQTIZtNFmgXm7be/wwg/b+D26WI1IuB/UJjxRi4fMbdLXPHusJQeg/nx18fGlfCCPIvZhkbGF1r8srvZ7CFhiZNpvnFev6kwp9d/Mky8MisMQ1nHyVo5/ex/o0zcreeBLT9O2YiY/dbMJhhtPEBowPVzLUqEk00AeWOZ1Tbb+DXdpKl5ucB6sSKJ+sZgSv4/pCzFyUKS2/syQJlDzV+jgbdOgktkeOhAph5c6B8nfjk6JGJAzP2KF1yYFWm2nXrWXF27bOVTimPYgpLjodfoQfJTTIgeJi2rFPpw+NOwiscnj6T1xn+TI0+pSNPDQO4Lnf7/Fg4f8OS89QwIPObHIjy44RCuygw+Bte2UN8RMzYKDqrq6NlESoBvKqqJOFroXHTUsDKT+t26R4VWei+FPt4bcPHtwfL3RfyRNzu6O9IG1SI186f0Y+qouLN+amzm61vZ2rjQ9omMkmg8/5vjxbylgwaRA2dOdfaOJB1j8twQexBRBWzTAMZAe6+OHMCbrnoX5Gl9XPxheWRkG6RSuYtVLoJL5emd7M6Ryw//VklY+9908oYkFZMIV1Fb/drROfA1kPdToKJyIh/X5pWgPQ0vLFzyz4JhHC7SXDM9VG6AykkpYoJeB/P+T7/rkZ6+KZ2iTlS3O392chPwtoRelTwjSbxQrP0DalGz/ZQKWGTXSkNKPQjM70M8Q47kjIkNdCiMChhEVYoHTtclcUN8P6YN0oP4iftb10SyHmhwZ3SWYgnl4dbyrgezSi2+h5ei/+oFTN+sF9GvprwP7ZhmCEjfctVzv3hzAj9cgbgVva4gGU54a/P3ZG1e8A+5I4/RBqP/wr6bT9CexspT2hlTkQ3wJpCNZOFyLc/DGdqsPNJ7MGUtLCKeCi72ibQzYNZwYYx2WLwy/8QlAAd7qsA8EVRZwaysvRjOBglsm8PcIQjT0AHOgKajnnL+szg/5UY47yp7pjudMzKxnmh8Auak8uI1kSCnKDyTk53qf9dG1yfK3SXzCv8HNApSNHanbnRcszr0BzWGZmger5QXtHnG+pVKcg6n/XDur96zhdPE6YTMglFD6BNvzZpKBxTRTJU62wakS8rvmE38aTYr/x5PvSM5GKJ3YclSmGovHnGATWUx/O4Z485WglEEjVcwh6D+mVvoNtW2FZ1HYUI/dX7SjRk4WOL7TBav3EC9NEl/tA2u7SOLc+a1bNEixTuTLNs39MhhhE+jd1pOSuaP2DSu9T7Vla761dtAKe4hFvEK8POdbkiB3EkPwKmgr/j1O2JONM+BsyVkjOMNa0afzT0a3Vu2M1DSiloS5ji01991x7phnHeru6tu0SXzqRdMDoSwVtDB8+0dCza7gWMBTIOCJWklEe3Rzui4o3QK/Pk8tBJelNvHHKEo7D8Z+fYyentNqJ8YlP0aH7MRvhrQ0XBaxAD/Jy+kCrUirjJizJhL4HaUZWb8v/dwArk4T9r44B9vNTos7DY44DS69C++6usdnXGEkHyrN4XlDntkso294PqMZ72cGxNG2Mfq7FGSqTCeh+ek0xYipl0nJIHkC5jJ9jIARH4DWwOF/2q64VU076N76x9XnjFYopf8HaatZBkWuMM3lCVhVx7JKcjAtH/csKqnMADywaSqfh/+/LUY3cPntHgidnZ+Jus4+Uo7LIwKa8Ax6FWWW61myUF8jXbOteOUb66o+L5pjt+m0YY+XbtdJGS9rKNL6LgySVR/iCElO0j8btwrTBvC/26YL45eQXhdNmyq9j+UU8LoI1Oza4gDxjr3r5fWjWXKdhLZGRCRmpSQprzimnnVpQdEN7czGxApmXlS11m6isDfiEzf1m/eAoXzAjl3+a/qEla0RfVasP6035C/WjFegriHAfJGhHJtCbxW/8ostoQ14sH92nZggx3X3hvE6f1VxerLt5OUYxNhziZSdlPi31SFs9MUXFSTJJuz/CXQ+xvtzQEh2mrA3jhe0j8kZB50rqLtmVmidj1WOjbRVlLdhyn5jhg8uMp72ijkC66JiaEkvyTmLx039yzAJPUhVvVfr5m1K/4JeYCGM4YJ7gELwUFXqIVhZGLwG/VKw/Ly2KNMt3k0xEAN5tK/jE3DXVoveJ0vqQHmoe0UAYSqyZne/9+viqGxvxRWAxxfBG860HQXeIPyupfWyOLJBb+yPh3Smsl/wEtaZmwe8QYYJKNqcdP3JergPrXpuFrg6IZVNwPXnW1SqXyDo/2rJgMGE1CJi37Mav1hymafE+1hRh2bgtP4J8tklwx5YXAZsjd48KEUcmVyGIbQSY1eygcYr1Vy/IblKkpEmj315MS03Kc410DkJ8DTU3VLRqmqI7QozwRgtXhpoqBdsuYsAFwNTTnvnX/FtuSLRiE8rjuvII52lP+timYjZUEqmW6woSbfw7PNEHH5yBcc7rZLQDG3FQH9LaSrNmg5VFn1NdWoOexFNYyPd0LIFtmT9BfUHrxxVj2B/GC93rw+eOtfrqXasUIVu1TIRvgvxV6UYkykK8KpstTKvCXkf6vxktSWOcMg+JnCwx+mePD2M6xmuDAMbnQujyfeLZlz5bwxSDaeY/a72cRVPTQ8bzf8wy8nPYD8XYyI4nPZXD4HI08pfnr2J4a7osny6msX1FBIB28tzmygtuRgVg0lsCzbhakLLRAIOzt9EpqbBYfkCwbd5hgcqJeUmb6WmJ3ed13SjdBjNEpA7EH7lEEzxvmrhL8gXTmZGG3mi18DKU/TcmSkuuWVxK1EvBOlMc/z/vphNzBkUMhv5XTtw5lj6vjbPDvxwUB7RHYxVWeKSP4i95ObAJxPgv9YlOiQbtV+iEeCUWvtGUIE8DfyQadMHZX2JOuqrs1GnPu1Dm66p8Fo4qonb65Z8y35Xe558+i5PjWIX8qJJyIBu8FX+qio=
`pragma protect end_data_block
`pragma protect digest_block
b5c73fa781fdfd5903892ea55241c773ba93221e51cfd76c6c920665b3770f65
`pragma protect end_digest_block
`pragma protect end_protected
