`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
LMXN6bJ6anCDaYtn1CIO4pqVbcnMOs/yzien4heVz4TRGfa2g8zwBVGoHGYDmgsjPbfG6V+r8yDWVGxczFLxTSqQf8meejzJ4eMHLfZCwROkXNTwSLZcQg9bF6oLbn6qQ8NBCELTQ8f8v+RBwwDKxotRZACO6VWdfPVns8W7fCyQz9wyNq+6uBzxrjoR3JCtDNyABAJt7BLeZzgMt9g5bV/938/eRMjEUOlHFm+DxtugZmhV2yXDQRvG0asVIco8awvknVvcx1QIHXsBaS4+8rwXc/FVf+TGkfsaMzcKXuUGIuIuDj2yIYr3r47m+bttiO8Px4CY+p2zfJwxW1d9GqMTS2naYMGVjkSI9DP4SSVwuR1lOJ0dB9rgBknfFUtUDByPmRlzf3F2OR+iYr3hM74pN4OJpYXfjQczlzAO5Zdof1ToXwcjCqDVY90wrAuBE4VXioM8R1SozPtpg0dDeNO6a4/1IJ78kk8+9unCvajFyac5sCCMfCQRJX1Bb75WKaHBXNuGhO6XHvRQy5IDpyfgBc9FhbliR21qe0Pe1KuB33fZgLGNEBW6QydcmU65l8f3k3pZkPlCUeuKL7BD1qsFR/C0P1o78L6tyqATJfkI35GuvUBt+AUmyGhU0HjX97r4C/GvR1I8TrxzgcEQVhwhHUnzEeegr7HMrIb4DzdMAHrYvF4cPllzzDqTrb3DA+ux/97OvOsf81l7yp1DEmQp1IOviAz1qc1rJr2KEtsH0B7eQhR4HHrPXzjPDLGtMvt56cNcjhnrGuF5qGmUKhViy167aMdhGNyAVlqD4dqOhF0D9SLo07Fr08NTqU9BvKrdQ7M+0dqkF/XMQLyGBff49DWDRZ2DQzchIEfNQpfgSPploweDczZYGhwzg1csNZ8tazEDWzacJlFQh4JbkPkyLXbmQB7+mUolGumalJiPoC01ZeHaTdVqN1L17tv+7GwT68Q4GSyeCD5wkOJMF+Kdq06sw9rNi4ZleaOJ+jGww1Q06yt/cD0iGa9vji7UAGkgGUtTnNd6S+Mza3DZXQd/n+N6v2yKDqrNwgED0kODcLFN5oCoQubRaWSW8+lbLJP5u0zZKogoFpOv6LW9MljvZ7FItv7uvva0g8d6kOZlEqfv46bMqp+XmphV24iCzHgx2VZd9ujE3AP3CTstV6s2zez6xyo/NKsM29VgxWFuRGwNFOyhKqOsKwfJkf0V332mzAtVQAFzYtqQYG5oI5Go8ThjkyMMJgaPdFQQB7m4kAZtymjUTr5cJ50o3GRniKip3XVqOa6yMs+Z6psbVhuai/798vITV5R0+uaawswUAyZSeLr4tJ6HaZ7GRnL0OONiHYL9pQX0///dVL8oa3dWcPxb5EQyePYQtTVEgH46gVfnqMJc0bJLWfzwNscQFhlW6FNEBJEkoEvd0aCQ7IBfz0Gsl3ZPnp/yQaQpLqJIpTlqxgZeIyGs8d7Q6UxvDxasQdlOkSpgzganI1eqkUB+hP++XCObaeDo6EqeqosxTGjvkfSW+CXfdLUqp7Zyr7X+HJlteu8+JC6Vfy16i0uwpnIVSO92Ts+u6zZuaGYEuDcBJn/vT3VCKlkTaYxWF8aFfprWlXopwslNFR2oK0HlJGuPvgyvu1B/eFpqe6+MBIjQvlfYyaqX+Shha7OvOoi/JMMT2+lRwAI4/LrSmznK/5FyC1iNd+rqgSPMGC0R0fLVfnumtfBa9iWWFmGlCeIAvYOGhkpywZRj4tjMAY3TVpQekY64ehB/LBP7tbH4DMgP/F1RvjJF6+72GlEA1qfpNCdVFhDrDywzUZVK3OqTOcq77P3s98n7TLsSOWQBw5G2yQKnY5iTnYpC701e8CypDgd0qevLP4JY+f/AOEA5ISZVrzhjlTP+6w2gJfZx4p6QeMlE2QOOdkWDTkQQC2UrGjbyVP5FWrEfHbDoJQ1J3spMIsLQGc27NhPD2R0yQTzL1H6Y8gbAsiB3WnwAsJgS3OE4Wr4XNm0LdzeXQ4x0Tf7eJ7higbIxjEIj/f8fcFgnZDr+5t+uSDS4jE8KSPAE67wRXJ2jgcWQuCxkkVjwerPaBzmNBjsPlHB/GeaY481bbXP56eyGDi5akTYg3SAmkguZF1ArURqZDoNQt6dSwwJ0vKoT1Wc8KdvtPcmsIPTHb7UVOXQsr8xO4cP1YEO7nphQNhPMOdSHvRK6DR8WuRSS5Ltkk/PK1+ERme3W0Z8YR9UQjnXhACfxGm+5uEpg5fcKfNgOnVTfXTmNZiNfnMrBiG4lxlmfdgWsdyqqLpLFebu/EcWdEPJnlwURNF1WO+DQe4NeUC3s93gIG0evZmIhIa1mmnfOhoE32QJPo3c9CieszHTrk1qpT4vfb0SOad1YGkCD38/sAwPmck9HrV2WIoHg3Lv4mbSz9YV5vYSWdCL35B+96ZI2PE6+GXvfF7kWxFnpXDIFUt7nADLyAqj1+NFJcUS1+ZFJ7V3z9OdoEuaSY34VZ7xwVOVMP2QcBdAiRPs118YX7iGB/BUStW7xTQS7PLn3aamVuedgNljruPJcJAfJpMomD3KhUnPZ4JLjI5FVogRxZiEe56SJlfxeGnJFaam8vllEcWu5m4iRbKeD8ZCdqbIWK2KaJqoPtLrRLHFMyPpZN4iFNN7Zwfb2ePIRUYFYXv5ydXhaDuCiRiz5nuBgtYmgK09MVva3CWZlQsc1qoRyNAJf7uS0+MTLpCPziSNYAGpKTrzwNxW2EXtf1QpBYSZ3aePPQepUx8EMK639YiH7aK0hKIgF8s94DVtmIXoT9U/vY3OaWqu34rk+b4AANZHv9WG04A/B04aiYORZmF0mWIC/BIcDRyCw/SPx1TvetS0Q80Oy+uN/b/+Qb03LxWAkScZzA+8XUqvzyqbGlZ1RblyezjgvYQ+wJynVUwGtUoaKVqzWDFnno/KRbaAVhb7Jtkh6BpsZcjmslKrLTjM3mjG1oyiy93bHHZ0v4NlcdvnX7nlptfA+D3QM2Jof6biAzi15N66aq5a30JmGAM0WGgbVC7odTpsW/ddZvZm9IyCuO5styo9N50+gU0dSPzJsfJzew25bKla8ZVy4iDlfJqPtm+YK/L1R7WgUUUOpmGoRldiLWjxbCI7hw9h3oz9NKKctGxzltl/kqlbQTbz5/pIHxTEuWjCUh2dkw82ofi2BP4aVKvDIhy3iqEnmUW8bA96U86Xz4XhIv55MBVyv50R72hsO1IQphWkMCls/UkOQ/CNZNgyVh0Z9CO/Jg9fVBz0LeNR1K22EKaH8o68N1nADSmg5361CwVv6aRG3hljbAClTzXD4mT/3dtSpWL4DihY4Fr0/bZyj9POPoZWCVI2iIt/7Rg+KolkIWbzs2cpkex4aoQkU9vZczHcEzMJNzC6l/T7RcNYa+y0+6pWTA7eHXtJ52RuarsB8fKfN7GWlwiHMQgJa9D2MjDywCiCD94ArNPMenaeJ1aAkEoaQ7RqLqTMD5nLgUq228tBaYeD4S2Y=
`pragma protect end_data_block
`pragma protect digest_block
e1aa09d7ce3cae265a07e283d19eb8c49c5cb8e54090d3ec3738ed515cb894e7
`pragma protect end_digest_block
`pragma protect end_protected
