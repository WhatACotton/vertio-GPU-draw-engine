`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
ssDjNbRBAT+K2mHJqoWznUC9b0cEmaNfaMrVETL4qtBRAruSNyttOIYMMA8+1RnzVN61AmHhrQTwfC2p3T1W0Lai4XnDZJJNKu5CnP9+LEH2f87gvK7FB+AnCzMZw16F+xsslKT3uC7tAkMwNqASTkwVl1caqXA11LmU+bTBcsR82RB9xh0x4KRKZm5S+9mUZBmLMdmW2dPVZcKiTE6AJYfJJ7awFJFlOdZmHvNNv9wVtpYODGWAuvuqUaabFFE0jS/4Zgwg46MTQUqSwqSG+7dAXQdQlh+sz9Pewg3Yj4JkthZ6aAfrkVIvVBEh3I+KUuUeGUReDv8kVLwaYnivDloSj5jwEr822vNgu+NVOqedBnsm0XBTkL3py06EtJarQl5XdpkQxClWWg5SSuVTHPViEKq4V1Qg2DimpF5SUowedJRqOSgHiSCWgbtnWzVnnqIVCb+nZAR1xLwIkwlzIi9bun3MplVnbXVzwE4h19Yk5qCSj5q/MN+GaUaKqjv4qMdXkxR/w3FjoXNZslHzG42YrrPpuAH+s/Oe/dIq/XOFID9jYkkTngUqXwivOxoj6YG/0AbP31vaqXJAO5qZmnAusH0aWRnpM44rW/+rnNfpMjcb/nE808QukrZXT21R5qxVEAch4CoqEMGdpvv0aCeIOHCLFS7y6InANb/hm1a6GlzVWTscCnaVhxtfnhOVYLbDXyuPSHYof2E3ZGssY0dxiqs/ef3e2lzOtudQaHCdPEiYnzk/KZU7tKut0/M9bkRVYnBVXKXLju7RbBecBSyac12aqRzCaQu+FBBaJabKcN+qCt4qCF28yTgkvXANfKjB/p3Nxngwj51EolvTf/NSxWzj55/YZgWDbaMHT+hYeMA8DTlO+huPseQ5LpFDfkS24Bf8MiRrFQ4lLXnhmDo29ZyoWpc51apbgD4hyj/c5nrkqpoc1LODcQl1cPffB91yj/NABZ8+VAwVY6d6VwDea0YJSjzlW4Aach3MFykPvfmq+q1ChrIV0fmq0jQgH9Uu8NnvagqTpbiTBmOkDzdQoLcGgpVDgOTBF+wVUsqJJNhiUe2nf4yRoGXJgwVT62lfdVNv3QOM47V/tz41A6jeuDulQ4fD2eleQKAgnoo+BSOhKTAhVZpOwlU5vZmR6pA/Z+Ad59tHEVCOY0DNTUrfVAcsnPDj+FBKbnO8BxBZeZw/fDMKiQwwvDvalQHAYbBfEPyqWZuWGGGwfyDyeJEnt/xXgfaV1H6pCF9Gbnu3mh20hrB+yoGpuHRmgYSFStHVWa3f5O/5dNvM1z9TmzwitxOVrtEGwiqyC2a2k2a/u/XVkmhhhZu5VDHAwVWLvyt+80dZrERvOb5C1yZGjguxw4oSOnL7YjNFpE2rgI8A1UlG4/2FQU+/BZvXKPnDbXOcRptQO8XX2+KGoWB1dVbzueVbRTticb36kzsy70qMzeBXmgOlB8opK0KaPX8X6IJgMxTmZ7aHc7v13P0EKbmK1XXbg/9CRXPLFcRo9hIQeg3pKWOzuO2Em12iQRlKMsSSXC8nDmaPI0sgeyHEyhI3Wpxvq4m/kUPfXWZz9S2RRhd3UKuJLCYwJub603FdbV7aOqJtsUS9A3D+o5R/HDC+KAj1sI8S4WYlSTYfYoO2Jc3ZbhoWCEJvgsZ3t7k9imPKV1tLjnV/Gi1JLjnfmHUkHRwcWkzDXtwHSx8CsRRbwowtzpzSl22oD6KUGvM7IWohW75veFdIfCFQOrQuuu3HwEp/FkccuCuy5+6Yz0LqrUf+SPxWIFbIsprPhZll+E01+wZoKnaJnE/t6ezXoiH7S6sEQiT6oJi+1wz4/V1ge8lByMdBzwQO+fZ0JUcK+FLrxH+q46eXg0RjB2EnlBToD3Vn4EjE9tIr2vTJrbDdq8gefJDHw3XQUCRjlzS0j9W6AKnhtqQJiaYyrMEiOMRhsGz+FWTKnnnBDhhm/gEKglUqxNUDetNnohu7OB4HQ02WXaIVLA4pysliws30nEt3Mcjzyhl6ZiGG2QSGbEJWxpKNFrt59GJsQCAZTzvttNhn9LQ4PQ/VAU04aIngwazUDjFxnIYTkhVoUzgvCoMmqvVi41I3AGZekS8XkNC4kgll9W0zssFfRG3ubeaDbBtWtaB3WYLwXhbvpb+a++O8JuU10w/KmhljB3yapl60o4adjXUFPJPG9s3qBcnYpDfb3743J4fjPidy5tqNIfS/UYMPnSyWZvCDRf7081+OCJfgGRe1m4BcQY9+Ozr4HGH7BrLeYKU9+3GswmcClE2EVaVKsIrGBBGAl++7OYi3uXECOT6v6CGD88vYF6JXyaVkgKe+6W0VcDvvekRmcBx3A/UPsibAl5gfgo6bEAGbx+VdyxH7EyHZt7iumkJoRjuAVwjN+uWnM+CrdyQkdKwC606tYjHuVbfOfqlqXcDQ7ckVr2alzTmKHcl5ShPE2KUv6rm2qXebfl4JEaVZ4i/tCFQuEbEaLFMsKdQ+jLLXVkInLOuZvGCFGpHtCSe6FzsByOvFXEHHb49Jclfb7DsbvKNKC+3tHFTmbj8KwSjqsfF/Z2GtEnELKKnBMzt7ntZVS3ApON06pfnuMC6aLJM320qQLhYz5G0FU6+lshvcnvmb+ba8z9Ib3pEW3DmzIYbsiJq5TMCsPeZFn6FFsGsdgSgDPw7+/grUK9M2bNbGNzbXBLUJN/WQ6SlnTwAAdDq/ZX7ZO39dk1tn2sIuyLRyrqQwq5BDNx+ZZiRrb0/ibSjvfNcmYbYlX5UpKIerz9FMxhB7W8w1UqM7IP5Sz5UscbZmPiXR8/RXIFoPe9qOsYNrqXIe5HT0499TPpL13kjReUb4twJQ3d1HJs9XIdL0J8Qasr8w4YrODjlm+vesFQC8j1WD9w7ca4Pf6SN0wCWalFWgtAI3XC5+GravQuyBnm+oQSgU8DduByOCre9jDv4/eszidpUl/m5FViPASY04MYjgxUw51ljdCoE9sbWPYj7CCp/m9KCYheLVLrmSmX4qTWuRLVX8Xgr4HDHvkjBCWnUKe7fW144Soeqcg3MzHaP5HVcuw8ENMjmpBOG6ww1t5u7sgRpqC4KsGdm7AjJhMz8/MhElkgEznYt8cXX8BQJE+MaKonydTg/JN8m1jguFqbVDyUi7u2nvm4jGavbo+X0QsvsRGFlVQ4a5H+FOWOwDXHK3GnGGhNLBFd4HMEtH4aSlOmL3PaLcKFFsiETHEO8DFKpRCg510HLUXlG/e+bcB79QAFyQJPbnxjtE2DOkhA8Xv60uCXzHh8P3rDm2ArtQy9VdQfEKcgGxDa1/cyr/fSb4WDghS55CmJEOkN1N4sMYO618ABO6JZ8OdISmTUzcEEf0/UxfoHqKu0Ry+AxURK1gpcXc/nOIqLO6augnHSSimPY1ZM1IJukUWDlZlat8Uf2UWo7+2dwfUdZ2hxqDy06cOZ5a7kuJz3XyNLuUpy8XxBpna11zfxPZCfG/8xniOxihuOoEXmsLpIIiRyLhMdiBhhaSA8AIPFSnxaihMFbEfVgFZIcV8fhbGjxZtj32Y1nZwDFLr1libUTnh7V1yLOgqz34xbSQw220YXd5xPH+cpqkXT8fT0asFgPzXREVhyBNiz0Gf7Xja0Uh19zwiQkPm3sBihGzwUN4VirxS3P1N9qf8er1mW41sGH/VcfagB54uHYcDiExUGKfL1lp8UwGtrC8re3r1C86kmcEd8KuHQaJAX62hZjLmbRs9P1S77Uywl0edE22AcfBPMU/nLDNAYv5UwjkU4p8J0hVRHvHYoFORC0S2JvHc1eiJA5LjoPGcp2Whx+lhZ+fl4fYp4sPPdLCYDIII4efZwEknX+MJRBguMH9dAG6sOLmrfayKXq8ZnwJwFMqz16RMjUUMEinf4QZUpnfZzHCihar5W0+Z6YBiByoXkGYUIOUx6PbjCo8s7NRHmcBsOVDkwdqfOi5sCbAU61G/lLbWdxdTHqfAuJ1cHCkCzvwH3FOSQ01b37HBntVHtFAO0KJ3EMmwIA2CzLfzkFLjRHQsEydNJrFGbaAuP47LoCD8qyjIQ1puOcewgVHlYtYaamphFccaQxizb9TOd91OxnyjGl3EqYgubTG/rRBgmon9f2HXcgTfytEQPOHngrpJsy99GTbfY3To/kdXXj6AcSKq0uZB4V43yxNmSajCAyLorlwzc822IkfZp9e43Y8NO3ZEoSJX1R5Vcb0+Hg/1lYoW8/0Hh1mCCQVegZy5TTIIIr+Wc4IOYGz1ENLQhAERMZU+ON0VpIM4BntYgfIsB/hAMdHjwbD8Njbpbr6LLf/MFfNDjue7vYezGm830WHpQS8R/HAu20GbohrBQ/ce8LUNKAk78wKdgcqJIoCzwEIPJ7eJUSatOYmgNtsXhidy0nUaATTUBgq5s3wOBmbPjmnze/GC6hE3LqyGvfzer2QLc4MuIiVSPMpSNwAk45+gCyl1tty4b0JmGTrMApLiis2FvgbcRqpmOhPhpcUcY1lNP8aco81VW4gvvX4UXyG7VaI6rbgaAH4+ckpcD9G6yLDJXhcjdaMQea7rCpLLTuhuIXwrttjRea9Tsek9crbY3E8/ZHpHrtv4WngYUnn0zXR3PBZMqoxqA+9BGowFxA3Lg3f/MgsCWc88guz2PvaTIilVT9Hwhsh7Vnlo6al1aJv+JkvqneX/7WhnH/rY5tfcv4jG8y7GgQKwKU28DGi0hLr90hkxcRIGw5QMAqKeVa1oQkvLA2nhiHGfJIkIKNsDl9FRt2ykSRqlLQPDNHso+1sBN09MlhVVz/rSovrAVtHsCNA7yf/Rg1P76vU99lOpBvN4jh2TUxKzjxCEFSAHSnekk7MN04TiOOJg7af6B7M8zNfkN3jOC2UDtsr/Q30j0Md/QGuvjuNFxbJ0h62OWoEBBSLpIxF0PziA5VHEbSSTjbTI8FFrGHioJBUJ8nnVqEjZam0+gPZu3g0FRDCMTKWxJ2mUI8zeN31hUgMgIS+pcB3uGhs05AUGc5AyR2B4Di5yeK+GghcS1cCjDXMnE0tMWVH3LQApPAIgGm4iWWCoUYtp+JeFxz07b4GrAmr2dzvEyrIIGktPcZ68JR0GWwlZawMFxOIopxw2+ITcsIVRPVNggAXXxPiaGTWTVjxFsl0JXx8A7Yp236Arzxt4QSkQIq/dFFK1OTLpQm8GALEpu4tdKySIfFnm9pVqDuxgiCd+aC/TXee7qykItLPaKZDRBT2LQYIjjRtNkSgrEXDcPvQrUkpBVXr197zc5mN7sshnwAjgjkqMIX/FewCDqECPCihLhYyoQ3uLEoAYsqfH74XBACA52mF5JKIR2EwDX8D4VhC8+7avb0GVMGk/epGumYiM6lgPmySBVxMgm1VnXFnr9JLItcWA6R3JecNZwg5hhJLlhhc2t2Zpf+sl7Xi+os0qNaf9JCCN0cWsLs0flTwg16NEGRJGIgHXmpslsoRxI2RyM7TF0eROH7Qo07s2Ipip9J+1MYQ177ejqdFJOhTbuAiPLUuUz9F+YRDqZ/8oD6rGi1rJc7/g3LPYR8j87yYT/mibhKSdNGdcsr5gztwN34PpYCGd/RCFFm2Ubx4IGToOR1K3OdikR+kUrxx6L0j+8TZhuBpa1i/jYC/vmTQoWt7iA0Aspovpe4IWH4HzEmdru5x64MCptrOyCVvGg8sofDPvrz/MB+8ZEhwJO0GbCkwU3C4R+GQ0q0g580RsH2HNtJuCI4w6x+ygqny4VGPMHTW6EqFHXnJYSfwRpag4aM/ASV8stpogrxPIZQhTYdNWQWlT3XqgBWqvdRfphYPxJFS3RD/kUUNZigMty37+m/okS9Fh4ZhdRG7GolWmN4a8GVKXFZvHcvlqp7H/zdkQJsbDzqJUxnNqS8rapMeDr3pwS7qx7r04emTVSZc4FYtdlgL/veM1TpOpazuW2xQCML2bqK7sq/+AFABEex/gmmPC4JX8TLdC2QwB8ZZnugXc9+yxNssbVta/zG5qli+6RApQLDokyhcx8hF+GihreMNJaL/IjSAvSyIhFouCt/ozwB44pusWaQhsh+BUc7xojGMGMR9mv8zWxc4bB9nTKfekJcncK9XKtDs4K+9SobDoh2BbhNyzvWmXYCg9pmfwYuFv3MqXZtkj8yeukQ/4QKYacXNu9MnlIzu0tdkmYa96CLNyc9CmhZ/1Fd078E7s9mkLgslmAt1NSuALuIY5M8k2pBVnWHMimimEmW+vYHdSrIxsSD3b6rOGnvplRsTiTUifOMXTwcTQxgdawIyq4P+KcRX4v3GykfLdRHhk2fJ3VwMKwdM6fHYEZnhlStaQu9I7gVOfz7s7mMyDIAyuPfLXiGV1l4nv77QnkPQbrHhoYSrUoOwGQW50zso2S3Lp9lg8jkN5pTqjQy8jgSZI3glmLhG8EWA58BbWf4xL+fyxFN9DMQtb8oKKKBERxDf+JojXvtcgFXaiBdHFHJo5JsDLDVRn5+pI8uDGXd6qlDexFaZIleXmomACwrp8pxrZ/gpf9FzK2YY4VZ3NZycnTwZeKHxwKdROaN0Ckpx/zOt5vLrF9dKC3cPcjsY9CgvBHrapoWpnyJmBszUgS/a8/SvSEzTyZDekSvcGG4xrlhf3kAybwbuu/COJnETjPUBAJfQizWnuT6ILBvr/f1mJsr56ha9Z+6cI5Rf+buLQCycrEbdn9Md1jRli2vekWIwCUkfvKCiXGvaVbbVVCSh6fhLgmn7gBHCNuYNXJkATNdbd+TKhKu+p5L8fZPNZ82yZyRmcbhXs5xjt/GlwzczacE9WI2JZkudqoN4RE3mHGEEp7EDA5w8y6D3rX/6Z5ib0tdutMrRSipmWhZ3YqYdi6z5kCEldIFFrhISArpbPXyRY3ug8WQKjtFEwPMvumsdCEZOp6NJDh3+td4U0Ep3mHPdB/V1bH8uAEUaarfQb6P8Y8BwSzpMua+IKQFbmSzUABrK/YpjRfTTkejTlkt+VeS5xMnYQ+Ce4Mb7e2dfchXm7OPGC3UfaOY1FleiMRfn4j0oF7GofF0zxTf3WNq1FjbuKdblsNryBlQ3NApkcJ5E9ByFbU9+CpUIiiAP4jmv3co/hCfN6j4tznu9l10Xy9K+fE+rGesxshamR01B1wAvpMNT4cGVOn11m+/ZUDDswnItpGbmReVwM8KktVHnC1I8prfE2OrBTHTEMn4tccm0Yb3gOTBfCEfUNwXvTfYXEcHweaBoyKF/uc692pHUp6JWDFQRxswXoN8nnRcc7EYH3EOBavT29+Nu26Cd9mEKZZaTEuQzo69MFLI46A0AtVBo10wvzAAhsgDIexSfUIjzLxB64XgON0cy8eTC9fty7SemD2gIJ680WR5tFn8VYSRTsUs9tlfzWBYpQNiu5y5q3I+ZN2qr6BIkgPf/dnsZs4fEKF2rMd6o2szhoLDP999LxmQ1WBHcs6xVF479cUigl2TpqBNbXRro8zoR7sRjSf7YWfLHDBflyOeNeKPM6S4licaz55e6zFPUqBNdTHVw1kma3nD8GLA3x0QivZLhqwcXA5zsg4ykJJEK+xhsnBcww2u7ZijfR6UTue+Cxn0RaXlDud75VW7TABgOXPux/ZWNE+w0Zo+yOBV2/xXD8ttq8dakGjPR+UJOUClzk4qelEihzOmBnHwu5CAh1vhXBYlXpYZOdXRyq272Nz3aILvKhq3FCoukW9i/tIAUl2KTxtBSWXYPn3L+9QQAzWxF41EXKo7k9rusO0VJkflZEyL04czCKRtNWvbbJYZe9YjtT9W+k7KAR/GJeXxNBj4UWJ/FsM5MVxngTazOd3x0pU13RpNTfm9ZbJ10UJa/d8Uhnb1cqa728O++tMq0cChsN5vyfkjWiObYLQFW6vLWDhaaNnyAUTzfLdNjxLEWLBRlF3FvJlhszFZR2ClKc80hI+16ZafPygE7xitgseAm4/TjFpturnQ4/b7ooa9/ptjlbeNNkD5V+bO6WLaWf+yiFN6Di5lsZw0jV5+DQ8tWlmq4j23j+9tivtsydAh2Ra+dlgpdrZV84mb1mNawOr07g/8ocikl/oAZJTTzySFpUUjljRZaNUQ+e+0aOi837BkTCTrboNPYwOMVkY1PDREUjfowwjDwx3wMtjU/ZNlXYcQpsYG4XoqEDs2B81RzVuQMQE6cvOqD3SZ4A6rH5piEr15gdFi+UJ6R8wgqVXX5EfU3hLxKHz91bYifj8hVm7umBK3eyBnVLgpxsYF95ytLeWypSb4zkRH1aTfY9WlBPIF8WbukrCHmcxNdTfqjpP+sVIefTIbX4nUNIBQqI7lfw2lfpxT95L1pPGUDiny5AGEBjuEyaRNsG8VWVn5h3ozdujSLlG0tcBXb7DhlN8UEOHwH7ZuvmhSs+YK2RKFfWrzYit5Bqy+/Ek7VX+91U6/NtMmy89V0fC/8zfKmAMcsbaZGjooilO9QctxWgy0iI2K/r1qC43LMeU2OYxV4vDLdW98FDtRiNZiiki6sugqifBnaDkYSdiG1eOpRxYTcLLjIiEoQbQyjI5saaq6UNUq+0RAlhyEU6yDLubVyVPe9nlonpN5g5B0NSmfl0oSn+Ipum+N7zEIs3BfpPSsm6jwTaR3Qdql21SSTs6fGoBExePCZa8delRM7zt9UgfcyIWq/CjudsGKhX4MNzMebqV23/6+fNwaH1NTYEAWjdP2dVwE0hrbFHhiBWq/cVbXu9SAdCoBA8r0UKBCHZWN9YDGlflN6AvTJXDxNiSZkUvGB5j+pHBOgqeP7STyIRsaZ57e7GA8c6gQ0vMzX5E/Bj+gvKkr9o6p7xhMwKswjbWlAkJzgMtElG/j6w9KA/G1UJ/i7dpFXra7vyC1N5QoJQe3leSZoG4fkcHH7fWBJITVjIOuuc7mT6XRQkw7/RO6Y6fkl2/pFLZ3Y+/ghVVG7thL2+lXGh2kHrxknq2ZdDbxjTQktiGJVLz1ayAiYv4/xGAL0D3BewtFLnGifs8F5wv9odFU0a6hwcnQAY9CyvSP0GeptLIZH+qabGbJehNbMo8JIShJZwPcCqJrnxt/9UR64toFCWT5yVxlIGylNgOMdZ74d6c8r2vVRru5QsAKF4IL/2jFWdvBwTfFE9rOnblVPYD6kKUgLC5QbN7pa5QoHuBxZpGA1mu2AaNiny0LG3ekQ5PxwPLr2TLBHpIjcdGhW0wRxUx3XiC4YJqQ5SgvZhTVexqR6OTXzDC6vrJnfCSvXMTIcH6K+vnWrLSjDeSkiOY4Db+QiKU4UiOeaf2OrAhP7Y2YWCOaUy8R0tiIhwkZrYrQWMYEs22JqIiQsla/7MRBOVepItdrXfH5U/xjwDbbZFe4IdavwI0ACa61Q8E9EXgDt5PybdPYLjeRBw0BlktLo9h9evnON/+2++zX1v9rIZPoI9HFT5vnOnoFNLRTGteKx2dQy6JtNaAWWrCLWfpZEweCWV23/3Mzsz8VZIuYX7fwwMVsWoKBhb86BCIMeh8Tq8S3VzJQckLVVLxMfFjaUkVJyps70S6qk3by84xjrVppdwbOYtO5+nGn8BADYAmg2NYrxWB8JUCxa74VO1+sSBm2AzTauveZIrqIYnbgZlPrn9g5uVQAjARKDP1UGiA1qs7T66xTFXnYYG4AGz1WjfU5DsJlvMAdHAJRUIaFVb9V1BGI48FMgUVBPhrjMvU6QTSepNjtnR1/flp9WcwWhF5Gcr+QmHNLOFwd+d61fw/RnZk3qw28etCBCxbwlRrqybnx1G6yS4DEWOl+G5ClLpdlwj7I37xr4pRmRjeMe2sXMjxfkinhiBLyZQW1Yvvn4kWr7M3r2nUvd8rnrsEluQg7CAuUBwJlRc7Ucfm6sJmui2/M3RSGowbXLgK/1z8G+ipQvtd9oUSlpT/BJxoYS0t0NL3bPuANyKWFYDmq1pOXGhUXWCq7e11RURH+tJ3kpBQqELbVrZhVy2qKiQplVmCNCQoWKnvE74ehx2uNcy4i8wxZIIMSQN4qEfkDYElmhM6xlzFEzNhNfE45P0hCy9NXt2QYUmC8/y/JNA89KW2fxdOt1fKFxZ30jO8UdJacNOkTlnOPxE8LUNg2G+5OEHCmSkDOo8S8Am8VKelXuqWjY3njMOTTjdSlhMx33L0U8/h/GOEkKxWbwV/61V8GW0MeTS+cMF6nCKhoZBuRCfZkrRrEgYMncsvWSCplNth+8gbbJMIK6zR7ElIAvjPYBXaKnb1hqdc3+WL8l6uV7xJuk7cqhcxS/Ro4WdyDXRqy+7s8vUFvPIYRArGaH3WQxXoZ9jHZp30NkE//633t9Vy9TGloGts9nU626LjLiC6/3OGCPGO7gdbMuPhrLSTab3BE6CUI6tBDUljBtPlLNh9ZLW/3DjQCYMvJkNNlbEM/UmhanyQsogswWws/iDOocyXvus4YI3iYsU/LZk2FbcIsSKCZHO8eNam7NC+CJx9fKl4AhO9TWgcovJOx4bZnW4+Sgymbjgc0LmfRAbDXQwpvptMJmB/cj8lqR8tCotygr7+oXSCY8/pAVvm4mZUAEPnpQBugC1+NoEO66Jq+UqNQ3vXV3kw7zLbLfurP+HtWqUgr8YqKE5F0OzQBKyqp4wNMyo9Rp3lQg0/7LuG3FUc1+VUuz1mscNbOkrhaq7bGg8ycDjjD9R73TVp4fPHhsdQ35ubOL5hxeoiEky8r5EpXxAPE9NLpnZwvJHy3qaErm3xqNpIsgMh9GfIqxiM+pX9J736xmk9t1xa6OUfJRLzcEoj7qAKb6OeWR1aIWLZO9f4nWX6LZbeIbZZRUeiIk8t5xKSgYcO/Z5uagtoiSlYYJfdu3AENaQRXd7FH39p3OY70GHz730Hu5PebhRae2SYEGx6wv/+V9wS6RJEt6AoEcQyHf8uA9wXIW6RpQURGnVCkzjCea9e9V4hlY4y4ZBgbi73MHDgzTgFhJwu78Y/CI/PpkO74DjmKiTr1USzLyRHZ4hPnOGOr2k1we0R121ig2B2I5VYGRQ3vjAJBSS4j7Vyi5jI3mYZwvHSYcFvzEYwovntbSYy0JLUq+q9owAFlJWPNn1TNKgU/zIhxlSdW4u0+kRGTBXHY2ow8KH5Dsn+PTOfDLwb/N7l7T+7QgyG/55sOYoOolK2rqLDSp7SwZQ3nsyMJoYfzqn1093bXosEV/ziOS34Qc11e5LjNdyhZCnbgYG7ZbI0VR/6ObEGfG9E0Iv+8vpHAiRQJRXYth0H4rICABWHQ/7UPiZ11zsMgnPpqtApMNJXh9hprGGflI3YPITy7UljN7OoKFbMO3B9NICIAC2Eu2FxmFZMGn05/anjnjmvJilNZjUaxE1LIg3iVjAhXq5bPELcvKsVCKvNy5cgJEb0elwmctt8qiOfuFo6LkR99YpqYC1OQmvbQCajR1Ab2e4ePWit95ZGk83c4bs1uEcfwFZsx4SYSSzrrsn5BvaHIOujIOeJL3Ck3Em90BYphYnTP2vKL3KJ6r8NohuZ7WKnjiPfgmtbmDYvHYI789PFfWLLcs3gsNVI6yts97e4kYV3xPe5qLf5cz/nZG7KZ07T+zoA7W3b1iSks3/viaCB+TfCFXEgzh/X3wML00SrLvUMDtS5LI5bJXY8nEpN3pjiFgOA9kJrp7ryb9vrWw/66oU0ioQbR+Gk2RJPNGdbqkwm0A7eE9tjihC43+vovsReORm2VuuTJXINFT+LAOdVsq3lzEI9xpwzWPc/goYtxGReJOMy1fDaZZP5W6StjOTsUCH5482+d1LtNbtD6RDRCzs/KJrOI/y0LEOJ6U58XYUfnTCp3h2ajOdQ5WauQ3z2XGBEdso2fO3la5bnhy+avRcTWX7bSdzQtPtnPWKmUyKZlMrByCpuZlI0ZSEc1iVVHJd/5mnwNBpGPFMyuddXU/wIgVX/YEav6UKmLKtOo4h/nIGKgRXx7uK37esQVs/njF+cnxP+E0CE+/bdtFqBBCkRRE+QvoHgSmA3Q4Ir19Q6r9IXJSu/M5sx/czg7W7nyERzlUiMXrYVe4Wj1l7MtTEy73foGFqq0eIqlrhf7JHSgEeYeIvUT/+UX6Uttsd7LZuldIBo0dt6qItlQc3VCnJbnww8Au8DgPGZOHQbg3Fe6SWeqqHb08PcUvLE9GWcIJRfZ4uE+1UtTvvCV83F8o7jkyg/KVA8OJ3H84xWeI1mK9Ev00VBLxKU/xNrklJPARDuZlMooLyy5ydNPf10VFEwiGtTw7I93jg5K+Qxlw3MVBeu1uOgFEb0b2amXsf9LUWF9iJVR0CGuDvi9oSNg+ieyUlyXjPj26M9/im6s5DB+o1Uf6ruY25mEovrlhv/7dGE6HDIGd+uywFBL400lWG6Fho4lXSjR5ocH2/a3NwkJ6q0QxTn/a70tY7z5Xbs/H6AgOvYKKmenXF2IuJnqNkIE8Q6+hiDAxJZMesbjoDYKcAAt0nLbDsijK4tlQOYW6sMobxQk66obV0TFk6ailVKp5GgLatB4yDZ4rtRnhsDmYvnBogMmgXmiBs7xMjVU0Z1uzg4K66P8XJ9ChgBujQSCJDse+o9AFP3zoFIL/5IUjpDu6MSPa3mNbGcACLeTwbiYk6UClNGIoJM7MRpVHcNErwLsTuw/JQ5GTKKa79Nu6yHZU/6pQIlaLZ8Tiecikhb0kRrn3fncN20IKo7h3uWwhs2IVoZJ39BcXXQ71XMXJZJinMK0fSw5x/sNuqpTamabvW0QTx3a5xxMavrhMr2C4eDNfcjAsOl0LNDn/4wxI4jrXGrdCVS4kWsVxCJ6cS6eRdoZAiu9rkVSH1hS+Lr4QRxeTukQBllPJ5fa4FPukMG6E46mpqF0qHU5zlhFZUJSrZGzf5NQDLs8ClJShTY8tbldczc17bEyE982/Q+Vv9heFp3zTdWtAiyiXB6S4kGyw6ZQ3+rpZnV4YJthC0HGqit7uWa3WknWKH/GzrbfDJAAB4vHF9BDSxvWl8w3ReLsEYfS7lx7pvoTyw5OY3z6+xI93SlSGvO0aTXSP3eWHd4sQ8zn0xEVDuoCpwDbIQ3Gz30nBL6guH+zFHeGXZBn8PJ58Q/56NQIFKXjlUMdJSGz4I/VvDc9JyZ6Vup82iRM1Y4AKiAastHrYToUxAtgW7erCF9WNTh1JFj0exlC9qGXr1HNMZsKMyTMnjLfsXrgWf35vg2X63eSw5S1BUeG4pX3cBZo+AHkTPmbz0AtLX/QWgCAehzdtQiSDI6vHp8XMdmkLn8NksGT2ZPNNcooUVX+Xe00H/i2HwPHQl+DvtklYDTIG1esXBtQyCBfSXk2+/xAr7I74ZwRncVuQfz8mqelCaYWc8cTaBT5VWIDIDGEL3IUcM/B0bYVLJkNktOCGS7finNct4KSen4etlvLCtiC9w1Chn89VY0S6v/FbIkn0tZmXS+vKeiA23CqgAq+j//udVc/38PFIwL13RsJxbbLDZfVrrGq2keIymKzvjd7qiM3znx39EO7AHI7KHF5Nz1CRkwGVBx4ne18yi3uUZoeWLHkqioz4erD7aBGhIPy8IfTtxEIrfr7q22bo1vVocddLA5PcFI8OEB6SYQw30jiDIm8txzuLQqJ2zxLoYPc9tWXd3Yjs6Gy/WDkWxD4zHbTT4I9a71yzMj6vX1SlZA6jmjEIaLNEf0tSEXH0aw454o9eYoB1lBCjs7kz4JKvhgSn9h7gEhopiW8Fi/tt1A/iX+VBObxaiSx+VXbr6Rg5N50RBVZV2IVjI1SxK3K/TUO+0MIGxnNtoW2yHcUyLasjgC646riaeT9/rFesN9XG7RauRosyq42aH1pss9HIEiHvG3JaH9EdBsdXx28xrGg17uSDNcnM+c22b4+i92Iq8YsDOOt0D6A7aKfhMyoVRTPavTvlMgkxzSBg2ThPM5tUnvw6KhBS0TCWROglZGgj8rD8VuJhmJirHowj7wopW0JyvKMA/ZBFVXKrZ5z6l6fPtYpKs/bgbn2q7EvVrkKf/2McWGBsZeIgf0gUsRrJqI/JsMJcYyjxtvebn6BJzTqZWhLPPFol7FjdjMk1YYi8NXVA/6LwUY8edadyty/3/GEhM5LjPExvRsl3IFcJuZ8l48XdQH0eWPlu4Tio9Bze+o2WdVWRzYOr6nGXNA4gE+EP2QrnKlqAwsa1Rc1USBeXswOrm9343Dx2X5EhDIDl5DzKF4O77oMt9O9yRNynmAOiC9fk6x9dzgkeBy+Ht9Uc85nf6g7eim3sh7FIlZwIF92wmKkRI0z4fXuwPFbGGkQ7bCaLisbvia+nyrps9OdlOouKw8yWl1Eft0Vvq4vKec84c7BkV3HUKZPRkA1d028wI5KkozWgHLSQhePT+0aGRAR36DBJ/d0anaa4clpwDElwwi4g0uj/0skYE1/pyRPDYfDqd7WzIONnQRIGEJJQ35d6GHGpRVfoxacbW8Q61Ihr+jJQspVMTAj51/YnKk4IU/1jQlOXvGt+6E92brLz9knVP2Vwr2/y3cQHGeGpEKYuX9yP/0dhV6LYSlM0Nsaa77tmv7lPRWdu1AQdMPY/mCczQnUbnNPCwnWGyCkVTT33u9lFUyb9aVA3tvh9oUiDYtBf7Z6HEH57yqGnOulLIr+eY7Xn77k/mc2rKCtyKhWTX0HIA9lNMhc+oC9fPSsf5vJUhRRlFnEWjsSasZTetZjuJqSfxRuMcZMjbocuXlR7CwUJfmIACfjnjnOiHRVypKMj0xVQCwIksueTbsPah8HBHOsD6j7CTPnQe1kWGICa4Lm0W/rDAsca2g7XTHjle97AsmaWu6MLjN3XFmgoem2Na5soNvnlmnrgS0o+xdY46d84e0PLI0haXB9XOyc7viMGJSK1fNudaY6c/5iQhGsu+Nt11UenJ4djEmHBGTtJixrXDaQTOh2j1iXFhaRYMWks1e7GndGJzx9qC5WhcN5kJJX6VWvymhhPMV/nwr1cTF5mbprDcegKNrh7MleSJCmWUqCuTqI4Lq6Af34F33SemY+SGDWZAidCvPBdHdhX2m6p8j8TA01p7n5MXQXW56CtALh8kC5o8uUFe6pDhlZFeEVrpdq/b1hwluwtdzxHXIE8qqns84XidHgaqUCz1gf0+/KVDMz01fn2WG+GKQ3U0NKeAyTToIGOG1J8KIYt0N9mBTkIKVBTAs67wIITmmRB9D0AI89nnpfe4Eybw27J0j3qFD5tMkex4UdrC8rjvRHJtkVyaWl7NG98Ttxx3XUgiEp3pGQTGZRPVpYGdJUZGrVvK3V0TSh7oycFXQQl/r0Y8ANZgMpzfzFA3Y+RF+erUX9O0P0hmDNn7k5+uElZOBrXIpf6pBTsAW7OmSEgLrJss18mmKpQzGr20fIDmfLWwyTacsEkjSP/spVrC8e/NxHqicxSlcoFEvecyiNrMk3n8TLSPCQWCPZIQgQPCXjN9LYqsyr93EVAWqP+6/Xw1Vwn9oV1AWnKTTmyTiyWHfYjj+XkMU4SvG7ny4nqty1SN6rVHx3nptGxVkopZ5sn+aaxBhWELKQ7YYfH03CPn/jS8Rwx6Ip48G9XYprL1HGYSk1mWvDED1uqq6UocEmbCHN9598NDAn2UhlrMl6PUZRfDVHwdWKhvptZmTUMDNLh1pzXkN/VxLAnhbXeFqTFyhh4HbkfJJMghpYuqxGr5CNGwsPconyE9v6gL/O7taIK3i4+ewl2NbtTQaP65m7jkiR7veFIyHGSJ9Vlk+UC3IKao5r+9AvGNwfKqMwx0YEnVio8SV6UhY3YdY5cEs/Tx/nM1NG30PoUw4JZnjq/BG2DO1E99OdrCZkv7VGvIUt151rO/deZL61pVZARBQ6kI5H3MWasiioPigygR9jqtOlvEIPR3RkXcwOMT3nO/ZLobE8HkJKNSxctom5jxh5Yh9m93I+SW6skjBAWEGgtc/KlHEiguRRz5fQwrkKm7SUwvofoBXPgfRdShNJS47O/1Y1Mmn6zupMbCqWwyli4aFqj9E1hpKsFbFyJmmwakEu/7xWSO33hVdI0+J/BhIbKxe/teP6MYyxLxqniigZ0oIpRRkU6knnMfO/vGglmOWFwBuKX6uJUpaP+umKKCsI3xebV2kYAZkzOUQciHgKU5j9BZYsDeoKDuqNkO8tvS15/gmORHmi9qR03TChUxS2hOsssdC4HzbS5c20gX0J4TOY8t49nqDu8x2N8dr80SClKHnr/CgtCoLqeBdVDIUFhwEVizxID0RYRRBQ/TxckCvIBQ/5bZxMU5OIN/sEAmqiNK2Lj3dEitSx4Ms1xqn2sjA1UAOXxN3j/JjHqg/WWmZ7gr9PVqe2fifP1n8JJLnC2uAl4/Z3I+sMHNN6B2J8MLWMYzhahpXrWIOQPONxTXGWJ2d0pit8tTI2nQcTMwEhovr+7cHdvsmkiE5p+uJPZ1g2KPR4Rmoz60X4VOpvqBId+tQ/mAMkLnYSR/FuvlP/RB1KhaPwAFS3VrnDpYx99P2eEhOdMjl7yKOEkYH3GzQz3MB7dltfpE0Hj1VryCdovDNtqC8C/8jCrKAJc9y8UgJ4qDZBLnR3m2OV6I7IupVAMn+8HK0Hdi8UsP6gNiBc8FmMx1Ijyx/7fkYRWitaU1ht9TBQaZaiI9fJupjuyp9AmlojxrTaPAUAcV5Fy+//1aCGU8QmgzZWeeSds8vYErC+Y4ll09DJxFz2ilMIBzD8QPHEiT7lECLKTHB8oov6EjVhywJ6QTtXKcrenBWlPE9mzYqaNK7qyYt+j2uPqUBXKTiB/o+bM+0x7iZBovXyZRLSpsrJnJB/BqKJG71QhY41hAdCBeiLuk6px3N2AKuwnIIv3Oa5Of4siYyyg1Rd0UH9j42WMthJwJuL+OfT+0viZq7wDlfIJiGUJkqve5c4d6wuI+3ErzCrbQhmBlJbBrJEWIkiqrDlZZByV+Qpzg9s1Q+D7ajF+r3dnatiXqQvk/PPxUxDZTxk1R0hMGcyimoY5V4rKM80Ant9QnTcQXCDoHClGyjb3x17dSYhmNWR352u9aNThxGcUlDoTfqALl9uXAa9naSQLskAJHpNY2+fO3PPwglHxwBgfJwnDQJXPGiizb9IDIwZaW7BzWztLgmF0Db6zkltS7/vqqz+XfA7SCjsXuUpM1fqK3SBwqnRmyCzFl+UTskQoAoNzViss/0BTjW96/WIa558fr8h9MbsnSRE85HaQtjn/LJi1GFxHt6pQRs5k2HEcSiTSW7HNXmdHUOc9izthHMj4Tv0fU+pH5Vyl0zNrbcFzFeR3lbZ4ojOUtfF8qup0HSwogwgzfadE7iM9PLRbfeohnDjCsZG6LYGjiddOmmg8iWhp8r155lLJX/naDdzUVtDooG1+NY/kfL2NvYd3imtIcVIyG0GqZB5IclZ9G5h0MFc9b8apXmB2sbWngu0Az+ZRSDFsNwceqD2V7p6DmUpG8uzVK7rf3WuL6uyq9owyqHOPE+OCWdh5edGHvbW5mXackn+6QWq8+GCC+5So7UQbbjmi+UA35J7WYornF4lbbXAvaqBqJ3DEVLlevZN3kO7x7KsU0zgCxsAKrj+8jGSFHHBSVFs1/G03lst7oghoHMPCjGkLwoJPJQNW8QeRKWeki/6js8l6LMltHN+yPwDPqVTzfbNHlTuD8KA9z4H3ztuig5D6nW4kY882b7XrC7NVeA4qL2thGBvVLpiCWlSoAeB7Y5GJdcj8cb9/OhZUInolrBwYBdIAFADpQYI1mfK94YG4qEftRf6WgZFleR4JbQEtmrwd26A3ptnn23XYjaMoxiQFskALL9dlXLuhFyRJOYa9NgdTO1ZwDOVOtr25cI2ZpdzsXZ/4Xxyq2ikX6wFgn6sKgzizTaJUYEr7zoBvj5yu6TKVbqRjl+A1cMbBxlEq8iUE4JPWTwEy3UiQI/UP59tTnkzmKkZaRhZnOEc+0GOg1kWZYsVT/5U3PSKuaRYWtn78d8gn76uABslx85TVfDQezRkvDwkikdgmwEruui8Z7yKFCtLvG2taOZDtYzwNqga8On+YVJTj8n4e33XlGutkbGlv7jGf/GiPilVuElLRPJgzjvpc2WxvMYUUVORE7nN0Tkou4MNZY0aQxZIU99YTtSy4nYE5VTN9YTjA59Myp8eWg/8JIXRHDIqJcs+bf7A0T4TMDKhd4G7NzRWIem5mDNKkRrKj+WONOCzSQiwYOpCEXrCMODsB0lhnQmroCRXG9PVka4d767LOpHQX/fvnRZEWUJumgWp1AwwPJe0rV9vhne72joIESxHTq/ogS9rRYPHfEyLtNQ0Y+i7kCrJLldgBEmSzzvWBHwM2qWyeLShVHW15hHCVoMZSiYHL/zxubVjHTmITsjTuXbINp0oihW7K2Yca5Pyx8bI6z+/FSASTR2JoenSpnc7gMK1UNFiGUeejCYbkCpDM2paCDQMw0MKdxtfpY4h9aTkEBOPIqowBmoX67o0ym1D4xwd35X734GGWyOKwh9ABPrcx8KXZBmvW7GS1BuY4Ji0vu6H9fgvIRRCsf4Nbw7IQYbcWCgcrgUMZZaayHmjupdMZU2rloNEoYMncuQN01qT945Tw2VBgIJt0SquaNV2TdzGAY2FivxnHALCyh8jXYl+I/q/cdOsYhEv8uBckWncKfEYx9vMeG9MXzaE+G3b594FBFEvXdXHLXGJ6+O/ClMBC/GsbQ7vR6Lh3odUEEkWn9+9FePqJaNCrHzrqbQkaXyYP1NcHyCZFOjmzC0oJ/pfXqKR9PU9blSwCWnt6st2nqy3FQIY/rMkIxwLYm8l+Btb9sIePLGJJx0x7nI1NS1/AE6JtFhfc6AasLu113ISGJtC5+ccIbYLJGsnxCkn42qzieKdgTPthhJ/hMtNxcWjqLXatN9rR5pDYibdkQBI+GKGhRiEeKx6LxB+EDGOY7H839fmOgxzIjN0q+kfwmQfebDIiU35THPDFA08izzLJPj7lSlKwT7V4orcdSlQPKanjg4BicF7/aOAlQAaFpj4fIgxZ6AAmI0lFvlzjlqsQqjxjZ5uRzmbypvGzPTkBgCR/dfc1ojRuftmz0439jg8S4zyF0DxlyMeMV0kInS882ZGnxKIRc499fwDVUqqu+049g/hedmqioXuN3vEOC+tyNby+i8I3OPs4MQPBuVITx4N2LKY/ib39VazLqXhLxtWjGjZOiEo5BK1hjq9H91A0dTPoMy1fVz1FIAZbUIfACfUMgonDOlfX+Hcpbj1+xOQQSyOFsrCHiANZcfD5QrswuUy5xVAjoPm1U378rBuRIuU3T2MapGp1QqJhgRzDebjEkfemGtYt9LWS+i2rPkoZMMUN64OyjXHMahhCWawRmr1CGcLohE27xwDdkJXF7iddHReVbRepx7ZySoQv5SZqUNxeJBSmRALP+f9NURePv7sozY9STSokMggt43RKc7Nm8yUg7BO7aKi7zvkz2yZ3lMP3/SCFZHD1XN254fJTI+tqAipU1go2avNctG6ivw7oyh6mSW03W6FkCLCwBiyg/Dd8bNk/WDYDMJdUpyOsBhrA6fUq+qePOysaKvcJ/srVglwtAE3SPwt3DsS4y6XntdCvlnj6dP0Q4EEopVFxDgGEYOVT0VQb0nsajhq75zuk9MDe9Godjmb1c//wkWUdvp2OF7zfoLQu1Bsq+Mx+29mMdtS48px26H4C10LbyzwY4hUHbJWfkPLo73iqMPZNh5G7XZO1vpDMQ09a3arz5qrfpH7RgwuDjMc387o8gCYOt7+4ssGFS0e3UUr2UBcir4cey3aniWLoTHYa+0KprqdM/FwyaAwZbUYF/L0fOxVK3DIfDhRy0YBSKUswRkjorOPM47nksq7iKmF2k9QMXHCNxq+Fcy3NaesBNPW3cRnaEiS/f4GFqXGFGoqaNR8LG17CsvI3pYCma27S+Z7ULUXvO6a3IEtElcRZ+iLTAJ/vFLztwW2ufUrYBsynLoR6HPn5ab+zU0bvqBd039nOh7bIa+h01fa/OhJejcFiwVcsXJS5a1MnLlVP3voWQZVxGicJ/i0vqmozTfYtZQqJ0CzvdprLA97yWttFyBcM1TjkwBztpovlkv/+OMeIdwoTm/HSg9ECEj21btqcimt+jmDQdftKwuZbaa9+uqQq3EaVoZXilLdjJqAsGOnVNYUPjaBKJ/TUkNvzQ7MIgaSs4AM6+nRuZcx62sw/ENuA+eyjQ5h764G2pveZMuKtZQxfDm0ypqNfRmawGwctfS7DgOt26yX/PTiUim2VYemJm+HTwCN8ODpGZYEPfjfMv723ZB6h0k9X+ZmtNApmFawQYyF0FDlRxDl/9ckBvHZeMOF2T4bXiROJekG+taZ629s3rih9MQDCX4paiKL8pyXxiaNqFCclMtov0lXAipRSZgReTrphd3d9qbgpCCcbfYOMUz2b1/LXFil0sxvKem8IIGof6xajEbof3hLWsv3mEoSnFrFzBigzc/ombpfqmhz6uFBYTr4x0+5Z0wX+sN3kRTqul53Vn1vPbCN57ab/jHzHjZQ3LlvQTxOXxBxXIZOzVT8KubGnvGg7h8ktucF2YfGKHVcLNnfZa0wPT5rQmQApRussU371TAkEm6ueECWNJ0lAIVkWC/tUFR57XUnP14NCySvV2xKEWPeDv4/XughLsb6wFQiQS5rIOF2C00kWWToh9OZ6kAd//twNE3zCvjIuk+m8uvLVYMtqjIH1Vizdmxu3dCBYTM++YzDV6miGOznrViIGsajdfW6Z11MG9mmYybOKOo57cNds/VsutIHsfRiA9iPcSD18SG7Cl+LraA7bGPXN2VtHLLIbDAg45ST+CT6qAkDtOTWgsNuG1iwkiMRAMNeP3nrkbKhyV4gbXT//1xZ7trZ+DKH7EK+8Hr9/IRz7s8pYp9lhtXy+VyqjlLEr+pxn3PzBHdZ6Q4ZVenj8HDxGIfj1P/FsFn6xSTGB/pUYju3UXkmhobk5Y4uQMIMGXl6/B3cjU1NCrsPJcjLOTo6Bbfb0YzIFbEIKRz7QMbSXDGMwaeP1HpAjskb/qCZockPTXBxWDwd1tiNdgIipdMV5j9YKb/38bH0yCSEzoRhp5j//akjTwi2bmM+r/uN4woQwsXF4jf0HcjeZDLZDWvGCfosq+B2256u8XMfb2KvXP/V6sRHZjwCbUnNHFZRqtgTJGThh2Ic/rO+DmMqf0e8oJj+nfTI2kM0vshgrWILMGq29oIscljvuZ53Ejf7S/1z65cK9cchAhyEdtWAH2etQdQksoRGRO2wRbAjoFYshMtlmzPKQkSAMeCZ4hbcO2BVRdrpXLS+zJkzFuEz+0/POtiGM45J3oWxgbhH753A7yO8yS9UxK7dNw61toZ5YlP1R/VBeR80odfr3QDkKa2L061il8bmgcCF1NCXeoCO5W6F+rrNUb3/WUPth7AoPLtxHDqZQRNnNQeGjdMUOjnoD2Gu5NydFk6kJUoc80pDjV26fknseZG607Bn33SOEkDUDfMSejh7kMr2y8KhocREaw+AzbLrqZbHpf72rTZT08I+ITTtx7kBikoWusMK+V4pQqcdL+MiaoCYdvYR3ZN+Iz/bqiGKE1QdTyeDOHSGBxB2kKZiKA3+MP2NxBYDgZbXjoTcySnd89UREA5bscqhWekes5ZEE3X64wC/csr8JI0C95B8CDJYAtn/y93ddPmq2J//4pPYdx2fZvgSHuD4eTXFJMq/vAfZ8Azr4BV/BLt0uzerDm1M7YaEH9SeSr1PYYuD1ALa3bbauxGiPmN/V/dsgSxVd11ivRr7S//kztANq8ppzw8ciHKO7MhUo4kVIWGlNW8gcgSfKu9990uDIBwYayNy4mkZoFupKAnwGxTzowiInc/2EgEkhENqa/IA3pVtYFSP8I/vJl/V1U6heJ1yWv3U4orE83f3NXtivXmc41XKyKxMPhAgBlZRd5d9mPMHWzvM5ddlU1WYPXbgWmohYuxP7tZaLYXT9U9izIATX6PsW6XTx0suWqKyBbh5DE4fAyzAonRVC0j+S0KsB/QSOYwzUAcz/SeHcWtfLItySrJoBl2Z7LW7vmYBYkRt7AzFQreJntkAj/9bl4ULJDxSdwkkloCdA9Bc6QsWPofpyCbkz+13GRNyKCN7DJwb7AiRHxR8YdfVxGZaCWZwRdUWCcLswr8KDYgTTFQls6Y8Rfsb6BNjE/6wW+tqGfd+nAtn6q2sBcV3WI123M39iv2T6Uo+iuL3x0Evik1oGNBwnDkwrrXGbsAdq3SSOssfGX55N4EsHBA8rO8mC9Zsx1xHtVwWBAdwfoqJcG/1Ihq2zjhFIb5M92ZfGcUwwBTZUCGCyYciPftBRAhqEbyyL3fw7tBY1JTCAek7UxTTbXNx7IYCKBL7ZbnBo/cSC/Kk2H4+ltL+Ef6kVJ7SxgWf7Ay7zVKHj+6uqLzP6qf0q2ssTCEhqsKkI/xututcbHLYFdpIA7z8CeC35lDn4RV5noTsZjfi58dyxJxYpOdIQO4pipTYzWwPY6ijP0p76jJQuFITveP4x05hbfvIWynYmD/c6spNRWXPcYcBvt52FA7rLquR+TItKV7t9764uqU7DOU+RUBznMDilBSxlY089CCTEIvvtLnj5BprA+v9enLq6SEsRQqllKwc+5BODe0dRAU939BjhiS73ZTmldUnY5bNc45EX8W2CGfm/Od9sWX6wVX96S3vSbcGDYxmdGVU5szsN2JcHvFyygYMwvt0alnlE+YL1mv54lRvtf/zL9GUIUrXqQ+nSGzDyt1hzfyxMtoXHakR/aGhhj+zDhinCy9WrH4Ja2bfVrJEM1lYoh4Jru6L8xWCHTvxLOMqXxVA2ByyQ+Pkn2RX0RKMPt7N3CwCN5PjlBt2YV5kopG0ZyBcdKMmgBn2/kOppFzAzCr+NY6U8R3zj9io0wT/nMzRGvg10wKixX7tP8ZDpFFwywVDIdvVpzqdlfe9Mg5pOxThLZLsR5uVmEUZBZ5iTbuR4iD2XAIYJgQ6kJGuhBBg/1UltzTKE58zTG+h4UvFObjc9XsF5WvOvdP/YCg6ZLC1RaX1faPlBPsHNiCanMz3xXt78scEydaO59MdvVhXgJTTW90Hy8rLbvUYGHhRt4lArX2q3BJD/CIBA2TRTPRJED+D8yBledwa3b0LQ0CqzrhBN8Mz+FXHZTf3YmB/z0o5/oGKSq8QiKSGfypF8T8bRyW3zvloolynvTFdoWpW25R7AYgc7cMNhWSkj7nN7lnSgcOmBh0Z8uurQmSlASeSlz74Wdn7TYNbOwVvuBlL9uDGzFPsFGMtzGmtoApVZtY+0+YSLdpqVN/44a3Nv42IqzNNDOwWmTq0kTHr8wn4uXR7/rmRgG2rBfm2igVOe2G+obufLh87oh05AGSKhiAMWxFWKZ4O0aS3NLraJiG5KqxqY2AMrYd+hcCiEWiZehY203SsexLbELQiDGYHFbXx+3dDx6kz6mvVMCB8hNESaF8lotISfyvi4py2SZeuopko8hJLsWNzRdTHvxupJNqZMTG0OFaY4w8LKZoAKyeJEmW3eRuwU5umQgp2mSEiFyaK7lGtLcmdd5KZlSYWN0CYu0KloonYoaaVWsTu2ckRuKGLt/ziSpza2x0G1Qk7SFT0KnUmLfGaAspKKJtZ8V9OOE8VsbOGct3K8uWZmFLfdPVUXOSzRBsb8yjSYRywlJmhXI1vMerLFa/m+T1fuvIB+S09TKvfxlrM+RK9UD1rnRwXk+qEz8Cypd8Dm0+35WyoMyL1j7WICz7RKXeclvYgAx3o=
`pragma protect end_data_block
`pragma protect digest_block
a5647e1044ca46e64b736674b35fcf3df88c2e100294dd913d0e69f7c2603201
`pragma protect end_digest_block
`pragma protect end_protected
