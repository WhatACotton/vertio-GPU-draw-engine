`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
oLJQVa38TGwdWy+BCvD6I7harMzTNVOz6WOkEH2PEo1fUOXaPDdl0bUuUq6rOC22bMN12/ErfGtg841XJwxFwbCDQqILGZRBf82y4W20lOVM5JkxjlJngU2FzjWAqLMZQ96WsRSHPdTX08v6eCQDTWvdk1l0Q+LPByot+CEE40KoYtyu8L32L14TI/SDTNob1ubB7U3z+o6/hAb1sRSqXAu/RJPOObQEhrpiMD9SZawIdum96JQqa2iBFp/oukJ/O9PPFrN9mZ+/V99ffafRiCsJx1IxpJOuNv9V2gWc+lta73D+ysJVhIPt3loUjQAoTjKR0+e5lwzD6GOUlDpSA1oxsZMwtZwnJyYqJLsMZj4XG8RqSwrCUmc5S40Z07u02Jdf27q+kDrH/cOEU3DvqZNtBmmtLL57CjguB0VJ6VG+1fYAkzP7ktrHL02Xx6HkUsAnpyml/TJqbAuwi8axJUUO4OIPc0BfuBIZbZt3+qjlWXjJ4lDsH6IBizkAZMt6KT3MEL6iH6jVuXW15vOgIqEAUq4BlkgomjqTdMuQAwm/LrQV64/dt+YT1JpMTpIQoLCGCEgSxYsnjjpYRPtrk3sFc0mqJpXTDNSCclt4hqZJQKCSiLjE5rYywJC91TFedJfQ9iPyrTgNGBQLHXhcwmBN9l4P0+NIee3dOuIGWR9bZ2jKVdSnGUj9LnfIhzLpfaKQK7FbCAFIobf+l5bnxVZAkX9DydUymstTa1c/cMluBD0jSeeba4kZIlqTLdA/tQ3I+JVmXimBEtkIJ1vVZHrT1HNAvq+4vx0SkIfLxlKTwM1jKh1mrq6AyB0i6Fx4l4BwEV3/KYJu68Kcy6p3HLmVeWZTUt2IZ3invxMLD4N8XsS6HYnW4zCd5vPrK5zNHDXYtq0TUDWWAtRoDmyUu3s1Eq83F70+Z17IZv5ICIBZEk2cIaqyPKrnkS1jiw9f4MOnGy/JufWIJ9LB7+gAlsMJ4vao25WiFCgGK5g7hLXcQOhLSMfaPA1zKL3ab3Cw4wR4TevTgkGvEcQpc+KyklI/Vn7+yBOh22yH4HlrQ2OOIdxo2yIu/+BKOc7KhYPiPqZJPzlKmhKVNzltF7VX1YA6Z0H1fnJeu+N5e3QzphzOG+UnyqWv/zhnSz6ilBfDNN+Fo1++Gr1GMGqvrbQXd3POuZHtvIc1SiwIsu6MZKiC9wAjjZ2j3iDg3EnwsC3TdXHEgSZLhhhiUbLmWMStTMopUx1wB5gyNsPwsg7tyE5aa9+9eFl/AMBmMJ2OMfKljQS8xz+HaubANODSNwMNLtl3le/kJCNO8iGbZe8cU5thW5vakjsDTPKFn6K3mPxNiZv25vMXcU1N2stQRPG2DcU5CSK6PIpjGfWVPu4nxgbJES9Br/VsNOb9oXtxS1erOLN4cwrYCGgje2d8OtHarqLKCjwSQzZ+R3ei9zMY9634dCVUUBQCzSAzPw3RMy8q7b4q4yf7YU4aDTSx39XsYKUrVcawuluUIZwbinvWPJaLofp2k20b3mKxMsJQ/8uG/vMATAXIBslcKDYPMwAXSp2TDu5X1FBiJazcxU9Mo9hrV2CH7CB3y5ikhYWdJhPehtb6guZiyxIvToqc45sCELC9ZK6EzAdMsNFQapVjMB6nKO2b51ZStj/y1s83dwgxgzn6Z8s80+f3qsrNOxN6EZiOhfbgNXyXrX2dGOI59GE7AOuoNmJJE+2X7Rkw5hrQpiRmJgg5YevW8ipgLUKdx+pHSlHOsDuPa+YtWwklYf/LDTgL4w8tb3R9bx65osTzdA9KBsMPyrlCFBxvVyMpep6x3iPKCkG15inZV2FTmUpf/tUEjUqN/599zzFWrgjW4K9lxX+UeMh4itz6u4EgoqeikJKybiLdxXVHQULHZ8MWb8MFp6oUgaNoSqwRDcksAbnSDSF8NYyGyzPIDJEkCmzuiy2qV94kLcWDNQkBC10v3Q/YI0+jjPzspXSJdlfofsZQYEImic70nMZa0GcvlB6n1neRs/yjOOrsbXW/AgIcodeVyf3h2ki8gITCVe6tZUxNtiICvhMzCzLRVn9Ogw4qItkYdfwVWp1feFK+S/V6wh9shiOVNDCG7PhQsxAbi8PibBmdlB3Bp9I46Edg/yazTaKh2CH0OhaCM47kB4ghJ/zkGplCnTgYm6lT1sAIU4N+1fdgaYZq//yxLVdhIiYP8lE8D+f63j6yOMwWS4/M2I0SkKt2osZOZe6GJ7Dne6B9qvKQmqu+GCsnWl/PhLFBtXneKnnQaO1J/CodivKmzkVIvsUirwm5rFBk2kDKiqhjT61ugKMYIWG1G/h24SxzEPMQ3o8YyDvRuh296r/UvDGreWqSNnaTLxxwyYiaDh5ZsA/djLp/DvS8QNBcP7eP3TZ2dprKBzGSDMOEyAXHlTVzZat97puIaXvTQWjFqkU5uzKFee3fBXrFCh7TyuACp6gGJnF9LJRAYNoD8apf/dRny5+6uFZA2z99z+sf1H3H1Zds0G0A//lv3fYwJ1PdJLI13kiyU0jbj8QDg8b/4jMt7jBfhqhYv4o2zIjuv/Qu/L/78ESQLftoiphDlqgbMie/2FaKG9m1SnHgu56ZNOW8yTYtilM++R71I7yg0OCm+nE1SG50aNmLC/orxhucK6gk8G48C4lA6u2WUpaW3zsBIp/Ss0Jwn6kILiiFIPBTMYPp6fhJMkvuOovphExJkFyom3ok4X8edeSEVxFPNftTPCGb9hVG/cwG8k9bLxJlLsfNcTSxWUjisJ9Z7m2vc5EYkjc8OlcDvjr6dqcOqNp+WiH3bLnm3z2uu2wErFpN9c6872KYDFRNIjYs8ZGwIQz64thu5g/yWDF8Rq0bHKbGtZUtfEksnNAO++xjc1qMlJctdT6x9FH2ChNwM5+8MKS1e6b+EX+u9zp0/cO5kJZRWK8CPYu5ly119tQmSwr2woQ0lRyH4oUztNsqLwLqIqXHahJBl4xzezADSzexd+BLr4M48lb45uZFKr4ck8erB2Z5JtNTIMzUaWwBH67PgN4gKnvS22lW/qpX/6yc1yLSqE7RpX0zqvLLl3Xq/nQlSRGeZu+wLIeEbalHjLy2A3ufzKmSw47qSugyrJQwP/QpzF3bNQOnXWOlqsVgPVHF8lFZhfiqjroxh/To42nuDw8ts4BHkwYfSIImLudm6kAlZVq8DTLSyPf1X1LNiHrzeysjY1+5NpClozFBqR6hMv2JcvjuChIYsFxF01JmWTKmiivpvPxdvt7x44VUM7LIkYfwShy2gvLPEH/Ygw3tJhrnjFdzBHE2aqhhTJZiEkmeCEuqC0n5fFr5Ay9Hu5p3d28YOPqYC22ufCOidr2IfcVf/1ZrL3MMW041Os3yGaPmtO8Xh22k0HNuOywQsT+JD6bu2qR55MJWYCH2OK/2F/XY7bt6tuobJrXRxf1ZrfhKOh6bnbn5y1Gw980CVAHagv94enmenhws1aQbixdn9uF72nWPV0gjloBQZSnsOU7yVKcE0uw4uCxgPayeSGwIXwREA5ln32Gu5dVQNTzX4E7oDDrzjRrD5JqCrrx6bv7065sjmm+6RKoxa6g7H9EONVROEKBl6LTC5EHz35u4/XPk4rwpGfZYl60L2UKIKB2dx7UEIKfM9NuNpML88ipt3FtmR9+5r1KkLDyLcvgdzBRt2bsQX/qBdfbR7EvqH/B+AUenTgxqaJ0puScX+Z0ogEz/l6t1XS0WgZsUJeB0FZFtz+8qYPkQyMWbmyawtjIfMiffVxvn/DuTb5dDuDTHo7w/F35U2iAYdUr0ydLpbC2yl4LeRAipoAz00+6vXXUT1DlYOyhaUC7dje8/exNS+C+myBlVTL9DNgnnCS3Q30GnuTSE0mOm3uv/42ECPERotYkrusuCJ5YKV6TQP1srJwr4/7CN9dRAVdQp05QN24J9zBqIZdul43d+cd6/ig+dppfFt9JV6VfWKz/OajOh1OtigfPN7ljAtl5j3ULnsh8WbD/96900oCpTrR9DSetoYg5Vrw2xYo0QikGUWxa6VQ9RLwib5WJNKulvy4DbjKioLjVzuFkVghVSEF90M0wS1/GKzM0i7I36rgjGGYhOpfF4IzOtCA9/zT/t7X0KbHVBJ6z70Ys3+/JRcDFMljn8UDxS8qnAdFPmS9kMq95Tb6wgt3tG1fE++sqtQ71Fem6M4K+cOk6UG7Kol/iz0JjcpaU5XSjwx7awZRabbzvkHjEU+0tp266+Ed/PuU0TUo031OdtDC402Igts3TCLf2QQ+E+KqG0eW5S8jxGd8/ckUEjbSU8kVQMMtLEBpFe94XcYAc5k6zQjvoXFKHRjssMWBq7zYvXUymD0PSFaR15l9GtVW86tFtBNCruJxkpCbR8dHcxYgH92ISXNejt+nk2QQlO9tNpxMK13oH3R0z5QlTBt01uKbuJcWMjwZOeOLY658y5bv7DB0ZCDoDdegHdJCkGp9d+DCUfbYj6l/hdLfNoTRe5YN78qU3w4SFtpNWI1owW2obVGhPKhIjn1/btSlM6c1Obyt97zwbNhkm+mh+rjV6iOQerSt+CJy1eT7WRpyKXT1IsxA5wHkbCJT5ZeYhm4fvOC5iIJwgHouqg/75ncy9DpuzNHm02LeJ/ytJySo+FxZ0HtoOk4WsZS0gz3GjKsD3MWzxmnNd59dbfOLbx9QdvkCrshfzZ1aHrvhes4Ap7bb/Jl7/QQN6O3m4vI4jV/TT9qokvdh6sJ6mKWtSVVg00W2qYasJuwIH21QUj/AWbZ2eiPAjpl/uPoFcXNBLqqA7cFaB2ni3SI1lTb1asuSN3LSG0S+Fi8GPyF/K6leDmwfqu23jNyBHGNiF66d6KfkD4rpxCidVH1kfeWKCNKNfXywm43fspRsWScnRYI0pG3x3sbENPMabUykpOLrQVXP9UD0RG6pDO8mrN3Zb+1Z9j3mOdrHwEpM6sgCafgT88x1+dNLquo2vmJGBODxaOvlgeWj1O8rEcok0WGRUxkmx99+YFo0/9PIkaK5/rfVf6d4nGc9nOwx/tDUTl44GfgtrxIpJn+f0SmobhuZA+6mCAeOtPGjT7numeBkL6xRMmJKzCCEHFqrdt46iThq/GT2x6z1tRcn2ZbyRddD5mm+2v6DHsgN+35fZxzczAi4j+lcD0upzBQGo/kLnVVM40LwSJnTbIFn4jLzinuE3ZIv03VUe+LoZOWyHnUIaDTo1Pc26re6CCz2WODafIBZ2iBTC+iZ0ImfR2tqpOIc0/oSYA1/fW2Zj8dOAVlvaNfpQK3vWsaEbjfH2wfWY7es6ZSeF1tK2OcKQgd496t246aydUnewm7G5ONjiIrrqx1LdICarDKn/EM9p+YLmSmZQCdGxIf45hgmETxGcg+MbGp1qwnzbBAquZObtreuWeSF1TLovpzazXKe0xMW3OySERBf+lkEQw6xKuMzv+7GB2KMwzxbxeEUf9h22DYHMjvKxkJAjil6iEFwKv9KZ7SYQulZJAcIb9Wq7x9avT84r24ebj69XqGs/a1jesk12kBdR97sGb09sx09LhHtdKgegnGWNyLuoJUzuk0qfdJXhgmtXYcJSjC2ZKDNnZTpE6rWKhCMbmtDQoODBgm54NYU3DHKCYdvWth/ol1l8M7BvZH61yot5n4xh+Y1Oo74lG5k4c3kv8zIrEA8S1BrTXjg4okqIImAtRUSIMjaUSix1PMik1jimyudlvQs2C04rVswaVBDl2St6utTVo2QtrjHlD12pLcleZBysGSVIEPhhC6PLh3h2BerCSUUYmP67mirRXrz4IC6G5eiVqtL6qcqSBprr1h1SmS7JYp7waGBkEasR3PDJDB+C9zEggqGFWMxl5Vbvmf+4+5+QQqyAZFVu/b6Bq1UHPRQA4+gYexKZgI9gImthglR9MIPkLOC4fGF2LMapYz9RpZxCaGIFNfqYDBSnF5WnO5aVoUik7vforV3DU22itWL5dPKpJ9IfJSbHkkyb22d4x94/uz0iIWdSj2AlFCaUmUa5qEvZGVgv+5zCEwL7R/+WduHe2L0NhCoqUfL12Y+X/OzSLb+za/9p0CSSmQAu6KQzIAhTmtmeAiiFJO04wEd6+txlqbsKUePVzsj3P9AKEl9fsiYgfvuH8l5+Uzs81vNA6vRcuC3NCqj9XaRmdQfyNy6vmOGzbzCLBTh9e6Yh3drG1kT9WBTO/mYq+boQ7I12wsmLefDkafke7oahuxMY2PShhlkWq0hW8Q7mQ93ROn+OESKOS8xuTqHkorKryu1Y8yQ0ID0rm2yksLcalpHV3qsJ9Vfm0MMtGQ+FTywpR483ibeNCMbHeJq/hJmxY7IDWv3apmuXbW4MyIFGAU5oP84XvYewqbf+efRPkV1m1LPOiDMGA9TyAD0NjjYwyyYjj1VohbqnFzbugklbt5pBx5VSMsYk4QgYg1LpW5DGqyvSeGJkF/ku8PdMpQ7eQQr3xtpcdEwa4UibPxO7sMB4oZ9P3z5DDS5Fq/tSHBouk+9kyzIL4F1prathNtpWzJ8bZgbpCETMPWsnoV5rq7XNn0x0bPT3mgB9HR5ONVgebLOBpEPdlUQdE3mDVyl09NhJUCNfjPkR0wuCn9PhQd6Li/PpCjEO2HZwONN9i6i91Dmp9NoYDzyy5PN6o2pMQ8SUbZhJV6hTfrLdLLzwFXP6JVT3MqvtOcGsNCpMPefuakj5HnPC7/fwvBgm0LFlEhfqqLT9XOTQJCMwkvbKCMnx55QEcuQ2IMWMDtL/4hnX7kuFYryhO6CuRoivRwob1K3WKKlZ8+zwx4xJifdTz1hq4xjaA/zAjZ9Lx0egtqlil0f9qMK90x5CaF29SyierNu/4SHD/qCeJhjufj/WdGjfHGy6auFoDVHo5GY6UWquq7eSsSuEL5mUlRAKcwzSceQWkN6e5UMb2U4+TnSA/o+X94J592pom+4Kj7AE8qvdfJC0j6m9gGeMJNArvkdifZfzqCydb70wPM44VIH2MuXjG2hup16mudWNST52Yr1LeXBtptwjMAPlt6Ig/10McdAZtmhEUyWn4Q1NjpWcetuEaKWPMGwtkWjmPJTF47TGH0nds1qicQkugc6R4aJij/vXQZv8WEfVdZSHx7zqB6rXlzCjCAJj8Q8EV525GvxBAjaIMVqJzFELy4s6vJk9mm0b1lwyZXVj7Q4NilzrQNCQKkVqFIwoZG0hao6ggZlsteMTAsC6Ac8RRfQhyQrR7KbNw7yu0REz0ewpp9T4v36vTwOC5hASQev3C7JwdKChyJgBPghooUa44HFOWa4Rx/HSAtCkxHTyE9Y7wjmWEc3WxFjeLXGjsDUkf5LAH3RLYauYhqsazW/gvz+lmOs/y3WHYeqwKnRnsCE/6pStEh6U2gojmcST/+rUpI1K8X3+BWzSjH12/kyt81xVO/afqieEnqPXf0WBioe0sdItJREImQX5Ukig6jJJ6qXXahJqEhT/15mYqxPah1x9SAWS0MWtomOr9nbVYl/gffm9pBW9VoW0FOKs8hUvAxMJ/TXUbfu7JVKG7eV9mYxK2oYxO61kk/BZIu/9eEaTabptIX9YkQ8tOyeSYZQs7tJ3BxHbDpWkHa39H1CmTjbt6jio76Zg7/YsBSYLyuP26vKj35+w24sHKw0rFAxRUyRaCrLeV9JAymSxqmpo+uKMATg7nygcYAR0RvbnxVbEcF41EQdvX7BgfkpY/4kvhbaXJUfv8yvznE1OkXqDbtGWlmqCe0vYbOBgTe0kMU3COSPEV3ZsV3bz6KCj+23fcjzJOPDEtHu9Ao9lOUqAdjPUTRNiy57KsoXuascHADSbc7SnPYgo3X0NEGC4zDJ0edX6NxktU5m3VIpginSldC2WA7/f3afWcjn/IAKT+00CBz+/4PnITsgJxXfOB2yEb9gRpO7NTL9pG8eLohtsS+CsoMZMl1Kv9xU4kNESCqqYhm2rdEww4xRALhBCuDxtiLgE601aoKJDGw2BYUrL2uovM8n9jCSyJ6zpvrGLFDX2AqZbytmFIDWIZZlnr463EDNh0V5Jy+OBrcL3TCjpShGkellcjzpcDv2/7n1B0ZciinxfvsyJvluW84sPxpIYaL1G9918i9ziYybLzd71RiQZE/oyhPL1UVl5Fg1Fs+Pxcx/XrFkzdSUSxkKZPtbyu+vaFN5RIA1BHxQTC68eOCPSCNglw00kDkS68nByFg9ygvg9Tu19miY/yjthyGrhIw6S8kiMCfvT1SnEXDQ9C93Q52P9BasU7WNVZoEUHz+l4EVujeE7XwFP7QNNxo3ClF7U03LePLhByGVRah/80em4zUqt4WZl/g6ff7uNsWdH7Aqd1BKsWnTSv5SfNaTSoY8EQbgNNBnllYlI0CuE1oKsbCY6cgfBHu2J9Lcz+ALbJNzeFDPOcXHMy6FQKogO71yUsuWfv8iM3tb2sJrxOFy9AfzI6CreXOzs92+CUKl5rSEY/O4paOGuaHF2P4T93DPvQ3doyhm3A03apLEZguwynaVJEb6ZUBduieH+PGl4D7HHEYTfMQLjGpahW2TqKe56XT6qM+8NfQBeSVHV/HpDhEq+v6VObemF+t6UBYt7nYLyBpTwWhcKru3qQ7mZCccsn5BZP7JjeIFuIx/NVLhdGt1ukx+ryKxHpIG3nrBubmlQL7ZlFYUwGkUseE/NUdwSBRCm8fQXnZ4uYUWdoURLWKI8C0T2aIE4Da1piZhJINGMe61Of3yeRJSh9i7DVuZiEjvwiqyolVbVV6l4+ePEYKi5hYY5BcvfZYh/zKHnHEb9pyFMpwz+cpYAL7DsxeieOg6rA+WlsR8xVAznOJhQje0NiF7x+BeLqSZXNh+5x5NwRffbF4E+cNERE2CptZpQSJpf8xLy5bG6e9agnYmFipvFQwL0Ne1aeP6b1RgvhN9f+WkkrIlsA36da+SZrc3TSf3wbZudvHmnym/LgH/HMYA9/yRH75wLXA5ZBwZOZr1Wrq4nsISjriQ5PFV9QGAVgMLGWa/eduQ/ndIMnRDX2xIWcr4ckPQf/7XibAZEIEsu2wqfplQUb/G+VGsP7/DuWnqofawzqijfZVfhrou3mJdZB49DlwHjvVj05wGJY5zulyXnYP8LsDfHYqy13JBqm1CgJ+GfyuNYt+NyKmD5uHKR080S5XQZCwgBttPJe3egfYuksAMIdXd2nH1S1861ji7uM1CLEvKtKi4u8HxQtJ9RlIGbZIkvXf94NFdP8iw+zLPLQd9OZU2+w/Hvdubog67q2jviefekREx7B1cbclnrkVdtXpi0Kp2veVxR1YvmduHATQEGwB+WV9Wz8eBdb/5hD2KmF/l7S1zRVQR/8ony73GnmQoCD/JkbetGUP3GcuAW8D6EIROLDXWI/febRZw84iHtr0sVcbltE+CZn/hW95vLOAJEWa1oUQox83qoa4GwX6206ocAXQpgpVjMx6BTnv5ZyQ0TsKBrGqThGuId1FhWrasRCM+NdWaGcoYtaBmNI8e/oYL63GyqQOSA2QnBfrG05lViFHVMguGd2iIhoARuqCOnp10fA0webOkX+IRSh2xFCU9CI/bXMZYgF/IvhjuE4uoWUUTZlk4WU+OWTfwHSF0gV6nuSL5n+fvXiR+TIZskP49ZKyAYlPiX8uJfgri8wfveyWFOHx98cK7udq6bgRNrB8nWbmjXI93xBbfwAfvheTLZTWhUcBmk45VyXTqklLjUzYqXyrhaHhCRVCBsqzdEFG9wideTwbEidlGuuRCyt6T//+m2ZutlZ8Wc/m9THtstkx3WZ4RKA6ftPH+ND4BWKd7PzAnj3XooOoKyI7ktXZWNIzKT++KXzxaHeLZFEU6yYv04CC/Dd4hdoXntaPCXSkI+IIiiMGJLgYqjaTAGdpWu+7InaYFTycNDYCEDbmBq6erHhvrY55AvjKm+Dqlv1+Om7/AaaB9L0Oz6MGSQywErwEYwX35HwzLWitXDS5REm9kGlmo8z3J9oQMLfCdtRSY2m/yRHvVxY59ekeVxIs8y4LsrGgn9FLJP7LlF8WnFoWCh86bsjcA3Wk2WZDuvBOGrVVWr2wytScqq3JMO/YcXk581c61uCQummCQMX1E8thfzypygaid6VpX0UHNpLickOGvcOcPl5zD270/P7yGsZ+ANt4VSt1bEV57c0wcQF16+ACWRH4Vcws3thPfXVN+XROeYy5PJuc7K7WLr7W2TFXj2Vcyzou9K7DkH+NaAyXco/XUiCYflzlFgMlZdjk8np7qlO9yE6DE6XroV5Txr/l7bBnEQlkaDqdhykNzr1DDEY8Rhkggg4JWANA72ii/npsxODvBxQJtgVZ9ALaofThvWwBrB8BaeGfFKMcfMqr28ub1K7BqagctY1YlMpbZbBfPAfTuEKEY+EJMIZ5AmWbZVC7qZTJsxixfnZ9s8bvTp5Ko+Oznup39Z6zWEYTts+6b4pu8lCcKfnEzjCQUn8dBIzrwn3Fg6ek46qqeU8z0FB5CKA1zdIeOTJmPFG81YGO4U72CVh3t84+DuwnPQl9185G82duBaB2Pf8nYXKvpQOYPVrA6WeXnCnFjPV7NRk2ePwT1RsyZw5v84DWMVMdTJbGKfq5w5/AzxtpwNQ4B2VbQCAFrmWZc90WfzCb8W3b3mL9z5a+o+l090mxHzLN/lECSqDiJSnqey+W6BhLs6kcopdbNBCmXo/lQwdy6VKAzzoCmWaN+QZtYZGzE8XSE4e5uf7hECHTNtt+WxUJUvVtQdK+xiqokTmk0q5TUW75E34OHVk94Z0W/+sQjPLHuKN66gDuqWP3hhGQx/wijYmLSNC86HeBzwZ+D3ElVQfB8Sz5Z/JFfhV3GeQMY6UlqQVoI0oSA/g2T+JRKHJDpCpZWKxvNazR5pu2ooqHtRt6PInQW1FXjShyWLQHBaOg0VGajO2NEOHoc7XWWNOLL7wTVRqP9TA8QX2/XaZx6LWygDfAkWIlhmrXJRornMYPpOHYukWJDAOh8BpwjDojYn4sIGaEvgkbo/mYR6JVf+ocqkZcMFwdTdILD+2NKshKpvEr3KY8Nj8O6+9SpQiDIG7/AgaYC9PErGg+u2ZlpvPdDJjA8CeC0wWXHUwfDdRvjaWkEK+Tu1+4aO/jTX+suSWHj4Cdtk50AlgG9jUX1FixwnCX3APLGXgwEdVqbmhXPXDOdujFfUgEkm320shY8EjVKF0aksGxLafdyYx99XvtdV+IPC3dxGRRCZBO5m7vFEn9fSMr4M3w3AMFplHsJPtzv8MF+EbqE2SrJYuaOxr+KgGG1rXIjTyV5xllOOfG7EsiqltcLvyi3zgtO4mv7n8qHFHAzSWNd2xth+aQcurzIcQbhR7H+2PGrYHHOpl4BI4I95sNQbXBKqwhQpjGoVSZqGdrwL0+2jgv4sSWIi/2QH3dhxcmn7GlYwRt7Jppwimx+rqvE0MfOxN5uCiIevwlS42ZGNADPhwwKX/OtIhCQu28FNgGaiS1261FeAVs97zJLwOHhl49xPUmmLz3JzMznvqhnvtIIKB4Kg9QtM4l+TXQ/YQxWGgCOWIrWzI6iK1evs0tkqjowdGkD/r02W2hCJvTRAyRWcC4zaToAEmzNrycRi/Hl8KT6BiQw3PNRacXosU2M8GnvG8rSBocQXpD7K8GdLkERELaUxpsVYEHrPwzRq6chEjwNo5SHXeSGIOUt/dlmCLFHjJt/w+wc+CHTSpHcxOJcUxL9aw7uoOfZwAOOE6NoZ9oVaokuLMBpDm7vo9pVYjTPBUbQD9tEoGTs84P2nCnE7Nllb5lFWGsrRYZ0b4pK2sPVq1QIJvO24CwjBNGykB/2jkjicsgMNb5Y2RNKc5UuTX0YFZ/QI0IA7BKTnTFfiTYznboqPJtCF5/iH5UHSaj3I2TrEBCgjSFUymhu5yjMSu8Y304XC/9KU/sUOr4J7pFpLddWwsF8om2KHjFL1jie8Ug65a2n/FsEM6YYfTVYsXjxxu6wiU7X5RuoIJwINutDaLb6LSBy+eI8orL6/jvYMZjZG5qkvibsKM4DFvUvtt12wV39IvMQzbRLFQz6lejKIAs9muLlum46hdSk35eNAcg2q1G4CZXCz6UZAEa8QObWfoCxX+hzZ+7CSRGsh/5VIub4JQgcYI+FSGJGkrQdmCPDR6G/xAZqvmWHlKiVamGAm7ksuelOKoj4IJJDduMXMRSqrnUNc0/o4J0MQdvyVs0Cfg2pMel5K1pq87nlOnJtNT4OwKPebIxzbtZu0W/UeIRjcLkeHs05MUcHi4KTuLDtkQG4oops4Fu85B9kqm2tX0sm76DuXHVqRdCL/KuxllSGkGjCMf+f0n/xKBgXlhJnT5KMlo6TE5IGdLLMDSZMca7HrtTHuUcQKich5oHSZLegk1nO5E/De5ANdjUhUqJ9tCaC4XuGsGIUTYDA9BfIaA9nz+2UcffczZOcv2Q+fEpsv2I3/dL1/OjLzDMiiv0052I4PAjd5CJvji0pEBALYN0isu/r858Sp15CGbVnmNcUsxp16XIZd/0KBI8OUdKn0SQQi3yMUqVMRLsBn+lF/2bcTTQI53Jxe8ya2nPKKaRaQ3VXTS4Lk5o6LBCAdcN6UCianzSIjDwefMFNscy0U+c8d9OS7A8fVuNzaW0S2N4b61Gd+1k33hTypvzBZFofKq3VqAOyLLdUdN2aY6TngLz6PxYLkri9miNaz6jyEXyZLUl/keCAYpdxbcOxxLNLc6NOz4TgLUICRSyxKCHNIXha4tjLUNiYWg/kr+NjpORv8tiMArk1n2uOcTgkJMo17NIyDVfO5pB0BWEgSJ/yCHuaR9OKWg/kDDX+sGUiuHPs0jI0QAAYaJAx4IdQPlb28eJkdheoc7f0FkaiQv6NYt9e/ihrM/XPJneUMSva736KjwGkbr2NuI2W5ONvScAL6v5lYWcQB39BiPbWPuzqSSRrPARwyGZeh6SpXrO9RSAvJWaRxqYvil6JxhUSgMjdZ08EOp3ywMjZJx6inUyddRy6nAA/wNXSudnMV20dQMax2Odtr8GU7YmX2pfKs+Knm5+N6tHlHI7iN52D3QOksSN9XPeZXcSt7dN1TNlwXJnsjMjK7DHiC9ppbM7FqNjTsVaX7xcsoNU3WG5GXr58eNd2FRT13sFnA+JASmlwarFuZj5nl8NPkSDhX4RMIiRs2HnGDVrL18DBg+/whnzFGoqkkGzrkO/bUHmlYbk6uyW5rWZvylPmyjm3KsGjsi9Vc7ZxgVjlwKUrVXXSxNoUVkQN6wpsJvbKeo2xA5ONgaATebahgonOEx3r0k1ZoZES29aDs6rwM9v7FL18XJD6RYegmtlx92HeK+L0veZ0KjGhxbNj5bv7wrGBqCXG8ifs2Kjr9UOwLpx/4Sc3RXjDzg4VetclG8bWFcpRzlf5pHFnOdNh5qquC17ouskifEMga5EJ+D9AnVgtPnQqZuKNb9fjJaCyMKXT7+lPYNrVGR+KvGy3RH76v0AFew9ORmAnshNFCc/GO+lStpZN1MBTtWIzbOsckvhBkG7QnAalWmB+qHTBjnan/HIy28dq6TjJ9SsKTmCdoj2oq91sNy7x1UU6z/5zhXVmzkf81ycHfVVzOobagNpveQyRo6uWbYs9A1SA1me10/DRZsUYr8kbE+Lq5HMWohkOYlPCHlj6YjiFw/p4nuag0Fha4EQsT3JuNhaUl84BORzaIRarJh8Ki27FJ0SBMaVxEJol5c2WxYVdN0tyyLrO3wZZo6mRBxNxIwMjAVSq9F7UhgRZf6IvbFPWJl98KQI0wA8fd2jhXiopyYGxlMsFmBf9q1GW3VYe2TMY+rI89qCqQw18MAQsM0oqsOxJFCRHpNzctqIwVqsVy+5deypU0V+W7jcT/dLjglE6NKF03mTm+0SE5nJoxK+wTh9blP42wlWYQcQpCdoIkyCqHNBWMf7swc+W6GliDoQ9tsM+FDmRwAOQmqFsi3ijc1vpvlLm5irSqRMbHrnVSLKDRc8Uxpa/cSyLqUXWJTC1TguPynOMsjfMenXS2mlptII8AVeC9+sGZWgW18y+IBBokvTADvYB2yQB0otuK1+hjHYDKJPjhZZZXJ6fP9IvjufjYvbo9PUpIFQrB25fSb3z2pzxVX90qjZiBVgwoGQRUkQecRqul5HHuvl9QzJoMP7/kXgMHpR2sU3jusO6mZdBlFW3GbcS+LjG9KkbNCIWah/DcpSVn+TsCvue6TbqREk+2drzvhpxuysPRC9j5g7hkxIU+lQ+irO8xaXNKoKRUxyVGKLE2EUdeSUh6o01imHiA5cboRZ06eZP5jyu3y1vESbCP37rVIPxyNpp2NPFjnGC10yQlr7KIihqwrn/tRyUmq3SACQkarnuFZxwVqFmVH7extV0ceQU9NI/4OdkTkvoGYLT/KesmETwjjHtcGbpLl7dx7WBDcUACsF4WzfmDP7IBDvHzmpfC11HONuDeBfci64tvX5X0GotTcIGcufCQlBRYtJlrftD0+J7+JzrWyuIrb1uf+uPu82nNidhL4DtvbSmWoM9+7QsjUJgSYI6FHtQgvg+QwQlB24YyL+aVs07QLlC++uw9QUOgAl/Y91jt64aw1dBM4y5fA+qN/jLBVKBiwHnLrTBemeDkd8rhw3/vxSe+TvQpQaGGBeYXoMSX49903ZiS71jMipgMjM9nkKm+pMhIx7zGSvxFv/LXJ+arEo7m3E+C2qwOMt6ZUj0SCIB/tEEUdmKGhO6UUSQssEAvP6VO8SSPH1Ipnwg955vyJDKpUISHJj2+wmbaPGEzCKJv8hp/Dm3tTr1lZ42Q67lODrwHD9X4x7QLnv+AP7bCs527uBkOa3tpDfyJdHoXFXAsHP1geY+xkwC7UW2lsLN1Gx4LkRzgJijgFBuNeWbuCcXe8qOhRY1Mz9iVtnAIPcR9okalXMaYmXSr3ZQqRGmF1bZJFJi4+QMTbHyOvKsmHC+wnhjOTjnPxywcXub6r07gSjVPxotufUaWpPLH7HZJT7UPIIUnwmKZF9NTRVOFteul/OklF3Vu8+/EpGSYxK19lzv4Nv8wRUEeZlH/O2zXoOfb1WHlht3o3hdysD0rwK2MZ5GUr1O19zRreH6AICy7cwPwmB0Q3KphC+v0t1yAohW2HqYaPYIAravWKVkyMty+TyAxeAteWJ8ggwnI8RUh2U7nRizkcK+l3CM+mv9Xz/1YznN2xTcrbwTKGXevTLoPavr8E4+Vi1nkviThss4IT9skKfZAx6k2nRWbObdaOhH4bvJAPUkdqnCdgKw6dAP4jQZTIIX5YZvuxliof9Fl0oVI58BZVPuRBNAUOUQ1hAmMJ1VZfZCOPMfFZDSWWku4GtOF/rYY3ZRETkcHjZEbcNS+0YetLd0UZYDwy/1xofdawZ1Vfel97n3rCX2H5UiAY7ifIZCmOlbiwK34m3WdRkB6rYprFLYsm459AqX7GBHS/9oMrKZ4VZidcAKgLQSHTWHLxgYeheKaWTnMfXlY+zG96E4h/OnFhGeRl+pjR3wrvxhOtXh+K5NYmuPjv+D/SmqTkXQSX937jfhUjQfQs65vbgeKbn7bWSc63r8G401KZ9p9BPZYN8e1vIxYz60l/QU9sbP1NjqDuGvv91g0OY/VC3XHAECPm1z+gTgyEVUE+iSAp7hA7Q+pVVw4Vnnp2n6u9Y6Yg164u8tmzB3o5yOG/AOyF9t5S3JkWoOHf/EpLQ/X3AFioNNHDOJrfIvfJ6sKYQH/LDoQe1S3fclc/mRp6u1mRQ+H2NnPfOnfffvGYcGPoBoa3xj898teMsbY0zwRhboCZgRCpsUf45t4Pyz1QB9RiJZ3yR1prF9cutmriY7Gwk57hzkZfjC8kDfYXeNvdzr0mmj5/7D6j0I6B5j5U8eX/k0E4FKtMZ288kxijYYury93rKwCHrQkR2ELoPDdP46/231VD3+WgUF5c8D4ioto3dVOqvxKqjGheOZv7cmAJHTqb++4rorz1h5rVvMIHsVkaqF9AsDJ0jBuJn//F+mzA8Yvr0WLM6VF61xe4ZVP8p1sNMMLywZwuJEqHU8aYswbeDlos0Lr5vBqZd1IS6VQhBEeoVp2p4OweE5fZj2f/M71MYErc0j9pWDtdXuBq8dPhIRTSJRyXFNk0kbptnqAQI6D4lsGzP8lOJn9GbwgSdpBEU88v16pW+tGfZTe1vDG7qNOwa7a3ZO385BLHzVOVeqZu0F/kaZOxDS5yj9G1uhypgzEwa5fdxNjPWGHl9fzl4BCivME4CQH5T6yGdzeH3yb3R4Qs1xPJyiyhDjGH5/RkBACEwZBbGH/RW5kFzqkgAzoC2N8OGlOeGfJomZNqzI7eJd7Ikog6RxjdIDmFbFPgYLi/9ZeIV6A7MRtW8wSZl9MYgsnKBeXu0r8VUqG5P/vmJQzgAdpRNfYtEvCWM+QzGlq04WbnzC0ltVkS3T+rv5/ZpLXvJG2R0upD2iazAaWE7yoUqJhwvJS+SULJqXkrs0Ct6431Tz0Ly8jOF4jzpnbm57j9cPIjqDIus8LCuZJhKnBdNXq8imSiZjMV9U2GoMvrH+O7V5NPfq0bM3sdBO67oHvX9EaeEudot3crCNh0htHAOiaudr+eqmqObw+HHWubvCa/Ng3Gvg0kU7QAzbdNafeR+mRU4mGVDY/u0mUv1iyZd5WfJkTagIVLjhKNxUNlhc/8oMl3muCMf+VuFJnkTm0fJJzMXtbr0cga/mbYAcpi3jSx57GzZ9D2dcga6He2R6M7y+g9TJ4NcW0RJS+zVIn6Kwh4Rjg0l0NsSEApIJd707nXBlAn0yxTjJwBAjZBAmPw2deH/TyT1j4DbeagYUC4fiCtCRBAY8Shr3DTp4pIUTRpkNCbZPYONhLJh6NPagOZQIWPZuRCxw5EehkD1DlGi5hF0mLgf+EBijPSS1pNw1gEsZk0ML9TB5hZdqqbRomH9zn5caYT9+2v83uuwb4NsFUvud0GcbPUagQJ6HQvrasUq/Mw/ImHdzaerd5KINDnWYbhTWIrK/lSZKwB+xQ1bSY+Zw4SJllz22ZiIu8m/HTOX0NqaZdOJAVjMxqvx/qWEeVQLbF809JLM28R5inkNz1yyxN6WoEKpllLvRD4xREpQgqNsxxL5Bik+wjPCJqQAaCs/HkqVeVm8h352VLqOKpEAiEHy3Y3eC0pNZNVEb5nPsgpVlpgG/XLc+H9VXZXrYsTzXqZ1CTcfmTESdzrGtThesIu1nNv88wvZBtz3aOjOlHj9QYXZU2gWKyybl/VaO7jWqaesXa5olzS3eAtXKApql7YR56wuU3at5qs+Y7hlV2pWZYf5WO6zYWe1A/Klzm4sIvDWl+EsN/nuAhechcdKaEKZ6OfIuuPRUsU0LuZOz+xrX6v9tqu8vALRgTbpDjDxdypvadmeQz979donfbq4FVCe3hjegklakr6AW1WOa9X1bC6T65/pnjjJSB/aB3eP7nttPM+eSGbrveVvYppXl7EUYjScfCn3PnruP9rHSp3NB2+Jck44N/YFHD/PqgY1cxQxHR2RSfVEdGToTpbA+FYQt6abBbCgDAnExesTNDhpz7XrAzDFS1h58XAQ4NfEeA0Se1HLasmd3tzWdjqZhYaTtr/g0x0ZNmYYz8RwqX8zNgvx7jRny5oaqbvVxCRsgu0p86+rLXLstbRgVlKRKTXP9M/1zXug9AXWQEOr1KZMABB1xS/YeaXyFhBpHEP8Oi7352mVZiR6izVO+1afTHnKv15D0/bPmEJb869/XjL/r5TxoEx7b0Zbt7zmPFcW26mGzK0kC9YN8yrgmj2VZAYZgavRSobzzxtLOWnBiGUB4emDbJRMfBOH4aHMxaR55Z0Y2sCYJTwHbBewvqWyJSMEjtfuenIbNiA59rjQTpbYkAhCPkRNTQDxNRB9LwOkh27dcFX82S/s+5NqrKoLEhvcZaKjtzKXaQJAheV12GDpfuprFf4/NlYjE72YvLo9t4z94ctfnO0ydlP6g8rVicEm8ECjH7DGJlSIE8CUY8JiuhsMutX5nQps97wdzceJS0rYdTSIBqjUH6eXGUt5RGEv5WhYTBLzm4EZtbmkMjRFsOgFApyRfVyenx8MIVhdBfDXAar64qZbbXM/0MhSc9lRo/aetlEj5AnqigZM0ZV6Nckf9MvVyif82iFrIqo1WBePwGNr4d688z/v7Xr5mQjfkYGpL5MNmFdr6gAu1vpi6JS5DdOM6nf2ekntX8+lDbN2qvkoTVXRcXfY8qbCmd38A+CfBVcYTikHA/P+85Vu6Xn9mDQ/jTLkmCPxIdcikfjvNEAS68HK5Q2KZQY+YdsL4Rz2vuoxsnmSPS/fZ9RMJo1I5GaM7w9uV8Y/kC0mFkyup/uL9+GOh16ArqIP10yY8ACx72mfOuiWrIr2Fm6YK0fxr/p3C4r3y9Gl5MPHrDJtGXj/GZj5MAqTOISrQnb/e4d0tenQGf2HtjEKq4fFymsr2ooVnDw6Hdvfsnao8t/JTiYvSLwJQvYZu18MDyiqE/61xqW/llOvvLd6zsJ7rO+klakhDDIhenqghfVjoyXWd/34iDsZxRpBwpYlZLwK0f8o0npEE6Pk2uZprKZsmZLWHOefLeReiW4pUu/AKtdkpTw0Xt28uj3LaNprQAOfXOZ1kr1fQ2VyczK4jGv+3pqSznAltmtLGuhMLtvT391YWg4HP2mJEi1Ac9VeIevkhsRDmzpwjHQ5qCdgKloLrmA+I+kyA4YkhTZWWoicfHHX1/I+DxBXTaSNx9oIa0+XVTdHld8uN+VhZnOJFQW8Ttno9PuljMSgbVVNQzND/Lb4bL+HgiVEop0155DuPa3aJF33NR+Zyzm6LkVKCxdbUwkGzoUhmoHNt/R6QdpKk2ux/0vlJr+7gtuh9uCogjljjt0xEofDG5nZ1bVmgFvkCePOLxfa3oalPFI8fdkG+W3c9cFDmPtmZJS0N85pzpAH9OkHXHogJCahSeAzVysrfeu9Horfr72KGA8tg9r7XyEndk6yQ7aUyFJUtp2/OwsVQc7hVRfo0gpN2xKFOCowYN/aa5uhvgrw1+ll00zEijZS8SrrsBldy0oAjnaP0MWBornjXnCfpmL/SrK6THd4jUovTouPfNK4IjFYOMRExm/Nbi2Hm12BtbnSdXhNC0yF5uYQDVg2eZTmyTzwzEf/34CCeHbn5HnKIzH4yWd85y/NyiNljKLpcQgHEcgrGQyqjHQH1iIAmas7vTScmtvXawoIPxGaucIz+Lte0KXdb0Q0FwWw/2vAOwi07D6CiOFnsr+2II4ukaXAVEH+vxalJLiBZqJ3dJzEpQYsK7BiAlmn/jegP1+qTVR5ATFuRz5jlBukcmtzrdUwqRkzlr4if4t3To5D9aPT0FwJU4ak9u5j2d8yWi44cW4ftR63HYSfNvIJ5pBkl3xIaHJ0Vm2c43qx5DE0ls0QW4yEBw6nHbS0zfFe1gw6euk7EsvJOJrq0hIpoh9qOo4CpAjVcBE+wpjcwcweMlAmiuj1azr7SOd9HHw6HzSQOJGqwPb7BZbf/4CyqkmYRwwObAvgqEKRtD2sF/TdLkcTEwKiIHHApQuZUg7OPR6J14lw0hianIZg27A2YMuaiSlLGdxAyuZtCmjoLnlrstQJxLcNxvZNZtWFoVj+UiGzJ3tpVMJtOT0YrAgoOhM1QFPCVe0JUH3SGztOPWym4Xae7KHiikUfukb6hrbPqd8TyCOwMklLzBCdMMrCIXXt0LdfKOcMaohlIh76DIQHsiK1oEkmj/dhAxKKtjdKKsPJzw89sjuiqJAhUBuCOML4wwBDh636GGrxFKxIS5SMVMSUdecOWMtalHJJ+RDnX0LFInAaXArdD5hfVzFdn/lskYcACspnfeqo5YQMttUcEoltqXsbrK6PHwaMem5TpozxyxwBwk+GiKMqoEjyaVnIZC8nu/RvdsA8Lb4bp0yr2GHYSS/MKK75wBhFphwAYyCZIHvzvk3KShD10WvvGDAD/WKTTqWrLbRisfCRDLf3/1+qXctTvivVcA=
`pragma protect end_data_block
`pragma protect digest_block
b7dd82347172c1a69a31592f9a86d7914b2ec531f51124a36a43fef5013f7835
`pragma protect end_digest_block
`pragma protect end_protected
