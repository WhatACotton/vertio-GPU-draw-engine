`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
8WEExVKS92kSkgoR7l1UXxAPeUYc5Cj2jalqlFxgOLtwwwIz/CT8ZabMujepBG6Wk0Dp3TtJPXiVrQmcXNHwapJwOgOj7wJ+syGnDTbe1EFNTCBHBGv6KZDmqTyYuXRoLDzcMOQ8SORs+TjSx9GM4uyx9RfEOwdA6+qW4lcivBHpaT6WClQ8urVHsAHJAKhO4ZKpHZzmX/8neiAgdqpYa0ISyHbG7k0E+p3+3O1faSClzQsn1bTtRSxmElHJfAvormjoa9Rc/LOcm1hVmOAcbikcFJh20g5wF45bfezn37albDyxkdWIWSzgybf4DbpFz/ixLPnVL7MU6XQUPSFQCC3RnI8O/h/cxEV+crEDpt7sL/+YJrM/CUiToBjUqThm4wzfnSjql6CA8w9z83k1x9CIQb5vofye2nu3g53W7G3+u5Gx06eqK/VPVpFJoQfm3/7S3W+t8CEZ4xVRfIK3ffonRLSezaQRq2LWJjgpQEQv737DD1cgNNsUcE6ZzzJAhZJrust3jbsJGVU+oTyZbZW6H38ArjkaxoQ8sEXrzQJf4IU/XDFack9gqOkmm4xXG+9+EWXx3K4NlzaTqwh0OEDtXZ9UaI8Xc0mSaSnUERYdjIsnSQiWZ6tLs1QWGVUcVdKVD6K/svHEOK1VaVHfSDsaPnVVf/rF+uHT1b5SGMTN8vHzjgT0mWkOihIwWK867T1G/QEeIuhj2FeHkzJa2vN/KVTMDGuK1lxHHq5R3D0og7n6QeKec/equ5dhYOY2HU7kzvYMQ99dui2/6+y+IOSvpgznFWznjEKjwKyLtHHL+qbwQtHbI3NuJXP3DEQU6GqhVCIhMZ//qIHkV7BTsqhLc1jxGVoTbAvMcjzwSjx7rm/q5kNh5BU93E+qI8SVRJODPFPeX0xZkHmVfcTFR/l/qiPP+21LDxI+wmuxJhiBc8spEkY/Dk04Ocsg1kTyFi/Bix3xPNvFoHiI/7ME6s/WWxxvUc/iDMNzMdfRjtmYh80N3+6OkNmk7tLIekcW1xUe/Y3NQT6Q5Slp8jXYShWjqtGcrngkFZRnwFaae6J/kiXNDX0Lvo8HuDY90NFe3h311odP3uUP5OE/m5OnRiQxNCcrqKaAIHByZu4aG2Rm9ksJBSQ/PRIqqs9dsVdIGXVpPZ+xg1S+utQhkg192KeBp2TEpaU2VwJItOM90DllpMBTtMeLJpEX8RY/GZGfuXzAJ02Hs+XD9AnDdVfhQVhINg6uOToI4zJMPMwZjD2sMM471yjCJE8/05bGLAa9XnI7wJ3XHwAdgfxxyiGZPuAcT5RWFIDWc2jXgLSBRZWe6TdjlBChNwtaKDc8xF7ZIeuIv/gxbolUP/1IY5mE9JfjPENXqBWncNxI2LkDYG0b6OlfbK/82cuFRiKfYRJOO+u3Z+6t5ipV48YryNlyo2ipnUvgkpQiP8ZRmzXT8eHB+yFh68RYvksiX4PfieWXpI4iUPbqed4nGqjB/mmtFmJrSeTjLqyDeVHPHxQw7vVWsD/BO46ql1Ctv23oZfNHvAAkhaV87zmlkUWwe0qQBB8Gp3UcSNTDdI9Oy9115MhU9N/bpv5CdD7Kjohlby8LiqsDoLad5s394+l8+mOqSKZ2+4/4OWZ5i+YGN9vuHe3LtJXPy0TesIn5R5xFbyEMMb4r313p/4M/kyzXeBBfNk2f+90zHFAAxDsWayO9o1ylBOUoxDpVvAcH4RAE3XPb2GkK0R/2++CSCTkQIj1q26bcsXFs7RcpdMvZ34YR2jjhwFtzlxby4e6TQdVjwlCZOOQsBBgP0j0D+dnzqbqeeSaHmEPrUPSB5ShiNNxwz8o8k59k+OZIyQKAHuEg3z/QcbM7qisoqC5tB364wnuwMlSFXq94zdK4RBgbLyfE4lwMPaTROqIuqoXrjIqvHHbrMW2y49MrvpisEPq1ZDL3PyNOl1FMsAyiHZ/YUEAeEKljIOHg58kOyYDpkVqIYVvLdFcxLMNEO82Rn/LXIYXXBAVD6+e/rdhUoRur+4f9fp50wV0nUVEx7NazY1ZnOimxXy7zrfTb6MR3HcEhRzj4QAfJvX3z+3Coh0UixgvuqfgH2+p4YWp/pPiwrstzhgsMVEGHmAthopGVhLRset6jxTa/a5oyzZenpsske70Jxw2xVhfSjrFObDDx5O6mU97QOwzEwvF+oEh4z7Y/1SqnCoLdaUe3dYYV8z4wNpRWElcN5oir84ehGdQVwpaLrIif30x7BIsScYU738y2RPCxhEx8YJxzGN2LNnxyMAkNAe0hRkt1h9M5kWGegQYt5polKi6ncsT3wOen93QDlVa2ACrQzArmslPn53g4XELEtXB1KmWMZIlTSxbGZwP240Vmlxob3gaPPUfERNPN+gGGOoCpybDYbGXf9I1+W5SDHAN2zEKkikFXjC06FPRrv7Pl0lDMPPdki4fatiIHeBnvLvB4SklIAd17WhLVpb/UEO2iNHj9mOskhERIuXk6hVLk0+54xWPSmnWNaS/KGkbFBVX4EA/ceu1vAlejq0+YJZWRIbymOljZ5+gxQb2SoawEwwro2RqwzPhvkWaKu9o/XBrgSPewqVEm3enWsASw43fKDDfTZR4V3AbQzqnLG0KefaSEcMG8qaG3bQk1h0spkHf+lQ25B640rBtcc5TenWHTrv6aOlinqBphUcLr1VJ4iyv0A4+0YtedxC6lguTH5a1Lc+va+8QjqAlbkYewjisythFnLgkfHbx/CJiHDiB9HXHgvkxmit3xggpSj0dyAmox8YxhS/p3Ahk+PDEzNDPpMiTofo6668+loodc96veNr6NVuWfDIMSPuP2qbN4uM9mHurVMv59yC14fvhQnUzjRhkCLZ/baZR5nJg7RJYShibLW7g5Qk/FCQwBOuIxZacKYF/ks2pAJ/DqmM/70Af/lYAqy0njNqKawZ2Dk6XMi+BFSscPxRMws+4c4wyggU+HWtflraUtTCI3AR72WflCykyZrPrysCKY0iB8BWROpcB5XcpedraVEgXNqY6ffSZC7nPymBeHX8HLYsZqZsPHHMJCuPog3o1cjocwulP8dhvqpqI4MCGPTPb2V1x6XginT/Fksz/O6Gl29w3Mdc7CtodAhPKreHPw339keeE9cwQ6lvzGPaTE3ocoYujTMBW5YQCltSzmXhf8YGMnf9BSynfPtf69x8H7WB5uc2mm8fAV71sx+8wEX23lzFBJZuoa0vusITqk58JS6uDrFjRFFDZnqiHQA0oW2alUoewUpSH8joNyKhG+qZKi3eXOjpHtjSNKMUeX68CsHsBeCI8VFlR0XDudtLxgotqlx6Rzn5//BdfTJK3iZ1abtzV8WrqNKWkvSfEWFNMNRXzgu1jalYaEm/TJskIcHY0EeTmTuEVXVQGuAUvKQFTdTEwfco/ra+ktmMovuNZr7c/WL/B7gDUR5MP9HemFGa3qnumM6bQgFpxibsiaiwUltQT/wIXKzRrTtdo9Dt4N+qwAHCu2mBxJlpOddRdGU2SPpkN7x2ufc1FWLaM1hHfCMLStRxBmXSyplhKPr507jVqAbkISQOO2zhHIxsk2S+STLFK031PSiiYLuDoFoXOoUaKXBCAbaWBFZ6GLlSKpEtzVAQFu4US7o24RDwWgISzmIee9arjlG5GYkuIBAEpMmtULipULECLbGJXHCTPbjEE+rKzGHuCKuWPorsZ4P3phLg1861Xev+pXUDO0ELOdMRYCkOzx66MMsHdvZl0neuKvEghfAz0YscQXuWOn+G4pBVslmx0gcwCT/R58kDxUEtWBfyeNzJ19PuRiedlNf9bxPZ8Gyje8P3LnzwmqllmXM9FGxVszqqAv93RjaukklUXbtVlsAtqEKCSI6ItAfEV/f46issvU/BQx3G7bpjR9yK+UcuQxL0CmCYy/ba12BTlelVtgLqJWAzx1izyufXIX0QX8ifA/sDNALYKsn52LF3OSBgozBpom9PweuBNU7z1x6QsWsN8BfVtDHN2t5y17btp+ZWirqyfVKeolDFhnm4qK0z5u2gwtTP64yp3pER50vM8QFdy1qKRDIgRz3/iGP46OP/tj2mMu/0+PWm3mAr5H+WxjxvJGri8EA+AgDiQ89n7pht+6Jj7HfVDMbyeRwb/HsZg4dIdfIDhlxc58pettiSS4Lu+2JMhuvXIaVly8Y4qU4VX1cCSNm3/Z7sSJJtwl67WqLqje0eGHivrecsHDC24SPPYDxV4DruUyzB3pNqa0ClRqzfvUOta7c64eTIZYyTOjamHrU5k6zUczxhE7JYHWBO8ixzj391f86tTSfrS0+5NadUKj1A22CVS3IxzNa5tQSNrnluXJi0HIsYzRJxExQorHrBr7XjRrueaw82dAoX2IwX50yfivmOXvPTuutvcTVrXJp7nTWsrARyGObrtd/5HGs2/ICxQLW1UUf3o52hrzA51apO0i8RHifxybVL7zjsW7IWmR+YLGvVhwUdIbdGpYqRdaJgXIvnIgSKDoXMDE5Mi4RkzXdBqM9/oslPQCfyNyKUsJgAxqcrPVhbj/3qwDF7zn0bKrBYJOPb640IJjXXagKAO2k/N0LluuWJwvW03kdNGFjSJ2rERhfia1G+ndL7IBS/p9/gJeq5RbKGy4rbVhjfUrjvqMXYyAsKZd+wj58/+acySC7Euow//juWB6Idg+ps8FvXJtq9DMVcO4U+RcKvuVwpnKVS4q3b+JzyqaWsvBgap0h9EhwxkWXQRpL2t59oc8P67pr0mkGTTYYtwbRQRApivEIuz8miRS2gk7WkORIA0mhVUZC9bipMLTO5h+woo7aBRmm9r6kVB8qYT9JYrwm6sANif1lxaSGG18Gw9Oiu8l/6iaapDAcWFReoGqVqgvZYcsoo4Wq6n4emNR3FEG3LT9gHVAQ4IXhlnq5xTobTtkgi6pfwC1JWIPoMTA0mil0p1NMzfcsAgGYCbcC0fgEs8nDJp+UYwwaouqhPTXlq+ohoOXUkds8kvfbAHqGhbb4eOoMatwJO4OMgqgrMyGrBuB9/KvvltfuATQ1y6Ow/0OcnnIx75GJ1CIyIpMkg7Ymt54+owPmJEHMZ6R2I7G17S7pguPWWPlIZqlsczpciFbQ5fOZ2O5YdDqmSl3bsZ8SIdjJVHodkywjKUPHJ3myCIDkvXn24JOqHwFT2vf55+wd+ViyEooN8E0nTP3rlXpneZ62aPD3HOONum1Rxf+Sxj9RlNXImdnnnASGcG0C/K24nYdjRflfkxWAeuBL16s0lZZ6V6ZCT8r8QhBOy0sj86iRQa2cgZJDwALERhhk1qCFbGGWgWTYpELDEy0HaybbJaNZbJrical6n+/IZmJ7AghN6+31PhwxJBwyYg6FWwi65PtFDz4icOgG7u8ml14CsAcaQwwV7CQe0/nnBR0zL+v5qG3NU+bZw9nX8TAD2UahgQmD7xKFe/Wrs9DXtcOLVuuaHDpp2nPRQRvcx+tj4ORVoZFJLp+LheIlT8FMPiPVLlx23eaIZFbRu+r2au3+dlC5Cg4/9uP3jQbFFfDxC/QaRgaUO1SKnfZ4PXj24+uTa6exV0YOO2hlymvRhaYUEDltUTOKhwU6d2vZaWHyKximqVZ5QUDAN/X+dgenvdxU/xp2d3a+fDenMaQWm8Ffc8a1+fSKY2JWmy0cbOM2JAeVd5fL4YCWkQhaY5kk+Cm4mk9ifYHAEXzp2iIB6EE4W+M2Q1q3iYnERFpWYm+Y7rtohqmKhdCXgt3ZffNakwfE1TaIgLZriCimWWUXYQxi6CGBOsE2vJBfDWx/iQA85MgKosFwk2X7ozcSC6uR/EQWNnZgZdGKavPUferl5P4eH00ETEwfvGyd97uFn8zXUlSDCh73GEdtJdoN8qi7An7+FjAPT2xFcMR0Bd9fIwXtKSnNfNDks9HJMxIrVYp7J+2Gq3/xu75HcwBrTDW8W4ZDD6Ae5DN5KuokdnO/Iq6CXwAKaTrObKm0oefZlAx8ZUagSRuZVBi8jwRjj3MWbfOdU3YInve3Uq3SfY6ZfHcPH+16BbrNvvtZkMAKK31GFQ2CgQC9FDV3xeg0KahCcsX0IcHGVdzI0TnSOZKGirWnO+gU1Mbx1b7rj6ikP2HXBH3aPleUHw593KvB4iuxi6YHVDLoTnOdIoOo2CYtMziFh5/ubGLQ7EIdJVd1DSi0DWP0lu+yDAu//I7oDRHmdjpa+BA2ZVM+Mx1tTiMeiHSB+P5vhioacv7n2qtx6d0AkQ8Kw+hw5/zTxKom1lhTK/CAQOqhIwg9+lgdqv2UGi7f56TcdX10lSEb1bvLDQgG5MGcYpms6B+IZzKaRDh+BDRFaRFVfhvCNca5HCg0Ya/V0R9ddIhp9SdQJ1m6V5M2S2vuTXoGSdvtmSriPlDCs9+GthWRznP0nj9j0YLhtzb9wMbv4SlpObnuON35BWG8o8JJfLO5XIWYgosBTV+b6zVJMrMKlqGsfVCPtzyPbC22NtgYtX8a/B+B+cLo8GIheSutE1d8yglW3aOV/nkr39KuqcyX5Q5BRz2KcgGIBPqixcyesW31e7kQnXSM1eghGZ1ZFx8UQP+hKE4KeH/1eViBDAn/PNfw+UgL9WmHSButTXUSTHbdeq62tkPxFhZ6dqq1IM6VhJ0KncE38ZVmyE2m+JjT8DJe9lDleUEAxqE6MiS9On79qZDex3/e4UTymHggiV+IEynYu/eUQxgblA3SdEs/Lcsl2yNMnEtmXIojUM+uLsxtG/3s0SfBx5ll9SojLGG/pHK939oxs+gLxdIYHjt09rWz7GavzjKovwLJH7L5XVh1k2Q1IUH6pbB9ebuUhkSTJ7ypOown5z9oQoT19n/OC1u3pJBttsk79GotL4aTkhqx8zX1pC6LkKe82SKY9WcJUJ9x9fmPUpoZKdXvkSPSAeA+ybD07cNLt43eOyTEmVbjna+pH+x17o1mvU+j9aXjB566GzGdoyemjTtYde4MWWCFJKiU/FbRwIW/OaPiMKk6TMhAcy9lvagb9dZpfnbCETfisg2SJoD8ELIm9vzEEerwXewwhf9tAFAU9t6c283AwAMHTOrSxa8XI0pocxOD5y9rx6f5/9Y18ybXtkSdcGUHytqTZNLPlwkjjqs9tCUDw8uH+3gGKiQZMMt0aZPSR3NJU9153K5wg+mZBvq+Z1dedGSJbVIqPcC8km6eUC5bHivH5FO8We6JvJVR12hWyQITWCM2l8fJHZCFaJG+XCs+BnqbVHsVjZEYHw3fByzhTWicg8/i+1w6aWVhVIVP8tYJWUJaVIk0+MuR7UwBSdU/39DDqzdukz3mQ+E1NSIXs/yZyJSC3qvU0Q4JUAXYR0WaJ2qOF96/mPFUpJBti49wj/K8JNtI2c72x4KCAqyu6Hbpk+OaB/iN0kpc0c+HXq69qpXt2V5c5rT4b4Ya7dV446tsff58MDoOGIu6wtbFhQhCMX94GlOFsfLZ5xW9ArmoyW7gQ6yM6ubqse6iiHSKVdHA23Z0VrZG94icA0ffARk8LM2UymMhWwQy3Vn1w5SAZ94Q8voBNQ0m6/LcqxaWhyuhXK+qvfm5+fiV5aSSt3GQo/l4t55CCW15C23CmkDSNCPDifksYF9RYQLPFiZd1k4KJUkSnJtWcVWLuSn8Jv0mDDllWq0NpvPfaZrmMYLJdSIWoUeQ8ii5b72j4pG0oadU3D5H/M/zsH6LcAGjOoqy/F0JevbBL40K2/6je3fwYdddyOHCvhjFqR+jju4fN8L4WcQ03MFVuRsndIhYV+x1OQNE266c49+O2I19VYzo/AAOKHPOrzppMvRrviyxtebqFS/A6g6uwQuqJHLsLvzya0DVVZHk5bpoI6WYySWM13nm80f/F+sJ9I/4Oa/4gxo+o4z0r6vYVyu7KUOdJFYGLAriqXiekojq78cGxccXQozQ6QclcFmpbw0lzz9owNA77pNMeDJ5DzqUZtdT7peJ6iN633yoLiAVPRxF2WZQVCAys5IH6WDWJN6d8bx/pJElQn1C28bl63LMgUTqjkOCoFq6cKxzYps5k9ZJvypSfaEtWIDiWbhl5uO92gQ2OgBaaVVB7Iz+f/DrSoQ9F9VPslJfRh2XOACDlOdGhOY7d1NykIQOKVTGT2fnNzRjdpHv7ZqQuoxh94J3eAB9euQp6/8Ks8Y625sD+gHX2nIZ6TDH8y4zfspUeh45a/AMnSW3SS5FByNvO2eEj4QcJMGClBmiZkKiQvJDLibLGbYhmjaY0HWxMQ+cuUYrQ+Rd2+sOoRFruQsBghi88TZ9gfL/HsQSTg7HWH0q7FBzA4AUYxecEa6BIT4oZMJFJA20Og7r7+vYlYpQ5cNlBZo/G+dKR7IEh1mvg0oXV01A9B06g/cXQWqlCPl7QwV1ay5i7J468F/LUxG9EmL05TRjePjUCOByjIfFspe3T3yJ36pzqq9N+k42mmypcc3QjPBc32XBxsHCowK3v228t1YONdGs6ac5f0gv/AXY+NoOQyxdzhxA2lGMEoP/BSvV1E+FcvP0EKYadxBuQWdb/3Zy60KLg/95MjIzSao12M4roSHrNpkPCuEEyQbcidUXfX3I0Ub9DmXiDNJMMOffvMuxZ5XIcIl4NFsI85NnLiHqTIJ8oC1w0dEnjP/8A86u1jfLa5eq/EMl/eK83bE0zf9QF0pqUDlqV5JQY7ZTdMLP3w+ujfWv1Jg+egKHQijmMIwuHFX+gZyU76bIn/gaF4gRVevEjIJbiJfGDrfIXrDpCahMQ5iRiNEXwQ2OMNif2AlTTA8VYqWCdvPqrDSTSusuqRIDdATnYDjMAqEiwDng5YC6IPIqQg7N3XojRT8/23vIP0j2iJUI45fjlLw598BKj5TsrGhU/5zROGhdadkvxGmr/xAuXkYHzKh/FaWJukhDIpyaKaXEfrfXoGY59GejM9LDvIDiJm/kUp2x11SRtxfFbN5rlDhKeqXagozLwqr2nMbAGwbSPe7aIxTdqc3fR/zT/L10ak2otOL8eh4NVN7KWGhfhwDKc5DkrTcSohGYoDP3SdBrDltKS66cBnqcvNN348t/YLovNbsElUxspVBZUq+9Htj7TgoSIgerWmBYSBy9UHpmlJrhkB/+heVWfV1rdcAEcjgXon+wA2xi76UbqmWV25N5RkDY6sP8dghX6oWaOVQj1IVGgpcieEQ5D/sEGdZv6hK5qXdwtec72G9aiiolgmRelvNyZLYYKR1aL09AkW1cgu4YXxpXRxo6tuM/F8541SJdUgQUDkkKoGuu2B++QF/6VmnuxlNp1RMJu8zHB2nFiP51qlJ6ROpsL87pPEUP6QueyKdIrBmW4SwddbhUsL+JtxJjstxN4Mqw6NLP7nHOeshBfZNH9Utvqs1fPSLuPuots5voJPrvhsTAAK3swl8LYYT8Pf+plZbq72mZaJ4k85sj/7bRrBtT7OQymiuxzaRI/Km+RhAgAUncQggT9gc9lYVSQJWDreEGTi/cZg/6LNc6VzQWmdEOfA5J50ywF3KtHcCANpow710i3XCyxfndGPGcvWCl14My9hyFsq4hVaFNBb+jeeCAJa+vh1yvTNhDu0Ib0/sJ6yT+GZHmFtkB5YYWZxcql13bNzszEdZEtLGnotN4HiJQjWfwceo2Hnwj8AFG1qYgw/l52WnBoYw8GJeMsAQKXzqfus0ooZaA5zJF/NzyHYuro3fUQIGg/lHqVta0SCrJffxuQsphf+ppWNZYggwjwJimaiISaLgtacWHem8lJXEplD1AAkg0K7b+6wgYKodby8veDiB4ULwNuDKihnNHv3YQz9IpV+ZfG3iVZ8jzPO/+/Ti/7p8Rxhs7ouZn9tQfIrVI+1vQ5LdyngsOnIJOj4Zs3k1VWh132Gj7ehCD4ECH8JeojHRsWGbcOuC4cP7AZgrXve7k2zdYcJMZ5m7LqARfOdjOmzEC+PO6Qto5LXgDpZL4OHW+d79/6N8DMQdUam/BeJccoM4v77s8PGembyweMFiEcgoe3mNSB/U94zPrhVeoo45WjsgmFhrtdwycVCp7Mlkqfcj8EoJACt7iP+lkEG9sQC6wqyU0m4lq/V9oc5P1HsWqneMQsIsTATLbVo41F2Js2A8mG5rXKBqfChfu9Ro+gzxYdWWr0hNGjUe2Hc8JygnfZ0ifJ47myjGw6lzwyjQoODhwkqnYpN4K7u6ovhVihBuP7qXV7dq2EyG/e3Z7HrH4leMQszR4eFCP+HeCneY+zpR8FkheUB2N+qoABLmIMpaYXs9Bp6xLgrc0OWO1KTHutBsZVbRb2gIBHcoS5nq7eKYKzO+/jcGiPM8vgit5z3oB38d4seOTZ7Nwwmhe03m+j9js5Y8nK8bEiOJy1hI/Z8cg2YjsgtUjGaLRZBctEDX6QRK8U0q2tIPjHhXJcpCa8at/EkEv788BhFr74sYb7ZnBttd77KjSQGwGDet48am0EAYEc8rfteS7tpQ5gd5y3QWIPOOofvkWe7sLc3hGPyGloIPWBFQbNuEAKL4NSEJG8BdK4bF6sab/KskexdkbayhsPLFxs5cBgUilRvdECOUBh0f32/jCJmvZ0La6gwg58eLTu2cuEXQ4n/HuJ1caUrOwhrPlVOWX/JWDoDrlWkhSFGRcjvgRBEtn/T32Xqh/E9YFvgZJA2TBrYQ7Cade1q2ie2aAFysttBUXQ8rSHs2lZfRU0EWZ1xCNlNGgH510J95rPeiS1E7dOiPIRPq7pWGwUXpuGiK5zX0d6GxHhrTN7CzJVgwUnRZyFQVRlGYdXP7wKJqTVXtYpxyUuEFR+m1teJ4KELIA5jlgS7AqKxO8a3OKx8+cQpF7dNeosouabGk8qQbbPBQRqGTbFxcdpYy8P4CymUF4L9Fe3nG/OEZngD1tJtB4UzLQWDXAv2JSeA2bTY2CZ8pGvQxdh3XHesHPIB9wuKNVVDKK+JfQJ3D8vZxeEyMbsrhUdt5BFT4aCa1OWYBgwFy91rZK9xO7tPGDagYjnxke3eidrsYXwzyvXlOXqy9HQX+wMoqNq/VGKBICbYPW+QDu/gKqra6x0z9JMRb/gKBEqO27HWdYEzfkhVOINV9W+qG4iHAV/iecKdOLMfBNzNRB+TD87D+FNCf9lWp1sU5ehblLadOKWQfIZBsjDauDpTZOW1NnIq99dpdgQ2P90QXWWLtmd1ri5bbcZPKS/m2/giuskzEiArGKs0ryapC5qVPRPUC/yzP7J7EjUtNha2+XK2Pv5rHgkzVkFcSZlZPiHNCBQ9a7Ygn6yhWkr6qORJtR9TMVuqDMezSr463OKGepivcafBzNExMc2vunzOv7E/+4MXzlV3QZdNECyVjdOzhg+JarwQYBiJusNn0h63xdBvKjVm2bbjX/+rTGXNPBW2i1pPNaF+v8Z7ih3nGFZx/SMMOKrlUExyymkBn7JZ5807SdUXfNeAi7ljwiR5BeQZMGcr7akcSoC5mLUy1dJVdqWRsM6sJgdsTsxdFruDHtJgVgEF0GMBZB6RzA1fsUHGzUUp+m3YT+g7vqRdO+IvATRGNUGoN36sdHsaCRCb8mOEUy1z+abeCLmkkEOWj3R1v3GSYA73Xz74C27ypjeEYVKqJAiCEbO+QDyTTmtPP2uhGdlwAaYuKYGLwOLZWllTRXevVwlh9rArhbk7jVbgTS+3u5pDMAt7wbU9LzRGym6YEXnTYIAVphcfmfxytvYmvfrgC6p9q8XtosZTF6MpmMVgWavv/mF2CWU2Uv4F7o64yhdgl0ZqatPA0LEGTFh5LlZJ+wz9EJ2RnKaq3E+S2uFW2LF2hZyTKHyZHUKUaeZBmNtjqgONur0/xjDzQtSbPxOigdHGkh/HVB4OgPUu/ystBohiPbc2mktl6wf8s04gTsJd08AW9Hl5HQ/P4G60+S3o5StCAg6n0pW02NlPYAqgYlHxAyLxWqCn/L9wXaRlQgOUsQFguRRoBvmWhUjpcx0hoFdp9KnFrNeihZiD+JrVnoKHCS1ml4i1YlCijCWxjCdIja7Il8GRp4jvO10SENx42KHSOFjlanzCbTZtowsngLWx8ttkzxQ/QIc+saRzvtl4pxLVrZmvdECrNm5uH348vgJHy6z5Nosqrl/95+xgoskQDhkjU3CCPw7VTeRc0ZALj+2ci7Uxl6AnXItF+5QZxPJunLu9ht22+zxITaRCgwrAsRjfr0jJ9WTQ14+cIKahAepD7wGIp8p+fLQSJRE4ZSExPxXoRMUhcOvBoySF/bvRG8jVA9yUOFmGPlgZBgA8hfFSCyB7QbfpDEYAo0ail1keGKYMLZ7cmnKuZLBz1eDKBukVfHOU5ziNQkTykFKl+CLGhyIjANrN7POrn3o2qA9y7Qjze/OaRrlMcdIxfUqK6ujBBEloBgwdtKV4ryU8vDRtuskHDtUjKuur1ygKChRjgNLPLUntKVfYxQSFaal7znuoUL+8G3djojy7Fgy7ijqJPA4oB8GNVfOfGscTsB4/xnOv7me/QLfGsGS0kCYtw5VurPuCQo6fiGQh4A2CQ9jVXSBRXF4BwSUqOFgg3AOM/rmooTqTN1zhfDD6B3RPt9TWhhtAAZ63o/sJmb9c653ytjPBmGKOrbcUZM89lfx1bHe3aGKfLOP9TI6aClzf0J1SrwI9Jmj8GF2Mnzu+aPshjLJ562bDMnD+taIFVKpM5h5Mqr1jruAlZ5SIIIzxWXPzFT+iEEJfCnNgmVpzRTT8/owMhBXb8pidT5IgkKq8XmGmrVvZzwXF3vlOnb011hkTiS/Y2FJngBwXCaLReRohQVKAq3jmSyMnbwbhMFGJFKDsEoEwgl3sy9AB+AvM35VTQDbRFK054JSjkbcD0d7cc3Z5wMI5NqmQa7u7yCn+iHhBMp/4wBAErBZX0Ji9wCExhe8KzHPRNEn6kFAV/hfjlP8JDXqGGjgEVr2cm9Z0DmaNPgj8rHOR2cuJyowF8E0eia59/EMQn9w5R5oXOJnYSTX38gch6K8HbPsTYSkBDhB6KjvvtFnTv56jURt4NhapeONg/9pYGnaVx24Pce3jyLUwlQ487oJZ/l6Ty/04LwATw4vKJwzsJ9P0Tutiz4gWxQpGW2eelRE8I9HPF+rh6AB8cM11d44rpmlKRh59KX0onQwq8YEZy6wz2Resyp1I/HaR/2AFoHqKWHUBlnIYkFofl9YQLw1As+U2aQqexzaRokWrnKgCWdW+xdZBi5axpZzifh63MxxHR+4sAsRNd+qKaFWFCS7lDiW2d0jLUOYBvrANecYBFEjyiVi5g3u36dMfTUSrVMzEIn/IPnANqVYHofiwTbAImuOwd2PJDsWol5ekgMXxE0yv+yEVAzfKOi+ErIHXmBcG9jQmQ/NYLfzbOQTMdFMQGG4ZmStmptiIUMW8IluSn5OZAJUdszKOXteGwKdRufLnsGNTxGzZwmtv6XqLwm2Ikz77Ygn2FFAbuGyaIvLhCC49n3QwmVbHX5Yrd4tNLqNcMwkDNRw/JN5ymwXzDvoHScDjy5T+Y5IHM8IwIsPSy5mDE9ihWjloFexOV31HKL+Y13MC62+QhEXgfFX51fPoxV/lzY2tXGWPZm0atSixYwE+3ZlxDacdpp0Yt61nWuXoeHUgA94WO/QskK+ui8ENmjI0IzIGnWGZVTQUAiQFAMYS/pa33DpAMqpRzPfBK6q81vWxO7oA7AG2F/oZ0gSfUFXznNAHRJJKlZntc4mT9QqtXrdYL4h1uYaYNyExbFnW8TLhWIfWLQvKozOVj2un+A/nWMLHRkRsYAWrto4tAprJprKmIbtknZE/YTMar3EblGf7d5+wAquig+Ib2y+sgyJGvpjP2ev9f0cWKQD1xao16OQU63SA7WM2knf/wZCxG699pMnifNUH+rrIAGV7mpKcjYWT4iCPOOgDmzKsLgdCOezBk93q7tm9FPvWsl+VbAS/WbtrjK5rm8404MRy4gTATGX7GotlKHq/pfMxA2RyQn7nON9nf7GJCaVEdtnGHPoU8AcgiskoBffOO+kWj+cwVk+vxZxS0FUVKbKwaN0icM3pQ9Yty23T0gTVp2vZs5BB7mitj4H0/fCx+colqVdWb6ZMXdmDBHPH5lAy6VYwNmIRlAra2GeFX4SNR6O86fxDfhnGQh0YafD0y1qLH4zjfhlK9kAI9lmlTbhC4uouMvUVNYipN4c5J+ZXM7ZtUeJGT2E7P0p/OOgrLAKhdvVcpC6Ts8eo7vpuNHii0qGu7BZlBsZ3Oqna03aFUDE9hyYQSP8FSCWu0IKEm/bYKK2VG97yKmzAMemlz2izxI7TPDbKoILvXr9UfkRRtSWZjcB4OWqD7S+bLpnvWa6Bkio/x4FYLoyfQQFWpd2QCj8EsLCXMiREyVfc8ev16nrNH15iqbgUItmjkTrCvQqnFCP79yfnNJquFtX2eGfccaCKA0SlUmXCLk7XGdxeuzc2v8SDaNS/FwN+JHkKJQMe0S9guerg/X/7O6k1iSn3M6zWWp2tqZS4a1EjOh4ta4w00KTkaL2ItMPc5bJ7QMknKz92Hhb2sn/G5jUna5LWM0lwPVMmJeyUeTaWfTid5+NqOo7PO+LMGV/FpETs9kbUkKOoC3NqAGymjqTcBpSLYUxp2DV+lvNaMt5jZfDikCm4K5q6DklXPxt/Jj74T7hZX0N0qhofJvRIIRRFadFbBIbZP00+zs8i98ZqxlXGPUq+wuzW/txqmXM+/QubaQNirqUXkHQBHKNLrIlokT0OnMLVsmGnGpQEcFbwnXbVAKPpBDcqsYnE2prfHon/d0sTLLoXCxjmqovMyk8oWaVCEQKM1aEbsT5AeLooiGXpkT+X3kFeMH/q+Nq2frnawzEBfCMpPou9Om7ghdk3+ks4tlIlBQZx2a8dUOnVeLDZc45uH3SkwbAR/ALjQg1m0PyWTiv/sTraUuKELFhIsojNU+jCzraMlf1d8vBTPpANW60iGQpIapGz9AcDK91hrl4L9xU3go/k8NwP3FjRaNnQzTmX94uO0RvFUd/JM+ahrIykxnIjhkKHqWDIsrzNV1lx1BUcmztkd8xYrifRWkm5f99DjWlM/637Vi47HB3xsyPCJKafdbIeXuvLGSOzb1vVRwwgTZFfaw2AkQa0nZG9cIR2VQ0oKvsFQJe5/Hfdt/OrUeDo5Eey+AF7O/PE5RexIXKCiPyxsvSnfp3mrM34vvMBpvHZhA0fAqwypzLNAnoYmx5Ru8dCgVuXHGGCm086QyThXP4ojzOmrCoxf/jyyOftLolzvF3C+y3IKUR7DeR+k4xwD8pZ7580pMsip5qqpqU4TTaCfin/ESFEwXkbhkMXCOSmka+deNpOmiCCGQmug2i4JuLO/t4s1yzWh8DhzjUNgcDtLQH1REuWBT1oz9Y66eiEjBgLm+Aah+cL0fzxUrojUKfYCaOiDMvWeMce3IIA7V5oiIBE0qbTLXnnREr+oTOT6zNhq/CO0NO6kGMzuc8wHkpkT/JAJZSI/d/i3xCOs4IRMPES7cw5PiqTYV4/wZSFSwa9wY+TaLxRReWukK4YeMZxl27kUiT/VriXFAL5cn+Wa/na+3Mq4qzjovjryCIaBA4R9CYrdy0TJGOTR0pG50dLr+WxLXrPeslq7fUVH1SEtEI135R1adoqlGPZC1l/9HbJjt4eqGzLjKKSD/zPPAOzwk7C/XiWRhXhfglZMixO5YCg+8dmIE2T5nhgzMUxDrQaBeHLqqw0rgI8HB0fAye8Fxu39yXVObiKesHKZrDsYfYknpG3ISrXa6YXOP9hH/a/bm0girGaEsDTHO/APbxKQfombcw+/s0bVsFBvv09cm+6cyXlBWWwxRD/UXh2CvRdD1tzg3h8pzoR6Q+Iy7nlwplFqRoOq05Ofnw3ziFURkIpwQw/OdcjETRkAEhREm74DTKmp9Wthn7nUrXTSgHgkGmyMw75hkUdosX7UXtOZIJK54wLLaISzOsuoDVdmDftpiK9pxc1LVwetCv/Jp7oNtWKXsb6NNF0Gb2JwkHjRnU5NwIdaIr78kHcrpyrKiS1aSHhWyPuHUGWI5uX9oiSjRaZzLhVJG/3L3RMNhDU/wQcVv9MUG2EcUjzzSrjjseOX3f+SB1KpOljN866Ra64kfXo9saKVylR4u1JDS9KJSqxXJQZX3rVxBJchWxcEBbjF58GkX7cm71HfGsaGI9sekGyLZc2fKuO7mf6JcfawTJnQB2LxDkz+9km1LN8Nwn4QxxCUr28PJ/AQWJqMkP5IL1AFbdEiPBFUGLSwN8QkQjILERnCjv1qgpSoCWcCqRW1YczEvAqWGcXic8LbCZp53F8sz3uw5UZSdxr/+0CsZpozVfeLQqsS+8CrkWK9BzSIaaPTrzSE/l3CvtVM/dHQlQlUc6adeziXBZ21+1hokv45NnWY7GUj95uP6tojCrxeQzg5xJKkZ0kQGkHSNC6juSoW0NYvxeexNniWNGBRKTlJAQiuvTamN/Wx0PDJ9BXFhbFvXT3gHbOHeYZgsiY7tLws7mSMYXrhAUrdFRoqY/HCZdb+609g2sBrYMvbcOBAQZTsWxc/iYOV+tckE5yeW8PaOky0yZMlwNhilnBDG1uBGWF1/UGV3iRWnZs17OAQrkAn9WQAlv8rwA9zHAFR7uaVnmxYKJRS/OfjdZgBCPlMRCcjDvn5Bok3JhqDeRk3q7vGRXs7iTxPDVp1wNebiQMTgvv1lcTqrQvNWwuXIJL+18VeBWVpI1WHb/4jfzcM88s2Tda7DyScDmiOPA2BE8WAkp9MKczYeYNhKKTo9y760zdt7ANzp1oMS4gbpStBPva2HsHwCdQuCEYcADYoTgwTwBwrviKmSQTH7Cg0f7HSzVTVPc/eUxkQCkAm9qm0oKDfKcfW1hsOizN/g2x5kLRuvz7S8Jq9NcPWxHxqtI3vcpmNgXI6PyrmkrvmyGltuavSEY2I2a/Ih8Eq8euRIFuK1BDSxatVWuA+9rMd1o62Ybsvk1O82LcvsUowWlE+l442pEj5wdodfZJ4251+UUT3HdohksFJLl+eX1iqPYpKvLKBK6+MhRrb9q+/V4MmkpxpO9frUnYijnJlmzoWDl5q1Bz1s2n66qlzRV27leMgRyi/lL+yS9kDwwGe0rMrmHWP0F8I01knQa5neZHubiZvJDtUPaYw099PVWnRbY2MGYaIkGaJth2NuYwmQC01mKhAw9xSYZoBgNgdnd9UBxdKMtpr3lXbQL6DeNNwGh0NcPu7tpY2r7RMghHXY0KTeqtcR7tkZ5xSHyJO7RHki34lYjn0/zb6OnegtXqvFYIB7RtfiJTIixqxBmSDjDOpadEelOjNMkfPb5KW/mudQVSNmEVfWVcCOhu9yJMAxODLgnZqety+7d9jr0+n1z1ruf4LA83vKuSQSPEvqhYNhOTwKJ6fzAmHGLeTy5rhdnkhpmpp7oAVQhpDXPNNWQGfJp0c8SwoQ04YxOfSfIVAQ5kngA0CtxriX8Ly4GR5UVaIx0B+Jaud4HyeQq2Oz5OgPIhF/s9s3vJj+HTQYL0s/qayMVk76B8o/1aVXMDEfuwGDIOpAi4DTLrPaG4OKvN2Ie1rp4JH8O5pAl3mjNAsgLfPb7XfOC0iawrr+6EonOluKAfMoHEFn2/0+IygbgJLqL14H4Hi7x8G9uUYHRUM2rsSjhvq24X0zdFIEdki1oIljV/a6L3OqDWqHd8aGZwaP4OjGUvw8TqzX/SkwkIB2p5gLI24d1WXNtsTEi73oSiYJm+AX+jgR1JR8BXclsmq113/5G6jE4zXmkSo0TKbrRD8NBJJ+coVWahrcgXdsbPC57+sei7JojGvtCmN2YbSYPWHSTSZ3pxtt5y6s+FB3tjF2xucoQnl28rMiTjdW/3RyI1WnReUzPckgeKs/NKuWI8V1SNsiJTk0bWCknWh7fB0uvkeL24y6QiusbiI7nDnyiGv7M88UQts77AHD8c9dez9ZF+5SkyLl4U2Mhntw6D3G4f/4Rzv9y8cW1KN04OUb14Hh71UBm0cVo5GjFzefgdaDAYfzDTQDrFFtXDfCftBkjrVUntTSSyVPuQ9pBMedA3FPODHl6VYmIAA3T3xVH5CZ8Ko95t5qiPxvd2proXJYuVkfymebM8NPerv8unuySq3cJDRLer47fwuaYYvbNXu0oyYnJanV4nBd2JWDR6bNxY/3SVbT3mzmx5ywFoiQn6wDA43d2U8Wa98YoZaUtvxNrW+m96Qq91I7hMi++QhSErtrqcjOGHQUaMxbFnnf+Oq2gUKVsGdocftOp9fUnb5oclQxBj9nxlLnPp2JInvGhqrOHwvKQpJQeix0ovhMxzH52MSUbERvd6uX09Mian56yM1Gg6JMWCkMJj1hljumU8P3VguWQWBGcVqg/cLxqGfx7hLBr2KTnL9SJS+1eDRScVJUtTyPPLjzD5jXjZMk993pab728MuEUI18o5wXSEFof+NreFBMlmJNIvqxJ0VJoRMg5a7RxoDdzsL2WdNZrzE7ZeIBHdJFBVayvPViUUIW2uubwg506oYZzk7nlH190Q4VofeHqJmWROh4FHQSonov4RmT0cGeHUNyzDO8dBqE+xl0fHcNQiVj93eUp6fP58zDaU3241kWjANx7GsP0HfctNgXVcace0/qIycC7rZmgsj53RfJ920vBVrjt5GVfCxp6aBKMMCS7nV7StQKVrrEPo64Pwoq1NitTPBMoQZ0JOZGEzjWm0TT8gLEY7rEPUFgd7kArTnQO0NMcj8pZAjBGVK2vw2j45k8ylS7TMFPEU6C4Yi+TVmMZpWIYFldMtzNmXYkfIVVi1dfGMvdXEIK7Gx3ZdrvqhLKjZQjm8f33uuxhdA3jf1XT2SWRWVu97aqcl+4w85305fJO3H5zAHYfhB8JKJySoBuMOJICqXNzqLW04T/RFXWkMyFRRY5wEqZRpgf6+3a6j4inZVhoEYvNofoVAGp3AG7inoCQEHRxLyaXxnMg2Lvh5d641WvXjP2txL6nV2BjntSUMqpHaab5XmpQ5jejx1iGs4DEia6jGfzsMAK/Hu3TXyf6l0vj5C8cOwbg5MgL+sfar5SlWTQMmUHOKZ7OPIudUH6Nh9sbWjCc9Z5vv0dCa3i9KxRaupnK4iY8DRwjt/WK7JYkbJ9K0SHpMEZErTuTAyTq3D99Z9u1ok0CLmMAiBcMR7rUi45Fjdms83HGs4yPS+6luxq3zsICR+/3WYdCm32CX+tN+JZwVPZG2kZ5ghtgehAiqOUJDV3en3XQOwM+02mBT97HtpZkg16sxmV2oCuXGCnSibuMJ52s/Dm3B8V5C/Ii5zejoCsxlfrrqnr4cFQnqG7zjLx/5gZ9mK3a7emzEkvRvhpuL2sqwFsGMBfKL8UFISAuQf6P4AC0nA6u6PN2Alz6r8/zg57gy8qBmUiA/5ttNybUQYcf24cMwkXRwLFtoVqfWirmJoaSZTrR9/VWY/ZjM//LI2j8LEZaAQ7OQgS6YZjhn3KFwO9jqY82dsw/3uHb0hyTnfVR9ZuX8psxU9JRe0G1shQSHjdv2oEP8sRxjqSzy1aI199xTJzbXgjlJdRi3W+sSA2HSy8GcoS7bGnsPRHu0WTg0t8gFmSdnAWiSNFcTar+dj/8EZEQURHpt+4IbdT2UJaexxT1fzvY2Z5Twq7mqEvYtiIBYFYRUQrf4aAl/BmVybW3MVGKtWd5WgjHA7ri5P813759kEUMqoIm+GHkbj/t93IwE0oZYRXSPCRA8gaGE3SJyH4AeiTeF98YEUZ7eFCoz17xRS+VfdBJBKhEjxevaR3EkZzs8M7NfOsJ7JTB2BnDwek5I1Urt0XVVTS7te5rBDwwaGRnoZCo5ONk/sa/mIcob6RLNT1EdGoCe05vzj4UEl8hFJKy/a0Xm8AViaFMd8YQUnaeqkXmMf/Kq3WybwC7j4yxs8UavN8BXu8jzt9zGNnB3QPUNaO4tGUu7hdselGbfytWUg2XWJ8rGmwCuLeyXkXG2Ss/YzSyJW5J8+qH9OPuTd7qF2fX5UKQIBmipdtqVEVOsQgY/6fNNXbtDlrqIY1hgBysbchAFZUmZTUIb8g9BnvBBav7TDXCq5ZimfnQaqMo8uDeK/1qYaeeVLz51p2sZLOdvp2T5lpjUWRi/RyAidxnPQX+mV+aifyRh0P9qrslOptoUQoLJddxGquWtrDhPsuq4ayGJnQvsqtE468RxxSjR6nwUKsqYF0h7IYWrQByVzI+nattSobw3LcR3lMO/ywWtOupnlgCA4o/k9fSYG2VcrTtDwouG70BcP0s6/LXg2Ig3O2282y2Qq3GApHbrV8/veNO9oKsEsRs8iOl1y3DaTN3MV19FRx4Syv/u9nLBIItb2gDQhgwU0QLSEMtFJtLP9GuMqxeLDnPREsBCO9U378IGZBI5yxMCEHvaSt65Ob4Gt8lYaNK0MTGNxPGS7hegC0w9sRr3grlFx82leSCLv87RJacQjzWGQy4/nezQpUe6zt8xo13dy4brwdgKZJvhIRzUSJiVsXP6hQmlnnWiMlhtp8yV/XHmH+9KIPgweRK0KzzagI0V6hN6W3nWA+minxT6/V/0XxB1DP2XJ4xzfrLzPz3d5JS7VaiDNPjoFQ+ZURfxVu5xwxBhZScNdY+eWL31AHrT268jT2BhmClshBfELPCvKNbbcA9FvFH0Id8iYW5RZ7P8zsnf7YSrstI8+0rAFngosnSJaAIRhEoGuXF6ZPhlMn1cGyH5EE8RNG7mx1uJwihDaooubpZ0liy3HXiHGwDOJila5crR0LJMfPOFxIKpNTqYK72ULbrtrRE/HYaU9PLWBMNe7LHwo6bIHXh+S1QJEMCjxBBvxYFEH+3QSPqSu25FYlt/ha/Sz0E3f9nBQ/c9XAGEgdh4fXnEMVInJ2YfQ44uO6ra/9xCccwlEnj9ng4mYj3WC5pzHYN8RZRqGhUFVCX56ubPpweC3NkSKb4PWX9V4m9HjY52fGUWmFtI/orF/XvQcFD4rtOqxEtUEeN6INhSehGRsbzhfHV0683MwpingCIYNrNVBXpe7csuJxyLlnSLULAm7f+IczRophohIqo/cjv0qLuiynOMqGiIDb752SzGXmP64leC0jSU1rNtMzB7NHGlJ/YSu9urLk6YOjF/AmszPjJPyEGUEUn0iSXiKwSfdK6MYUSob3ApMXIFsksMwsyXC4o+KqcHOcPK+yyTOUc3FsOYSY1QD34NMZplPPttzZYFildN35CB1C9RACq/O+7YdRqQoJy/4db9Dt9X3XoZgwTgdviPL3Ewfm9HcChutcALc2Q1gRRRKnRj6QPujPOJvebpbRZVoJMU7J03vNtPMIPEFvaAOtltx9zHT11Nbhgb1wpjvv0ylFRDQGDjQtuwhCkwB3NyTjz0DAAFTRBUR127iyMHpEOO6gz9U+7aiIuDTRR8+Sn9WiPogL+iBnq2V3ITAegt2NtdPcuXh/JC9c3WtDAVDP9nOMYrsuSmiN5i6SJ+aKBk4nonQ1WA2rbnnWwfu6tdDE3+hUsFvDsM8Ia59wkCYpIQ/yUIj8cfib3THDc1VZzzibB9CSphr4poDX/715tXOcrc0gn52RVPAjlM9qSG2iEhLRfh6P4FHgDKvgOYoUaqMLbJRvaE7WgyfhRfWgoq0yS4BitokBPdLHl5rCtsvTEtETmYME3aIIIm4Mezc8QrqtBWr215M78LPPPdnfIVSAyGp8H09ilu/GVd7jZNQzJ3Tscx8k7Sco0ym6ag5U0z4rwAiDSjDDCRgRS3Lp5p1zBlUrf2cyg8dT7ImQsp2kkuUkXTh6KFteq+BILRVNvqXdTtLxmGsidP3jq8U12X+ZJXxl8lHcmkyjAKNj3FhCAclx9uzCPJjYFYeKAJkCHb8pfFZ1veuh0ZAZdI1QCE18NYO5heB6z2jDgMoh5D5bf9FOtJJROfxszYuONDcdAJh320my0HB0923TcA9ViEWMD1CDzxmtZmh+bjSTeVOJxqn02dStldACYXidzQL8XYWILxphEZKVpykXRB5DsSyTb8kih3K3dI2w86UiBMV0peYyvw+j7pWEU4qy1mLTMWKjYBVjC7Z4xZUK6sVqH4paH/ND9MkG8iQ8fNMXKpKoCcmS+Nsmpwn1PyRM6Zkf29Jl3JVZUWRthyyNq91g/z0sCcQQoENNrjeKRtJqQFZ7DH+1xv8qOqqrq6/UIWPg9emmXJX8VxkiNoIkMkwyjNKe+7qeQy132zvijrRZgk5sGrtOLvutrGu9K7rBw882eb16544UDldvwTR9AVa7IVkN8NUgivWvAJgup0pM/TNL2fPZTTfSxH2Hf1W8pAp8gQn/CLYK3co76GsgsszqL9VyVYgLb1F0z1bo9/oSE/1EEiwKFt7nLrHz7jV5G3ov1GR4nOlqlaDBBhKFaADhClpHezik/UvxWoh9PTgbhe6aD/jM55VqL/cdkniaMv0W92uDAw4Kzijyt8xrGvIqnRTEXShXMKAsM8Am3wXevxv+TJepG72/FTwGfUKfZrfVZ0rwXqdOO9LS34rRp22PZ69MEMA5HFL4AVdzF0O9fCgKzXNQGka3tqqSV+VBJI8C3U/LtJ4KSJ9dvR5qhBzLxc+dYrEDeA8BjAYnr9CLbukgER13/AuvobSpwP1xi2oDhKKqKsGRkKRkDEKqC4fdZpyLjjEn7utB+5p5SyLO/NdRxTkuPbJ2lPlNnn18j+ji8xSVzUGMTD3Y06z1lhatYNyfGbGZCppPDFqOq5/ujhPgLtZ/XOp3IG4OjcNQecB0bkQg3YCDpPlVUO87SHJncvpSRvwVtJoID7LtKnHpOBQSnRgihTXQ8LeZju0u+JeJrbAfGTKYOHAwJYNZIEgK28yR+vhOZ5rbfqVXPnQosRHLPEjw9EYmKcMmULD3czAZ1UG15wO0IiMJizCFQFgwDjQNPEiNudwIZFEw96bt85kRcCqsM9wdjBPfoxhreCGvthlxs4mjUU98bQ/r3C2SO5gd40WOWtDpg/V5zOEOBfS0FvP+1h0OPRDduTrR5q7+uyuQnBWq/9cR1Jvgl3mw2z/mywjy/P6M4YHBz+EWV4qlrsjgTSApbIeJNg7bGitxgnYOWivSRPcsWGqk0e09rHQzTxFogVTikojNPAS49yEh/54Tc4GhbyFsLl24FxVasLbjQlLyENWreX6O4Qn0GFonQjO7FDuYcMA0YANzxCiACuYKOpPXtYAmhRvLK8WzcYPOETpnQJY2vV4WIwxFRtenu5V3fMumZZORwlyc1hKb5i0jCSJ0vcMFAfBLWHUkxqS9v2pd/vgcoo9N8n7K+dDdgmqSilcgNfsL1SzaUSKKifdcewP+lgyp/wyKjwdHQ42z76DZmOqe7x0/D7cZa5sidPDVE4jfEwSj0jrjRK+mPI1AsM1qdxkPWGlWoAZn0Ng4PwOxvLUnTiVAV+u2YQw3Idt6FYPxA/yH0MA/nwF8Zo1L2oUhtbw/EfE3nsm35hAlAkDyH23RP5E9ZzXGNtNZpheqWuWNp62W1m5sfdLdLV4z5JMPM1WxOoLzKBonShrW3EJ1+Ek11vzvZV4fazKpYbXANPLQkOCWyW6pLHn21pkq8owEVO5T5O7rWc075YUlGv1iKfmQx8LG1O7X1ACKolnTCXJhUjEbPA9TSCoqDmPHGccH3hyIoiOofTeSdIYn/bZBA4eZxyA5dvcxhwfxsOUPs3apq8uxOE+AAF3CmEEYNAes6f+sNhZu+e2mD9GBA2eYTqYiiRkLozwNrSWebXM0GODO0VhV85Dvfa8mKmAObInTANdGZYbPk7KtVXMvnrIkKqtsB+p9f3dNfnsQWrd4+2XqfAu/sS9vuxXdNOZqHWAGvUXJ8TtFCWCCm2e7jne1EXlRCvKD3VAnKKz4VYP0lXOLD2JNQNBPxsWse9FQpkWxD3251rF8Zn5TL1Hf2510/0wZFg6ofcQ+6tDBwjThLA6SLDgUzBa3XpPdLwox5nIUh+zsyTG2ZzVw7Bg+pPMvr5jOCaPrcmkIiSeCGAF5jZ4/Pu0Cy8SBB2aYT0kyLhWayHpZbFSF4I85FMlaVpqNIW88Mc5IYXO1VOq0l9gDque19ffQgcjGCzHM8VnvaivWPl1nYi3BA9MvgupGgZyBbEjSZ1osM0nb6LABczdIUCL9UaxdA9sPBec38c5p+Mf9pagi3EZA+3R7WjzLSvXS0Pa9LvqZ8XFSfDIt8Gsb6KR5yibnT0kTIaDi/wkzcj73VSgPhQKqZQ1desm1H9/lZ7V18eEsl5vTjVNcQDnoa3D7wy7Lx/vGG/GNzL84ayaBX49nDiNESc1M04p6ID7Li4+sAJLkAyaq7heZJ0ykf0+5CeFbngaNctQlNX0dPodgV+F7mvBxelqp01QPASlwUES67ZGdY6oaeHco+Vc0zFAj8T2BFTFPyLaWVaRnmI8EZZagRlhkqqk7H8KvFKemO793B56dMmxi6ttsgl5EF0+Vb+dVUM0Dp0xgkj9TwY5HVvwPmBGEJ3dI9mjkmWQKX4iHdMw2ztLFsyK1Qn48qEblcTz7ZPETS839cf0fAC3Ix/99eIyP595i+56ZsB886PNhYIL1/t1cfKj+mAlp4F56+hWkMzsRWXcFC2tThwQ3RhB3fJx+uCmMRy+d3veQfI0ABIl7ibDqO5vDfP0mYN8dqLKma9ocI5E/OxMtmvqrcCfzj0hKi7fJszQld1u0QjLjEaEv/VmXQOCe1C0ENv2rMYvDdM4qMkw6e3sFWbcVTmXwn43iVRnISw30B1jIbxLk/tpUlMpBOV6sJeOKVQTHv+RG+/7XwQqjyLd+7tnsL4SqHzxyf4MvoE72KEhRCPAXtwbCK/DvkRLHcBGOv3/SralNrnZaqUH5z0EqxySPfuHGzVhPwk4GAzq/reiuSb/evZTrayP6QmLcY/uBoW+/MOGhsbDTks5awdZUivSL0hTTTWwBNEZDQq3Y3NVb8YbT93Bq2B2thSv7sDftu4vTiK8olNr8zFOl42fPbfMo1FyZd/BdCeSp3pvgRConBP5bLlipypagRMAA3x7XgAYjti+qE1aeqdKpnb7wmptB1pY5IZDePtGYX36DcHPOT/mMyDfd7uqK5HU7yDqWNV8NZGuEAxMOhKAUPcZAL39ukLPFLS7UKuXTqma589Mcv4JFILuct37VfrzFjUWHVNHf7ZWD4aSKvS0rOGft5i1DKXV6VOSvV6WVqZx+w/9o0c1HwYRuD7BJDBpK4N8y+O3DJn4iLjQ42Z6HY+3QVRCSXhYDKR1Rq24R8GOwOOG4LeTkUdK+Er02irbSXVuPQ4jqv6nua72PpMUk4N3Me+gT4Wt7Fuco1dtnQWz4HR5H18mtEZRPfzGFUMgjSnEdnTBEd6mTfHGe4NiAqkCIqnDlyNZVkd/ZEL3D+atC8FYaXFxvwKnpDfk/CfM+i2MJe1ns4hY33YZFDlHOxygu0eZGYJxqJWWmhytWwKOo66iik0VLo8GHpcxiTdHlteIMAtKqKSTOeLRl1S+19ZhVFK4Db4wIt7Cn4mEmBwEdK4qi3vl60DILJdN93Aqky5Lvgi+o3UrZxio/71i1Ql52UNPw1GCkd7Y34qn615qgXWKivF+9WUzUI2++8sbvQv+Z65jLmup0XTAaXNil7kpaj/mkjdo9ZJJftvM07kf9sl5hKWCK9pOWmYOvAlLG3BZft9M0mRlRs4pQCZW5+OU98u7GSCxsC/Hv+epBNJGjF69FO/jIHMDn6E42/W2yKBrxVhns+HtGIorXAZLobHcZZdCLgmStz7LNoA7LvNrlrOzv1K7YRWVyWSZz2XMH3S+Qx+BXwiUBRCBkCyAiNUChU5fasnPEDNx+AZ/431UmR7qofN0nv9LjcXB/jfDR33FTIcMl9jSCZoyc5B+Gq2obfxTWQnjHY1HTfCDqWVhv9ekoQyof6GkzQBus0yX+6AaaUkDOkMEYmU0rlg9gQJ3xNOUkjofvrLxjIo5oO9s+Za3E4NfM1aX3Uvh3er8n5EXBwFB+DD5DCaIck9N9F3O9fkALm0mX4whuAHPbBPlrcs6lbtyzxw4kUB/J3ACjlTbVASxCzbUHas4lrwcN/BhlS+t5iZ1lHOMMLpqfTsEChmJpDqOGjnc0UqYa2AXs5raZ7o/bw3pyk6qXKNvRsgn6RnhInX/3HaXU7WfAr7T6+S+nEu8oLGKvpm7joqbaFLtuGq5BxsBa0DeQrrIaCGR8O1Ezz8u8h5nNSxC+zNWXIX3Z4vDr89mGnropWL17wQ4cVFVn4AMbCZ3Is/MRXweD4jUI3/8nGMMCpRYY9ozK54dpLDJhsnEOETdv5Ce7vNNpj4qQcSbkTjZXP8HUXN21E4iiTGyec9ZpWVz3BzqS0jtKhDTvaMNdvQbZj7b0mRQGHkP/rjbyN+dj9qJJ2VCyhSTJAMcsitLcvPflY3yufg/JyNkL55GyJRzqtszHr8olml8s8es3l3kblTrjXFwuK7+03PFqC+ktel919RtLSJ/K8euS9wzHa8gd2VkUe0eYyiGeirJxy7w3TP74UZ6PWQBGIsQumaCYHwyZjO2qFquaHcX/uE0Tbc3lHj/FMBt7pEUa7dTuW/GiFvkV2RxG7l6YZQ9cg0aqXBESJAYfOXrRasqTkel4DHSVWxtNC/zrvLfOhnxJDXF38sKnY+0DqB5PUk46elst1kw2on0TUH6EV/X+F1REVpQIb3+5xMe+x9hpqDpPmN+4B216j8t11cRd1kEA/19wHVxcjcHFNcPV4EUAjC5Fq5Ge4oFT1tHLYcPZoxc8au0ChdQahdlPKz0prEEFrJMv4GoB9h7nZypuj+GSEXdMMXfm3RuFbcFWLO4bR6BL6jOWyVerAXYSgz6MPhOk4pD4k77XQVfvkkNLJPu890kcnu1H3aNsr3S8lZIrALBplszuolnGwcRhxALgn4Qodj/b6Eib4Hb59JgKmhFeRkLfpbLxkL8gAEHAnLXcdnkEGTPR0LAnZGIWZiR+j2xNorqhtUb5c+oCmD/xA4XcgftTxL8lIbEikglmMQ2gT3RfF7Ox4TuUi1kfJ/AqYk5eIFLTK8Fk9PMWfenqkfsL68luchs22/n8LOYsEsfFK8ST0xOR5rBBpZN2iNu/MWbTQ/vPLwVUdnnmgzkDDoiPc48tzQJnDgfSUMxAtDuiLt9G+Fw5wZSx5/gKq5jgQwCRyciUAvC5GunBgA6y2/yO3r0JQ2wHLUsNePBLawIF0Z9Vp55o7iaAPtLRX2fU3LCzz5/LdTXImqfdcKcBrxObbf9KVSnh7udSzmlGm2/3INA0SEzC8QbNSidtUNox+tHGSLOWAXfweFZR+TOGxpBwaBktTWePDSPJX+yRNrc5Mb35A8fsTJ5J8Cd1OFjXl8BlWOK7GrtH3XF4/Rdkr9QYE+4bI1vc10IHmqlEcDpCY5HM582GusaoKcB+twVANggP1Yi1jZ+8cghSr4LHSTFmk4r5Cfwnj9MOU203hi/KvRybzRx1lxyQD2/u4DhDhXN3ssbQ8C387/H0ngHK+WkLhNyoftKoSIV0Lqvjy8QuBkiaXOuW5aaSW7d0nFoNM5QnXoYE4m8w03AhzBr4NO3+qU6dAicjKNv8n5MKY/Z0dYwwpZPCzJp79KnRN9rH+wQWV1MvLBodYK1N4jEqRNFWGCuixBwM7MzgPTCxfx/djuxtF1jKl2guWpMLU6GRJRp96JP8/HomBPEUo+nlQXlF30gk90YM6ouaCgiBhQitBFhetFn/uF5IYLUm/GOp036TLliyoJFqzf2lnLGzOuYFVxrMQgvhT2ECyQDWN9EUy6rTZU0+Y7YeKWsZbhaevBT8J96WfefCPr2E89ZY/zyZuR5uPCczHYyne+UPdeMJni+zrd3eLuaU/NaEIp1wyQyBd/cuOeP7j37QTQ5YgM6zas2NODL2VGOKpUQ80SvP2676cgOj/dzkOVm7xexGBtWCJjH71AqdXeDB9/m4uSQJOMy9GV0q9G7zX5y3hXxh57QY2+TzGxtEBC9PF4bu0MtoWukhJnO/gU5zjJl7DDTEnFmNJtV0d41DcClEfVwyXwKrnFA5Uy5XXiXlhcOM6anJ/1Drkn/G7gM+IbekPJwLGjRi8RLYHZgahi17HrScW3AIogIXesRSWcLoVez38R865SY6jG+tjFTuxuH39oRyyRT2t8sc5hZLU0FvS+tOnBKm652o9nrDqlYdaiVwNoZeFoX2MT4gZkvalyIibQpA217q0vrIGdbaXAoz6jlvP9rRDN581VG5JjQ2z+wtfucsr1n4cnmP67e/KmevVi5ZdfQcH5sKbfj9v8/Q1/JMLp86Uq7WhBsM7nwe008DT9x/a5YLo0zDM3mnClnRoL9EI3P0tDEL5vm07twef3ibNtLC4P/VvBqLxAmmO6GeW9WBToKirdWbxaGLZ1jV8Zlwhg2oREmPcXrmyyU8tktvm9KwpTTV7XcvWi0dGIt6dr/hTA4Aan3jawBd5SMlLEkPV49hWi65NqmOpGne9xZIDjo+zrHwsXcTNl2QtUxgNmOq9cG7/2DYwE9Muut8V3kyzfHl9A/egdt85VIrb+vq6NpEtu6zDjcwM/+VPlLgzIdPX3EcvGsKE/zLkcYOmOUj1iQ5e0ZkmvEaf3VKdUSVxVCEw/i+YJLfRxFTAZVi7+Q5mf+oUKi0yXUDAryfM/aId5fQG0SvDdPodndf7gU2Idqm0RrSGqeKvZoTH+0w2/1HbBPXZTvCE1B6fHsH8QmhFkLPmild9cZLM4jotoCmVKEzFi4n6h7GVuqM91nFHZ4wMv0s7xE5GjjIW4a/MG758gh7XBYpYromWLyMHLXDgxTHi9doV9W03vVYEmhYFQdrl5HiNAa5MnaYDCxw8X3GEeqY/PWDQ/qmTZoCsa1sLAJYK1jgImDCKem+Fst+TkI5xm/B6u3vh1Ls2jTNVmlXT0iA+OPCeVLF+94Dn93105ilm/oT+lt331ElsylHgP2RB/ulU8StVy/w8PoaR5SeC6SF5JAq69RrcL5oNkyAJMZ3V8CExKEHIVP9UYiaphYFoVkQFQbjGlM1h5t/eoXIcpHrRmX5v5HdgprPwWC4xMmVYCS9drfHo+60XD+uB6z1LBEC5V8/qZAjzB7x3HlcY1wHuHWsf+lUf9r3ECgfTbqG6qSyBXWI6QHq0oJgtLzcJtpP0yDt4e3UKZXnB2oVp/tbad9SuzpIMo2UHTXzmlesFFANZVMsU/ZEPSdJCiQmIQKthgXyRZDYMI1gnqD0pWGkDbCGjjbec5+O4dfPONdokTkeTCBiB+hmrMKDD1Cpn3x/1xGa5O0SDfyuSlF1TWLcyn9Tkj9dPD+inEQxGmEqMa8opBaVVyYyXE4HJkCZdgUKg/F32V6pdKuthrwZoRDy2Dm+lO4hcA450ISHFJNxJMEFnMZcwYb6giGkeUQGNJ3ubCXIy58SbOl+PTNeT4ayAvjYvS4e4sK2z0bkFcOrsVEkG4DpBRDCkYgquvrXL0NMibeuZruKdZJ2wdOcewb9WwMz4zuxj36n/7U60f2hdPt6DKtnTCXvUcfwUIm9BAHrtfItyI8w0pOjcqTfU2WkJ1HF7kW5IarsH66s/OqlBR2m5fYcCSA1FV1FZWifh2OqZrJBMRHbKI29eCmTn1iIPOcVECAwXbI/Hu8vBedaqykJJZ0PhHJ3kywl7CYJOIYAtABnwSlM4/tWIX9bMk0gx75PWvDfRrGL2AiwIinoPXf7oE1Z1i4pCUOAHUE/5c76Yl5A5/XUyETIMn5eY0G7/6w4bxzqp9QaO5HOHJxhCuZix8uDW18b3Xjzod/o33DkBDGN6xB4fD/hxtR6qo9NmDu//JRCNxe8X4sFLdFZ7dQ7HIX67UXEaIZtUAVt81BQtEUgCVOAnbnmMnN08uArSPf2GiqCb/5odKux4eK+qJT6+LGiylSu71SKHtzX/AEiJgOEQdsUEHDPuCSyVsXuth0J68Jnz1M8QIYTzO9mpdJXxHOIa3VN8RpJpncknOfdNHdpl9skEwL+6HR84eugIRDyW9rsqSrC7DRmGpmYFTcXjYNOVxFP8fpUHygeRzk40Okn4MdZ77opwfwbm4QtZRg70JUA+22e8insc1ySanjzpnKLGmA/hROFzKe6dNgDbb9dyOW6XsgxybtkhMANnUBvnUKMFKDAH3E0eQut8+BR7Azt6v5KCHhZTyAbfojIaTmuQUXxJnOX6/SAqrUcz1PILd3PPcU+/OXf/7UHJ1VeFyejB6v9FKDSz8NgloRnPccylH17fsgfwhkeegmB4xZMkBOrgr0k6G4a9hVwcjGFrgdAIoyM0iZAvrJDd+u8uOEXqsVNk8q3+ZnLmSFwNV+pT4RbiriJIY8IHolda0jg3PEdrdXHw+IHbMm13x7p8K6IAtMfpWjLahUJkb2sIYIsxIGK9U590GXXi3b5Yv8s8yIt3G2vLlxirhE2rklVhH+SjZFPvP+OWhrSjuGmnxzgTfAphHpcoC9q1wTrxqJNKsOZ2+JNlE+ZVZU93JX2SL0niHutvkH0AUf7it5AdUqBjEagXL0hE/7JwrLSRj1g3EVk8vAhtUaR0oMTWeZpucoCx5L9DnSovCUt4MEzkGG/T3fXcVOHlWnOsbuNqtLzgN0ZKE6YAytYd52hrVkf/nFKsvg2Zo1gJnoUC88ATq5dTT0rXNZaYz0i73eRfjCcp38i8R+ew/Ne6/tSDmbpqOqlnKW8veQQwG3easQNTM+1LRzDVxj2XU/uFcLcxlwMxgA4RZJVMIPXU2x8j+/+L8Mt5BKhJwJs5kimkcoeTYDiHOzD//9NbM6fo4DBkf5DIaltzb7MHk7C1jOYiYBZrMGW+GPhBRBj77BABFvg5wcT6PBqF3NCy+Zy95VhDepZhLIBeD/3FA++w3w+vx3r1CSAwRJaUFCrf9wiGjIjN7tFMu1qmKy8r/k9lzciAWjCy7i/nsiUdYFpuvThRqumV0e+quX/ZRVSa1G6cJ3KhTJ6eFHCSnL+KrAc8QzhRiv7Vi0850sHU9MHruA7d/aYqlYZvLMnaqgdwYMnQLY45cQowRz6gIBK1Uxkcj3KTiC2ro9zm9CwkIsJLHSuO0062r3fJMtXNYFwLRIvqXKMj3cGvlcrtpEnsLeoYh2SFUsiAnFM27NclJK6WsNOF5YvvbfdQROiQTh0h+hZ2RRUWEESTAWLzytd71jjWMYQNk0NzrlJnpQOE4jLwTm0rP7wphBl9ly+ahWOJsencuhhnY8rLfjQIRgbl9A6osc72mIuRRhLq4F2pYaa1D9PxstxNHB+pDyGGoQ37jaUZFBwxqKuFhXjnSZ0lf+MO/f4ofsM2ai00IfEOTix5OvMXMa1bDKard7ipxWk8Uz5z84wgP6Gj+HTmxvJBNvxyvc+fCcr5FgUUlNGlqQmI2WbNQ85q3HAOz5aU0eZ8AvLl7/TQm1FuP7L/qJVC1+P0MOVE0btGiaWIRU64bMU+PJ8Mhyn1vsnksNa+cK8qejW0N+EWW/sSEgrvUoknuY/qupRQdr5pR7RvF9dLBEZ690Ihz9WDYM1yGSrNxoHFm/sYTNU5FETJ4rH5daZydVN0oi7fJfD/yldQm/2tf+zMrxALUxZlJgfLFMDp+8/Fh2DghxHs/TxG/88GfjZcMgIF8PIRbD4Ah6CIUC0lbCd59ORkY8PghbZOt5250lGmuxOxe7K8GiaS+QIcoe5bRt4+ACya6iy5+t2Qx9mtra1ZWQWQp0FjtpASM9uc3xCeggRfg0g2rDkbrvbfuQ0rkndP3Bf11oas8WsWVLeLxip55XVxKNluWYmwoMePoXQeIBjb10hdlLqw+jEQwwwIsHYWpRHvpeuhc+3/DnYs4GzGMqAj81cX9M5H6HI2I5zokGmTDwLgWetnMc5DH9G7+jW2vIDv9IrUY4NpEvL1bM2rSg9BTD87v+FGzmI3rNeY47ANYIEsuQ0nbfdjmk232gyYNv+uUMV6/OhIdHxqZ5aISDxtK9PMyfTUFTHXmzy3Hik8fszOIqiSMEx2tCR+fREqGUgj9aHYq6dZXNpOUL3VgQJSg+VN0vYu1qqiRa6mmz019UPRwTJEQpZvfsmv/LzLfsQuJMDqOtVmHoc4YP5Z6AiMrxb8V2zCkBUz4Q7C4e6kgpoQGlT/p/T5ph2L0vaJp8+eUe8S6E+Xpqp7qyrp0B0E33jZyZdnFbwEnFs4aB88xqFcVOH+fNPDmTV1PyR75wsdPPMHMUIHq01HBxmmej9jXaoM+Jtw12HWgJFn3u8IFgGprqRBIcEw8zFcbq5cdVxNJrYQn0DT9bfhFAXl/DBXQ3HSfKGvg4H7VQULa1IUMCIpnxlj05TJmuX5jiChvQqcJH/empG3KoY1WGGC4ANMNk5ZT5M2ZBaLclvhiEseeyuZ5NVqHjumwk2B7C5pf2v6eAgePSnWndNohd42zXPTMjyiKNG6hURP8wfSTMvPk7afjdCP5bj5RyKW+lURL8AEYCDRg9oeO9HG9n5vvlOQePCRYT0GnY+6tXlEFf0EQpz4SMJosQO1EOW3xIxErqoh2ECkmR1RfAcWYZ/LuldM2oZ+XyOZcluLMHyFH8TJv2VuN/o/EnGQtK3LztZ8ZlgYfkCY03BK/ZlZz4zhBRP4A5JelukAuGOuiVG9jJINTXw2ac3a4RdUcHtLazPNUW8IKTuTJZYNIkSqmCvNLA/gPPSdo0zI+uk2kPY53OprGijLllGWlNtx4LtAs2Dgc4B1ndeIraGideEIGOl5075NT+fhFPZtxX8leg1YgTgeQ1V00WL12vRtdynKKkZNiYelvZIZe2uI3VFU50a+R28k3ajcRvu9MYeHZD+nPpOvAQd1IZJ/XIzBo3VGjZpFNAAOSpwuSO4vl4Es3RkhoCzLBTTekXBtcnxkFZ1XPloKL69il9Cs2PhhIN8sHpVs6XyjWMJV2Fs3aW4ZOMoGjcyton1u3a/D98yEODGPjlEKJwoABY37EkfMUcqltXwywz5TmSPzz9EjNODQy0qNmBlRsYnvEQ4EPW9c4YjBwd3mWN7WgFwNBaTdBTwwNWUaHovwqs72gyCF5mBMv0NkC4Et7J+5IfqzYAuCNHetWTHsLbtBr6WYtw1QC08CQ5VaXFyLQMywBt+MWuOKCxxQLsLbweJ8znY6BoRj8hrLt2ANzTlYi5ZJitFEFoQLR/eNCCrGYlc8mVNMOghFCM/8c0gRUzbI1D4Gq1T+w25+w7GMXnZjO7NBF7vl1bLXjYVHnnJYEkJCLKfDVOdG3eCvxoXlDDSTz66evmQ6ajhzFZsVj7tgV2tcnFMLPVUTNVW3/KnoXWAEXp1OgM97joFv+4g9WrClkohdC+V4EDQcvfTpP+p+yb4wVq11zcS6V7BAMzz9iRCBgQEGEyrr25jMA53vrIe69HUk0LHfsI5kqh0/Af7BSUJLS5Pqzskq/oJY0gbkWuCJyfG1GW6ldqYWwtDa1RoZIxK2wMv8z4q9MCZY5pBJaeLQKZErZlekC3z8vGL1wd2sZHuOD9dX4LL7rGQn/W2A3JcY35dZTB7tWDfshnVg5zvxy42EwzMZsBXTCktzsyMycTcT2xzLyqStz5/wNZ6bjDhn4v4EVNSqBrY/6Zxn4kBngFdA+Hx76vMxpkJGRipK8zBE3cjiYM0yWlSa91p8jt3irHHNcKLBNE7Jku9SRzug83zR/WnzCqsqc2cyknTsRyXDMEH1xMjSEAW2hVbycIrauXAxmGV0C3XuL+RKB+NzAKeeFdfVp7sQciABxv46P1lloWwhFPTK+wfz2gYbTXpMZ3WJJhAMt5DNCvfY81NWf9bvzkJ6b/R4kgwH3zrKg8JMnuDR1NA5aNIAOimHTcrTDufRKyJwVVyhHj4nnDWt5MX9WdJAD9D1w0m9F0dTkO8y+2WEmnTTH0E+7quIFmcE215D23K5afXVyZHd6Cdsp7cSZgPWH4Sv/9ZcF72Kl7GCgP3z6HQkosgoxQFQNz4zAZjkswkqJdmOFyS4Z6v6nSMHL4tBP/LFBKzEDUIWlEi4xGiWkYqVZRsDivjzC/nB7yKNZBIOsgMtRcgMprztrKigTISlcLICDIEJtBQtI1lUVoTKD2620vwFwotyLri4j8PgDDQWK2HGJx3/nrXBrjuLVWo9OBt4Z/12mwGOz2tnn6GLeAjUR3WgvSafRuQj8KGdlob1sbe3j37OFcZRdLv8FbtPHLpCJpCRXGBHbq6FrsLLYIVhY5bH+/vSa9DlHz/5LtPxJu/tLo57vOOoj+Ae0BhHYbyOccjJrgZs69N+waTNx6zoXWrjPOWEhjV87x15LhDLNKCXhjaCTudmFtXzqQ8vKlYfC2r2h9fSrAQtrzgcwbOqmaE1L7YGVEW99YD6VyNwDAFTDgILjJDzGZ4sw4sV8WDb6yaGvZn1EbXuDlfICYQ2tKNELYCt++XJxVQMVgdeE/FkzfhDS6Mjhc5gVqU0CAKYtTji2uqUTk0vTqpCqJ70ed+xIbmcbVFEOyH255IstMYHPLvhoOeehdj0v1BpsH0RUdIPEIftPxUUvK5fGM5+NfIzS7dBZO5nUl6rlyG/rGNV6h0dXm+GV6Thl86UvUgyxKpw0XRtJJ9KU3ghOn1J3j+m4MvVP8t4yEkiKBtIANZlTxE334klGPU5yjH5iMa2coCTWoOCVwjb54AmSQI2zm0cCgVL3kTqwXkHpy/fHMwxbZ5StTYMZHG3hHEc67pxheeCjoYunpvRHqMTrH0D4qZ1SgK8YwWvIrEPRapGxOFa3Oy73+zjBgWwz3Mvy1AXe/Jng2KtujuVMz6wl4vwgQyWXKQImhRR1TxAoalVqwNClu5gnVhdSPsg+JORT37FOfn9SsUIlP2go/EZ784+LePVpRWL5GlDkNSAfSt+Bgw9XFju2ycX716BHEJhGY/M4Kqp+6Z1cRfAY98YNz0LAoXkUlDUb+osfOhIiTbrswzZlE0B+BRjL8gLHi0f9oaAEevifMCRKZQrSpMJP80srRyjevbSngk8AKWgyNR1Dej+kcQGRfyx6cyGBQdW8YAkr2PHlb8ra5MFdIhhxgbCCXP21QZzHJ+0L5UfpHwWYhLPHPQp/brEQE6/fXHhxjJ3kmKTBvDJ7q9NvnK0GZFNGy20EFocU8bhqe3ApfWmdyPoUvXZop/AeqzyUHYBgCHLjlsGcH++O2mTJ3qD71ipigPJGgoP+0n2+1aXVbaDH3A3yMePz2StQPZjmB4Uv6AIc7BdyMdPjNEhULI8YzyjE4eNBOkOoNWHCJ35sHy/piHDPDoBvNqGol1EikRdfKkBuxZflA/HhhxPsdyF7QR+QvY+AaN5MwART8PLuvM96oor1xQHCc0t/3atjraGAp6h52XNRCHldKfqSHVlTiUUCJOM4GVdDDmsKDjtosaoiexMh6dYa2lUEUDrXZGc5J0ftn8MxJcaf3G97/z2PKRbWSK/t1J/za/CQvkKKR//oqRCWTwwBde5PMsiPNRHLKefJSloVP+lF5wVsOeQ5I5e4icyrhnZYzGO81qu3E9y8pcx9ZlNUGWQvyFM12ZdM/Qa4S0iidfy4HyU71C5RAFKbpgGI5re4KKW5NRtf+su4xWzKIP/gYwFbVB/8FQm29pqLunz6PwiKSUnZ8b20DJWN2cdIa1/OAbglGRjVUWTm54kzhT+8gZy6VFRVzv2rzPPhO/ZDox91eFQXcXkK2CtZo/glIq4J9UWkxwdah87DNmJn6PcpdcN8nGBpgNWhNrqwwHs6x831DlFQTFjcx2P+/gXrRe3y0uNLrInCotrYTx8p7RZcRwu9XHtGueBZSJDNHPIeuob/YImttUqQcXO7vaf05aGY9+7f54mqVxU8QprqTNkW2JI9xD7YlmqfSIV/TZcsDFGMhCYeDRBiGtp2QIbeeT6BgGwtZWZUILEPesdIfBPlHlYGLrACnpks5nFvN4Vh4t6avG1cspnyLlEIpmpJ34dTDS3bP3iW2F3z4GeA6ZuuGxP7OiIzRnAHo61Vs40MT+NJy3CtgK/OJiZM1Aov+H8Jqh5M9Cxvo4yys3QbSF8FWJGnXWiESFcsHjsukq9lNbpCIsSWO/JXS6ZtOW/07cB7I/BaMGIn0uKQh/kfSoM044dG0GTtlX8nY6HlM7S69eGTMUHWg2P0HhiFPGzlY38kURyIGEOR4x6XoLKgajni/xnOitL40Q8JZr++rRyzjYSVQtIEw1j1W0HpdysKoIA8D4Yh+Duo94/CzN/dk/fn0FTk7sm9e98uxOrAZ3M8kQWxreL0ERnMWRNN4uZ/6HA6Dpm7UFTt7GdWk6LGrhxp4R17stcid8MBZA4Hery6q7dHGHnhgX6MvaSZkRXLHAMU+gqxHGK4PuGvRzVfT3CdH1THvtrKVdbC/Vx2jtld8d6scnyuhFuhALm4CZwXcKFmJSsdongG/1jYRQwaC5GD6djBKgvtzEOjbp4Ldz90AtCg8g4pSHqWS9Fu3sr7qHgVVoI3H1pIyjTwA6i+awOrkwrBz1kYbDxOf7cWG0XW8kR+gUw5oXi7j+KjD4gHPyuZZXyTIDGPwrS8tETfOIM9hdM40gFpW6gpHq7XBY/JGSGDtcn9ooVkEZCqHdsICO/X50mQvBJPllECJ0pplxiY5LF+vuosYny4CXJp0M0wp5wgg9Ulu/be0ZlfSsPlOUZBQB4SWg+5WBVL8lkkE8qP39E3IN4BECSaUMmNyHuj8zojWmljxJXizg9dVHA8ccRZ/HbOlDVf0zv6psA8bXJalslw2Rq3WThv9Lmdlbmb++bVGTvAmHgWiXZU5xJBovRNKg16AO0utR6xiQlFsta9pLdYwi8PioFGr2o+QHrsQoMFRQ/HXh7LTl6ethmku/WkA8oQ6Q4D3FM0K8r39WkBkoR0REzQvVp8wRudAQuW97Wdg1eouoP+WiV0BIVxwNBMpcuWGnxTpO39hzkvyVVnr/sZ1Ccxa8UKIR7GYrPtNolYhzGE+JKRSFc8xkk+xNUoI+rYnzwCwHUlePTtE97CMqybmxV2nZeHn7nFWnJyXFx7OovGEUopA38pFlBRiVGSi5dHCrWw1Eh38nrgT8spPB0Ak4/Y9uhcjoKBQj5xlVlpVEXyh+RM4/UIaM96WHrxgPU/kqyoCTlTBNJHrSsPwGAr0WHSl37C+qRkeOTNAkDn09yumreZO0m0lSKKpPoFLPY/edm+Bhu9LaT/QX4w3pNGuDdAE9o7NY6Z6E8Ahnx5awtGI8UcnSu4Bs+JPYx+FzAWjSKwmJf/Np6WbIuAO43IvOMBktoqrc1kCa9jqROTlCU9Vj1nFzBAX3KO/wplvkUNemuL0D5ji8447lcyIb3XKf4jjnnNxh/Cf8BytUmtkR0SpCpVElRyvVbIbMMg8JTDaV0H9ROg/OTJ7CVLPjtxqqmqX22wXsCr7oA03yVjCdYPsDnZHGNgNq68g40QjmBPQz5EGHHtnp/iPCYQLvodD6uQ6U6C6jZclSbVuxnaJ/Lb7BljCSZBbETUvgx99uHVGPnQl2XZJsAPyr9iF2UEFaucllhzYziSZgDgLqW5C4WAmSPTbwYXsMVpX9rjIFT76IYvFOnDS3FfIGtuYNFSSlV7sVvMgAmxjPNSaT8VgtdjOJiBhYR7vypQGHqhvM3kvgZIHWOtRQKOF+3PtpFq3Qmm3cpVdTsCBlWofst63hwugGudFqiRJZtRyrHpzGGPu45Nw2tpWYllOfYtoZRcvDAwACr1OgLD/De58AFMefdqEg32TaHXaG8IKw+mqXA5rrA9OwBM7d5Y20lT/1p2H2q8NBs7vi6X2Xap8Mt9aFcRVFbo9HjvvQvXRGi5ZYmwVC2Nssc02Vj3P49/nYV6p3qqTcB6CnsM03OIdtwagYEBB5IxvAIDoByO5f3qkI1xiiLyomPWGSbw8SzMccnjFOGYXo4hbsHGyHPIDDLloPCgPtj2+SqVf6KjTIstQvcd7si+DynfINPbRftall0bE6H+3GlbDNUIWQgrUg2UnC9sf6J8TDnZagaxetXzXEhY8RW1HVMiIcnTtR8pc5rNveYDr0kd/BQHkxVjx1I+yUXWvEcmTd8HM1Rc5gLc9Cdg7WlLZixbIFuse0gvSsQBIWJuRBrxFL5UbselaLjo8x6k5CRY6Ew+VCJ8ALrdlq6pau9pdH2HRIO/z7v5U90wLYEQfBeOcZecO/O5WrjUJGh2lyW9HmRTu1K5ObcQP7Z28bdVqObXPMQCx/XKGqU7NnXiQ61dAr3V8epn9Gn5pdG4I9680tmsfDRHuHwNhqQ4ntjHyvIpWzNuRhmB3cU1dwB42O9KcF6DCZuYXirl1F3y97wUeJPJUJawj2FHLesgTcOnjx7lqFrUx7GHSR4BcKqg67ho+EZ5Fr9p+IiirYkxEiQV8y2GEzAlH8x5sFphr2DjZxMEiKgh/K49wuglosUZ4P9UFYJP+kcojFNJIFNWlOhDFU6YWSPlW6OAub1plLVFGKJ7bY/sx4woFjTfNda4yYXhvgsp1g3PT+ix4dVgULEcC+ZGd9cQgjsz6qS8f4PTZnWJ7xfVoiBATKPLxY6DMQMS0rMKwvdcfMJrFDm/dGGBKf1oGOu6cna0hFsb9/MgfLeFWXdawfXhbKoFsQGGnmbyHVmZ0Sc8XKyC1JB/331ioQ4dNT1XKWyVD1wEch8rXjOkG3R7qDWGZKwwsURyCFTsFfxaHnoWp1+HrwuGofU0s+tvbN1siCgr0c1KszLpcncV1VgPIpsbaFnkKYH/cPh4LzzL4Z7nxCs7EAZl2+rgnQhgtKA/LS5fZqAK/veJEsvfKntkZcDNqsyNkj7mpKqQ5ELhjXhQx0Cu0+N09OhsLp4T2jV7fv+oCKPZcnaPoG3LDg4w2DARU9DjQmB6PBgorKfxD+bxU3cKruiyv7/VyeqEVn8mktIvbC+L9nwt6o//4IAGqFSYRJ4209ltmv0MyH1eAXrGNsHwp9cEl1OjEBK+l0YgGFysKn+DD0gEbCBuU1aYiUJhPm4P/kUIKwr1TiG/q73TsZTJsxlFtgQR8bSZKPszRAFX48P2GvVMkzLW72FweDLWbrl3Ow5ob+CrBouwk6JnErtHfyEvc/gKp8n16C4ceez10CwP38blwgU17WEiIS+A6RyvBt71ngQ0qH+9zInsdjtHteZg027Q/yqewqwvlcWuBtWGpw4YpJvKlUXgQzICaZFw6Nuyu2eRoZEZc6WTKsDQiJ41c8WDbqNFDm+0n1qnd1nRuqBE0Rym0FnRIm125LJyotKdoARykvwVLs3/FOnG/etoTZ0IdMedMjrq4fSV1oz2KVTl7SCkNehQlvo33oYPvMv69JtEtRUb1VCddigJ2bkiy/Qr3vtJXCXRfGHuhRS4VPp3q4Vvh78LoiexLIqtJOcCPyGqvfv8QnR+fX/aHRldywMJeLaam4nTWnKQsZrNedFYK80fE+oUMRKgRwlSBXSP+esiRwssCQA80iwNuPtUPdOdBQdbc982BlGwFhi8BUaTuOtOcFCdZuctd82t4h4REOojfoeDsCW0NA/flxE4Z6vIParXYYUfwkX00UzVK281uuAPLp7hiBRv16t+GLJqHRFmfIaTfdhb28kvA0iS04/TNgPKpD9aoAntpS838RfxyoMp+JD0ssdD14BQistZhgXlcNKfKMGZkhXLLK+jftw9+g6kEZjZoYM10/jO0sVQ3kQ1pwYOJLg6ZcvWOCD9e2AjGzZkBV6FBpJAgII1HYkZ797dFU9DcErNESN2MFguumVSoHvqni6UKZNkvAyvNLtbrDEBwIUzVrDWXvZWeOP6AqeB/DnDDMKdiAeVEWxiDhDZsjO/80Ej1t53XJVY644XNg/6Ddo5/qsTA5x2PYzS0mOSMEsEeVSbGh1+40YlhcoycPvxv9TTSdnW4VNIBYi/pBLsCnwrRLc+2h4kc3eoqclqm6jCjztIv9Vo1+04u9gHCVnX1HP9xatPxn3l79aLJSVd4o/7eQJUQsrH6VnPqsjTAAs0/zapkY9YwWJij27Yz2sa4bq3qBI7ALiOKHOGwbe925nW9c2pcUI/MBcQPJ+TRWqteMM0pTBt9NcCdVH2uuJBafgJ/enaC9c1/pgYuu4KIMwXje1Xr/jdT55Gc++DSQAIQSgXaqloPKhVPSr7sQVFEYJkiM1fYKSSBXCAnMO7mUM6W00izELuJRsosOOjhecbh/HYWMtFruerRaeHqcEKosmf76v0gSrc2OkB595cZp+wk2i04tFiVoeBCuxj5ZNC9Z9kLbmCCZgslL7JBMxEn8nzw+29P+I2W+OaCyZAwqpdDdSmtD4ZTkeo+tcArXUYV3DUPfAzcdbOUzdN89uQz+dQRhJQu1jZOncfryWfnFhvhygvx0mzpySj6zk+DNzWRRPQOjtFzojK57ls9kA+FszTEK2gY6WggpKL0mrMSzPl/STcAISOZoFnqCFceWq349kix7g5EoeXHUqOfeL4nx0T7E0KZ2WHN1Q2RcRIoMNwvj9SMszJu75aMS81s2kqCXHO6ayzFaSCw/VSDUTXyVoiTQnD4cBe55fww0DG84IUA+x8HZroNh85s5jjDycnf3N19F/u3XxPgOwG5vMytzQNAwarBOxD7ZYi92iou+wrRiVfaF6ika8LiK9jKsFVUbw4TpEMdgJ1YXWv6AepfnW7JEmquke3y4lVq7MgJ3NccY35YSkHUEMa7Ny1gOEt+Sv1gFuk2Bm8dsfSssC0=
`pragma protect end_data_block
`pragma protect digest_block
f9015c89104805d99ca00373b3d14c1ab732d045517d673ca628aa0aef9d26c9
`pragma protect end_digest_block
`pragma protect end_protected
