`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
l+uRB+15aNJrqxd8bOsncjXMICtcOpkT3JbBUF8K1BCKraw/yETl5cZP2ymU1qQ/52WVS6LyZ8S1o/aio5xNl+77CMzdWEZ5e5fVattnwrLxIRMWKYp/TIBycudNJcpxoc5BrNaSRgxPiZ2Mgn019Lyn9YjYlyS2kXkyqFgQyD71RT7MQ8dox3n7X0LOOEswY4nPTCj+lnFYt8YdN+Iablgajfe74bE5Vn7YF0KfH9a8pAHm90VlVyRuU7JIV+nAqBFYDsQA0a5DoS33WOwzvg5oOg5/x+C4eNFQM4eWNhblpevaFg6greW1TZAV4jAR9UNy8nBgXFXHrxtoy0qblZRyiK4nSYfmTQ4SU0URUplCqqrM1aI8NzAI+Y0Ok7jwblCjtzS+bgKVac+2fYTks8F7puOtP0opvLAAiWf6RHyHcj3paniPdBKqxnSovoPLiSCjyaoOgiBcK1peynl/UIhq5L2alczGRx043pW4k7fIGf6tlVGtRErhu7XF/9+Mch8oPFccgZ7AJHAGyH9GmOadDm3G//f6257krc6Yw6WE7B2/HbSyHSlqp1Xmz86/jGj+iPENK9TRze5CmQ/aUoa9OGzGzswhGh4MxeW75o0WsO9KJqrP/SWJVLkLAZnBSEJVwl8Wep9ysLGvHeogIJBv7euhShQEhQwakyX8MDbp+5rvHrNcDwonrqI1eMBowfrtWngn/lo5BY3GXcy/SwXLx5fMH3Jwve/J6GNkuNWcGvvPVEj+GJkPvx6VH/w3LpiXoKRXEM1Vrm+zwdKKQyJFwsivwSc8exQOae85dhgsH64RvWmo0UUxDyGCpx0It4kWYJlVY6zuxhCH3ZjGBhIctkcInpPuSbmwx0YWKD7t1rc5cWDlF2wi6Tqg+rga2XfP0O6XbBuXHI4DxibBkyM5Js5YqhHFzPj3RdslUNHylKzopCuXOVM0LpT3DRklz8skoXV0ZZEL6iaHPCE2C3e2bYM3UoZSmRDSRQUTWuFPyAzaGs8eRbim2VkJPcMvVXpUVMzzknz9VQGDtQz2NHSlkO1dvgQkFsn9+uDZJ+ye8os4h4V9aeyg1rSNMNjAXTcN3NML0ZpCsobOVHXirWZESXzqK5NwbnWfyDf0O0SOkWFhcwD9/MpJJ2e3lgbWkLIrTQityhElBhf/jYQjcs4fJs6LAJxmKjRtJ1TJXRXDylr/aPyjREZaa1d/elA74Y8uFELK9s/1QWU0PBCq4byLvQ75tiIdN8lD4DoTVFpnJ+EyJDU95kiRYyr5lDNRS1zqu5j8lF1/a+XBk3MitrCZJTh8ihq799LpcLeN97cpxEkZ2xCb8RPSfiL0yrjmHImCeHB+GCJKf7gOz6Q1lhpPVT+6NAu8egVOCpyTB4HS1xI9bs59O4SokLhRSK41m855f7AxXoblOoSC6cDj9wmAkYl6PqmiArxVImqvXe3rtFcUGhGsvCw2gEeA96/8zel/E9q93paMrvqar93kBfybHaH1Usj6EylLkSy/OkoLl+2UUqDvjljz2iltUxggMSjtDjl6GdHr5T1HEzRbugt/96h+pMBlNyQHSTThykO5obFMUtlYwveJpHXU4ldzy+4UiNMRG5KFXeduJlZ1Iq2W7da6QxElYBPstiU5OdZVSSy1IbQilg0C/p9iLCCwIoRaJ+L3N44K1oZu9537rbc5WgE2Xg7CpaJkfbOZiUKwWhvvgUqrDAMAHwnWmBgi/Rd5GufhryoqML3JmIek95TqQ/rs7if8YCDrv8MyycL9wFxFg8UqNGEsCyTSJT6xafmYY+QBYJ/NurYtZzewr31lf3d4554YNMQncmYXE2CNvTQWhe70QexYxJYy7MCjjXARcPRLxz/og8oADVv/q6tn2Aa44KLE5/QQIRCEBgpKfMhy1g0PvLsKz/CPFpcG/8ySJFiMvgO1Jat3Nu5M1XsKYrir6MOYT1r86nOtIYgNs2/89+rWIGYpOqiL/Yu2g1wyiMB+nUGvjtSBWqA9eVk2DIKGLw8SgVziEqujutKj6nYkmjucrQwuo3bCpRMiTK/sHTkodm9i6DLMecdm9g/7nh7C8TQVMYJtUjnja1dYCUerjL4csOthyNoCKHb6yAhlZcS7mIUMhrTJLk+HoG9EX7zndcCRsd8btmsGrpmbf0/UnuAkQ4MMjkWx2e3wpXTYbWirfd/46C9sqFoKeyHOs/svWI9EJgqXyARXjBoaw8oclxXEvtxqaHz90dIw7Nb9/PxyYfbkYhgsRRyzHvhhBWsm3FZKIk3iB2rGg5Xhm5+CJLWBqx57BCIWo9Rb6GkRUpPIxdVbEWuHOI8grtNq2SEZ8F8e/cXeJ7F0oGzchC142btEQwoTaDnlYZGRGdG0z8vtOO23TbsK1Bn9KAeqlfstT98sZq5ehGSWhLvrJHUlinAycYi8znhpm4Of+4ZzlPS/SaVe7UEUa5qIxCHnYYRZ5dfffxh2mZwJgxxO58Qx6Retd36EiZJJh29Cb225h27Dufnq6+1BpY1qMY/Bq/PSS70sNF14iMRfl0oircuaOBv2uCRx2UC92Id0yw2TAmYdjJf/ov8lS3ewmK37e01eKYFMIA2ZnkJWxw/D6bUlJAqnsQtPckx+YelpUZf7LKn5UpJXi64FnwlPu+MleWE7fxoob4fqwKQif8vPlI8/hGhB3UfheFW87TOzpH5Vwkf7nuRFsbp2TU5NPgYAfSCbH20EiRF7dWQ19fUBAYMgYZevbs5V2rIKNgJqSU7A546UySSRlmRSlKd4D/Ek47XX3s9w0WFujzHZFhPaDtSCBZey7L2LG78MsUwidRs/m8eAo6d29RQLK4V1f+hPTqnfULb9C5oveg29rEUBM0JiDrx29jI57CN7AhJHKRa4VOMjKt8IfTppYNdQi1Kre9REBK0WKwTKx3R7P6SRz1UaOGSZf7w9XX3GJAhqDpDLxgFXDvMEJBw+Jc+ZDHDRcDFzb3oPQcBMqTH57+nPv7ACKAHOGUDxlGgmw3O/IgK4QyvSae0cOCJoMVaJcpqCOWlXzDAyePtZsG72fQZXY3PnYMR3KCNmSC3X2LCqCr1al6LYpzl6wgD1+A1cRfwgSoifV3xVZqrPNCfPETKhyg3mP7L1pxcQ37PhN1V7ZU83NirHpihBRIZWo2QJbmn82fGZMJNvtzIvJhAUlbl7696HQ2Sz21KPz8gfRD+C/lggZlhdE9C8zveaytt1+D/iISwAGPow3r3kFK4RYJGyjSgm7sv7u9eTR5v+0rakFtMbAVHzQLN0tQY/YAgIPJpu4JRGg/Kr+JU74PXwnNRmnOK5PutFr6CzvaCuXQZbzQBCboBTUOvyRtWkdKWnBJQETF44ZZ+5XL8lmx9YUiVohdnmgsRkwjC4OMu3FhTy9+fezaGKqUljYWeIZd+KvcBqb3JxvBqjPR/T+dhCsmHqlbyjFm7RehGSJ1R7wdkOUxRupm1W/dsBq1Qn7pqHdU5NmITw/6z2XbOkSrHFsqIAgZNgiIwI4HLM3QQBnXidh6JJ4ID1GPYSiMaVXBTIGzJGYmZGCViMLSyclUmL4DqkQ8yiv2B8dNbCziGhH+gpDUBqmFbpPRzj0nkTjpo/4q+GbLaS/ddAUVPYSdJpv01D3Ycy3ssgp/5HtKNwjAbeAko30I+NCds35fhj3v5oheNowMiuOKYBu7kJblCyX3XARcIEhUrP8ZrB8Mwo1ys9YXL7sZ2YEQoHY9Jac0mGIskkBd2Twa85RYNnFuoAtY/DQIZ7RPWvdFlpvHoAETATwBlZ3JhE8aqhHZWt5N0myRhWMH/Yf7lf1OkmN6lw4ccmT1Ure6Ckz2ST0auUZ/a9wQoYOQ8VMpR0MtiBMZ4enagq23k9MKJM98b6qKdZ5u1etfI5KggzmWsgQnKK3lK1xCrKhZ5l+hAsdwXHwx2ZZL/EwWoHLvVqFoazrPiCfA/bIQ1rxrXpY4W+F8RttfV5OURRJ2h/Kudab+3kRCPn1VxCZIHnvi6ziozwWrJwG8l7sK/Uy61LO/pGBLDbm4YmHw+EBB0Ab2uLLSjdg7BMg/aVkolQivxtJUl+4oTv0zpgYAT8N5zn9qSbeJZB+m2Qu0Ma8SqiOav5xvXb1SAYSMaN7tSYxw2eT5A23T7NqfRzM3mYEG3JcR20PzauP/W2akY+kQV9MyMlMiQrbaoM9tYzL3OT8diLTNxz2kBCRIw50X/WAI8HVkjAVgUg8B6k3XhkTxTJ1p3oY1ZCjT+GDBdxPFnKQzohz590wfvpLPgSpM8khljSIqFlat0djKxTm5XFT9JqvfhmUgRVeONgSGjHNaW+diBYETxsCQn9gg4++k0WFKZuNj62n79mgj3vbChU7Q8ivzf44diQEAitXUJKtnM/6H3NAZZj5OX5kwdCdFLtxLtfSqR//DTxz9ySmZscrwX+ahVyMPRBS3V3EkDtc8ZkDu5RKisZvdnxqn0VvjeiXGVGVzSwOSt9TKDD1xfsSf6tWjKfh3dKVAUNIpSL7G9GYk70EbatnYj9qunvEU4pqeQwt97a+USGdrcOCK9PdRTDX8W4q9hOdXE6bxvvwwDgJIEogYDT3rOzW+9FUahjb9ygfMtm/f7iYxFRiIl1AHoLz7ikvrlSYORSYWjsYT5pT4ITYLU6N/e76faNG3PiChDHALsd8h28uLiSpjIfbB7u2gh3tspICxcZW8tMtZdtcjt1l/FcOO0ueBfI1cZ2TnsalhPT6W9Dr8N1IfmviZf8M2pKdB5zF869ox4+dOz97q4+2uCuyaJzDxli2A8PKUqZClxPkqrPQtQcMK0lnL7Ayl4cxrl9EycpfGPYjXc81yKXgoWpxthVl7XBr+647W+sXlLAWIWb0KNWBxaPs2WQfQCQJCozBbUVyk9PBwt6JBMIn2CdFM++abvDrw+Z8kXAKIcLVR0AbJtDnCogv/O8lDDk8WGkQC73NLGrKNjJE4SO9MXjesm2BFGpGDCtSnpfEu/5S+XZxvUzxvRQ2FoyOEidZEQxE/nNlF/w3nc33rYIpvnaEoEdRnPnu5j9lV69FwbdEFwab6jm1jwI9V++JFdD3Ir9lupn0xeKjkgrzxoLT8nqAJtvgmqYsiw/J5Xt7pPQK9ieUAW6E9RQsiLjd/bJwoMPX+vTHSCPxsvjQXS2dg2HhNqfL7PCXsvw7ZnxoGoFdM4JrtMvlNZ2wbhNFxavk+FM440/vh8et1mdt/+dDUMENPnsY8Gatcrycmk+KzBVGeJG8f3i8cOHuzwAmEHsTKM7JzjoLh5zKTQAcfDqbOOql+T0NqGjZR2fPVOuw4bWol8mXqXhk+Ev9kAy7x9XSpSZIkwMfDynSr1buPpz5UoWNbylxoYmPa6iliHZ1mvM5fLwyIXPvAXU7rnIFKd35dxOWAJnPPvUHvR0O+TzLeQt1Ge3P0r248o+nWfWwNK87V9pT57lhRdG2hGK+upingxT76qCpRNalWhquQ39Z5+mVSKm+JVc0vMeqLuIMMgW7zuGYY3Iif6FnI2gq3fwJCq1IKcqBE63TcXF2NwXITOTkjM8wiJzQTe2RxRpTMgxMZZMLXk8o6skjA1gRvtaT5uWgymSAP8aezq3Od+zqBAR89xpxhDls8litQma9No4YI7UTaaYZEk5pTB4u88K/NwW/VbNclDNMO4ydiGEfqswhD+aKI0dwAZ+MgI1OXki+GkG/PxB81N72c7toMOQ2BeiJw1KJkx8iQJ0v8cZnNCKFof0qrLy1XBe8/7qNpiu+eu3SOSy3bxv/9DDj5jJK2tbpO/5BqpvkcjAPvXmeJWq3DALyxMDkAyxLJenko2MDUYWIBpnnn9adS8ZXsg6AAbRECz67uPE613dWkoscc1aONKXs9rXLaZF3G7z3nIPeBd28urAV21lCVBoikGzaoP4xs1NGnu3QiTAwdQjhs9uFl9EgW5gbw3CqG4rBVqaVNAS8GiLOBDJkn5w5Uu7XW49KHqLXlHafvv4mcXlEV3b7Nh2HdIEvJAIY/sYCgSbKLck1JXC6yg6fl0TzjHmWiN1rMb2nbXhAqBDmzBBz7ZNcBsKvimG7hPNu1lAF/ICY2sl52vsJ71cRHpCxJc4f8mECwiAVn03fOfZITZ1tm+Ut9ekxpcdAy9FckZOOsBrBMqog9XaIrRZ9z3xVlqwFFCQHrdefxRVGkYVwp6L0AMabyYTNtbi39/fcbBIHzsvfYq4unPPYmLCBoDhmRmTV9/b1A6rHMGS+HF7rp2DPNSFF0iaOYfSR172HGqYfGz+osAWhWt5srFyk9UsKSf6oy1vTVAxbK9b5V4HdtybYNcLIBiR3jXUk9iXBuHCeTjVNhmDamEKlauLuLbQf0Fj5+3l02Su53szo4n4ss82tU73mVUAsHj41xZ1e2BeEyQJC+VAf6MQ9WgqDuGiQilxFg4Rl5p6ZWuphR962Ise0LgPMV6Quohpctw7IIPyflEXDMGSQUXgcMWA9dUVtAIAqpqhfZ3ECPtq7Zk7+hTLSVEHCkUSWf2om3sc6QqWqCGHrEAwJDgZLGuJAV8Wz+haAXtb98bqbtELGUIbpq4h+4vOC0dAnNPlzFSMGBIfqqekMn0n/RxUSe218q4/v1q5d9itbPGORQnmDI205P3JyNOiCWvGOzLeVi6KjFIWOIzqgvCK3Gah94t5DvRvjOE7inlxtNrvIVYCdJt2XHmlmWfaSIANKf7CsG3hWl3O0iKEK6RHV79+1egXL+IEGVEeISrr7OHW8Ts89wOCE3rpm9Q8Ia7sc+G8AACuGBGyK5dapGYT6Odja/PabKBkWaoVMChuNbWjgYknvej+j7JpgGlPhBc8BsDDkCK5+k/z2qBsj6p7gBfSrdfjOClThTtgeN5eFkigvAssi0Nak5KoHsyxiheoTjZAmBtCa8x9TVeohotWktYwjWKv67Ih9lCaHRvkuCc/Btbk8iSX6YAUpnLHSKvpVBtmIkSzMyTb50JBQJcdTThx0k1vrwWp3iDF9Z+d6i1gIaQXqlywNo1UXJILpI0n8C0Nsc8o7Z9LAVvbQmpJ6b3kDTdCXP/TfoLlzKa40rO6gpD4gKMijfqGMTPDlXSzxM9rMGDOfDX3T8XcRpMJHwCtZTgep5HWypHo19nkTYR+wSF57EakkiMsJicMRMBJGjVK2jWQXh1XQofbxNhLPHzU/mAUsECaw2gyXydbZ1e8M/Doc6gp6T8aZ9CjH/bBy7Lu93/vPjW4j0HA9ICYAWbd/2IfpJkGgVXzHUv61lMjLLYWclDovgA2R29U3Imm39u/ie4NBEgTQziEpt8QgbpMVlApCw8+WfD8qF1rK69HYQDA0CK2ipC7WTun0xryG1gG+wAoJNJGhqULSN3UsLQJ3+Q53PsppOjHhnvgPIFtLJi2osh80G25NGWUl+ag6ZuhzncCX1Ns8OEKf73UZyEbDduaKwFantd5cEyyFuQ54C/SPx8BYDPOZrakPS20+42SQ0RXT9oaLVVbX13Lytk6XA14cKCjLCTBnbsNnYiCKUW33x5Hk+QetUA9eGY821xm0kyCZs82K1JBORfbJ3Qp9/bFPoipGnkcGG7V2Z2sI0j+TXduV/0+j8mUIIRxp1nWcrfWVxY9EQUmsKJ9mmz4KhN335iyZjv8BBBmuqKA3k4tER5Uu4QoCec4PQmlOZT4kJRKFUv+MDHFdYrxIA2ArNrwGqdDAUKwyaa3Pw4i9QrXz/8q+4hUf4gTpnwvEWTqjr/2IXlooO3FYKsQPrBanGV1xxqnpVBkD+yTh5G/j9VI9+C4rCPVSpA6pXb2zB6H0g78d0xIWfN8cXyWz8376rk7X64lhKXTCITZzo89QW3fNKrKe4p76Qpw3RA118QHSn3eeu3rFo+QPs2nblpcE7YEizPn6hipwENqALDYR2cRJh+WarefO3TdrIVa4v34jaJFFhsEgXeQdwGwTxshOePA2fWYugXTOIv1X6UA65QXvCCK719xRk2KhCqpE2vlcZSDAd8J87B6A64c+cIeLHVk4QY6IzC1EOgBwQF+nkayGDoAji4CD44LaB9QMV572MMUVW8SticHE7PVrEUjn6TMSZJL12sy2c7WlZc2hNvEhYdy5Nnk5MdTtb/4AGmoFsdbNj4do7XVvBqsyml28zbOnqzUCTt2o1LVMlGvAmGesajp3eEmV3/N2SEwji7Y/IcrJZby6nrnBtbyJFR5Uw/u1mpoG9bbdaXqAKVBd7rcPbf81Sb5u7qVGGXtnAe18+5fjY9yHn1YN1bo5gmHopRwbuPj7j734AyyRwQJ/ZjW4KNeJRembVo8UVsjFl8HtespwLVZi+jRbXnqmu2pQoe5nRsCv79b6UTdKofGMQNt5Y3Ovm6bGLAyXTh8wMd8mM0qZvt7akfM04NuyMxrpBxfrDV0abfRaYEf3u34dD/2SgwFxMakbPpO6BNtddFrehev4KLjuEuE1e68bmGEsjI/j6O40O9N8lVw5o0q7vOs+xQdHT5xb8TBv6kJ/dBcveijwuHDBf7YQg+BBfoIa8kg/oh+Z2e52LAP7hTMfFIWKSzIZ1A6lPAekVQ7CflsPT7GjHO8IgwSZ5uY5XSBU2h75/taqxYuCpijt2JfEtDMTL3zk5CQmv30Vc6O8uekHN/w/8eAkeRhxPIZs85altzc/Mby/HYghXRTKIo8rJn8SZOHMi5u7YM2DbzVdO/8VEQ97Y+JjAoLVHLuBvZ/2WXEbBMm+0uwasRPR13hYkrBHaPj8Y7LNnbzbH2eaEsX7G/RMKnKrTcwgH9Z8+zEKRnVr3VSAknig/v2nR21wujwFUavnrjiZ+0dXZnaWWbnfJ/ArzJGL+hydGmNVyA9JuW/LPhh0J9fTxnYGEPjWfkFFI1ogx9YPUcvic7jhcCXc0ccue1dFTTJmvA9ImpvXUHIZT4IdQvsNri1v6JjI0rMcKjNMjPZoCc4PL9acKcjpCR4tD4xEhLUkqhoDR9F8+MSBEkPgWqpLuqIvGpptpsiAFgQjKrdLyLoP8XWeN15AbkJIu3nG3s2PQ81SmKzApZ9xWt60S2LPX/rqxfZALZnymk/63P+OA6kuwXLw4XmSH5cmxwolc393SSCGpNShYgyTBPd+KhUOg6KlBz9+n5UQp76HWQSjJMKs92g7DKhd0kkw/ugOVFW7IedreNIE++wZV3Zifu7MkwF7nSgTXqWwVGpm6h9ojEibu18iQNggJx4gC0QwcNZo5RloMvLkkwFC3VjGKbK5CXamxjkdy3Z/VEKwl3/Bh9DVWUmUDdpycBdnT38yt0Ns+DEZICb/M+wuFEexp5Pv35WoCuhpGpViTB42XezIHA0CnkknMgTSG/t+W8QRXJlkcGjW0tg9hKG2bHCat6TyXNDIis4Bdgwmxwmv1JmFUBrmZJrGOLDV44lvvtqqM3OcvUlxbGbqKIpnhVGdZ4emEZZlDRUKB1v4HWPCJ9FmWW+IpsZfpGfksbEoheIeg2/jBr2zAJVyHfpwxvXv6DwX4NlbTQXRIxVr9x60EWipUJ+n67XEtq28K9zXv1IGhKNIMtrkwO229R/u+VRN+lsOTYC1ogj84Go5mnSkJjEmqYCupYCmy2WgAtdfwtjNAyZiFGo0u+UjneOHf5e9klGm5nmIQZK3iB0hS9tWZqTb8V7vzsxza6Br3q00emdgdByhKqmwc1hUtQRowCheJqTRxpq1EH69a06QENKrERbBOs16UAIXczupCEFz6BvJU3PoNuZJQnQ129HrsburBhXRqrHEYIdJyvtABlds+Zg/AhyXuNS6vizrdavPTP6evMJQaZsw5Y6sA+b+p1BFA8FvDjRyyC76HTbuFmd4mAPwKl3C26SvYaesTBIOLl5YOSpJ3HNTa0WCO9VXJ46pnaMS7kshVRf+NkIpXFNFYg6FcaxcSxECdmAzzIuvF3D2YMYeyDPh9cakwCDOPEnzLtnzf+i6lqxL4nNztH9lwg2iYZ+sQPcq7O65Q4i0kxOpma4pClvcspQ/aSbRwT76v8P7YnTlMHzCY2n4sn+XU39qNLzLQgdLrqzGTOEx52SDOOjzim1esNmIH5b7C3JzWGMbxvmNhN3PP5DtRPuYYPsQM3/SjRYRf/yqQV81Y7Gi/MgNLMFGcwyhcGKPK7IVYWolxFTI48x495MZiR6Mv0c4HhInVtEnBo57R3pTZpFF3aadQaijdZvY2SBPnxTWpNW5ZXEKep1NBraKeFA2D230oT/a0D8SfZFSAVT8u/gv0kWE6BghQqQawMk++12r/v7jtg1D3AKn2JRYGasKPnJkSZElVWZcuTAAt1tCSrcgAzfqwc01ALU3P2lTALEkG2gQ7vGNj/Iz/BLqTQX5vMfH6a+xSuA8I1xmb77vK7FqQj5PaecbEdtvl94r5rWAWK8AiTJvH0il280Dm7ZqsBw8py0W9CWhCWiuGjNqWMyBhUs7xM++tiZbntEy+H4NFuQ40UDGus7+bpOGzsCpPP2UmAG+glDXxqe2tp2wFYQNGJOqATOrHjm5EzlXRSTfUNSSPrtejJiJyBsRqNZjCunSX1plGyPQw2sejtCTX7RGqaH1j+CsO2UJh8ccOTeCgmTk1QHqhLjT5x5Csemvc5aKVvF20RMRvZjUDD5brKmXTrAXeBISz5zTdNVjCEw95VovQCbzANrL6k9rmXXyZqmti48392IviiUO7lnwVyvA1L+QzHByNOHyBJbnW08ILSMSS/z9bNQPeSk7DRe3Eny63IbiTnRvC//hFEEmmDsYLOPVdtEDJjZuiwn8ucNCIB1T4YiVSZRt+8h5qJ1spamtQtEGHaLUrtwBTZFWFS48LN8UwhypNE9Ip2ZZkrQTK96p1NfgXLLEgp0uPIp0jY7+8J66tFtvWSDEoedEd1sCZIVtG0L0Npy+59ZfOBM2Ul8TojTd9rjh+FTQIbHscOut7yMwKp80lW38jGbFMCvhUTyLep8cnsdMDpAyE4+sIUL20XTNvYoFn1gWex+baCsglzPCrVhoDHK81V5mll/YFL3CgRsk6jlkKsv9jwuOhcz7FRkMldYkldQSJO4PqGNixK9tTwT0zvDhKOt8O3JnTg6jqt/mQepT1EjEzkHkrAog+8fmdTxdQ38Ye8GmcnlMo71NHSeHr3rtuaL5jd8J+CAhH8BlNpMoOvLvIBKJL/Ex+/731ix0KKCuSKtWiTCsDGs37uJxjY0ScPZ02WzvfWhjbrDmRvKnLAHUmotv14SEnk9DwzBtMyMfCJzRf4YfhoFwPxGHEz3WepTh7IszMuS5+SmUuXVLQmOSlBg7+b7SS930XMeffeg47GD2Ln0IHT+FP33pmg6lW01ds8k14tZ+Ny5IkUO1qeYN+Z0yxq2I6wjKfiC6ELYTXsmy0dKmLR1pxqXZ4nlBhJglnB+ZE/J4c2lgluFP1K6/uTjsxCDXUosMzuNABEGgZMH6+xGh8p8mBrvplqOIA/s1ku55Elxv7b3webMriEWju0EKBZ/h8TNYWrlJocf0Bmay4P2OovAEQd7iDZNteNm7HZsdfwALzaybofvr6qSOWhTpqneMQ/CtOFUXspUjZ7fPlFU6UAb53z4yJXbgIHqbIPpFnu9vAhZnvRQkInycrCANpXFC9o4MpEZlLjrALPisJXlpH9dFV8NT/w63D1mAgzvK0yOmsqdpCJJr2Z9cnuw2HKaC15docydmIfp62gOjIitcfVX6Gb71Emu3pi2f4Rlm6HlatNISNEMFPKX+8MuDFB3vsq8t2ZnN06ZXL2duh6fqiVcpBjZqrHRB1JyMbQUKyKResiWVh5Njr4b9TNSfVdTSXgnoakERP+SSOJuPF2NvoYS959bUWfJovAzm/bVG6u0nq3Ex5YpUFLqmhS9VytVgzBE86jjI/O9ZlwrizMcd6/xKE+DB4vran35yQmEQNxY5k+kkR1Io3r/sUUnqWfvBbVKNL1RN+iEx7vIRht8agH4w0v47kqHKBnIJN8TJ/Ni1c4KEVHs2PEeiBzuq4wbyh62Tc0TJjn8ITRTLCTykr/+aIINSFKp5P12RtH9Cqhxbzdxtf3ulw0ZMWbudQ1byCXpnQTSO//Yno98yCSBLWpXzM9CuaMo2+kYOBav0vI5BhQIXWg57y2ps20ZPGvnnKkwsNCDuqjkl0I7/z/yLBk1ftpq2L4UOYya3xOp3w58uwRCIDIM0uhQwtew4YmJhsFCH6tzAhnLkcfrUihHcXOEnRE8yvA0Igi6DGhjLEDEg8fQJAGx2H/b58wRrB3Gzd4RO/Nd5WCM8FVV1NgY851Gn/s9q6/8wMpKn8K2pqmNQl5n3DsHbSHp5ICK5OjGWktiEiJR7p8KofniWBIOjV4fBG0GAIrVURK3GQdfIsgKoGlpw7t1AF/QA+n5gs+zOOu/ZvzNCosuzxwqm0UbAQLvBXpVbl1CXdgcjKcSDeSZeLdgHLpNeVl4idNd9dHsEWtcWEN9U3aBOfr2Ej4RDvhoZaN43EDcIXbdxgV3sUsrnZFjQOdwdiqxeuDZkYy1GatkTpbd4IhK5ENnKxpcI9e5HcMy5mG8PZjLcu6yE2QXpMGWrxTu6oTjogwiWoOYOthbCNcj+0+GI1eS/0xw2Ky04Okr4BMoHvlKmELPjfV1IwLf1MxeuOG+CL332FzkHvIRXHx8xnW077wsfqvn89nTmYJyczkwmFbtkAafv9nJX9vHy1KhmK4W9FO+Z7uNLxEIdoTpCz9/2zfkFTYA/3sQzkTrHlcCf/GLgaIFk1d2fweJwZ0d4s6DzhL188Z0ZqTknKSCbkCvDbOwprAZTNBSVWH3r9UxrJa6u0DOsg1tRQbg6dtgKbMAgPcQFOD/oOVUyO6v3OIMkhQVEs/mPNsGn74+m6beSvfnbq0cKoQFX1k+XOmskHAS3K0dcvy2Y403r3/n1/lxU+0hAOnPiOR/Az0BLIoMAPLRfUY/R9COp0MtVggxd6dw4rV6nT7mKsKYpdL2t95gtXrFbALgn9QjQFfbNNORC47jq8wKEyYTPzUc2lsSTUFiVzoOh1oBexQYgXVni8pYEWDqcI2E1X1MrjrVkq55RD2y6X5z7CW9PkpSoJEOL8sMTwEJIi9EsHVmMaYVOdK0YZAAPHdw8+otApr5bpeUcLu2YnqkPZBGIRbEy8whaPYEZudLw71VX/v6XqTPjGMZUur3sRW104in45jXvTMuo8ZMld673ZGFkdO5rrP9ggCw7TSQxfKAEqKNntylBUiOAUjxiyJ0MNpVGB3PYYSf6qzdIe5Ooq6OyrumQ5KEq39xgQYXp7NsTItvz5D77cp9PMJQnyE4jvFS6MLu5sdMzfRV4YZ9zgQRFubHG+QfqXZqrQfJXS1r4RnnEtFyo5J9SG8J+AnamJBcCZa19eabWLXL3LP+C8KgaGz++6HBX3/GYFG1wvXnaM0WwJFWZeeXXy7D1USa/sY/prOjoE8v+WmiVeICLOGXrb2waX2Zuiy1T/MuJRTzjgJS9oWv9SXn4MBPiWnUTY0iNA0pWC4I68KdG43PPDnxgPXhBIh26QyXVCFcq49XoSCP0afHWSiSNyT5aj6waGLzAJKiSf/d3FHOZj7PX6PkGLqIzWro69G7WG9/rjPow8+qAeTECJ7sUEu0VyqjLcUmTNBcHHsdnGPZRB21H0ZL5mX67BqI/a1wwRUymsII+5AT9fRLa8tEkGrKc5asAneAEtOKHgpeyPy+s+LdzpIg6s/hh6Pdola45eJK1t69tRUGBMpRDnBwWbKtBlu5TeDxUw8C6lVkoEdm+BFiWEtEtCYcOXDfKcDWFHJ1TvTATo3vrqjoMGz6Nigj8A+yIXCRnyEtJlOU4oTiomJ9qUfn2YqpthRJLdetja88EFA0vHvF1MQ1M4S5WXape/P+4XyNu2lmbQXsQd0fea5YAesuCbDq7HBr+BFKV9lG3x2q/UaH1JhvMPlUgllx9ix75ZeVUkg9iRJRk9PyDNwDOR7jTkvbC6u+H79uGXQVe7Hiet+i93YmeVMhdksvtDEqz5YcGNUX8Wzhahy95SWHWPclqFWnIkQbdsODKwLx4+tsdi3wi6zyBmDQwsfinTCE7t0uR/QmbuvVZ3LjXcztzhZDmN1G37hu2Z5pJXYwPkMITwwtHFiWiOM+xgCWqUj5nTX4oI7rEPHyqMCJqExRcyGPVZ2/s0On4253dkUR4W5NDK7JLJcEOPF1YD444SuObcfvoCbQ76wW4T355PG9p/d9nIMnxoyeLjxrdCC92r/uBaKaUTdzSOe5PE5o2Bapdk07PDVBTJuzrkEszxDnxc950vql3pmPqpTOw60F7s0EOmrRWyvnftGEjLZFJbnHPnsRHt1pBpaHSMh2AoM5R1zk8fsvnwMqyFM8Cipj0xJzCStofMDxJAu2ffysrPh9ZzMGX0kSr8Jacyy417GoJr5yvn0JF3b1vT0EBxxfjx069OTKdHuk9g2Np0A2t8PzpudVZI0QlvdkovrkZAfHpyeYlJyPdrZf3a5Gr6n4I4u+Swas7YhbOZ2jduHIZSanmTMXTVu0qvbzto8RM5ijNKEyEoAKX6ybz/Yl8NC1D8LXM5OcnUE+gvmAh1wJ07wuIkaHvyjB+T1PZZo5HNIRUubfU1PcwAHABVcuCsQg9K+dcRXdUDrGCkxYAJrn3hWP+xlbBqK+5P4HZfL1Xx04v/D77F10WQpdIGOayYfOoHRUN5GmM2xT8PGPY+ErT2IJc5BqFGdgRZe8lK+XV45sAbSmThge1I562rwvDEcDycrL9uf5jcFgSromeECVpOrGNiiYu1M5kItB1XEo7CtxKQAtu4mTdKO9B0kUGOx7yYTL33Vv8tHvm1ILn6Y7l+Aexj0rmwaP+Y1Zvfh2098H0zMr0cY8snjuue4jlpL8PVogDh1Yj1Q96fs8aPlINj2zKYS4S7AcwBwQNymmTvgREHbjKKOjd+Eu9sRMk9CMR0r5L6FXenXXNjdtqsWHdJzwvUbB2tbIzCrR4GNluXE0UQzU3GdOE40QnC8KZ0d4R3u1si9jr3/8hAGWwmBvlYa9hYfSoudwZ2oybhKL4PatzKbTmHAqJxKaUjvWNw7px/pAqO/hx6rxKXTkT80Qd5uU3jUe2S9g06XVKlAA11GCZ99Wb+Y2HOdsQsoSqrQLaL4mHqLmuo3cQOHy82nPyC7lO6q5Lkcu+5FF0iMLF19cf1dbl57Z75F09izWc2AvE23N7GdNDDy1PO0Ai5/ED/hGUCDRLcZ0lhfhoDTJYTwDEWiiTrjubHAATVwUAl2RHisNMoxLS9W+9NClaOFI8iJkmgiPtw+tFw7b1SWxWIa3eOZSfqNwjny40YGtICEibs8Vf64pDwiFO+Wj8O3tLBUbW3SdHvppcnrXRxBoK+cNWi3Abh1rWlsfaFje0VLB7OZ1pJY++SdpX/GK9xWUTYPVJKjUvNQIGsa5hBs1MlxEWue+DOpqz1n6bnYbXdQ4VzBdCjlsGWa0XVAqigQOXV4a+CFasxQTnhlQ1XdtH8GWikyI3SSYGFO86+ow8eGUYBuIw6Rm6Q6pdiFtX4blNR59fVuhwdT5c6XLmtpD8kFS7O40bseS1P/yHTokVxq6eYOr3zASUdj+KL5tbiNaXs12KYERXRI564U+QoXl0AaZsut7rxDcejUrx+7IoRUqEC1MwCJ8B+VcAWActGgvKEENwc+HPWeC9/OkNzCLgfMkYHj2RhoTfI2IqP9d1rqkbkPgWq+vGS0QiN160piaa/8cm4YWFeMEPco+AhpkCllNuvUbk/uOc1NCWDq8u0T0NfNs9cb+mO6gJxZm603wCCIpvURdwOOiNW0PrT+cnCMbG+G09VU88pIi2STQZyhE35snYioyR6+beyHOUbd2MzeIgzh/HcJfqhaI/7fZFEoDksq9MFY2wtg3DE8E5RTfZG9hM7oPxW91lxeDywwE0055Bpy+Mh4hWFjLqRacppx7PTGTyLrDkDJJ2Y3uHTvW7QZHvvQ8AlJhrp17dBSFWNl72BjuqkoAabqy+LLT/0up6b9gbEBGopJULOD264VrLwPSifkvuu/39lbiBESbjYvN+jKQVrXgxhItZfi5G1DRjZf6lTVxGKBfYx0bul+3wC/8Xhh2WLv6wRSL7JZTvZs8Jy7fURNc7AuxfoJwfnkQVNBGLH9ffITnIc3+xZfY4I5i5oU2XedVZLk5x2gLLU0vWhbFVHyudoMqJ7b/9i1bFZVxydTb6AnAdkTFc4PsxnnGwiqakEak3TZzv+VlO03yI8ex+N5XcWC5NzziqoYwU5Y6x8UHn43wBNmdi8v5qBESAPj6oLZvD7YBV8lxCE9ieku+2NWUm/KfF/B7t1cCWcs/LuHJwV0V5D8LmHeNezgQ7wziT640nqEUeNW2+lDx0OqiOtdei3W9SgLFfh+0W30hmJvqQCf3FEsk0RJ/oXq0T+tz8CIqzwkIIpHw0JJ4DBxO/GtKfkiQG0eWNfPCl/6AihyYqLwYCSF++kuXoMHr93WJIL930sqxKglVD+gDEXfwcufL2WypGu0Jh8D/HLB1kejJweEx7Et7qk3Y3vHPjBnUaZ05GrW6QnuvMAsdfJ01yI5LXkFAlno2syszTl4KRuoUgrcFN2qEmFr94F2zMUUDNA9FxihqQG5MFBJKkY0YSO6XjpktN7opLvwLNIyTHKKbqs4mZNwzePo8N2/fDtvwSm6PnVE1DbOaZBMZWChEgVZvJ4EJ+QOQRv/wMCsK3VTLDgVusXH8EoosSW1UWsQIIilNMZ5tamFxU4Hy2vRJunOAiJdDqHRaFYnID+CCZcdqB263z5+NigIKwerB4vCPn5DZpgJAwZshMBlggHtPdzYZ70Pl8ZYLXBGSGsIdh7f5xYD88Tqh8J/FBfz2L566S5N391e69GlSOOr3+5tFti8zfjp9+MYKzHd8vuFkgwRGrGCxRekY7s/p6xYDH1L6mtrRp//gCTGBvwzxqUOcTdV2fdISAbZ19HD2OP0TshruT6692eBolKw8nMwXzJp2j8YQdQqP9WKCjFyAG8QOnKLgpLLCLNejACOgBo3hAX5mFqf83jDUEIJyy4CJx8V1twLu+OXnQpVyjR6h7GjBswritcWNdg37KxAYcJPNCGcg/klhfP7wn1WHZ9Cuiya/PDCsDvll/emsLNdbCM73Gos3TuTAfsXhA3KAneKD0UBZtQKok9YGOmOg418hqIzVNnc71NQuWIrJ6xD5fcq3qOGjx3Y7gXjMLTmptaM7VOLL3yKQbiIMQKDFmXdhnyX//ParMxnYlsqD6Zyc2ULw5e4/yPj39j+kDOn4sQOjG1C4BNJHWGfbsZ7/APqeSnOJooHqFXnFxucFQ9ln7+B5ufcXUhBmcOTQ7HhppHPzfJ420j2e4WC/S17PmPtjGko2ZK8Ozw/hlFl1PpL9EUq8VgxI+Z8DoNBU6VjJtD4nYEsDBu1yJ4PaVNefHdUbdc2Islu+Dk1tUGiUeVqbQcqjV4n37PNC336YDaze3unp5ATbHBa8iav/AR/MaIijl2wbNyFoThvfrMEjPV9f3rYtZOCZvht4pD5L8aIMu+YLyeOZzDoH/Lw2dh831TUcm+Raj5Ci6etM4ojBVxpBrGkStEvuhAc6IfAJx2YDtI9smy7P0OUWOY2esnfTWZNzX2IpsXOcw0zIoO7cI3THy/Fj59edBMzFHkKuwdLkw02KluqJ7qlCOdfxUVNv7wCOQvEtUW4x4I2rCL6Hc7K1MaePpaiUUfz3TJWWUag1l/g47hdf54CWs6IVAfL4BnetnvgCpWpDXf6Nig2RaGJ3oSwVWIF3/Kqgp6bBaNxt10uLKxP2fpW2/PEG3vGXMNbxAQrcbNNnXIwieO573s/8tn930vYfX5g6yfRBHAru1qBzAROcKSlZnXzliPGnoORLOezFocWA8xdyiARzYyboRYfRccj7AHDbOAhccU26X+HEUeObu0rzuAWUSlHyvIiOlce380P4vytaNxys4ZTcvJ34JSqROE3BX8hgIeSmFFNQYglQCK+F5nYMfVbeNRU4ToZAkmTomdGyGcW77oSK+EC9XGKV//ZLz+M2PjZtwC5tr80sdGhdyqp7L3QolSndUeNamYIDdg1GVrTd4cOM8jLJfG9y6VEKPv4xoe/3KqiLaoQ99y0CTYtWU5c1r4uacTXIGt+vtu9k+62/4VsSLGZ3MXxjaMmQlWy96wm27xuwKslFS4QriQUJ6jC6txlxSHeWgm/W4ECWut7tAnuJjzblhvkeVi2L+dbcD1ghWqZwYOAm48DysaUqYCWZijJbbbQ7wRXuR0A5IvlTHwnBtityIcYy66RPzmMQwSn8WGih46ABgua/xBCM9QHn2PvePZlbGj46PVNpMrNSFTxIhB9Yevt4j/1g/hy8E97JG9qmByR0yCWeUDigMWdJITjrQq+52XL3IytD0cFy7zp1vS9Eb2Gj0BbJMjnuL6akb5UveS1GVLihpza0eQHqpVvUSZ1F5KAw7hkwWSaVlZNlhRFoQ/aUZM3hih34jLfdnsN2ZC43pg8TNYb+AhUkUDKBFzUygRvSMjUKIEo+xaQ9qUyW36dpRsntF8IjcuXm3tJuP+VwMCI+/vuWstHKpRrFTdMbTlbS2MK3xwSGZS/N+2F+by+WUVroGrE2j8UyEs124G+qYpqjs7taycdFrlvjZoZBNRMRnYAprrHklTM7akvaO0rRG+GBM14y+J2coYnTf9/Q5DpmPOZPQbYN01y3pfNz9xYWYD6Y/8yPUGTXekg9BqtQ2hHMuwXn/wtTqulkfQY+YRZXdZDu311KPvnVbCYH3fdxD1IvOrl0RnceQsvBMG9F0l8v7H185fSSitpaMx6ywAPTPCo+00CjEAqRBR3MszNdHpHd67mmmLzDgkq4cYvXqn4n+x2g1gkgDlm09mTXM2HU/xveKBrdgEiK7XqJXIvTAGymgBbhpI+B0fuREuCRHElCZC2RcWJZFPv92B7jKAJe5gB+KyVkELb8bexebV+YUcGAZDoEItzvX/Qz0o02oiZdL8865rkmhUB0pdb3bhimxPPatwhl13D8UScvV0eKF932Tk/94LdxrgVPCTRZjSSc5UGFCWH6mVK7vT9wYKFkgxqTyUciqc/Anuc3ZK0CmMWtLdokpY+bxGfIxlv3Fv2dGZlbdYf1ekrQ7/fKwQqLbRGs1FRYYfXi+EkMMOiBKvyhD0P16tgYd8Gdk+gdkCbdzDrf79Gr0/RjaMHZLg7MPe/QiownuQXdVe/wvu4IJPWeO/XY8deICzTBB9bSJ3aGXIhjk0EXKW/D0dWO0qKCEVie7q/kUwFkAeajz6ex3P1iYVirluaRjJKeZzU24x6gvS7nOmwrU41eaB5tCRGtQwhGeq7wTBw9QIzcly1mkMPHZQgLjRgJTDHQy09U6uTgnBGwzSJM/EcdcyCDIGrmYORqN8pTONIyeqoEGIVAuu4DOreSY7RjEmtDje8Cl+laYhWXbDjj41nOwGTr17h497fpv0zfPr1yh14QuHMDz1NeC3wP59qbUGyde+JPB2zFW2hF0TwDwEYGnKfMY1sWp/JE3r03Nkq97ERXHHhTcl/ED66jY9MSX+e1NALljFoo05bNaKitSBIp8btJduIoyJSUu1uU7fdLhgLD5jQNUcjhdmmciXlxDRpl5B658oIsQRrutPfahs1IUyYDVEdxQGQJhuwhXs4BNTi/2LBo9caNp1+sQB1wWjqAGsJ3Ydrs1iW6rPEylSLP3wVT9bRKyMSY1eEBa2OyCEzweo8eEQKTl7sLX05285PJMS5dVC9tjJiQxwQSR6qYwb/w8a0kvWwQEg0Nh10FCrxnJ36MMAklhDVt5DDfy99UhcaheNPj9sc2P5JTgnAoEpkOUae6GNwbvJugz1COqW/GmsmSyPuEdAGPaEMGhr0MJCPg/m7UR/F47rY2HOupHZESsiukRIRBymvpvvcYycMUD78aLb1dBTTMkYvI4nDhjMV1ExJCpJNNsj7FVxmpy0zB9+Oo56EAv0DsQ1ox+ZwnyeH/8fSRlgwExFGoLNsglOzwDdnbzNpqf90gSisMHx40FJi/3FiV+atsqKmVbaWlu7qWObNgZi661rgxXMjvTNaK5gXM6jSeeEiEboTRmQxqJbLz/rM4BNPC1/DcpiUmGSxXIj74hKi6xdTVZvhJQ2pjggKn1MB+aeBizeBG0s3i61RDvE2kQgTtPMLsTVC4n7QVMiWhoklHTmAI7mufnxlV4m5iUM+mY2oAaAWOzPegBEt6TEwsqAm6bEkFDW4q2dP3wJdfIFIKBcSPe/7oJ43wqZOAWL6bxqEHSGTL/vBMT5YQhrwz+ixCDCF23LQQYFjVJP7+mFbSIP4AQ6ccoU2fAPzgQSl7OTtxvjGh/cdkv6RDzr/Ps1meBUhPiqKbWsy5eqTNzUD9oCB7Mte3YO2kmGGthUR/ok32ZbzLpOnSDCZw+2Fp7TPBdNAbVdstQPEXQ9dDiU2bD2+DnwjFGv6lxtFxzIUtnMrrDjtnDwkDZ2UVV4sj6ZWiPMEWdzOboPnozzMGF0vmTuAwMLqiq3AxS8aR66OBUgPpl92flTZXskZ4ATz1YEXXxjCZE6i0UH/Bu6vMDZeI565IWkuca1zatLm4ChRax9c6gBM0gN40Nc59Ay4XsAw/H3dPMgsHY9l+64Ov52PmZuKxT+9Og8SV9x0RPBlAOxLzSuXlfx5Gv6OMJRbYi+G4NdxJgl0UQAqFJhT+KRY3q+B6BzFvR9E51xN+1NHLhGFQYzTSq3c9ASgn9yl/eyDU1AZRd7LLKZqAcSJg24Y/LMGCmvdoTnG++PlBmkhRdD+cS7m4VwgWCjLCcOxssNq1ybAdpRfBKbR+kdDmoZrlmw4GXReUbjhtk7qmsZBp+Fvo+HlaPdNOBwrBFhUwy0QZWKG6N2ZLzm9fppwOFHQ0ZVDV88w24ElPzsMuK/nI3kgKaqiv9E9BAkeh2JfAYUSdNNcisnq1kvneprh6Y+Vk3KUanMirjxDWCropEBfJ43ekPIhE7DAiQiq5pZtt+oXULisab36kIZvMGUggJvn7K8oMcZ3M1rwMvXFHb/s45LiHJtdx3MY4MtsL4ZU6JdtGsQiEww9z80B68fTuk2wv9scEuISg0uCMQLx6NLjPxXl/yykkYgDK4HGx4CY9YQ86iaV8FCRrUKc6l11unmdeYfcicbhCD2g5s9vX+R5Hd7n33snQqIiRtTByXWBztdxe9i+jKkw5fCDRwI3a0rqCjJIgpMseEa9G1QF8Wc/4oDTmfoqM3bHsXLa9/fnml1Gcr8spd7oUivRkuA5ZCdb6fjLNX1nxabq4iwssdQnSqS0N3WfhWgqXzsfMmjdg2Ico2gVFgcgIn5Skjtr8/gfRBWwV3TbFdb5pD+F0LvoqqjTg/uu8VNFyF706toAJ1QNoM8F0wZg4tQkbXDw9F3V8BX9C2zWhrZf8/iJ/Prtu9VAZ5oRpzvCcucQHvU0XUinuWfcEeRg3rUbIYH4nUPgmEl7UV9Yx6D3wp6LOPcG5auy+MSzS0fipucMYQ6s1Mdq3s0E8/ehwjqDhED+vFk9Ft/Wbl381336zXnlQgB5sWf+/Xs6Z2D2xb5QlZj9YH1p0P2if62wJoDXLzkuej+X5uprMqI9VvxWbQ/8eKaxp7oq/n+V4YoqTZ/q1YZxk810mE9jF9iOF7goVG7qCm/KKkz593h1ED8UhG9unXX7o3PT+sfJJWNzqTpzwTyILg0noatnZUuUECehsJEWbODVEqIyknNJuacOkYkuPE0kOBQAjVcuVbJK8RM+etIVPM5ps2hgKGMZSZ1+orxO4tbCFSZGoaYp3PQ7J7LJ8qoQWk42e3mAEDmLdJGzIrjX/k/MblpMfm+OjFqO3CmEuLfUzuWTCO12CDCqkmASqyM8Sp3rnhhNrhb0SIaxNeX01Awvhhb6TrPzuHQ/z1UCGG+OSM/3eTT2VLQ1W5Uz7kEIEjhPR9pxMYaHKzpcNIHPTe3CPn0hlSHWcqDe6/E8rYBnuyvhUsyGZCwf83Hp+Ty1+n/Ih5j7pY4dxDcgm3RwF/uRoJj5pQpKiMpw6puny33jdjJZlqW5PtXciISDksOPONUFG0BdYMgR8RHzhZAjl7/A/zmJQfB6tvXdrijlmyc2VU5T752jlmffc8MQIl6thm+mvW0QryEYmIqGoRdH64cOQkVLn8tpJWTBKSMC9exqOETP6XMOYrrXj5sZyIjj5EWh12iOvafBrUFTk+sdwavHGutbFEFWRX7JZwfzkQc8el5h8bbrY5MwNSNB1zwF5JRVRSKoManhr2NF2svIJyy8JhWL9jBuZSvbqqT+DG5eM3+QishSndU1cif2+85g8qD/ON9ADd+ab/WQv8q90bIw9SXEsC9nyICbVp5kXo/qPJceSGVekhMopfU9lpx0ZEkVxA3rmvQ3Ifu9+n0zA5YnoWTB6jcRicep2gaF16y2GySoY1mQQDay3Bkt0is4wO1TLyaOyK0xQqJ/93Slk4nwWKZvvwxc6Q0vs1Jb9NL3oT12LsWetLxXJ/iCeBZ97PVfsVYKdnWUxRSKACog94In/nCXrMCCZ8S8Id5BBrpTPX1y4elxAsOt+LnmgUxqMvMWYqQTVWWxnd72BgufkLOyWG+iZn367tWYNRZivaTG40Ux7KQBJEOIAGw59Nt8DJogGjSHoO1BW/hVBg0QQguBw+BFcFuW2m7xECPgGvrKPqQRyrXLGiGUZ/yObPB+/NXpWUsqSPXv3xEtCibIPbiStjcvGTYzoCpcB5WYHVopVw/NhOLPLgZ0QG4cTnVKC+sXNpV9u1peRITsiZto228J9+GPO+pUKnjuMsUh8w5uyMGgJSIYHcS/IZdW7ROc7rW0z7/BYahlZlr5GEXZFvDRQ3olYsbrpWwe1SfB4d+yBskdaSmbx5TtoQoUI+gIkbEd8untWi3rTRgVK0Mympx7fRKL/ZGQP1795aqQaoeFfUpIP+3Vg+QM3haDHXUXGa/QOPih3FtKcRsTeThhtJziGqRsZknjfCzlyWMUPp2DQoXdFOCVfc5BR3wPwprCNro2AUYzlhODCYbp37g0bf4bMsHR+QfjdxFJyg3RAnzJQmcwXch59hRwYx2nUdf0GDew9IEODypUpQ8y+/ztBj0BNsLbr7ssIKrkTkPqx0Zh2x/Ve5WCXmve+7ui69GIzyIAbOX1eY5ccYAt04quwUBXFmaN942YSKUg8WDafeQiQca5rQ2MMjSs72K3L61EC0J/hsJXKyiUykqHigNI+GZWAJJNSIrBjEu9xeuVsx3uQQ2/hdQDdQ4SxjZVfwnelgrqugrCfAMIeL/0rbpiJuYvDJDZ4Bm7/1O7m5BJaAn6Z3r2qjPBj1E+IH1Dknjfie0eZvnEpb6ZebKTOFJ+zU/3xtdEPL9K7ltGvfBk4EunlZjs0T6idaPjfIxvc8WfhO9jWeJJ75xkvHLq68KRVD7XfUIWdNiCtv+lI52h7rcE/qO5wovqeNnf6unIKvPFoOh+X9QdWorm+dKCfxxJa/U7/tk/SpmE/BJ1i4O7YevOzSCXGx+UqQOzBib59Im6uRgO/K/bzQrz5GTpHNCLH/76ZJCJCwETVdamaRrQmQFkLeu0WsJ/c7jJOBd6MhMHGVAp71SXHaQBHixcZg0F2uaiWjYi/lVTjXOaZepGH++/MsZimsFj+UOUVjYNCAJwArEjhqD7Bv4zVq0JwAo+nXHjB4buXm9eoDo1jO36355YmGc7Z8LAnQFdJTJFFX2zi9I8KxYNkcI8aUBQQZWxcgJYx4bECi2Agj1Ns9md3ZLCx519hJJQP7RFX79hGl1h2ao1SWK4E1PIJJ35tcAGE1J3+sKZGmupG82B4YqyawZLDSoSSsXI7yUzmolWYSfU8z4qyelxQUE6RO+3g84KfRGMarRDqtVxnRWCRoUH8wPhCnN/9F8niUQ9azJE1TYNRZ84u1kw0deaJ6l0djmlMUyT9fRZvy1pixv6lBTjICGT9DmtE5v9bgcNRqM4aMdvudCxtSLilKl0jqRCEk0kudWqdqA7ycoHR3FgcWBm49mcrvLFIGYgvTNMCc9CwxxVoQQXVGwGc0+cRKVRqlNpun4b9G5YpitPQcWvInQakoN76fA+FApOCTJaWdr+9jYSyyzx63Z6rcjxPsxrsV23FOGDMKfOb7JvblnnVCFvdhs4SRCYHEs5dQBwJi7+Q28ra3WZGfUDrksleinUJnJkKW6xMkfTeKQ0MpWSwaQpQ+ILSB505qwgKcKRlpVPSQ37hjX9o4eq9qfUrVfhpjHzkHxSK5j4sgDbMF5WGsHT3nvL73848RJCtiDLeuFnA6+gKAIOOZYE3rYctqKp6nqTiuqkx0kKi9OyJ0Uzkiw8JPfijRkd3vhqSBJY4C1XEbwDi3vp5OkI8GrwFT4KWczwVwbY3XkPZHgnhZYka82CAcqZWwon4mXMhUcmEF6fM69LKpVRXRRDDLElUXMZ5mLZufIZyR8goL4NwKBDDgZHcbUa1BRXiG3gm8LsQx4AnZGfCufhXw9zMwySuM5sdb0kMMAueC5gF3f0TR8hRjTeeZzKJ8CQMz5jrY4mJ4+l8TuDrlj86ZnnqgT4ezDEXeIwHAxr8OGp0McKCxXNMA8HDHL9Zf6hLwJj4IrQ28uBdAJZqbj9Ki4Ra33gbsJyYvyiDwZuJuyB5NhxxLjpN1dWmEgOzpNuP+WB4Oy1evw6edxPvD46mCJQMITdiMNpzycHXOPPYNAloaHu4MbhzSKpeZI/IsPCHKsXY1CVbqnoCTOK14kHOBQv+pF3NSFX4ncRnUExrCvv3zPjqI0jF+WJ0UGYuNCVRalkiPyXY5syMT4f44o4ajMjQxcAGVz+WPetKiDqvyEQ1NVqo9HTrMflZlsH+/2bhl2FVkF9b1jqwk/+8YWWgQX56U6+hxfdwpoNICsMCdKNb7xx8RC/BUtetdnpTxU93pNVfwWxCTsqtrVyfXjj/kYE589jhrowCGzpLnBG8k9DLm3AbkSHXpJTQKwm2Gg3gucsfhRtDQ0tf3vQHADYD5qq6PQEIqxDLTOH59+3Vg2u3mGQrLGpZ1gTjEtDW5sB8FhsxfVsb1q0cM+eFxE6goLqHYqPYuuou2r+dKYHO7XuowTy3+I1g+fZlABsqDNkV4LVpijWfeVHzheqHBAXUEBHyP6xyOSmhU2RpmoWI4AmugWi/uLY5qZIlIjVvG9FgZBFjHLFFPngd++M2EvuZvI/ugBaWHN7KXfdasCqB7cfXq05a690EEzivRS0lSqx9pyyIvkZ3ljmETW9LvUXDz9eZT334+FHsXLnrh2omKKF4r4VVCp4uLNwAdluFKR1z2qLz3fsiR+ERmp2pjTxWMfo7omVACwiYJPVw/sPS8x0JSsWG/o2nutaN/33pi8BbrO0gY0n3yH8L/8W23OgJ8Zf7ZVyouhZRjOmkip5bHt42EXB/z2QtxfhpWHtoKgzVHwfJsgZ2aBbhs+pinxodIb+KdwApzKaPYbEUAzcGrGjMjxuxSztkP8iFlSJZfoeqhKAKTeLfOtAywKiaHiowv/dMEUsE39c3W3T+Fyiu7AWHLn+Bm/rwG6BJdYmu3abZ7C8rN1yMJVT4fYBxqmdZDVMVhndLtC6t6LuyE2t6mbvHbnhhLYnPAZyq+abAqLJyjwMxgAyvHGVgl4nq8YekGT9v8BweRX2xLNyZPgqvrJvPpMk0CAYYYuQy5gFzO7OHNoJA5QASTSeCToniRHfySpJMd0lYQ6tloBSdDkQgg9/41EP7UNSl+1ZdkoEiabfz2KnJyyhK3pjp86DveSXc0lb3ZpqYUF5VNjdd7KDYJ10GLwLFeXpDVFneDOxKEyuxYHH6GSmGEyeXbQ4iKj3BYPGl1H73xVmAiOE59t9hKuhIMpsKWg35ZaPWEi6GzDFJf9Qw809+G+iPEvh6VNCDd89DQMv/iwGKvIxQ7LqSGMwjK8e28Co7PcKuSBzXXSokYr/v1a8qajAOIPKzB/yZUusCLFPpXRrsIF1OnccbP8BHHMF2tn6oVKYqRbftg0Z/J4/1Q9epghbBbBoXrmRNjZCVZTvjC85h6WnUXa4a6TwWT3dcOAGhZ5wRoq1fbKm7+T3RF07UeeQ9JcmDaw3ZuBwK5/ZFadUQuxjvnkxkFIQkXii9v/UhKwZF2usSBeOeeI4LAvWTLihr+iecGjweL/bGrex1VWB9GH8P0hW15cvlaYdVrdXdIHX2XL7muR7BLepZexaEY/6tFS+9pPWXWdbzidYRqGUz7efzLhkqaaYVP9qvFiekoC7K9vRVzajvpUMyhd8+BPDFVDpUuVub/TV7AnC1/eThzbL96hdBivylZQU8cMcugmOX/KZp4r95AVDztZYF9J25j1AJJfg/5AOmTK9wnpwi39b9NH9fHvCMy+7zvp+kNOsx6ZqUwFrhNQR58xHBMl9fEcwEFqtOAeT7OAPb1rk0xQ2giopYqzDHEZ+Cz+63tcQ1bfLzfG1zjVy2zvEoxYpdo+WItSRLoxihr/3qTwSxQIB8SyBMJAvvHp2631vfaFu9kDRQ2jCh1b1GYLN7+m9uYICmeE5riLfXDUEaAdm/oNkYo0o8rKW+gY9JQaC7BRnbAriwocbexGz8JV8jcrjCd/7DpFYGAazEjhPz+9x9aseuTLpziNz4EU+Y4gfC1MvzIuZ9pxJZOWc/wTztCaRTFV93UpccdFeG/xa0iwFPMh5MeH4wiJXfGyauvmTx72JBCpnQ/d8MwAMg4V7a+RtawKImgVKQU9UGW5ysCinJTEQVHB8stCk3iAXjeMeAd4Pdfqx2KyVf8kxgR4X8Q1IQB7ZdCV2SexxGDhWq1Su881V2sbDDc5ubA8a96gpxDsggDy/0rf4wpw6I/ROdEpNyvOQEHAK3CkyFVDMvjrhRsU4fIu8EEkESfiPju6neWE7n7SCZZ6tDvBNPqZfToKDIInSvhzU7mTlhHb5iPGwq9TS+3njHZtXwSmOdbGb0AlsvJROnuM5/9D0x6pQ7acg33E1xie7OxcnBlcugnSgybec/fpwh/3l8KFGZuaptneoIbKHQ/a7cZ5Jx71Br3Pw8ZL6SU0rHvHrAcO/fUaGLNo8NMEeSjaUdOB+EYt2ZTQxUBg/5FpDeHq2fqDrcEIfUzaUs+fyMfA6rDs/aEMnEojgInA55qTgsJEbZ7p8Ftvy2a1RI9MoEuROGqcwuYWZY1Gi/YpzCXVF7CC5TQ99I961nB7/NM4B8VpOmiomIJP7a+iMpv5V8ynAUNTNZYuJyNOK/nYwRMooc2iJnrmkM34rrlaxIz8l8C+jsT+nbl+hvvzpHD8t1x7C8f7oTkCI91PeLwf3sLdd8BNwRKlI9R1LKUotRSenoUkzHveoqvD3+hK5AgYUtAPDL8Ow+2wmmPGUZoHZ99lqUWUJa2u6hCkru++y2OF5tL+sBBFOTFVxJ8WZW382MwuOjeGcQUPsJ6KBfh7sxAe211SaGA5/0u6jV7M5ccRjfPVpAWcepkSXjh6+e0/pPULcEzefOrYQJmItQsu4l0DJRx1UFHKxdu0K7fx5g4VTFMCf9iZlzKEfGjYP+OdDjQ7JWa1qwzJ7M+zx1h+qA5gV2NXwtAmY0RNdZfl3CSTpW1ayU0iCivMTwp+CI5aM44qCWO3mlcOi6WzKp/cO6bLX7UGCbx8azZV2Xg2hXUfVVTqiwya3IATaHMXR+p/+eHxs3eP6MO7glBlL8DFl3M7DUYc5nc/W1T8u4gTvgOHkjLfjl+RPsL5HI6y9qYl5JFo2hmBx2y5cNDfD1hsFZi1OA/tgvfbAU/weXgTEKHlrbjjzgSfsqCHgm2wkAGI7xz7Nkb4BYqarP+N6GKQDVIuT44lLyN/Yl1TknauuFg0/lDBeBBlgqRfndViAK8yNjAV6Aa5YPIFBCwsAKz4XEYuLlux5DkZyMMsCahFuIZDDGunyB9muvFPR1kJqWUpsurXWTQKnocwsWQxquZKjuT7nl4zNjqWU5tz+ifuJaGWilefn1L/P+R4rHt8c9P068WrUtwBoKSBabJ6jOvH2fqcGYp8PqnNDYQXOFcUAjH3KYcN1IdgFhwdBj6RdcSaa0EWyNcVX77OiIGv1K6ZvG97On5UdLv+o7eGg1powNDyAyb3RPSCUK5URtMu6Mvs8DtiFxo6MDMXNzfehgemEQzVSK3CDtWxOm1esMkp3aIt9KJ+2WTi4ogbei7m/JIc/JYQJMHrbZaojHYVc7jrCoQU2lLDjGRlHpd3cUftsgj7xVV1PJjJ0ZQ5D9YdeJrbFvkKjOggMtoBcGFqIxXrHXblRVMDr6OovRvbnOP6pu1VfZBoXxCvWHaKxVhd0PmnIKi+d+MYg8Qrie4CcG1Vjelurb8kSI7S1QSv2+DJ96nzlxjM2xI9L6jZu+ugHu7PseMqWakVfAHAb6rJ2qJRF6udZMX/+GHSkk0R4518yO4fgEKvMJ4CDhAAu9svZFHcomsoGHRigzoJ/46sMkRIc5Rn2stGBQ5I/7xb+0bfbO+KXRvagN7YF7SUY9zKWvn6QDhQCF7WanP2YnEhDmP3pHdsebb99XK9CCdXxL4jB43bazymFaaMuw/M4XSaFkxVUPegYQnBgY2zhOyVKmjRAuwxTnWdhmmn6Svd5VMMsge21RcCSKPHTixJPlq6JeD+/WFi8GnQW6hUvx2OqQOUxExVQlPifo3M+LDSbnwSxopnN+Z2JKjb8s5W6b/SSIW7CE5quO8Ug1Dr1JuLkkO9FyGTuZGXvl4ubm7Doat+KpgyHdQQeGYWeWA0sUXDManPMPGanc2x3BzVBtV15WFZNADoNHLOjAOz+hNOIJ4iKRme8OjllWj5YFdCH7yATsm/ZTLYaMr9oVGA6FjWcwJsO0oudi1gI3qhL0VPcjR0UcOFbPtxcnQcjJbYu/VYCA22S2KCBb8s/xEDAykZ9L6MnswL/y8AUvH0ZNozxzgJ1LJNSCu+ZH+S1gUagisIwqLbg+syzHRB+xuMNn2tF6IUF0j+weIb7MxS3z5nCXCiQSJD+Y2gRtazqLp/Kbwj61nnpGOTtwlcijr5ZVphi0MfDXJdcfyOvuwWG2SKxsVWus7+jSVoea6gSkYhamrXjNK7J0mQoaQrgODpNPbLrpMdVVYI2KQ4h1zpYuaflndWj9r/VXFwiNOLiyWcgBRcafjzH9zUhEgkbhqI0U6elFDvKU6Tq83sg8/tRzh5QD8KeRHfnl0vyEK8cCqLM7Icftosac6ZNlXKhFiuvpKPRESBQMJIl+gYMEgfEYroqt/x9dj+FTEkgRdj05oTnEM1y4FCfHi8ksH9x0WZAcwoJwdQdEjN+MBPGcWdcHZYeyhreZAvcjzFsznxUlSrFUcag/V1hXD/hfQcu1xbFrG2EUvF1gHr4agYEkBFxkJwi3qC7b4w4pQAGDZppDvjECy4SaD2ERJGvF9pZwQkd5I5H1kIkWzBgduKnPdZ7XeV5hcG1CeZsI8emhRJJH8PEJrSF7vv/2gQrXicG0GsVMWlzBjqIsJsr3bunCrlWU8G/UYZyIoj2ab2eKcNSodypxHaJqxtvDdFPoUFPi9uhiAOndlwTz/kvb90QQIGjxUYnZkGXd+HWFFnMD+qG+loRqkMC/yyD/o2cCRifFuKQTkKkR2QtPr2JT/k0PsyTJx9jgiFI5MJbvM2suUCfgIQJjPuXSiM8OwEi3ejOi6UfBxKb+Z6jRlZJ8C3s7KVwGZ4oBQXnJRRkHtUbCr36DLE4kNiCrTebV+FSkf2Iip0kn/0dMHNJbc3vujLfSeOfKqNeBBTgV/GEv6vm8e7rhDZD3Mm8smBjiuHxhhu+V2iZcHDEGnOx+l8yxk14AKj0CLBu4ptwqL3ryROCwle4uyeQvJ838hVKh0xnzyqFLDtdSpeHNwR/RP0EUt+twvTiWgOTZfbQjdhHahQd06O6YRIWKwF9XtwaqIFnelSVD2AF4QTqQOtO4QV5vdF8fjC4CjpGh3H6u2EKHz/0410HD9Ttz76paHXdXqwaPoraZKtIfiGI1BPv3iuX3Q3yHbB71d/poFV173yIyFIx3C3H3LxNo3ctRC9TPL61XH7Gr2C+uvkLr6qqQbnD/CcTEEg9KxRRMomtt2lozxxukMk/HFE2epjSXdPVbaFLHeOm7ju2TRf+CUHUMAs5RrPu8HDwQTp8qlZ3M+dqQvUfv0ubCPQ91ytKyuxhvxdlZSnnN9v4Q80H3jjuDvu6M1LHsMEOvfJgUTeURdbSFD5j/RIyoA4nB7zf04rkUtKP6Md2piu1rRB6thAI5/l9rSnSjo3sEBCOHKSU6L5zRhm2270z+tcNhcZEcaG7wqP6ebf3IZ+Pj1VlDA4qRHgBtdFKHsAVkB8uVPzxSeYRUomj5kTYMaK41i+HCXpRIleDImgAOlU42IRVV8zwIpqL8RVEipYxgRBN/98WK8Ndq1Mn4TAFa+jBCeUWV55IkLsTwp3H7kzywrIQnh8sF4tYtqzPKkK+YItlO56SJghuAUSmASREQM+DvZ3EjbKfOajGrqYhyZN3Xsvriemz8WJeAujxBXs8mnTHVdpi62Kaf5eHUSQo5OxVT3sxxXxzn3QfTAlRVD6MIhtPehT3G7ob5xwEDTsjinh8VPvWjoYGQ7H+DCkqtwHtMx50tlo7cMGhQjrg1QqT4EIQ7YkWgbge4SvNPuwNL3jS3ehVDKOLfztWS0mHf+QGTCYGLXnCud2h73fs6Mim1XpgF+wpNd2HtwIfJTHMW79rRs5IYLgc8suSW0oxFcZYFmvyj55zxliIYvLgpU6iLFf6YZUTprwdam9aSuRts9mhSaDMhaS2TrEyzxyVZiP0TffJWoofjtNZQ/LogAT77HmmoX5uVwNwt0ZtPwTbba4NMM0srA0o+2QRn90qxJnthsbzh4yMayENbJJzZJc1i6L674+0BATKet/8XwwAoKtjaS7TC5+hRsA6Db12lB5nGxxkvywaUOwH4a57a8lTScuoDT98DWumM+8YpRGjrfG03E7txVv5ybVneOi2quAxuneE0oTo0ZY4g43wnkvu2znvW1zfehqi+FCRTSvr+PF47AVLCmKqgCaQRif1hKNBeb6cEcbXeT89NYHVXhZtkOVy9NuZgNTfLVJX0sb64iQ9Hxf6giWaaUzXzGQhU0wQ6dqmFsD1ILgzhy2xfJ9GR3aTVjaLzviDyPYFSUNVaMxYSU+D2uhcEl88+JJffPkZdCFWOokCaDTLAZBjcUNnkacNTSFCtavP7QIQs+CYiQFPCoBvin6JjkWBLUXutaKSEpfiOmicux2B9TfACjLA1a53Hx7OgoowWip54g5+NbNl9zB5Vx1VGOXd84JjQaJqm7kojE0YHmKxsF3cYu+/Wx83YUVPxYecUwislbpTLGscIrL5ZAKen0pLbv62RmCV3WXibSLxg0TSs62qXzrIep3+CYDYGyhkuFpJHE5LWy5iS8kHwRSIPQEDx0EmIbmyBDOk8vNJCfbyP1zNkfpFsMJl4eeL53F0y64HyV5yxs0/y8JtSpsI/7VCx23i4wyaqRu1eznQfeQl5l1QQM8Z8EgYatdmJXdfewKP7kUQbXTT7gCqLX73a8Y4ATJ0btchJzBb8KIr5UmMgpkpw+bIEjrIGJ4CPy2TNfXa5DGkXX5wgiA2kO1EuL7YmWH8H9Vdj6AC9a/mQLDciZYcgWS5LCRoE4pQO9E3+Fx8gTC6Y8NKAfClL1JhEmiSW+95ec/Vb2koxP4BCJ2YnY8iW3+6G7wk47oXyXupVvpegTmJe550KIVk7hUFUAca+evu9r5bSEbTb+WTCTgI1vzt0mSYtVYmQ1T0csbdkjUXrhoMia1AuJ6P1aiTNVemxBLWler5oXU72Pw4O6fHlgGXyJZCtlocuIhnnKYLSt1nHtVxNNWhvNwsLB2MGO9UVoJnqf+duJJ0JINH+6i239nbGMqQNS2aUxGQgx20+IeFKc2j7whNWSSJ8wcKKEevsKHCCIi4qP5xUYWIe9e8HaKqSqaoXtLv7n3AmmN4RsLFUlqzwyAkgxgzES0134wqT26MpF6T9/8ZudOZ48vi1Qdl99fLbNXN7Z0ttKLzxisfYR/NfviOyRJ1D2sFqhF8x+j3B1C/yQT3PuMg4LzEAMorZYgScK/Myqcd6lyFXP/CBEE0VV14Ku2nF0DvPQ1LJoBa2dEW4alpneDZRl7wiK+XAov/v8STlGNbW5M2PfoMdEAiPp3FQFCMRDQ0tjEWvLzZEas6fIpWwrD1OUj43f+fMuZecQGMExwMJ/eDm5Shd0YXzgKW/pFD5YNDhpfNV/LNaRO206n+mQvU9OVQ8A5PxwDYeFITVv9MqJYd1T5gTaE46E19QJ8fQgmJNPZqjAIS6XuYAudDXkLuZCk8fvOQx1YImYSdOGQ6pMOeJAK5yV2GbVzqhWuvoCJVW9hxNe8hvyHIGYeuL+2YojGUdk/A8ZOvw0J0sHDlf2Txwc53P8RN2GOvo1BzXJj2jjuDj9GjBiHVdM5E5WyXntDiYYgJW42kxXhmjNvSIp7F3UnXhTw/XRUYqdhsaFj1EQK0ge6Zc4+F2HKUJZOdlSBpzjFeji+L4ObTybQiiFPZgEa1ic4zLsLq3z4HSQOr+sVkiDRVehZJq9X1ll4uuOabDh6oZyYFGWCsGG82EfhYT7I4L/oegYH0Cc0WeG61os6D1/pKMtW53xNMLAGVN9fj0TM3OYMmzL1rDCUQ0nySKACgrYJFKncssXOi6BMnzeJHBqcFuNMFBEkfDUr9jsb/PJHB1vlZs9gJqC3bSgOPhA2riPYRvapheq6HUH/S+QtGMWgz/DzSitG4qycELRU8y/tMiXbZI6iOhvcuy04zPSD5G48QMCBsSCQtKGXhAdw02dCIFt3BWrYMswCtyw9hQpzSWd9lTzV5jL2raoLrcwIQQglRrlTcaZCo2NFn2x/uIQoDwtHJEFHksynkV7qthstTKXsAj7q2JqoSiDuuD+msCuhcosMfuNyU85ZhQC5yCRete+W8mivJXUsniwZO+M7MOks5g0K4W4I7U50Bb9/gEB+B/0hOitQ9UMy2GD/4W3iwSdYqTCxDnkgfzVDJt8kb3plAIXnclsDBxuqe4iSKkC12TjlYI5b0IH+uAFt+kpGb4DF+aoZAwwM3ER9Ep6h5jbhM+wvqkTFJgSey5P9+Rf46cH83qgcpHJovP/sOOCKItZdLAaCW8LRY4I26miw546ZkYtpCGkFnxfDYkd0NPfuGSaGSa9CZR/l/wcovYOK+aVwbKOq6SttIHy0n1uEK5RzttafWX6gwb++83Dj0RdgU3hddLGIzAY4RNnYOCqPhRH5wmQ13wG9yGxWpZevm4rRqyAw+gyJGBXcpemn27AIFIJiq0U13QYBppq58AA9JIw9jymlXNP2U/jpAhFYzlKtMvriNt7kecIVFcVv9HxA12CdljcQgPZ5pN1tIpnbvLWBTnuXb9J8BtOfWdXAUuLlGH0eX7NT4CM2mL92ghofDUMn1AZ0FzJu+gTY+tNEFxF7vehkkVSp+UafMsFLq+qC353W2jE9lKVw6zmNwhl1B6DCcFmNdtPouak0fs7k/VlgZie8amashdJ2jrJPZvcK0DZ9b4EDJWW38+rxAiyDYep9aebjxzQgDec0m0zHskSg5BTc1jZNT6w7D9joPwJ+A4fsMuwU+hNPeZk4cMF5fxdCDFBIbNZDWa/He4fzP39z0lSR+p3o5e8fpLsh7jEdF7wBRdjeab9RkcgLYhSOFjpFmvtJLeVz4in6IpkBI7Plp3LzSBks5qRW5Fjz6sD58oyKdh9AaKiJERok+yuyDIQ7+715hzxgRETtkGfUY1QKl7UL/8e/obb+kWoioO/1Xw62wX0wkaMXUN7as5CyETtpM2w/pb5a55lSMJmyfq1inMZAKIC0y93ZiXZ1iwuSXOQrmnGfLD2259qI8XHSwIIDZCkTOCWOCUDNZtDDrXrZBLZuptR/YdMHRpomAg/PGsVBW8PZJJvJhyATib+hIil2/qsrhnn+wuU26CKsPP5U2vOTWk/F4As5G/u376gBrWU8eTr+q4clD5Bl1Y1NbQsDCcl7xMXf3vVE3RHC+T19sAavHiqveaiS0hnTZlfxwG33VDYK2mq1EiZqcrXlHRD7KA3VmNePaKEjVVcOxK39H6NP0Z52S7wlXgly+aQ3TVooLUz1uJifC6A5vj/1DbVaI2ypQQwY2PortoVGRX8XrbIyx+NchZ02ZdSjxGcC3HiZlAt5cRPAZdfMLlnjrJJlvbi0H4mEP2n3VNrnQioA1Lte7xwg9h6Bxa30aoEhtA+NGnrs4ie9ay12octlSm/mlj/9NKnvrXNax6zGW36bWOLT5qrDNqSvbgSu0nwcwllePsOT0mSIbvoAQPgOB4Op9vigqhnNFoxc2tgraGnY/5DAnMiy9f0QRWIk+KfFQ/i9MMebDhs5TtscFjab81sRCdiUEjhuPoQedzFfq3u7PKAT6b/v+7riAhzd5QK7JN0e/TmhNwgIMAVo97TQCT307nG1XUTC78DfMA69OoelsfLsIlGYECy/UrwibolimO4ClTmXdkCAq4MzTAcSgmQN0PkcfcKQXt91f9T6LOrtMpdOjUn8j3K356OIDz9vRrVWvkGWvRr5rvX+7kEGhJ/umli8MvpBYt2PW2mJoIB04cB5aeQjMVN7haRjkkTUbVz4EoArAtG4o8AIiVUEiQI6owuOijtb/TJ1n5BSDWnrDP1oIXPbp28jkYKp92K/jT2b/ZTCXLxbl+c4RSabbImB545ilUNcpMmWG4mNnuXL5dzftlzS853+jO1gakyeJBoVzn9DHMT/d4DtZ1UeKPH0k2ZteCto6gzPCkJk7lem+XjiCrtvWFMKy6sqQ64KrrzirE7uO6CWzjmZ2fxbfs9mUDlJ1W6SOQYp2A15Sfk9P/o966WwmmNtCdVl9aAtj1dtf9X8NXpBSYRTVs2wOeCAimpsNnpy47AHYEolH+Z1zN80uHPIzEq9SBgoScn543+g2PHA6hSuaey6uPerQEYuqDKrIL4EpzsF2JdpMvQRtg1dF5IY3hemEemGBaXd3MJBQ751JSBnVwf7iX7UnwnsD2fQc37caC0v/LjxC3xeiVXOnsNqYSnndujv9F/DtcOrQV7R1qWLrOQ1lot7GlcAsP++gi63CDtlW13hRO3Xa8swa3P+gC0SVL2pFWfV80g6dBXYgWoaA5l6XQPahdOmyAvF3C3g66omGkWl7lBIW6RFN7yadvc+CpQc/cLY3srVzayPfKd76ERi31JREjtuWvrEYZy8Ex2goxoZ86UYJSWNaao6qzmIkho3+eyXgkm4NwobFPFX57X93rbcZk49MaOMXhHYwCWHGjSG6CXEWJ3fojVoUEXOhFqoMJfgeLXmxPST7ZjL3gLmo6Wk5GW5f+y4GXijfkjkMMEG7e7Q2VpxgiXmI9DmSvyA6xaLnX03wW4MTQzM3fGwUrM+vUkdOeZClWlh8K85YnmY8ZU9yHLnYWfkFEkxSI9KxTO/qts0neIJMsmyLXr3CGvP6xBuWz+21S0kHHdBXsboFqBtaQat7WNsgMO4hUQZKYOOvwBsxRsvhbhwxw+MnfwLYtDd2pSsnNpZ0qoqB5bdcRW4wIwJtgSc8ktqMzN7hK05Yc+S5zDZ1VUrSicsfd3KyR6hbfHttTazYmHsjCdfLe2KtAq05rokKr7D0yf3p7Jra9uE6sWow3KVKeen+zdAPHfLzFi6qh+20WjNlhKKVy8rzu9s+9rrwzSOjv1pIU+nt/oeu78LzeNLnVIWX1IRPif9rpQYVthyWCbXY/6PWyVSXp6mbQc4Xyv/GlEFp6uBVeHsCkeqWZS82cdRb5R9AKO/vERmC2qPItT+V/gz2hM1MvlDRHi8YfV1NT1foIQFaq90OjpfAvdtY9K/NSbqlRv2se69vb6DdcXUgUXuHVusQufUBDcHxlndP3TCX3YcvqZGODHT6JjYKgfmxZUmFSKSKRsuBBikM7poNHS1eWcFKGw79LNLUFhD4R1faiQP5p7kVPP61a5Fp/49KFAUDeim384f9NbrcnwVleQTWA2Ly7WFi4CHsuUzX5MsS6o/fCl0BxE9KwF21lS9pDvF4+6tT8qDCXhSfJN/ze5Cz0djvs9gsbjKhVMk3tfral2PG7mHYkvxEYh9JKDQApSRg+jsUm3DS/RezYleg5hvSqs624B3BXHsr8OiM+V3r/pbTEtBydm/hr+pGN2tykeD+4NLrquTmMHvKYuwUgmuz/IMQjyasuJA9YZFyUuFR7WtFVmsS3vIfG/gaDg+WGM7yp5mBUDYbShfkc7kvamADczgmwA9e79rUKaNbpiDJB0DTj2Q1DxVMmQxAFY+g2e0/jQ+i3DV+vuXhpPcbKVl5YebtYKtx4mmtxObfeaibw5UD30LSV0CkGVAaSf5XchT79Zg0BI4VfboPlosyQFzZGHIkX5IakN29srAlf6a+Bc/rSfqR3vFhpHdK6KG6ToZnx6n9iZwuVulSsqKsPqJ55EEVQX8zxXfTXbZLIaOuAS2ZJNbJDBguoG2DGsonN6Vgk4Vfo0icbsuUGCaN1Zd2CYViggmy88nYlt2lqNjXoq+yxzC4fqn+LY1DLlopNxXF9czjJ4UMAEhyMzf8IwDOpRp0tOLAAtcPNIfQyksYzow0GccImwYVDAgjMr0shWtvqyfLbmZLzBv7aVDZkZe8cQGRwMfo5tIK+3sGumuYJ9MFsOcx2jo6/Q8Nt4IaJpEozwAGRquGfn6oIpOdkYq7NXtkSVgmlEa/LidTtGaC8A+s0hve3k+MH62gSCdtSY1++cfH47t4o9m6oiH86yqZD9+BE1H+zQS4QRV1ztlkVuzQJrQPi6bV8pdG8fwzvfnzzk6o1NMoTvaP7PSTYn7WiwMEqQdj+Y2DLkY9u5Xx1kCXX6a50fGx/AkbhqklySTiWoxB7caqr1cQB+3BcNstup5hFldkU/4rkNYUDAImuaIsiHMReaR0dabaFbx0PHtQM8xrwTVkQQKENGmOCPHfqUi+CdJ5cXnPzjhWjPxbaGm1f2eRikVyPwmEhCdfAyuYfLpEkyrWb3ziWlRgEv78guG3G7+b9Pe5q4tjcoWs34UZs2Sg5zn79iQrCIt5XyW0as1kQ7r3r/MQzmfqxwRRY+0RKuRROEtehFxscYAH9CNW34qd+unro7awSzflQw38o+jyZLd1ZCKgrqsLSmgM6CNXGEEwenK87LXA577e5lgvHv+8NgwplcGgGSi18V2GsWtvY7qhzGrRqtEU1mHTC5Zb651RecXOZUWMmHs4suIh0sjNac5BwDIoe8vcllCe4pXT+O/Z6rkbcfWLx5d9WHh2MfH0H9sFmwihDyn57zJPCe3v8wZf3/028vwNUQMsVoiFU683APhRP1k0NaT/z8Upzl7JHnJzWA/PeukoiUy+5S7J13pJI1g9XtBfX0oo/ND81INHpFFBA5Af63MoP3x6c0iWrS/cta5VnFeqm4DXWnKNaowCzhL+xSYJ7n5yAfRoC6HRXjFQAUHrpzOFXolR+MiNY/L8wXRUYPMGvbJOzdlHVacvGGVIcPfbde+KsyDWXText7UKTZbO1+TM8yjbkwDjarHpmQW0Wpw2NG2aDmIf2clB0Iq3jcELHZZ+Z2Ryp66xXmRswTI8Bd9V4vK7toBU1AD7xtQIwXoE58WkI451+OYM0jCn4ckzn+wgu+34JFrjx+1ApQbmel3ANk9YwnqXIx2Fsv188YmYP364rD661sR5ZlIgBBKQxq1YMyFAeXWFtMBUNzEOOLgdUiKerNaYolcei0MrgoY/M6K31+e7gT8Fd76NC5X7R/THIhg4NZvwKJc3SRRpfgjblm5FpD54WBrfHZdelA+b/SGUJa2kAVxGM3+YN9FKkFtDN0FVWVhGVRFYKsBtw7IEuMxqEqrTL8i1hEY9IPbMATnPJMzsHs312E5rUyLTeism9QoFjKtOxL9QUDtHWR9A7QL9pqH8u1YInOUdr2zazg5f8WjYCiVWP0wIm6wqm2tXCq2te9h8uu4Vh6rKzpNpRla/y5m+rrFUxNQIbbl/Agxs0CpGkstdYqqpo0Tz499VbE56Pj937tk9hg7Sq5owv/BlMt+i68vi67zAaI4lNF6qGGFwxWm3Yz+Uiin+b89DTGiYt/wnPpM944/szxiI1O4uKSuYT5YGp9Ses/v5uJB/2LN4ktDZS2x/GsKDcXTTUZUindqNQFfXCch8pAMzAgHP3HXQzOlsfEoTxJxHXMq1IHwSf1Z0kkN91FunJxtUtuFtWwiBibvXxtn3yqpimjOM+Z8TaAwcNP8/qGTSbMSdGp3yhRNylNcRBdIkw41EavJDDImQYN8F1Z0bHCfXubo088YNyrVYO/nT7RkfuLEOstRRUvvz70snLhUdofgwNq+k7SFOVA4nAr4un0RNUU4Dzak/iXJ8aNIh2NITs6kbIQ7VDtvqObsGmgfVkecTDaCN+T0TaijFoAseUFcOH948CoX1la/ao6u5zYqfoeY06cQqZPEihtMTTuOTa1DujFx1XY0rSMYDlhHq1EROm69zn8dVQYBTD4WgTSvsZlLI4L8b7xljLbYygdqdnBCdpdlYzxVqwNjHDdQhlYVv0RhWvxN2CguUDUbYnOt5cH+JbHm0G9FSNlIY7u0JgHZuLjISUXzFHKBcTSHEGu9V26shz0sqpDjoMiZvPv6mKTJ5CyJGahz5NVZD1XZlzYA24SXMT/pgkklt7AklvP03eF1qHjSZWKR6phhXpv0EXsiEkpiZjzBr/OmPszGgwGfRcJgfF4rUCZ2ay4DGiUyKk1aTjM2sSkEQEJd91CcPhE59n9i3FEih42l0puf78BDJvu+SnpDoc8XhKDbuZKAEnZfI0pMFRs1hirRqh3XfotT19aTaGJCDJiFceNTZIgdM5YHweFUNA9gNpgB9fN8inbTJrMUYftZOuFpD3umY6/3kY4c5Mx/ShSIj88aIrc6VVjlRkqDdXE/4YyUM+clz5wrPMq6Hf4Gv5ueROsNTnLg5e5MlwtV7yQNcWS2Prbqo5llLtr8HiIWCKX6KDrCtfp5elNBXDmUzpqT58lZLizk3T22ejVSngHfNzIEvV25ZsvLwDBE5Pe1i3MRm9Q5HRRV4M4ydMuJrVUGdDGWlATG7TkBACqOAM/2fL4oD5i4Os0SiNQeEKzp8CMtsqgMCL1EOHOockxRGce4EAvPZwhvGyNB7n0z8HNKc3eGH326/4+ESLxOUjN/Y/sO1t4vzwc4RW/jcwnt4PUV3rsfowgho3NE1v69woZzYNqBLBwf8ntVH5XfzpCZjX9L3P5TKHJoErR+lpCkkxzuryIayY9h8ZBOT919ELNw6sOEoX77CClfoE5pM0wFr9DEw4m0HY2HMoM1R0UiEr5fxt8c/59Z3BZl6wTrsgzhdOv2pRkDan7P87blSUXRLO3dxDnu6WRNHlJ8z57yIBJYvOx2H6scnyuCe0DiDE+gzYNrZ3eHq3vEQrfwAeMuCTKZmWofkFfn3MSH690nAiHt6iS9YijGLHDy66YWFRTMaGL++Zlv2wiyzdRypHd/X7mP06vsF+064aE0SIakzAFLA0fCV4KPLPoqxYGuOY65pEVi463IX90rJ7Mqj9R+HZzzJnWASxLR3epqywEZ15ERTZqybjxf5Pa77xvKG6oSW+XDzo2RNsCrnNuQ/PUoMGHSAvDaK3VWL7UQfdKacfgPIWlA0C0iQkVUnSs76udlP6AGJDKj4azeTyESGG+BXHHI3u0YpaTdb8QSELf8VCxfULeY/HQc4JJscaIxodCADwDAV3oyWKVZ12Fx5n4/TzZBkXaDJ4rNGrhy7FJi3wr+02vDUJKmYziIHKhG98kqvmJuGOieER4ViQCLdmQx2Foh6u3njopPUC2qjUHqG7TOfhiL2BKDzMLgGfwZ+JmfQFVpeo+kKIl9hjczIKokvYkZT507Je/4CtLaiRQ/j28kYMcn4B/xSlE3caxxM1aQEqU21YImXGm52c0lc8weCr87I6QtJpfvMcn5DSELlWlJ1R4U70tZc0Y7izUT9WFxQqgMuzaD+df4N5PmA9E3PsQnUOUz8MmZSGPMP3+qgI0o9uxS3aATOR4Dg3f10XcJm3W4N+gTXlHabBomyGIZ4Rzm62zGV18MXOHA/8QxHe6D0Vc0KaMxtmnW9ymhEs7jt3k2GS075L
`pragma protect end_data_block
`pragma protect digest_block
98660535d95068c5daedb28c4660ed3d7599b4070e205ab32e51ee1acdd8023d
`pragma protect end_digest_block
`pragma protect end_protected
