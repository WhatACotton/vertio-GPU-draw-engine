`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
IQbX72FWdqG+wKy+ScnQjA6W2I0zqGWCRkUk29Bpk2Zj3VvZSGgsPnZnxFK9tCIijghkYsNTFO+njnhNaL+vxjprrZ8s7i5J/guLMD728o/HgH4x9vdE4pAEeTPiRyAY860YkEvSOLUDoW4VRfmwod86gwDIAj1372k6unf6gIPTWyQtz2xoY5wQhRLeSRogIkGjSlVcV1AciXfw2F/474RNDJf3cM2MRM0qGy4DujwzOWHs4LDW9RTx1QFjLKLKknq4gmQ4roz+AChqXsJQIRjJ5Odsu7ESTe4w4+1LeS4Bu8733M20zDEnLIb9hFAiU46NwBkMRQBv5nBvAviLp7Fqv64JMz03kQbthUhk8kqMWQx0EFCKC6WzbZyOkPPT9yT6+OE7G7tTzN82yn4AR/gDwoew+AaIAvXOwS7j1sgIYzhxjREhf3Q6APy0MSs9QlJdNvpCZVz6piT4DpQNQvIB8xJOB7KLhPRijza6sdkhgLfd+qzSuGNAdiA1BbQLot+X3R9glpLEjTxXEIM7/9XIY46MxKUFWlwsdESGZJKHVxUXHa2b74VTqklYwaRIbTdtQndDkrHpMoCN/uV9mUVuMcHq+TieKQ8xsIWxRBJA9iLNSVGTcBd27dSK3VIrhfGM1GHji/h1UkJhgXIE6AHGpoCjL3a4kaGgdsqM0gpx6ZmRgG/LelqXP979TcqYS/m/XIal/1zxsc+y6PAw/idbMkO+I42IxteysKd/aMzOT27BBeTLuTkYQQO7jS4zYOlGUnxNrefd7pmXaVuz0VEZmrIM+qwnFdf8Mg4qnOR3K2JhMp428aKqN86jh9+AC62R0aRa485cnCNDwmhIiTWG878WOgaEihBeTZfwuSsEq4UJZFGZS7SpK18IP10rR8Ws1hKqQ38L7WXmnjVyFvDEziUKkv4we4T7kMlRAAIQyCTMmQTnwe3GT/HSare496WQSNgA+vIv6x/irYPjPDwGYV8sEh/nCxcxap4H4sBiXVv8cK7LfezxVa3ZYEVuqEwm2S93RmNO25i89vhczovmbD2KCQiZCYjp/JV3K6TqYKST8SKXknHyQ3Day1Ay/WW2O2kLl2+MNlqWc90JUN19FzsSsi+jIMjsoQpprWZyNjpCBe/n3ieQ44v/Z6qY6RsvBdvnF3hCd/54GassO7k4mKIF7pJMad/Sm1UB3RJI8NWzxmHLiWzb7M68jaeA53+QImuRbAbXzG1esKCYSp9A98BYtuik+A6hox3+vDL6/q+XonyQs7YS0eEv7PQI6CyQ7WwrJEAf+BbaqqrJgOdLtyU+kW2UEKARwfVyW0BGes1mBlmolhTyEHH4WoSOdrOh9aQoqq+bR1a/5JxOOznHn9VWd56+AEmtexIhpVH8NwQv/zIHX7l5YIcvqvIpwrnnMf0fvSfywgLcwyu5SAZySjAW2DgKlUMLwv9+3CDqZJmkky3ds0BfJowXfRgAwswJV49nDqjmdAYZcfaKuyZCF8gdSW14QMlLY8+lm1I1qteegpq9g7L45qOmczf2WN2467TghCEP7XnIU4bcyHKpteu+4VtlfdkxC/CDwqiBeTAvZFly9pEK50VScmowhKoJM1LnjL6iL2RXd1RMBVpXntUtVRFADM8NQI9KSIO7WXMImfDfJcUWi38xTDEtB6BoYvbOHM7eZCTSNP4IWkO9Tyf5sOxdQmTd++fR1UVzqhOtB7IxIl8WDuwM9nzMBBd05MV3fZxndIEzb7M+Y5Qu5/SbhJCTAja10kr11v9navDK2LQ1kn/4F2VoBdhWT7emQjcPLPufGoLjSoQtS4HoRAC7HT3YicZh6a3xFnZCJIGUkX1CKP3jJAa3M3s/0fXr4+jgVrUGlTQKyb+39Vz3SoYlhL0K2CD5Pb4l8/iiEbswqmrypZaBoweEKxH43T5B5FU+Tj6DNm5MOe7Wg4yuLC2Z1rf4WtH3YFNNtUQKFP2wqavKEbyKsiGxziOp1688Sm+JesqV+DcJ/jMUV8aE37bS/DhURpktpNOR1kOFOERkUvjTNP2suCGB9ThnsUJniGvu4kRVjz6OfYj8IghueDOwvPCIHFJC0ZatFdhoz8KZ12u9/7H7hyzJewcbw/kiqJSTIecdZY6YQIIKpCMNyQtX8eUmJTdsfpch2CGUyNYiwgZeG6MNoPFj51JBZzzL1MPCcPS6DWQGu6kg9LyK2ogFP+CxP+WlnBwolRTQtavyK5ivr01LCy7wth+6krHRnBHe4Bs7hUMyPK2HAaC8/5xDlRm5DNG/WCVnX64c+0BeTj/XeUJoXK2e99M23aSvpBMuQs9O1SBR5iO18m0QbraVmjRlusnFP6jQ/DBQvhpRoIeHP4oZLV5sFZqi1MTfgJd4QLov8lpkl4wETwEPb3lhxJ1n0Q3iCfzMGFnf36ZVi1tO9MgRpX9d+Jx7/jqwAO4YsEoi6tv8X1PN/zwoLsRKtd1LAvB6tkeRqf0H+VgPYM2UIgnH9btFjbrfyOpJ1inzUIz3dS1U+kv8+9SDoLNEaqLG+AH4HI6mqx0EcK92cMOralV5aXTZf0xQdYzKykE/jdTatAQ1M1Sjby5+4of2rlIPAEiOt7vveaHaRskSDHYBKovECgGK7wJ82Ery4tGTGNSQdd7HGvx0EuasCOiD3o0De2PmoakjMJuyju1hbYyN6EmHVDJLyURJ/kkt7mdYHWosQtUr2nzIU9JXy18goLUh0KVtOjyihe1Vqm1o2zGO5exVIvxb44BLHGlOMYG+8hiLIMchnBvlh/l0ZdH1PCljG5hfSH12+D1lKAC1sCwTd8R0D5QJpDmzmqIcJTiFCBpAPZveGvwhpi1sQvqlp3EwniYTblR2elBOABvaaHgjlK5dR1gIHB81cj5F30Zf4PY4OINAu+h8cg3EyRv7P/7N+GkFocq8UBgP1BdhqcTLmktRJI22/n9JoAcFvvVh3WkpOTn8LNknp9P2S0XTsyl5kzZCDorT66lnpqW6qsOFsh/rV8zFbau6opIie7eO/uL7Z0lu/zFE0ERSFAkjcvU45o4AFCFuecUF9T+ZKS9cUNeIY1pwsbacRIF9T2ZEWySuJMhgOP+ROc75T+64RHBAKVpmgiK5W5lrhDihr9vmEIs+0i/lLFam9uMCPE4ubm0y3mLjhDW2EOR5sfkMXdGHmPx00XGjjuZRG/KOMoipN1nlVPs5O+CKKoZKf80SEhdA+i4Z4RwUyrCxxjoCwABsuJwYJgbADISEBqjKvMiW5UYItQQ3MTm+LKJ1TqQ3Gtl7jnRBhLw+Cfg0aajk7ZHwKhzxOjtbQ7nGdpRTHEfGrKyCXKIFFtyZYRwHWcONyiRXHTlWy6+KmLp2S8Jb3XYi58Vf7jQgywwYxwg8UNjw5WS8Of9Mj2AIj0Al957RHiauwhAl5Hq/meu4wKFiVJkYSN6raBRNeYu3VL/I/9EOMlmZitG/9aW/qQ69C5qhAIEvYnUYnbtIGrU63P4f+l7MiHiK/itLGlim0OZTbI/59fT/zhHccGwb08/dUvoRAk/cWhqHV2ygKMxTBUyDBR5Ftk9uCo/7nmFnBRt+W4xPwPzxjMaG/gxHxzAZw6+wELZQ6i1IxSyl0J9OEbusK0WPCwWlT3gCqSdq3erwMSrtniyiekJl5U4qlvZbiM4PEQTYs/S59IKowHIDlWXmRYyBGabTTdI2A/z8Ro3ntabXpdyCb3EqefYYbNpFCOYO2x2yeVFZ+eCNBgo0kIvmowqlvMBlntPr0nSLXki1szi5FxbLaJvy+GwVHRf9507pSje0FAhsmGOR7jEVUGPlmGTbTwZ/g9dRnYdtUowiZook208AWMsguoir/qo35VW2jYn3HhmJi/etIgwqv5Knqrtqc/oj8je41I0NBjuWCj6qjZ0l8ePdxIUayD6OAMU3oUl9nlLJfWX7Lg8S77nambrmAAaUriwvpujNdq5MZ9ADZyi5QqjSl+GijToitHRnlnkLA8F+2SH6bSGBBNhhCpiT50rZN0ZEteHgksyzr8lbKxAresyRTCsGbzd2ptADT7ZpvTDgQST59bl5EKQ35rqozBPO8WMjoUaN5u5+C8trq6En8PZE+2WgMmEGNnuUHwtGfUnqN71jYOd6ZvC+0vsu73ZxB59jwupBwbKK3o31Y1hO49h0eDJjpUV81DH/QBXhPilm/DQW4GbOWnaEW9zd863NTeOWYrLxt4Jl24NWt/qZsI43aYIaG1H0Y/j94RrGiIxEXM/YcRDT9Qu4KdV82Hd0GUBCMHON8flsBs9SRtJqsYZzKMZlr5rlTEEWDcxDbt8rhjgiPYk2jbBCQLgPLuN265JPVIVJ9ZV1ZLtpuUywJwytt/cpGREBrH1HkoP+mFfe/2EX41Ouzi+86q7oTGscZbXE+HE7hi3rPWBfbheoZNo+NZpuxmcvT/m2b2cPjzMWhSzhSuECeRmXgm2JqJntvuuJAPuphtfvai4ZnxNSe3DHyKjMuKOmLjp1GfzfosYUWhN7USG/hDxJDM7iiG//eH/mzdsUcZ2GpkCN0Qjmu4LXiokiTWVDqOmLyGNnENF/V0AEtZX4eXu30poZFbQ42lib6LMWN0hDhnM/UU7yXh5YI4RNOddXluLKeh4///SU2YDfjdXpt/NE+tw2UIRCWriyxLs48N78snMR6Xw1sEdYE6e5D1d3VWDWlJUUK3/+BIb0qYbCAnaygXZsSEHrgIZYri9msAqlCLMUztHEviOorBJDDa6Q3FFl9HnAyZTLrCZmWCZ/171eHRBA7HZ0iYYdZFfK05hSgTyTRoa4T5oDEAcWlEfmM7o51hTCLrOzBmGi/qeUJY9sB/mM2azKRAqexLqD32i5PreHj01KSfAXj8yIkWoLENJEcXLwvCOFjDftVfyQnws1kJ/pdXX49hE6EHKyIe10z/CKOCvqnHForGNO/PEX3l7jjFr99obTcGIFdaKQpzgirtD+mJuvXZxJkzwDFhsuIskeihSkbHFlXBlpdYgNUEuCWeeOw6YC4yuDgfdjzMCJJCC+I7y+WdGzSL1wxhWO6LcEOT32ucv4LuCRXbT5SpPXI5o8Ihqx9pOtxnkbJFBPied0lT5WWwHPtDcXf93qJ00McF7e/YShz9yiAsNxrmgSkpzZ6lNd7gbihZ9JWNoxg7h6/WFQZUJSLpVAXUytEPlGG820JSUG5l2Wpz6lDrKAgKrLnueQWnxSDwyKjzd2LqhjUqh4xDxs3y6a80cmu/tKaqxDDfE4dA1Q0ffdyo42z3lWcoel+YTH3dJmd5cmTWx6OKCZ1PyNdqv6huOTDQ26Vb2NXLlodtCqvVDM39zCtmCAxIsAC1no4vDR0ooETFAXx/I2I9RE0wpC9mGT4YN/vQUZoQj/8zAbeffFRqDVIpdplxKxE1vhn8ZT1m/F8fpGmG+POXthJ0XU+qFSciR9bK8YAOdxo406XnnL+sc7ZnUdoNfUHfTZhNjBbij+N/8KtOAFsSh9lNgVxPqhzjIDzUj3mp4x4w1LvGgXc9cdEwgmJbIshHw10yec4DX1Jl870bhFBQ+jP/cKoagHJpyE2oJejLd/0wwicnG0nIMKx6tDGYlU9wiOey9USDs+M7xsZg1M5eU7gGfyVNN3Mxu3S1ZjtG/NHTfhM3/elAOiEbx4QiBHFE0IdB9XHvRWzTSvGt84pih4hydR0pDBu+CjAQxv8o6A43VQV6Ifp/glUQtfk2iXqOo0kgwdPGlVHmLPRQ7quzVw+N6U/oHEqc5o3Fo1ZlbSKDda61vkmcjBa0eJIYsBHsyoMuC0FQ91PSSxSS5tAciH4+QTlxXNr4zDw3nTCfZyw5LM2/2JaKBm8jsjRaIf8e0igMQzT9aeO6VPT64Uyjv8pSHRJwQXmspdcljn2qeWgi5oHL69GMkNpTbFKqpda/oSWVb6gOnFGPGX3XRm3pu4VcmHJoCCyPHzkAfAI3YQ5hU8xLlB4x/qeMZo5BKxjiBet4z5FDAz8LAre1xdyBDafYbNOAeD8oVMTbMqaWNhl+4YSq3zni+iKF0bryKwOPIy3gK3eu4i2akNQPrAgdm9FAALFqy7C8s3msQuoXz/ivrowialnyKoBLCb659X673Zu4tfCHbKj7qXNPYEAnoh1XMA9Z/xb3EVhxMEPASg6/zJ7Vw/awoFBIIIDhxoQ14ksR62MeqA5nnvl3YkmfvDxrtNJyZtcWsKMpTLH6z0KyNZcPtcE88+NEEMwVHjLur/uTLUer8JQD5mj2Jgik5UPpCEm5mFIlPfcMnFg2P7wjjPtsjMbHkER25BhyYdDGXvaQxnAd56yx8wP7VomgUDd5H1fmwEwvE5xyc0KS0P+qptyUWe0uufk25wJMkM01HVYF0SYTmEFX1WVodNYLEtO7HMEj+Bp8REhGudfSJDvknQr99lYPS9oKMZrh7EpX+ER4SGNnZixUdsSUuWG3pCuLMDksS2kggQBYECfVziaIVDNnB4L67wVMWftt6QgdjAdS3LHzIp6rcSk/7yAQ6PY5UcqvP9aYCqo60pKu7F6suzIl1vN8fQlChI0uU+XkGBbcVSAWRCPsQLdWwMJcOZBsVcTPrFK+2MDZKUimupokyJMiTnxXK/Cj9sgpSPw6rAKqg2zlHnlf56OcUPZt3Lr1s1L5oKWJ6kz7pYe+pF5LUip9oInUCL3owwywjSb7K4NPQYkPGDwTAlLVUQiHrinnrY/kKwj4V/HswkIafte879gquKHzd0cgfIw6GlL+5y8AEYUpSDjjg+XgRq2K9n34QM911PAf3N9zmLTojTcwitnIZmDA///F38/24zo9QjIZliWDClGQ1OEQgtr5PIpPwgxYXxmyD4QiGfvkHRgiAznggraPCkFMofUfi6E8M641rk6KjbH+nXyAVuEeudiPoBdq2l0jzEXY8yA5oer8OkhLkhXgynlxlxOB/mrCZlWKJ4q0mA6awKbQo8r60ri2Xzwkf7Sg4fQ9nrUfrCxtaGz6YpluhoFqRMKcfQ7eE4/NgUPqBs/8LG/oXHN0iR+Vqca8z6WZQ7UCsj/3Id+MojMrdnU1FEAw96rEYuaDTBTAIRDtt+KsKib7cxonUPnFefyyAm22rehPLeCdxVjz1v4Yotp6LAsWb+eY8zCWQNR6ThzFasK9CRBz1gYSq95YJJ+RhXvRFybKck1pCVSjLf7AgjD5vV06T2y2y9WlnAhvBNHDdfx2BE1qMB0Ilz3//XyMUpeZvDD907e5RB2tWGwY8h9VTr8Rdq/8GD00l2rYhcmrmOspocMu2pvlcPuGWNUmDZJQRgbb6g8VfLOCl4okyZfJOeO1+9B2YRtPHt2S37DQ7Li741R0aR113sm9/fUBNXBfLWhNVU7RokxTfcwzklTAGXPfqr51eiukoXbkRkDirlY2nqPLQSYhX8VlRF0bGcX4o3EqLFUeECp/Z26+L1za7Y9pR9iOFWHNA5KL3gylIRLjqFlM76PvnIjkvCFkORMAO9PAqqP6fotI228piLC8p/3m1cxtvayDJazpMoMLb9p5/lyDIjCUF6wft+9zvsVypUDKvTJIr3iwxiXfxczlQuRgIAZJ0ikG7Pjs/YugZKsod8HLskznjVvd52neGfedssNk8a7xwt7FKHV9Z5ErsQNIlu8leoh632YHq7ERtafWDGiPTZbF7W4q8NIt+WZl7hMgqtvDbSKo4e/k9eky8iJEfO8GjzdcRXX7+zAfDS/EUOWfvi8DVxscr9GNGHofRFqv/xgf3tugfPKbp2pjw8K0VnbSRgWKz/eJDVgMQrxgax5qwJqoWhrLxg8szNCUvLQ5LmuD0DN2I26cOTMibGEiKobHBXOW1wZcpEDY1oFeqV6WRfl/WYDVP1iZOSAjYv+RxLibmTiLyEaotrlwRE0aCRb6CjyOdkndFzAgCsj5Sk+lnLYxry1RT+IrFQr8nbqBlMkN2obeg7nMI5wZr6yOU5FG6E2doAwWbqINJeRa/HKw6SseyujqNRqlSQWxpgUdv6Kp8xluthVJe37/ifFY/VkF5ef4h8gH6EnKpwURgctabGsY5d28vCG2MU+9Yz3jdT7p/z6XyHAX03Y4ITw2aO12685eD8P7sxpe+5HNlo/OgataiOHcnPzpzyO37lQWhYgFubpWGA5HbAWFOHx//0VBoIXE2d8pLxky26fgW345Wr3KiTuZ1EKSAyFWaqrOhckAgH7UiJD1H5zEw4b2e9Dw7rFr9zv1rGuHUKtkZH1A4uohUr5IyGKhe6P9/sRXnYzr9GbqooM5nNGDXEGY3ZdqKDtpT5BUyA21ZHZteYpE4wxPl2sGGqRRPjPvwcIBp8zgM0+YQobO1F9eWEpWNv9un2rr3YdDGnW95lXtzGrjND5+VopjeDc153AWsNHlwmAGQalx+H+xB4jbJqKC7xlypVOH/GmL7HH/El0vlxs9HIc8A6PggEQ3wBiI8pfCLWCsK6yxQI5vdTgPApbffKT7nVrhd468EQAVfYBZYwk4vkUvdkRLEVbtvSSYQn4T6FgHk8F91G2fI9Pl63ntP4L+w/vPqS3T7zP9wxD3BUENVRFHKopRT0l7gUNpe1ILznSR23Tfxugk7UnnhUWWKO10rtz5AAh/gitPtXreNr4VnkmDDMWCvezbsw1Z0YtRl+/f1fWsMI0sC3ImF2wllxkNCExxb6cRLXVfbJaZpMdzGy7kIUHlRyr3WAIOysu+SkPZYqtdPHxf16SW0g7y2Jqen3H9lNG2Ty0kCQHUlvnpsGz7uMrcTaS33LFBd63c2AozjqvAK1VDGEnTy3OKQzZ3RsevN3/Zopy9Lf1EKezKqf96J7w1YFPpm4aRm/RZcraVGY8h+pRk+pH2HDoVqm1NeUuvUiCB9910T1bVMt/wyd+4xsKq75i42n3KK0oVUigy1zSkkDQQG2P+JnyZ5bXrVcPw/AoCX45NaMd4A1lfTFnn1wwbv+19Ez8CkdkymYI+u3PLd5A4H8MZBJrahWiETMklN6vSKJ7Iv6EXZw48C8rsdV9LXWjbDwhL5C5gHKmznEGj2b1cOV6IdUe/sgLV0dqpTI/ntIg341n9o1e7CBlSANpsBxKlbqWJuInV8hX+dpVBB5j+yV4scO0XnaM5cNjWI3nxVvmjdxQT3YoOfSxbmZp/e939r2yh32M8LygXawVqvTx9XXbnjMcj7jW8F2W0RKMKBRMXv5y4t5CJf0PE4fCtx+7MareyMBkv/hgyxF2cGxnFLJdCMvH89yErUNHn7Eek2k7drF2X9pGfX04azUx7rttVZIVYtziBvpseXuG7LKPOEL10fg1HclAtxkHVqIpkprfR4T/fzI740+tqBLcTWf2pLuUQtzevHD42xiy9BsXbIMf5uP2z/TqhYoH1GobD2h4nr8gG4WYk6rptKk4wG7GQxhfV+z2Zf1XjMwe9WSOBx9Vv2zNpanYTwQMLoBNQBsmiExo65EUOCqyJhc0ou6yGrtJMI40240DcU6B0CgtIV4nEJU5oad2zmlet6GoQDQ4WDGeGdl7dT2d2Xm7J9Eh2fzeUbu+6+yvLfG0RrmBbRUDu2PJaCKQeUrs+Vm068IvL8T37TbP/xPI4+nWfVvTKQIW0jOqxJr2C+2nIX4fOsD1ykOxVFRp5zWQvlb2laPqOWvTgs5eTw0ebCGiDCRUU8G15vHww4LR+Ir28DEqfaUD6jBDVN9CwHyT/tfk+POavS1W9OWLYgBEbyvSxuh98U8+dqkmRXm2hbE3AZVbfDX6YLfz2FNT6w1bbPo8E0D5RllR/0foJj1Ad3nPLacpC7rhtvEpRpnFl4HQAxdoWoHM6MHiyXfnp7GqXzZjeOXRAqJ0xZ+9hoJxpo2JLtShtONGytmTCh51oUtuBKkUjYXkrZ+S9PhQooyltxo4H6a209HhZOf6ZU8G2x1ZiEPUnJQHPl10d4+V99pxXc0mpktSeqZnbe7ZtTMho5cCWyFs3c4BvJU0WFcl/W2QKMXO2NF6rEAAdibtOhxTZXQBLc0diultbLpGawLlHcSDvkwLcGG+KiEHTaczmTAWPGGQaAVh02MzKiGddCk4YiP9kdZytFH9mgJMYXQQrkOogRrxoqTKZPDxlCLqaJkxwwlZKQHrOiU9hNwsR6MlFVtdnJUVqowq4TiZtkcPyTOpCm0+zmeSTx8ptZdYPgI2gAr25QWCvpRY/IyiHLYX4+7h4sVG0ojtskgfConUSFdmXyNtd/e5syT8mLqCAW2kQvwZ2QWwkn3ZaOdoi+oTmCd60HTDhdKiFJxE+JxCBKEVcCO0Pr3GU8s9tmroXaJoDUJ0DGy/Ffib0dnwAj+l0JO4RqRNSgf3CEJHkaLdwURu80PoECUSHLq7iD4rVOCTJcZzElUy07p3y47TSrFt+8Xl7JF3M3dGboAygI7ghehSrztw3DQFkVlGsSpEAJl3kxD5UFJzgFSkycJAkCVO8723Pyjpo/Pu1fYpz5Wd+7i6WikmBv87yaCYJ16tLe325SPVFLPGnH0BKiv4/57y7UGT3zsCHBocHVeahf3Td9sMiZR85187Ib5xJD+qLyov2/9ahXZFp6xO2b2gW1IiGMqhjjLEZSlDKnapZlDak9iytqLXB+KTt/X43Q6wPzJcC8mCDMIdhpUqxKSkz8vSv1wkg2XJVMd6fD/pBhAkoeaSHat0PPtf0YDs+6gVTfoX+0XNGE0OpRPcanr3tiCXPvwo8IQHYQp6681wYGDkV66oosj3tnS3z3cfoe0Nv5/KgTTnFRge5wQWlQj4vAy8lFzitU12qei4XJAyp5CaeRjzfG2zTi8XJjl/v4laNrJ85uUo8hs5c8sApA2vtvzoI1G4t7VqZ162Vb+5QnZEVwWRKpnY6Sp5UG1hFTcyvlrGpnaU1+JuALENg1P/FA8E0okLCMuoeLPau/owxuzBuuOcuoWJDEs0707ZyVxxDWiX2AOygXN9WAEzpKtJiJiIXfX4hw9Who2Cl64ToJx9ZOsfONJhXITv1eJFF16I52BLAsJQDstMqo+Zl5aY4PJFdXHA8Xt/HdLtJDjy5s8FPEvh/cbbW4clLkVO8/1e3J5BNCVOC32d81o6mrxxmdG2TO/I+hBH5LM6tgkdPPObervUfhgArNchZtB3Uw70WsYQSTUtfYg6bwUehQgd5asO3AFpdFbakbo0BDm43HT3rbZ7uYcufpXgo+uFb5LsE+OPTUGv7xTjuOvJF9ZoAHNjKfYQwyO3o5MCG8SY6SbeBbEMPiz4Pda84T8mANtWqs9A8QVHtNkoEu9AwQnzSLe+q51HT3bNbxMS9Nk1jJ6MFlL+dgBCFv69qDTj9+VZX3BZsKnOLTdsDwDnowpZzrNbhQBJt5U7FYrAb56ag/KJriDfIi0iv7XG2OqehWUVlXb/KCZMfHpTx3fkPuEsM1oq2ar6RsS2R6Psw/+1dqZwLjIcFD7pE33SL9HLRUZRu+9mn2JNxmQDd/QGjsjcDn1SLyJlyoq9WVIPg3Y52T+Eb2HXe4FcAr3SDterYgZQFqSksdXPrCLoJfzlzNPSLTk6UrfwmocvjFizA7hxaRZraWH5AhYd5SrAnknOYUT/xqK04gqOAJUaMsH/WcAjS09wGZIcW5lwpsi718ip7LF04cD/VVXC8byeMILHCLDcIdwa6ZIJPLeTahFicXGzEkaf85b4mh7K+Xm9FFUjuQthdsLeiqiRKXAuSU6x/PxhSYkn/DqCxgKiragTPhGdyJrsFdhkytIKL4kHl3ry6QR+Cn0c0lZXLhnnld4haDmqmGtfXRSRTHmBDfT3A5Huq4sfuPUjrHhiVDrP6Ec8UdEFCFlPaDdfKZdHRuMhZr8g4p8Vu3HbNG8mtfkE4BFOMHU+4usprsKr1oAuqQRp5Jk4SrMBJ0QCw3fdilSKH9LXfHiEzFOxqMXA+alP+ca0D0iAIK50jMfDRFkIITSqVJFbwfHEVDUABUCiFY3cqx7s/j92aRQY9JIgZYoqlJbLRRJcOWl1Pw2aOCrBSC+UOJib/doMMZBTs8s4FhuPoqmwxnA1nGQ8o8zxtFSdqwJRpcz7krulCagZ+uufCVY5cMGDTDoo5Yg6VnT5sESy12qQ4FQcIJ6wrXhvqF2S0XcdHl5MaSVYAeqsrfZFpHBThL5U1T0qZSJd6iAPus51k53Gt3x0FXlu0XQsImFpvZL+UFOPtjQSzFXpbBnRjk8eP13z1TgWKr7iFbUJczUxe5wsGHS823r0JjVc0CjWHsQ5+8u1MXzAxAo/I9DJOxbBTqvAHbtG3zQYeCVsdX1eJlVXXBfN0GNaUp5xZaRnpeanrQCyhyyQJO0dMOsJlFeBJ3Rp/FtgRrIY8oYbuFNjIetv3WFV3tNPm8l3o0VSX8oIlFI8K9KljQw9VIMxM0k6/72b5ykWCTRtouOlHjzllXFMTCSV33dCOmzcfUuLFnF8+qhvUpRQyh9t8RfFdq5N9KhxQRQAA2SLh/+cAMnsr35FVyFFX6FBJr+G3kqgO335+bofWsK/mLUuMQDMBPEtHyPruxttI7p9jhIaNq2TarkEDgdqxb+SZG10X6hNuwsW5iJuhcLSUD93H7Ib6HtZ4+OZzOilSmoekQG/mqOFIZT5Ej1yywkmCHllZYxbjhG+zK/2iWMs5hrnxAYzfvU8kBGCw+H60uQloLLxUlpy6zJLDMXZU53naIOzGBysweJt/SzY4E12feqeDRn4sSGbUqoSkQbVmoHzfxEYLAJn83DxvXE3Qr39OJtnLi8YkoLw51lwPdim1Zh0iOXNYhZR3PfuqpumZDc3VoCohKaybPAKsVQ1p5gE3FntEvFyz/PR+QEMmIhJUNmfLbA3+wZpq6sg3qTaR2OZqqW1CMo2YI8sauZP/zamVP03CnHjpbGWPaIO+7xr53S4sSEhjAgUtVKS/QPcLuyasVj497ff9LBsyNgADW8PuTa7Cksza73WwZbOzn/+WuqT3Nyy8BWA6x545xGsMQP9TQIV0sX4HC7V9Wv3Teyx8LM1LFcktAK2lbLJQItsRyDyRvVnYb0CFtzg5CCWoLE7mJmhKLj4GUiCU1MrHxjSuIMgoKyR9nE+/TaJCfzrQIVQKbA9/GR0L1Id7380c/GnDkAGKJk3SYefVqsI1wFTFIwEL/TnOa2qmySe6+2WV1Et+XkK2TsE+PaEwgVp0y4M87dE8fvtG7/plH5s2kl5DTOCSDabIEwuDZeuP0FQqwifRXYgyiQqPcIHPTjinLCvb7euSjCab9v8u3Ezzw2afkG/qCR+oLqZ7Gf/nDR7qCBNfhTO4zuk5ipn4sDqArW5nIyZxw8Jj2Dygv2N1JUDF9NI0/h8YrgRkTNvco9435gt1DdwjSwmbCbXcnUCAUdUtW3U0Asjh7MKeY/vbNe94xfsfFkcD2PBS+ZarLZRU7nXLEe51mq8fIsTpGcyEF1MTlBIbT6nlldRsnoj2KqLl6NTkpvwpnlyFd9L5DBU6bVcB8Xhdxyh+fpsNnHaRJaUko81kFDPdcuA15mjGXA6TQ37yOIDHM+Tukukn6L76YRKNETFC3fvMc/kFGQPtlKROsk398eCJyzuqBwsOZ8lgJgl7WmXrjfMa0E3jzAuxCgr5NcCMyVjh9ErjREdTCZ6Q3vj+RlWy6BidluTPPQMkiQ3c19WBn/1h9smH1GTNN814jBjrDJGecbVgS30YGkC2Cv0QcQ7E0eUJ4ewGkscGS7gZiY42PPPneOo22BgDyrRMnSL46gnMBVv/pl8FH97A/NUsBHo3b698azqsepKXEqW8xD8A9xyQvkAHHADv4DYP9pCRnStHeiTyRlsyCspIGAWbFM3g4a7ZAMUfB6txEYF5yarC/Z4NHV0vKUcgYEY/b03GQsPBJVBkL7Ko5RhhL0weMOvaraGcRL25VvMQBhqjkbe6y0lyRDUHdiphzFFTxx+n4TBmxXB0YambMpQIGg16sZV0/AOrlPdb9Vm5J+Y3kjUjyV1a/9xwk3Ee00GFzOpeePjUWYmEipQ6uiMT7HcxKpNrU4NI9A6NvY5q5Lr9MB8AyEzI0j2qLsDRY3Ft6M+wI/kKB+DAIMXWSDUWPpMQ6RquoC8hNUc4fW+aLhsUXGng19Oi+U87qIPFaOqzwIYdnWERlnBU20wuM2J8HanN/Hgo1o9sHWGP0e7ZY9RcJqNF2D7gE0a7gn6x+9tW/QwM5PAAlAnxWgKqZd2MsRxOnaLNRAKVJfdy8jBIAlpmr6CvCdedKFyDPjsltbWb2nBVjfWLZ0T194YpGa9IL1l+pu1rfG9RpQOYdmDccX/ZG+eO3xW6u69d7SL05ebKsB8E/l35tlQXu5TUV5M/v8N6/fr7raaOITnrWZD88/YvvpPNMNLFlQhYBqaqjuRogTMAZExScAAA8DpSiZPF8hQY9YTQxRz1yz7Cegi+DXjvpUjc/jj7W13v08HbyQFV/kfzfH6ajE/JmSngdyksWW6wbJYwafNuPkEyzJ/FhF83TcW//Dm2Zm6o6XaO0dDovYmXaAHqD3ccOrYfub2hyloSaWNn8r/T6tnqNUWAoTixAgWvK3aTXHGnHsQd3WBGw40SkCuMTm6a3yd06e3Ncy7e7kwo01K+Fi/I6aO8xgpKo4qIrzjhibtVgHkc9TKloNNc0xxtzSFCl1vBx7aAURBSrmAN156juDjYPBcU0w70o+YbFebexgsfrcvHwTCsFbSIN0w/o9bFaxzqxTZrgNJZcWWhf8rXNtHNrFYIdw/glg3URXdriWXGJqJd4EDL0lGWl3Ke59g94dYtBN+YR5+NHmS8dAyYqyTW6G//8j6LCsQuXyGaQJU5lqw4V3l4JeO1PnIJG+NhKulHv4Ug4AewhlfjYQE2uUOQ9Khs0+QHtcRvFk76Ov5REda3m+PW7e7mKWheZP4gR5NwXh+cLfWUMyUPdlm8ErSeS8TtmneHdQ2DZEXM3SFAiui6OFShEeU7vho04bHR37+esdwfcoAmsdEcZ+s5GYLn9kM+dTVFrOfnyAD0ZrUEkmcKOE69KF6FIURzWt7enAWtswiWPcz4gxSqnk3FJyuM8NgC/nKwFb5PTAPqzj3jC3BBLC0522ei7c5DJmcJc5k1do7qtr+VrhfCzcZSk1YYt+x+1MUquBVlKL2LOI2x7olONbrvmEOH5JdA2azsoCOGR//CW/1NOjsp0FwnWv2/R1x+38pqFHJAkNq66f26hKjxXE7x/rT6wyofc+WNEnAHwDUcRII4OfNv/i0RZba91QWz1WEd/brCeNBi0gogG09B47ramSIwlMXaASS4GKi/EtkZJUDhAnuCNDHFwVE9Nv0Wfk8QjBe/TMJU49bkvY8PM2VXI8Vx1ldD6EH4LmBLLEftxZ0Qf+T4PMTNvoPrUKUfgeknBBkrZsULM+9Ti/WqSG9Zy8LDnKKRrhEi9FavQIn3kkezPRibrkW4BspI032sNVrf0Pn+L/3Ifl57qE5a2b29rN2NqUp9ruuNjxISHQJZ9BCrGVIUZw9vu6QjT8NcGqIHHJDieUHdB8ANUkquMRdi5kJaUOxoUX9klPigW41WV6NWnLIUOg+w2qWXZ7r64r/jCTqyMSSTHfMWdZWO3Q3CH+4RQ86Vn2UZRCk2luxDp2ZlHQwC9YPQL5Pq97Pwhs2mgGLb4G5ZM6InyZpTelRw+EWKxBN60uM3wraEgy/bzOntgmJUkco0T43lN0J0h8Utp6bL3Jbe6z06u7GP+MmjC2sFgw7gdM/Pb9aYNIVQmGLSMygXcsE3iWcuZLdVdF5rH4S+PoiUEWwUWNOCLxhbX7KAGMFy7WdYwuxv/JIdaEFq8Vfczt47UP57XQpU04QxArMHua4BADXR4R4agV8/gSfZNBLkbq3Dt0l//H+8raTPpNJxk7F5g9oEeAXBUSuEkdfFNZpg9NaeQmrCdRgL5XlPpGe7VVspht8XVrcQyLrTQpVp8PhrXqW73zIVA0oUgvT7CVl9q2Q+37MoLmH/0AqQHT3SmDHC6tcmhrbjQQ8QSee9o4z0j7nyzfdfbVfG/2Fr9mV/uMBfCuz+jYBnClCFSQ/JFJ8Nj47yppUyHw/H/xwG6OSfZNR01/hj8Wo4A/RykIMiFV9n67//hW9eTGo00eFsJ5e1HCEOWP6pQ6q57/yClBYu1D2Acq2EhBhze2oN43W7bcV5xWg9r2yU9uknObe343zDIGPx2BYN1FZpn26sIvCN0m/MvlJ8gijpuJ4bRYR5C6BWopsE6eY5CM5fmUAhBP3shiEtao0P4i2Vqp3BBedRjQert90O2fy7213v8dPUfg7fkvfBBBXD5EQM/+eh6jbSMrHdIX7VtdfoekZGNR0FLqCH/VTLXUoLFfqoMAjC9Bff4DfPFcI2sRcXh414oPaNEkgjv3jZ2d8+wjM/90NO+OS3M4x7dJDO+PD74ZbzSwWYOKAJNqZLD9qO3JtjdvA63czRdjY7HDw65DmoLa2lAU9xZoFRMxFV27bpW8DQbeDNeRjGON0bhPCZJYVgIggzBNUANDRydLxs0Ei5vBchtxYVOzbR3J1SBzfrPxUSnVfTOXWrZqm9dLZvFy1sFobvwvp1YGwoJYrir/FnJRfF4m+DetibLkT5dEEgG1UlWQQlVI3rbcpeczvl/IrMzCkmlWOClvlB6P8rYVsOhAGmEkGBtOWQgAkjujDJrHub2wKeUhNycdkCuSJlRmXGChDZ8XHEUHjnqQQcKNCYVDiUsxANQSGRgDQ4kj6PlGW4dDO98lMU5jVDr2O7yHCImPFc5FWVBkNCHmmmMMJS9VJq8q4ELdCxr19JX0bGd3uwpNtQ/VAX6FByrFVl1/VvWwev1v15oivYiPgGzAPIUeyz6epbJopehCVH47SJVVnmfI7QBYA9SX4lu9xYH0oZi5TSDcWCzZpdl33Xwr1SIqrm8+SLVlz9zpH7tDAOU1ndGTN5f+G6QWpvUfbjC4NMWXqPwTfAs35VHJHqxcSApxJitkAqNf6dRsUD3pxI6DlijiiZ4xm45eToeZwDbpLZ6xLvWvaAMZRaF9tTJoTIXgCgiFtjs9XA2mvylDnIYx1r52kY06EktKWT8cRidVyhpwQclsy58mKQnYbqotF2S4l39keaGAlbd0bkUzvTX6QxA8wgQre3LDUK2ubF1dZ5/814G/3eSEMuv/Dfzs59LvYjiN28g0xbE67xxsci2UApxJ+98ebImyP5SGjfe12cav0ANePGrrfsH5VkFBBM+KsZpCDgEfLsIuPGRdL2iqD8EC1q95/gWP5d/eVTxt2/y8UYKudp7HqNJz1z2UQ2yRpU035P53SMN+VBcnzyAc4PjHKKivJzrWs4wmVRM2F1wnU99ENyX6E162rn3m2UfXnGEkAMIegTM7FXqBfRHyY1JJ4/f+R1sIpHx7sJf0Efcppo38yQJn7Y5rmN4W1YKYDvz6/ZhJqwglNfRoyrYlaMTpWj22oxGSLbKNN48Z5PTAvus0JckcjYX2/NTq4l+1Hm/NXwmITP4LcOEvIn9FBXjW95/CHS8riHMeceZF5jLDUc55NwD3OoyGo7+GBVijVHsnPdSZ7codOFIA0YHl1JByuwQfTeUz4u9Ht+BvbATuMwb8VmEcfq6bFrdYCCEBERpdRuKmkBJWyJIsXajuxr9OdRe+pvQEX2vbzgRkOkRhU8MlqWpGsP8LQmeLz+b6DS2VC/WRMdBr/HTFYS5ru7/+vAdkTA4qaU8bwwdhLbk5nRjl2UQ6IfgDCLh0p1Gle0YQ86nEqQD9VTZzCjgP1zNQ/uMK3rswj5pkec5FuZv13vyDajuXgC1ZVrb07VJqBz6yRAw77ldLlTW9/JEbeqYpPnsnjJBoycnuXfQOT4v9cpcfRg+ZQEZTdmkg2+L9WXvRbsLgjIeeK5dcLwBI1plaEQIc7ob4A29nMZiULbnwDktbdFOSgObsAv0fyM2iN79EzuDsAxkmNQQE+vyDIBHexpNJwW59ug6xFMPPx3uDARAwsWY31qI6QZt1n/vUb1ThwPf3DxqBjSs+bD8K/A/pegFb/rtY+7GXxQ70DIdU3hAnVzi7tDavPfB4YzkN0FUT/GceCwNrbfIFr7Eq82AIEOzbPgSpmCpvN4t0aqLDhKY33yHsOiVfl3mXZizVPaGv5g6/YAk/i0713TnHqaONx72usC4SB0ZkGPhCDIX7VPd8uLaBtjiWiEN0XYTP5N0Pihc/7NhtH3wDK2O5PvVUPQOTzvq7RviHfJaMfu/PYG6K24KbMY2vBGzWWZrW4qwvo4ktlN6MUqW/iJGTbmiYKeKTwLi/kl8vmFGuWlmGpAvSqkSiBsLFzTKhV6AUQXoq16lPSXvD2NTht9A9YOlWkeBlpmGTpKJKRSif9xNHfBED9J9bszb8YQcmvZgnkbX9Ix/6UwYRTdXwdwxhuJM9HyuFv0rXUJNnYNfCt5vyBt1lEpZsxDD5m6reuz7qhQnJgeYtG3eMJXocPc6Xk9wN9yPM0mHF0N2G1Kf5OqhkDefg/0QDPluzff0hQD49mfSKQ1ZH14eCE49uIhrVIMnUTkic3ld3u1UFkxLRkscCFpfDN1U6xN/0LhHC1nxXpBD4KntCHVjSQamfVYATcgdWPq4C7AektTJql5FlKaUfTQvZYPd9OPUeFfPaKgkkYXvyLwJjIwOkMPtn847S3q5taCBtZ+6qwAEhbqFgabbWqckePa7+Z4nQK5e47HtuQrX9pWMmbpUZxwuEUGfJHlinfj7mzlWmYprggATZFW9ivgV7t+km396+RQmQHfW5oJVkmLb71gcKzH7q3uiORKZmfjjz47bHOya4upBT/NYpJF65b32mjFGbzOohVyt4p1IJz0uTPKilpYELH7HxH9Z3vwOQZoovoeiUPrxytER8ucLCCUu2JReP46uoVbxju2gdUEtbDWAWtnOmVUK2DnjbUY/PhzPuINoONnR/oas+LGaLL3239obqlw3K3TurerC0m06RKD2mt9EZPuCejGaw2jlzIJ7tBl4yOL2GtuoNfydYFZqY0BH2nzEK06Y4o3sTpBWJySxxTykr9ahLr+WPMf5zPx5C6h8Mqf9NVd9h0pYNpGGlz/ldAVnp6sEdsNbQefh48Yy63OVIr2v4iISrkmOd+qP1tVBLsgAzKjbQ/CBC8MQdnFvmg6KXWABM9v0kJ3KYMBd0xvoPzG9cI5HWRs7ZBjvW1ShDDPF8r8bqvktSDgxGTAxkWsHnawDPIsbr66/xaUGmPaO/ri411uKKzXX0AvTEz2yYWO5Hcuaz6bVg6G+vXQni7BPX3bUVIow8Csgp2MPGmZ6Zw1kRlPa2+LeJbJzyVHiaIyF2z1qM5JZcrX6lQ5vrc36gXpQQ7l0S+8sPeeY1GyRB1fiJqlJJoGjcE+bShuC1Z3gxJUZ0+KzKfv/wkkiL4WpOYfEL+gZvu7ZZjiYy4xSSBdkQpofxuqIETqMw7Wddg34YbvQaIGEsCgkan2bDjMeQEyk36GeHxVDqv0N4Bws4xYNL9/Im3bKtwVGQtpSgH+c/MkpcAFwD5Ip1gKpraD5tK4ejAKZvVolUmOl+rPJrtpRypGt4uBmTuPCGVN4D7ujkKR70G8h1frBB+QK3rzIzcLZl/Q3G1CuwduzT3ebrbUcHrmqebTC0sGxcLqg/EBySx0qNv345vGmY2jaYoP0dXDagFdc6XOF/QKShxC0zBDj45lDi4p3dkDDZoUVyI7YEERmHMtioyEs5tffhPYpF/NVn2VxpgP4tLN1YzvhhYP5ya0ezTNIIDOGSVgUSpZNV4ghJJ6k0vp9pU0pydPWnTgXKjTovM4cay152f09kmQlJGaANePNGRumpIOsyrQ66WiC/lkROVOS3PeOjvX72B8N8wLEavXS76CeyBFO9SsjotyZuQc/Sn8E/tCJH/65bhVEjwEXsyYsNbYHI4v8gxXGekY3C22YWJLOybz66DO8thf6UmaO2lwP16zh3Ke9R6LvltWV/UHE6I+hPXstMF48XOOCdeP9XASRGuN4lZFAii25C8zAHbFME1PjWaOVsKyuQxJZYzv140Tn9VrI8KbOPlo+dGGBlany6ANoQc/LUY/I0PAiHgbTYOCXRTlN75KF+vRwZC9yNkdATJs44IyzNZem5jXbUmhl7KEhtNWlKhAmyLQbhPPamOCheOflzLGwX5ylZfZXXG72+fPk3RSJZt43+MhUPQwJiTc5o49DRZ9vk/VAWdAtE3SRdbwGCNIW5Oe6FViOKYzvffNmtO0JURWRXwHT7ggffBibekZlYgZ4bZlVvHHDCow4sjmPM4JmMtZ/pR23f7l02FXVMZga1Qdh1hkJOtJjKOPTQBGkuBooTRoMMYnXj114y9+ogHJBDy+DvmGYJNvMGV4xiGO1qyZg7XTXA4vYJFPDbQIvSBFVbJ3MUC/BVAIhmN2V+jOBlncmkCJAhldg9ranEyPPNkrrb8DRtZyT/uwfebIiCaITxOMogxZPzTVlj/sxod7QZSl+OwZh82wnuKbsbE2JtnDlXIEyuNPktXYOV90nsMmUQRjJrF9VAN3acSwLYewxDH0z9gRaO/H6eySj3JEa1Scd4Xcj4tRpHAwjyjxBFjHhWC8ggWKnZX2l8uLNPG3Dypssupjd5jArHR5CnfcDpbGIOBqmX2H4LCO18HopIVkWu9H/TcnDRZgXjF/FrSMWr8BnfxnKBzgweggD0/vOiLkm56I3+9ZwK/Z99CesDOk3/6EB7H+zL6KLpDuYVUZy/T8AURmZWYDosnmsLqvMsWeRtRHBLj4JwtsCRLAiTGQ91CJYBsN1yeRW4eXVTaW7jc18cvAHMPNjKDcpLd7/p7Ewa2plHA+Nxy1pbaan211w2A1ECiiuDrKGuf1SKQjqF4mk350tN3QaYkpp14T+2Rl2oBT1LGJe80nWMMb5yCEMPJbh290APmwC23gAVjWkBYcmE88GRLTR5nId1FbjKI7JdI+cB3cqB19dVsUiSxCWvjUUQgUYq/vWRKaOZA0lyTk6hsxKDThNiTim3Cb8cJCD1zfGw/MGpXJNTRLk4UbfIHttaX8R7kca1KkK/PEXccZmPzmv5tPKsej4z1BYZlICgBGjHCFPYPqSxFn2/fs20aaaiDZqp0DtfOhBS/aPBRWKVz/NJm3WGmUvpXfoRkVF0Fk+RRklE52Y4YOfQlLrS6bxr/Rx+vjuUspPoE9EanNbwj8nhMTG10uTrVmFdfgQOY3yN8bm+CmNsskKxDTFn+MBtZ7ASRKJyL2NWRMKTgWln+B4CL3tym2FbSxr23NWy/LD2rED4A+65p4aPz4CrV0bzKruTst60tCVfnN35KXb8g0WRf8GbTEx7e5VhRISb2mdI0wghq9DcbubZIcwR/A6Gen3IhDMJU4z5M1jz4978wBnb2eABG7MQ7kSImGwXTa5pi7pTWA3MveP02IBJKeOfr5z+jV/GXSef5z6WMjR2DUsLCF41LUNNSLuZ8/SRkYtV1TqVz3cPZfA/RvM5O2z1UAK29q5OIXvPY4EdySNeRYWt1I0aG9hp4/SInF9qSU6p78NXciMt9Je57Xub5CJ19MnRGxj5qerKn1ZzSFH1gDBkiYVUMdyj9i3gx2+CQBKMyQURnquGfaibdr50lhDT5HdKY790AEHdDPHL1M53wNk22kb3DRIdJYqcmzUHTlknxFVVKp1y17Av43pBEKCMyIPuGZDRToX+VTPC6ll5ZAjK/TXxhy+tA0LpQHLeSpUIGE0BVtPXDlOUTojeN2ffEEWmXcZWvv159mZwIvYnZhu8S5xS4gFf7GmqIjjFQOPpFEp/WSuBFG1NMW6cVSiOEum0XWtRgzrYGEWwkq5xcMzbcQ5XzFtUL9X/7m8uTS8ZuBnGbeTNlT5uK5Chp4xyekGywg68dPyyZjj8qsj4Kl1do2t2ThY0uvdcFg50a9oLqyLCCazSkB6q1wKhOHQ0CNaY6Kmw4Nu7UBGOCn6bkRsWd9tVQ5gwql+tJWleGY2KrGWoEkelrTu1nnG3SQuPKcPxq29PmtzxO9ztF72wL+KXANxq5ZB9R7PYroEaZdBkNggIm6l1QYK5qWbM+Q2VfEmj5z8YxyI8AhCyTJNb0m/yg5D7ldMC3B7Stw28J02VqLsz8fGl/CkyRNKWyl2nd45jhqGIkA9TgzcWLpVU4xH0kWbfCG/qSuBLutOiCgt0P5Mk/a+4xRecaYxXwecyJ9gTFoOPz+kmXOj+bUyLppOEf1IFFxnxVSf4FZ/yIGDRKaXxd8HFNkjyNf5xxz7bbMZBtSBTTtCH34oITTSsP0McxldN421ER5kulEa/LWvIMNZtoS5nHfLFl1UeWeyk7bN+o8fLOy27LCNzs6azfwC4VkHpfSwaVH01c00Xn12iYO1tNCYTZYwc7u7Qopia+a6OWlVfU4L6zB5ZV8I85qY07F25QS+sATiU3CRW/WavOE0vVAJe6zvEkeVvEQTtC3v9jt/lk2Ko9gXAz+oYJwQHynC7oJyrGz9a6//jH8Im0XyVQHxTaydUS2KZizhHUP3eexzrRg+cJGNbTTp22GmltyKybQ70wNOz+hVmEqgWL5gdObCxNAAJ135rgvIs07B22Dsd8vquJUXhVJFG1cvFLyemwjBQv/l24o1e4TYRv7/syamQY1rx7OOgn1VtGMAM9N5radGBy7V5jqWciCbIjCMGzy5k+X310DmctVaLzCHgpwazFYCbnCKPs9EewwwMIRJ8zNfP+evS2glx/y4X8T9FScwV5IZTqcSGT3/VdjH6da83UZ44Mw900VvWbRwKBHxA4/eFl6wpy5NGWOJ4m27vJdFlV5xhL2FkVngmURDFZeOORwP+z2dJY1YcNehbuQGHMYKu474tlMAlqLscl2eDiEe63imVecppiC/0aj1zI9Bq7n6TiR9QWD8s4i3aIsYJpAtiGbsknT5p+NqaMwKkoAu1229ekDdp8QRrC+zuOrVKGwVCdEk5jfmZwfcUxJq5c3W8Spo35BwgWOrPiJOjq5nh+1ltbdZFgz+kDzs88IntGXwETCyGX4TzwNcNI5+YbMOes4HDOsa9q9nOmMuAniKVTQ9XO/sKDYhhc6ISzsYTtv9n0UvIbOJ48juv8TgHsR9AbYjTo+TYRFnhkyimOhcWkGrzZGMobF+0Gydl45LntJm+qpbs2X+Ku2q/zJ86lA4s1cfrecHMNUq8PHZtqhvSSpLypA1oQwEGA4FgQNyyz8zwVpA7UcGaO7RKVbr+JYwb+nxi3nAXO4adtXdK2VjTKXjSuvs7sXpSD5fQtawYRxZbPmXEXrbqi3s9YxnZ4GRVpUSVfO7yJTJLOJfDrv7B7tI3af0Wmrdh1uMeFw94CLjUQYZ0+Dd1X3m9Vp3LVwDzC2ObBze/fsnVp/KWJwIoTwbelmeszoMDc/oEQ6O1Zsius2X7IqHABUthf+o4564FuJgjry5PQJ6lTX04C72BOMRfGVWhVwra77enJcb6PSoW7FgLEGViHGhhxipCR3sx35tchzOFjAe7NoOmS11HNoqQX3xAL2+FKcEehxcES1tmVn5iLONEKoX/XFgueWo3XzQftYXOUrXM+/STzXR0huP4k9GvddKyoLAxhwX7IaZgRVlqs8giMre1WvDPpwRsNEM7CZlMbNE75qex1EUBrGQMf6wec+LJHsI+kGiIzCOd4D0PBZ83SsRggBbWP/tTFhoEAS0m/t5ho+F6mYiPYv4f2PuMLW6rsrvppHIINZibuYNwPdvqDJNGbpyLTHhIL89jfqfdlruUrJHQ2aEwU1LYvGbaZD7KOdswkONXaXinRiPwX+IFenqa7KH2p0UQS/XFGBu5ZAnLnUt6ZGuER1TUWwYQ1uBPfoMQlHOz4irjDmm76147/406/IKQf8Aci7GPv0ToRjwVuvE5whtFobWw9jJT2bOSnOgqJf5lmM9tE8w3hmmTRLy16XTF2pXwuP8KMeSSCTBdq0sICM/Nb16sfupvMocE2IunsxmwQVplyErcpHqL5WwkelI2D5Pgu3H1kYFKAHyCAmZ4nPhWxzpBMFyWr7qrBsEjW4htRIJJx171Kdo2Sbu+SCzkCA86sB9SVdb7L5iy/oZwRiSoA4fJt3gDvsmXDbivMNoy73EXtR48odfOUTj/NIznecG8+I2BwEKsJjD9CZGXln9aWNqeHMvBMQhatSQqBwMejBc+KI5lX0RwD4/Fy0MZUznUU4R+SJKQhZtiBFlaLB7aITCTyNdFSaWYQgrgtbJX9Nd8cwhS/dCfXJPC4/xYOocY+Y3zaqHcBLwDJXbZ1k2hwCGiRv8ilEejZJa16vUXyNt8/+PuUkIoyXDzehAfXZnMlyay/pGAtvO6Dq9OJPux7pd6A52ge3hJeZjdSNsM2pMgNvZ+7IAqUhKyFElm9nwCpYEjLsZMsuYbrTzIQQ84eUCiX8r1O4L/n9g5fMiRPXsItWA0BQX2IzHMaiscYr1OcZiWz6ZsDB4evF3ldaGUQEqkBAjdeWXYTLZvbyGH8cRO54xrs10Jec3wkopN9lSpsLSI6FtmbQdPfKJFgf7oLdsrcrGqGlZm+Mw893O4U4K5KNUV7qoAJ7FhbPz9Y+mgm6y+MRsOXjUj1JwfKvAJWAv6+Sq/aTH8gAf+eRvB0mvxCNsd9YTiP1ASmId5l1hbZKd+p1BUcMD4S8YHOCJvvyyQuQ2PfCe/UjS26uW7PnJwLyIncf3VapB+a4LECwPLk2FXEU+B75dNKHdqVZPiDD9/r+28w5sHPPCiQR2FRhnGpynxbOH/LDx59fosRi2O8xrTA5FbNSQV/8CNTctXnUs84vTz9c4txI3e3iTPXZonhrtIMzuJbAxHl3c0lnCHq06FnA4WACyKPJhoc8/v2JNPaRW7gVhj9SkUSBefgqY3Oi4t2qSLtxBiokc2XHRM4gIXOjMjGr//t5WVoe3eNcnuvCrCLr0nOcWLW76hreEBNfYYuHdkooK6hxfCMhevhBIHouoFqL0K7dxoj5Gj4LHi/1iJvjrsdbtPzM5vMzCiNIscnNVChT5K9MaTK0BMwN1kJT6q9xmgubXUgD0UhOuxU+v6C3I/MnfhxOFrNVAVrJ8lxJG0NoCwof7qXVSylX5G+IJmP2H71E8v08RkDXP1JNV1a/xW9NE79YPDASpRnmqsqnXm4S0x0fMvJvuiH4HLZJfLZjI+nQ7sXoFW7Mz1bElWri4INWTLggXBAIDCwDAv0O6EDkliqPeo+ni4NVANyEdeU623cDehlcWcwUFdz0GLmYLwwqAsQyVC36dTx5Sj+W4BjjA0EjrR4Omml5q+I/QXwj3QJ+gggZ/vWluZpU06gceUeBIcfjt+9DSAa2JAFv3d00/IENwpEtCOdzi/Xm3uktxdwX+huOJ8iqPkgkii7LLW1N0bF6wxTI2TX97CBfsPlAwBPhY/Zus23YOgB3QEO95PNgJjCUIkxqjLVJENXQx/FYf9KqfNdrERdjPVhTi9aPo1w55XFlE+sYmxsASKwe9Z8RXGJVFbb3Ry3fTjGEser1rVQHX8Pfcxf+5Cu5LdR2AtS74Un7m8J0QQ30B+eqFoPVQqzLWmKNdjBCHDa5RygeIo7nxf5NGcSvTbzwiLFer7QqWQVPWgWSO/hZxNQ4mfpJI/USFoo+EXjhy7WbGKypjGc7I9vOyRT01F1kzXU49Dim1wRB87fSbc1pDPkzFAz9g/VjXPgx8EFT+zshB92EzY5key2PP5m2ioAKa6qsAH0HPQCBBM+JoVmcmsRnAE4YtObUgAYBGrb9SNqdbvvM+OOcsFGqSdz5/x6xnlZFO7pfBtSHyJoRn5qkhOSpEs9IX79n3IMmQgNwJiqkh49WjwKsRkL1fjxmpNm21jIg+mu7DFrR8SItMH0GQIovt3On2lY/tJ6zZyQP9r6k3vDvkUfFmRxXjELY4Utw/kLe9AV/JSvDSZbmF+oJpoFhMz3ZqhPp7xU/1sxbaVbeNLZZEAXXXNH7Bk/KGafCl74sTtcUcboOxXhstuNKbGK0mgC+TQRTjBvED/o98Lc005T9i9HprLRf3kZK3X9KMG/TjPkoSX/8Y92Fqda5LlxMvFrbs1S4UvOS9yKCG2tNKW3x/A5FB/60xnfjO31s3gLFP3gDmZtOthwht32tu0fO4JAHdjwpQ1fgE6z/WUX+RNxv3SosvhheGizqMXE6dIx67tKaPBvHkFiHlfHNymEUxthYi+rK+jtsI4ueSPkZpLREKaheChLCLTCB/tIexyzx0v4S/b5edyPJd+CSXP5/+oTAFnFrxVmkrUs0EHaqzoMZqE4Bkv6A4LamQUTQVdQNPyxq2wcuKWy1FTIg8D9osm9SMQECn8hKQIiIdrcKVouaHNsFMwaLQFxJRXLOVoHJUDa1+o3lqH8aQeFji60ZkS5cMdZXTSRYPdjnKmqVmCsrb1ghUH9SjANPoYktPjVa4eb7cCaFpXINYHsoTUc9XclwOA+XRn6TctNROUipPxIKHYCuY8JbNjfvczchguPsjh7o7tpo3QQuXoqJuS4dqxekuf3AyOXMVyYtPrxJk1I6NAm4S4CEUoJsQXce1Q2SYmZizFXSz85E7uNoJSTjLn8TJXVchUjHzyrOANJpCAesfjNxhAqH6NsTBnU4GrGkmn7+1V/kj3puH7WLlgpTAFzsq+hbi/CgCAAaPZoTZ7t9lTn0+aR92tDQ8X7mI0kiHWhUQeVi1to66MSXhK5K9yJs9qlHP8PBueHijFcRGIp4sUYu3jUXKaYrpAHew4/l3sogDrW+y2Q/FoC/HfV4Ox0o0rz+4gD1yvwoE7WHI1rvpsyK8VpFBE1UsAaZJ6sPi/mrvqFV5hIdsjD0tXdJkE4/BIypusiAlGepnruM/jQipl5WNh2OoMbYgEQlVqFMeNlL5yn854JuP7rC1afeOx7xRABJ41Wz6YrhatnOkh+Q6AnRUWGVR+KI079lvWY/8bX8X1HHTvLUEiwXAMtAYNkyGPXqwu2/tItBhxocyEOe1pUT4gDYgUN3rSaSAipbt9y8wN/mEoSmya+u7Zbpf1KOdKFTI24WS5UyxQSHlKvr9euC9jyD2DOaGUEDgRvS5NwqkSG9LuRlI/vqbJIUovNnSQJCJOtE0IOBfdI3o01cPAM7Dp9Btp4UiLuTJQ+Vzq/MNBp/qaZuC2elt6oA9H8YyulOVvp6S2GbM8QlFQZVpEepsx7kOuEXUXBOkAIhVeS89JZsoslBJugvZnXTrXX7SIx3WR2j63IESit1cPc5HQ4nsxoI66GqZ7vgqi1v1D35u3LLTp07+6L1Py/yrZqnslD3Yl6EkBngyPXvSUbpS1YzbBZdbEn0fMI6T1xBvr+Fjf9mzXqbwRJPBL0dFaP4krA/VxT0fJn1eh96M510SJ8gdydY4VISd0HEM8WvGG3mHz9X3KcyudErjKUtzC7T25y4jb4ojPcR0/133oVVhvPNM7/d5pPlgYRg1lmtvNpkkM1INnlhFNiLD2KxB1PCM4j1UP8WP7a09QL4/VxPZjEif8AiM4/u3dRuBTqhBwf36A7nzMbbu5UgjqT4gOO27HvkGy84WCfaiwekeqcUtDWqAkeHq1jtbb0KDSw78M+YacwaRCQRMn3YG3DErVoocozX06hFIcQgNvJhVW/JMmN7tc0/+KA0snRLfTmaXGjNECPGOF0It1q+nprgVYI0rv+75M0dLn7tbcbLbtbB6JsFGLv+j2Twslh9SWGvdFkgVSIB6hOAVOF6RJ7hhYSBGu74Pa8AJozaQIOv2jDf3bJ0dA325Nh1/uyBMqb6nfHvZr6OgrFeDNYRCzEUvnDgpNc8JzNbYKssHJQOqYmLiJeqkzsi+MiYC5HLglJpNXhUbt/xJr697TOkpqY2rfBVUnqD/JokmDjpLR0ipm5/9opQZAfnCx1SqkZ5K2fchTsKZU2I4GBaQ9Po0udPkdTKFqRzOqUpI58py+GPT/ZJ9PtUyslWAFiRlO3/K6EkImmFmY2m7Y0x3R+vbyjpuRFjltCeeGSDyTkWp9m9VqyBLNpOJJa5etz6GAZiAqO2DqyrXZSzKYYC6QzrzU0Rl2SdBlmJxKKANicQ9XRfH4XHO7XBNNo12DdbYh+ygVVbNVU7JvSmN+EFRFxYDISx7C4FtAJ9VnqnEg+RN8fq1pvpoB+hJPXnfN9Lnh40A+dX4dAxQWfNo5SgT/yZBGVMKW6RNgvZj+Rg7I3rArl1hB2bx70C8AXc1qopqntS2ZSCmSTyFRimhuMyLvTYamxTnRMGwT7KglWOixdACCtKZoErpnK3jm3zaWFgVNOnPKwBFFCHp2EJmGcav7HNZv7lzyYC/dvu1qYr+SuoS40ZqBSziFWVLI9i8r7dO51/Emy+eeM1+MLoVetyoWbUscmy2/1RXSoYxGQOlQowBr+Lnm1dxSnYmV/gUgxDAp3+0HNe+XQT3jyGcoY7wZ0fDG3ufdyvW9TntXh8K+TWdRxckHE9dLzOPkVY/4A+ifMpUvPmG0V584X7mfRQMr8B661UCWbk9++dbx4qtmXfH50VhLFyPFkOYTXh6ybpBlju47qnEctzHkDWP0Hnn/rEl+05AH/+FHtR3L+GdmpiR6xapbL/qDOOeiSfNMnYCFgcmiwoY//rr8KUhGIJi9TDlEZvZSTupdZb1Q9OtFcPePQ01RkVlSjKN+aiYRXDnAhkyYxMQ1iltdxHW0h31AdNC7kWXhvO7bn7BjDOBuAajg8O9LM95830XsDeACgYswg6NegMxtjLwlgJIN5DxoxAi2kMX7avLc9GxREly2xcVIrii9xq1YFzD+2EYo06FewGl3sr4X87gPJfEd6XM5cYAjXRh1KYTTIpss4K3ZvRknYkAkdI6gy6VdY2TLXLFIlH37vxVHY8oZyee23Wx0n49yK9wnjFLzDKu2GVMtFTmUtU4sBf5SJtmaH93DZ73era5z/e0zdhlc5w2VsbuIy1SQsk2ewww4atLZcaL9mk1V+BrnXkV9tPBJn9c7igKIy9y41b5a9GgyDrWmtK7z3hLjSOS08n6FSR2UX2oyQv6k2jYElR9to9qfbMJFuwTHtthCIWnAUjG+THNv//N+JqRAiP8TILlJ4gX8WG73mlUJjXEiMLUQnOzcisyCjdHiM1+R5rSrLkj5hxeI7nZy33CpAbuaSMmCemFSndcWyEx1r8JdMNrhR7IvIW/NgeMthVWNz5zDJbMTcK5bmdIs0CpQgdIPSC+Ie4dUrtZBZ6eRYETbKb6KXr0quCx0269WW7Tlm0TbOqXTcviCG+89g3yKd5dDHcBhnD74jZ2SkkvUPDeMpLI2MyLpbyJDdo4lbM/e11Phk+fIafaqSoFO1dtVvpYet8uyetu1R8t7wnkN+kVw1EBCPSbbF/hxgEITtGorr1/hfudJO1vjxkQ27OwptROjPitY0sfcamwm3+cVtpplarYvCpPWI502k/GgnSlfLodDLgBKXmKnUUE6/ZXog5pONJ1EBbunde6+7IXoSLEAFnmKfiVrouqrHu12lgHlOuiuCGRgv6u7Hs8FK1JoZvGHiMevFlSQjwarAYgSZkb/6yRPC8ypt5kX8yQfHQknpG6h+idPWhVmv5g2WC084ZfiCeedsnKM8qZyvDJG/2eHFFbgCv5jPWdEYjbY0t1TyaE+d0Ct6AKMSnWJw+XP8ha3N74gJE1O1vdAHJMF2S6eSkJIDOYJJ4j3MvbShgzM4RJvZvYxUBfiqAIAhPnK5eucfh8D8eZ5rGQYSBlNJuoC3U1v2AH5DeSgIvJyS0J9hfUM+EUqhzRodvVmqB2NE5uE3lTvwtnmjvPnl3Rx1CMNQPDtxwkFmA+wSGqjLoFwBdjK72TzmDWCtw09Q0+Qq8FLj2IfZa6ii+o8Q7kx1gDrixMMPL07IDfBTm5wFjZ1S1LplyS89KXlecBPAN8j5+gQKwP5oE6Qx5qZk0sN57fmvwrAmAnIKPTp6pgNhIQD3xktYbjxcvPBUTaA0a7BAOruNEqI84y/KAq5uTSuvtRcJs6SgXFm/MsQTjoPcGXFvtlO/6Bl1jVwQYeeGUpTFy+uQQ76nN80MHXix8Akwtx65YKV3cU6n0w/voBSBlQeeqB+bykXq9fk5ANFvxVD6IlR5ImtWuj/i7GFgF6ytbIULsW/IyJTY0GCdul9AP8J19GFJPBdyqA9qz7p4bBJDXPAI7J4jIjj256McyDZXbhwSZapqZ6TLCybY4rmmgTyfaSV1m3DHRwwLdu8ihXAcWKOM4+KpsLF0GlUI996i+NAtPk0ofpNvDUCO7dcFO9ChHPJ+wxD5hEcWz3tKb2dslq52F7cwbbDzNOt+CipS00VIz/ZjXxnBj0pEBXxYz9hWTiilorkpq6u5BWx+IBjXr155AG1FxEyNBqjCM+IRquamBL8DrCh9fSYp53K+XGdRhYeoHSG/ELFqJERMoePLByAkhsJBr/qOE9RKCuf/MzYUo4XI0uraSM5K+QebcBTGkwuX6mQs9UmpcgTIXRKF2FFSw+jsCtRR9Sk6CyTY0EdSG93EX5/CwPwnmK23iY+71gdvOnveJqyu4OSZtfFcfBNp49s3rLGL8VdM0L71NJnRLZGQCCZVISKUCMjtRcYmmuGcUQSuGImPzYpHvYFa1bk3L0KKGDBpG13CjnGQ00/p4zgM/pkmrW3oYcDHGAqzRCRR+hPWvoy/rewAFimDlG8ONHsq1CEEsP3A/CEGoZSX+pW9qNWaG3XrGlkAwHfvOF0KD6aPQdBrkSRDrNMcYq/SEt1aybgv6lkFWCJU6k2lPU8Dm5lk5ZG4CvQmgD5lBoQmhe9f2qkaoEOUClwZrrSX7RGYmRgUtBLpaNjS+Ie5//LJLl9fCCN7lBfo1hIGhNX94X7+8v2Z6mZkqFLbbZ1RN7M+3UH/KIybkd3wO9ulttdbVpYz4Ykz4lDJ/xSeDCadj9nmFmO8Lmc/6ffxxD43VSuuUbLy2R5iu8eDpnjO7Lwx/hWM6Ye9Y1PFJq3MS16b6HfK/HI414LC9Us0BndP+8NDqz+u92SN/aZYimOG8Dxvb7qT94obvWN+4eADk9lq+AbgiRFuVT05Ysgf1PNS1uGREqzypDqp49Mo5M9LEMTUTjKy1XKl0Tm7vwJLEq9VLr0i20ebrb1urd9lMSvix2+MsSzVqOdG8dhxBN2eKdeTS25OuGlD99xyEr+yVUGm/ZWJ8/VT88J4PG8MXv0LQiDGu9rS53EulVEf4/W3FS/HLCCmrW6nvFLzTMSXfyIDsL4oCxe7Sz3A9m2r1YlBOyd4aVY71t/BIjBWwHCtOrENXIh2r/bN3z+X21sYBw4/h+E43CJXnsUHULBbIb+A1KuhA41Rk6rFFfgy7gkUvUSbmCSjFHqkuvbt/P+VPsTAIPRha0y0AiDVtUqV7dkTCybLVSDJoMUT4D/2WmBYZD2RTFV0Mpe/rucn/OeETlRcdlP4NZrm3eE241ssT4X02XMQnE27j16UcwmWqBr1YayzFhuYFBG7wBTiOdE6U25zdySYOPNA+/yQ3mi6wBIRSGT8hL5hFCPkQ+0/cai/BccA4bvJDIOqOfmeNCaUq+Nyo+9aLH+IqdUmBod99snTRUjwLgLCM3YIsSE2jg9cxFJgeQR14ZdpikYipaCdGcLw8tLHRRISo2m5OBlfXN6+FkKeEvAncOo6BqN/XG9mexkCJli+X8++W/kYpObveGh1hVM2NFPHdKOY/4poWT2/TVyo3WDCs0UbfSw3XYdv3KJYQSRGuAki+1SFD0mynabugbLCuMquXNsmhXyD7gakFZ2L00Ld9+kEQbNVDeqn3zyIu2AT227odBaSW6TcgoALrpzM/t50/FUNbWkLmQGMFz6ZxT2qj6s9ZIUJ1euUAtikpHBH1xLk2rGWqhX368gUBrNrPRaGViLK5KH/E1SdklGBn4R6f8gGXt6ZdoR4vXN+Q/BmRIbVaUiOEAZMOOQmCj471nYy+EfZ68Ha7WPLuW66UGrgRuq/VgDvkqOWYHXWQP23SQRbGsE/twHccqrWveIxqhXte7RN1OoWhhTz6Gax5n5wMXCqm4sC4HPUROjTa29LdbNT3rpoiKR0l0m9ZXEyofFRZfa4dK9K4smMVCWabG1V5ccdWXffhP9XjKAHoQxQOdTIwkoSlpKfRLE//ApcEyN0AAzIbwTDCZqnkGSNKeJVxtQK9yVT49bDKOTe2WxB0EVIP4mr5BPtuNldAT0Bsh+c029P8IK5mHqK/6QBT6z3gmkEPACoSdZtEyXoWFoay/jx0vtbMA6s8ljWob0Mjpk/QpMDpWuf7DwOFG3iXfOjUNJrdMFRYz7BGNRjF1yuiwGJO1zokasTuwWyqEHIOpS45I8eTdhywl2VJDerlBNXHQmnlc53B06ZCCNlESEZ67yGeT1YCVpOF/TYPlBX0iV9yZ+tcuImY/9Mb8d1iw7zEZl/eTNSL418NipZem9+2XLGA1nr8pp6XKl8Zcz0ytEIideiCORFIwDLeozmq93lSyA3dJoROJyw1HpTNhdo0Je6rqPhG8cmblw833zzEy/498lWQ47pjA6Ujx16okVgDMy6mp/zKVyR9SU8ko69j68uYfqwmwzc+nvb43VLH+kKRHiKgjaT86mduI2o5mqNA4Kd4loZjht2bbfr8KygPN0wNxBaCShdljGFi8gJ+UNG7BYhK3XFAdzSoCdtf4sUkmynKrj8S8WWzVjpbg+BVnce0U8Ir23ksr98dT1PjklSqX2l8zWDAq6IsDvDbLA2e2v6kYcY7CH1URdGBR4AgDJFS3llFUkTMRJSRAOxtp5r7LtZEOJNjYcuiA/p6Fo5Z5Pogizggffs1h7KfDfCsaYuczcvMurE63pVJ5L1k4e6s3ygoJK8TjnwCQzR8KffYjbjyre9dQqHbOsMV13ooXbyrE+O+iL4pNz2LXnrrxrwDKtgHCzLv1t7Foq5G1LmL0S4Uyx//UmInNowbvdEavkuaKLwcEut6YLqiz8PgD07obvP5HgpS914SrY8BEYRBzRqvux9adT/YNjinJmNPAUygJpd9mpdvabSKHHgtJFJwNVVpNQzn82+naDyf76hZgdDjQH//1gaNA0/M+7Ii3v61hgonF9PYWF4etYj5bdfA4Rv+4EHoXJSioGqbr1KCuJzEE0T2CN3vgH0A1D8byKgGjep5bDVhAqwtENyJoKKb91HtMb+pAPSqFEQyTuHZv56kQxSvh5FKCgw0Ihke0i/8a/YjS9OzvH10weFSFcF9eRryktI4qakxoeumewpHfWOfvbKUmaN7buYzjhUC39VZwVzrYiWA/BRnStvKinZ//WqTVAPU73FjWan3MyDSEIM0V7VXKM7qWkemOOewj5zo1UAAW9n3KNqlCUzFHz4X+QHrvyRLQ1K6rzh3IGvyjgrYZ6hHj063A8iWlVqKnMmyd4gLA2a/B3KS/TlqAO0ku61BQs+Rj6W712WRqZIVrPFvqNeKVqXCUUvl8bYDLtYphu/josP6t60MdETmdZOMagyu0bnrnkqZ+8iq0jeyU1xfIui46weqHhbfiJqaurXhDLCJtnQe9GiQR5GfCraZt6F8zynjnUoMvDNhA472MAwvlBXRmMwCNKpDWBtOn8MjRCZOjOIX7L7ljPlS9+tGLhp1cg5JIyJa6Ywr6zaAfJk1SSqhnOifwJ38W7GuxgME9Xd91U+MbswNh3n9d8ZAURAOdCfb7b+Y/aPjV8wrzJlxR1+GrwRm2rdI5UBowJSNyAYxqVJFDZwNmy2s/wXi8+ZnfSsDhJG843JhJxdVsatpGqR0JgA1Hk6xQ9VpQjOubJwtqmW0p3U1j8j43pluCJo6XCxQe8UWhCeOBmj7Cy3paR7hYutAHrwn9Tw7JKtVCg4X/06H8p4YFjJtqnx7v83Rcp8Rugb7o7jX7XDMMbRSkRHA2lqFFv7f01Dvai6dQFP3vMfDjzLlm/vOOECuzAXszPAs41PBseMoy+75T0ycZaoNYo0u3lWBrx23+JkiDdKqWTEvTGsm+4LdPDKc4fQz3TxJnBs2yT8OO5qfCe5/PsdTgzIBn3cowAXvQ7pNx5+Z+y17CPqCIBTLlz3NgJ7BXg0xHKvBNFveLnO8qXX9rPIZJxLVFYoxTNSjv/mEkEUsKz4vIAO6sy1QqOwIYTJWAHuEQ2la59wePcRyYclazDCezHZzE3IA8HU4yPlKR6ATWUH++Dq1/lPAeLsRw826T6EIwAnUJl1a3bEbfGEY3Mu2Ubr8a0jViIfv8ZVVPJVrPal4wXi7qm/cG5FUfVUdhR3SJ0W2BfOgzKemzPrpMB/Tq2dIYmR6lmyCQbQw1caSjEI+AFtQgLwjsX4kAIBQyZVu7O3GmCHnThXtHf0PNnHDklXdW6E5Fqpn1or68nv4pP7mICGiCREdn8aMwJh9vgfeYk+FIO3NmgCHxgC3l3ehSXvk9qr6wGLpM9FntO7wgrrDhq6RDjx5WdUvtXE7F6Eeqdlzg5qcgUG/W6t76xuX/WIfbA7M6SUJ5ZYw/8s2R7F7JWZ22wVO6PqyJawIiav6xNKI3CCfeA3MCzvzFe23GoJJQKJRoWc3PAFw9RYhwGpFN8q9cgR8CBbF9/69RN7VHVl6AuSinc5PTzkG+2Ym1HErR0hNov8IcghPd29ZdW0O0jf5kLqD2aPEqs6U0YB6WTMZio9L6QUKVBrWgMmEFAKE8gD8d1OG1SkmDGiyP8KCzMdAPx+SrgiKOgBk58Ay2ukefcIPoLGVSZ5DIlBmN2TBdSoSSk7gI6cYADtxaJuk3ESO4pIJ6dOMm/pVAy0lm6/kqyuLxrA+8VcDCd/Fa5CKa/c44LgkBsPnHi5x+MAmTH6Wm2/0wolNJzsJrR3VOfqrhM6q49WOahodA6q3Z9r/BGMw3p58YdjpLECCp7TGLhP7oEsn234zIXasUjj3vk8xgZEjMFWWbT05bzhZKiYQiHLzrewq8hDlzclruDmnH7wY2AN+3QA3iv40OFAblKbjWE7HBhJxiFesocFn2T2+gcewhGAzC/IhKetS42EdBh+uk9Ul20zp/JDIKO8JY6wU4XxBvmmlMkUGFFuFLVwQN7dJB1m3xGel1w1WDf8qfnkkxlhcFeflnC5S7NZWTZOcbeRoW2W7bOXfBmNcxG4yACY6GaYkCCOZAuDZ53ocZfleFPP3CwBiNn/Y1rV6WMJ+dTMKvwGvCAHYs2bFtxcjRL7jkeq8jo23ucnbqH+011gfjKarZUXAAG2rCjKq/DL4swr6FSuitjqUwA10VRil1SaDEy/1upR7x7CvJRuFyz316w6fWmZ92FNb7j+zdpmtgvsnLthveCzDOG9vwNbd6746RhNLmNImxnRaAhnffgW/9j/V/4O4nL0yQ+cheM+858pPi0HQEj31gPP09HTAm4g4azqBZrg+3TeobUEPvFoswxrVMe4cCCWaVxt8xkbSSCPQYcOUkK7YKlN1PaWaIh6eP7E8ZnqjjXrdb/Bhy5Qx4fZVWN45Ppv2S2GxKvSx8IjTFs+/WPOmsA3HvrQE6u6LsiwGyMXscjEQE1P2sWl29+7VUAq/KtSEM1ingo1atXlxShpjXkxbEwcmK13XiqcJ+ycrHUcuTzvBG8SgKGINEs+2O8Q1M397gQ/+EEu16oPkKABF6XYBLAKVMSZhQbD4jeVtBfU4mAhvgvWRWYDl+Dr9jAWxPQ3cgQHbQT34KzkNEngRvhJvBEKvyX4YTFqpJ8EOXrBQhn7ll3z1o/upvJ13a/rEqVBKGmV/YWzE7bDXvQu4pUHDwUt7roSXKCWNGPechJlWpYxyclDzlaWMpNXSUcKbhoV3WaxkOwT/WFLjLir5n4jrn/cdAM8uST4Gs/+wIPVhFFtxZLLLPK23x3gkc0PQ5agtJt6kOXpEw8UiPhpCutRbQOpCj9Z/1lWA0xwafADJ066SCWvpWbpYrmBcO9dOLAudY/J9iLKzN8S6ttgTRjfqLdqGYaIy6nVnjNgAPCAhDqP3ULLRnL2W51TE6vd7a4PSYgQmdQ5mA7KnFDKuTIXO5BG44RU4KcstUAdlJFb3cDjwRhukHAVk0GnHWQLZg/saEAZE5zrF6dXUjFCic4Z/k19D53Ui1ZqNuQaGb/HT4/2U52MGEYB7Hdss0tD0Wb7gcRXuJZrnH1DNGuRLmWWzvHoW/t2OmMyGPnJZ5deLpG92/3KL+iuOezb0ftv8B5clki7Crgc6QV5YB6m3pP+knRA8e6KFiXktBSCc5LnjAmY+RhOXOiSZizb7tzUcfblY0qWVECTLlGbvI+L8s4hBfU4CzhYlXmA4zMZBubqwPiF29rEUSmfnC5nB1oT7NKLfJMKfg50XleDg4U/+yv3YULnjlu44Se4kZ11X1932PgEnlxrdg1rKyBLl37sZWLvVcW4HwP6tejqNEfFrKwz73d0WKtyYsjHQZfeKPGu3gbObVGGeInO+1L7cTRjfveGX1H/ww2IN52I/sH8LfU20lQ1tI34eUhxeKxqS450L2SDi28WOA3jWUH06NSxP4vPiHfjqCKjSD752TF+yQ7QwevwjPYCU38lu78IIpUUi33hKOdpbY9sbUEx8kjd6K9Iukq0X/Z1fJ4TSX9hYaiWTlo7W3+wZTx0GhEOs/j3ZyxGzOonoWp5PVqi8QW835LxjZchefZ+7FJOBL65zJ1tOiyXNjJn1ibIO/jPHz0a6MljtVj1bXcxiDo+BqWErqlxzrOa4kDZeo3/sl7vBZYAP74ddBIpc9/Qnbl5gLpTFSANMXm9yVwLCic6BZf/Soich1LyqgRNSGG+JIgZHNLRscLVilZsbfaHPMGJPs2iB8RCtoEk6Wn/l4t21l/CanEhByeXk0ePATHfRnjJV2NS5xyNbGBYtF+MOk0M6SQ0HOhcqLH/gucFkWdTbrIP1hsr7KtCWc/d4KbsKXvQLVJAaeS7NHdPKgytUzdy6qwFWswopIoBRvmmg3lw+9uTJuIQdihAg8NhJycroKGggXCfVlmU7g4bdVF8fWZeTdN+0nzZQjLcLpLa1bToTUErwwxbgPFv8UC/ySLawksHtAnvDxe6C39yXSNdIHaR9VzFsGBOtKZapFXUdTCTrjgV10xt6XgJuB1kLvuGu2ucA9pRFk8HgryVuRS7yyLBpKUr+ymI2bg59UdcnPgYbfsCPo0Fg/Ob1evKypKHkrnu99WSnAGM4gXh1Wv/AoCwJnJRITLnkdviG/gKN8TMboEMawdaLORUQQw5y/5HgngNLfeevPoE+IFxTvLvhOmfwIESxSdHGoHs6/1tIWT5lBEX/kl1WoX/5UHMBU+av90BpabGE5CamZR8rQOoqsKaSgy53Wmm6n2AVcmabusAc4a2AZl6Y4bKzuy5jXzZ2lML/GprEgxzQm02/cVJV7YFLOfyClyj5u1zT3B+8bXwda1qKnCy0X2VdCc8yCwJEgJi4ORY3oxGEPdeha4Rtd+NevrXvdGdJznWkEIVx/SGRIrxXoHQ4lXZVwYaiRWc7xv5/AdBLyhRF9TX1fMcCyRAjcJI69Qy/V09QBN2sLMFrruhcS95NTeSVcAk7td261j/s4qwRZCf+DLYXVhn5oP3QJYihjxqdStH2daFlqZGWzzoaRKTpCEWq1bhchFIESwZH04xs/yshrCFC4yCSEBDuFM9xTdLZ1PRZPQ8ILx1rhPYk19zA3G1aUBce0BRiOmpM2Yc7jETXzt0gShuDRjhflryNESHIkPXLiJ+6k4RPNPs701zoAqNaDOgRjbwzRnV2K/Wl8hRxp+nlsn8b3eYkefpolNTKbS2/hKEGv37lozVffLIrUakfioANJz3moaeSECBpsYdR8w/T/UITk3y4iXw1OwgG2Q0R6ui/Szdn1isoZZRew8Y4b/HGpHSN6jRUdptM8nxaAcySzSahdaTEB6aC98g7Rwl4hRYLV+KoY/7x+uVE1L7KTxGOu0qQGnFuxc6crO+fpMwAzDTcnuaJAI7PDbIgD5JLywIjE+XLhZoFXPJiNxaVByU9JoQNXqLNYJ1bGs4fI/wm+Fa8HYzhWYxcws6RC8h4Yk937HtKDKMbJhRyahAFFiQ+f1NHVVFBRIw50o4WshUX50LCTZ/6nlWNDdvYUjFt+kTpOk9mE/UUyXFl2NBYiDwRZtKchnClLT/ISCxDlgt48jLR6WA6pdf9iMO4bINnKp7mJ4h6BwJFBNfEqja1M9z+9yU1ItQKSFAVmQyu571Jj4/23OKg31hm7HfBc7oF5CIX91oKcQxB+lzlVVYRgzzur+jDfzYCsMUkKsXLaW4yEBKiTUhKaHEqTgW+d4lXUS147dgQ0m2U86VDQfHjt5cIar0CBUCgWdbCrwbGU64OQuGjNzibozYRk+fpqhtsJevZ0ggzddhrmCJyhYgOBEuyf66EYxLyZnCQz3zLw8fkWIt5KjjjypJ0QbsM5tHJfR+DVak+3PbDpjQqVlBbINt45Rs6fwWb20cvrt69prj4g9APtUQgCyPyGFwplNFMyIpbKR1SSSeVrAfbwTTTjJ8pdmFAHK0AG883nBGeNmsmTNAMQe4E4QQvmLnZeVvobzwZzrRL8uUvGmRKZxWw/iBKHa6+9WLTOiY1jrihJIKFz4ZX0ygP84YlbTqBZ6c0raH/lmuVf9ccgdv44tvckyKQaNkXdTRtLn+SFvXu2Pm2kyZmV4lJIvt1a815QFy8njvXSOnjd3eDEAJQqOjV2gkZx2Hm/ne0roG0Uo6xK4bTA5FA9aKwMZMmtzcxaU2b14FmHnnYd/pME5cf4IJ0FuTlHEP7m6LfoHs3H26rsBhEOdBRRMXIkEaqKyqu/kyLT8SNoK6ZprS6nwwwxwpqpaDKj8BbYUmDJh7TlBo8ioXPwXdyb2ZmAM43WE1caoO7Q/N38s0VVncar0SuNDs800YAjntplLZ7bOtUkLUPwWU6pKbdrrv+gGeJ+K9ouhXichMdyanuI15OZt/TpT7Nk/8wvJbWOiDd3aV0+pl5gZ7C4bHgmfTiIQOzSAj4iyA+UFICwe1JTzvzvHev6Sib+8Mtm4mjy0MYDzWM075YUg3w6r/V4a6KEwsCIwLGiI2ALNfw5svLo2XwBvxTB0G8zYIegV8rEf/4GLk3A/jgyxVOCpvqUZAKG/yKcgIZlebcPJm0RLNhZ9uOR2+dQ9SqAAAebWJMuT/APavHKa+d6kt+y/AUAlNIJYb4raEee83qKRnkazFU3/ZC2ZFgklokKacQbrB83/So5i6G0coR51iq3T8mm1dJ7/xfwyzojJUgEMAju+z1MdW/IYznpHZH5DJn+sRb8UqeGObYryayZgjpR7/3xQuQiZbQZJG8IPoxSKfiwDM4EZ7x2/4QutWSX6brmiVF8nJyoKVi3zEKGUttWybTvZ/sU4V/kXm0s8VXSiwcKjOnRUWLWubBFhiKbk79PORYp1eYPXjRqUsKXReZT3InNqGPOD2Kp3GDVUW8PPvb1mt/5WxhAzyZ2MOmO9773OBHTnnQDesuOJuSzbOOZ4kuxYkZaLfwQaWqXxNl2A5xbE2Yd+hWr342uOD0pQuIJmCuZ/OH+M5oT2EZ7SnGpkwgcj/KaJ6hTcyHRjMjD+A7PXZlvCxj94Lcpj9sBqkRsSCeX3HdECopvhLnSWGZKGU/jTSJrk2OOcE8nb8TDeRk3+BGR5W63Py0TFgWnmQtnNpjo0oOAAljC0YAgD9r/6OQefYPaXV19yewM6Fcsckh1Bd7c+RLJtdjZhDngSAQfIeEVfvwwfhGe3G0Ub//rTiuNaIZpjpW2zUwg8JxNRdayFCEB6yJOLhGyWJjuG3tYaAv8nfgwvL7Jucm2teQQ+ghiB1tKBnLuRL4ywyk9MgF6if5ByQneEJihfKY1Tt4oV3MAwPdShmXfZDKDoTpPbdb6WPsn4uyZ1LYk8spuMyEMcNzt36w2KPkyQPKWNXXEpnMODfZ6EUrNBZhyCa0vPEbitYG7VyWssCyvWpqD96uCLTyBmO2Q6NfcbPhIDsRfuvx+BSk75v+Cmrs33Jj2IoEvBF19LqsLCm83Lmetbk/OJNcgnm/NdZC0DlBLkEbe2Ryo1zupOQMj+h2pd6pq/uVOkRvNa9h8jsBb8/0hip6Sdbnave/sxvwAeELyNtYbVWkdM3Le93UeuZ03DetsE4vchLFr9B0Chrs3ysBt8vMxs4JaDw3+XeoLSz902jAIuh4uZ+evoSb9njwUSysKCKcnlibez9FRxkI+VGdzaq/KpwkKmjeqZ/mhibZNe0DldZYSSMCqAL8uYFqJCdJyp05D2bM+y30kZOP1bgTyBCFyATaHgF1mlZK+gjUy7OmjUboD2Tj+tcWs0OeT5jHgYY6few5K7QXv7bkKs+RCd4g1EwEfCYIdayhiycAmHVn6ZwW75h22JqW8/jfH0pgqrNiEo0UAU6lbZ8mgTKVmaM4qCi0Ji1I6ujThwBfIbtr3nSqfj5WcuF06ZkfM39EcAxJGYmmbFRtJKPFiMJZAk7xMnsWf4lkrHrfgFTGxjQoJJdVn/n+g4JDbx4p3cdg5rCvI2XNbDT3RiG+yT5vw8+Z4LXDqd7UGP5m9zzPwmYYsqveH7VkhNnIr2PYsCLh985/P8lGQRKw0RBw3IXJ90LKc7Uyi8pwPiPJHXYSgsZtPARLo/1gLiYoL+yf0LQhdBEoDg2kHIUnVX3XARjfrly1WknsoB5FMWvGxL8Ah7yZ0eg4IiEwezuNKENoaqpcnfO8qNhbVVg8Luy7rl3fg/j6z7nbXvY3jAkXaoCDz9qoz2oWYmnHf/rzGHOQsNkWCJUREpMrJGb2WxFMr81hABFDB1pScGM/ZPAF7x29FSpBwcFy6ahh7mPpxM3O9951rvdbH3dVGwLxsh3HVA4ECZEcXKsfmoihh/uq1GLo0QrgrDxaulQfF7x84p1D5J5nBEDjsZODdGZfjQO5shi0ssUTJEAYOZS6IYjhwGXqEuYZTphdaCXLGShpdxnTdPNmIIsqZWbaWDwOD6QVpG+p01eNC1p+srjY+rB1OrpbglLDIwUEy8hZhRPyeEVbofWXaIRvKdRGWEwH9zqqMFXUWAn3PBT8GUVWVxTwlzbK7O/RMeoQZFeuGj1jcn9V+wy5RbwDdUEqXdnOqVfQnkNg5qVCKNzqoaB/2rz47+RoSiXHEW/u8X4NQYbQvCdhflTkdZ3BlggennZv9O0+edGCiO8WFvLtQgK6Ko+hgUZRNZOHNoD5tLS1i2xbJr9S2VGegPsgCfaVxiArWTiFYJH3F/xdNO6qEcDSeW+1ErJe8PPdedBhy7kOjiWtsZndRXLXYUQepBijXAp5PfQmnrVprRCKSuAa1QN7cAi9Q4t3U79I5YzvRE/XJQS6gHpWT6L8ak2Vkrqsd6pJQ/+n3UhIKGYDN0mz6ZjQkxgYCPhWOyUPq0XwKN7zQTYHZN7fUa9WzSA+WKtEmgu1UnYMa4UF78B/bPzRflf1doOE61GuNd2dW+jcEzKBLomWmF5BaiVRrWrK6NSGuBnefVoruXVmJu9L1bj73BjyI3f3NWrpa65G4S1ylIPJJbFfuShF970h9Eu7FDWTXgWbzW9UbaMiOQd+ZOHQq9Lu7fswFnnd6beWFg6YLNMl3y9O4t1ZiAdbJw58ihqt0QLLpe+B5fSF+ZNsHeIJfyC8/lJy8CzZLEo4XMUzDLFPWvRvB7D4YN6nHXtiMTJjdm04zhq5nRHgZjN1xiU8kGtRA9b2fc/IuC9U4JTTAFaIn1x8xTb9A6111llRRBObf+SxkJRvY5BAubWrWz5YHFrHP7x5Ow4j4mZKvbFpplrMn6iSW9hIicRXBNrXAltwwSQa7faD+Dr/VZz+5hhyWyiPGK0GiJ22XPZwB4rjxSbX+NSVDareyAZ/B2HiQNUnNhWTRSbwNh/iZRMcrUV8wrH0bkeuD5wv6FYTYTpO2HAmTPGiuhJlk42+9X7naezcmF7Sz7IzPyqz+jcTdtSrG/qdQ4mZgjIRO8gKmSHB2wa4ofwTvfwBKwWgUM1HUqLGPtwRE1g1If+jDGcAclSKyd89ltu9zuJ0nLd0arPWJrqiKQ55qvHK1mR1jP5sl5UesdziHhrraq1jacv25XYcIMwBJPgVMsXO2pcOIEU+YMsf/SbGfPiwRCz+rHXOHbNi+cr//GB9/qUR8Og8eSFRBrzbTSKyQNjeoFPr5bEchoXY2M6kCqpNsX4wn9BZ0GNdi7gN1zNA0ZgEoXrR5pk6OWjWJBuzewX+XfAix5At55pkGwcV+KdzeMsTK5i+SYt/aTC4TzMpotbVJ8l/WGn52ccP2sUmzj2kpg1i0gRK/xUK5VPmLl26auNFGL+1s54ysslwWz/W1sSGVOGKg1PALI9i73xAWeU5ixwLVzWz8/6R7YN7K+PTdoOV32Z4lJWnpP/g6S9xB6vThZNmrsCWTMwRnyJ5chUBpvS7DZPlqxvoifW/1C8a9JCfqoK+w7f7GrcdwrjXm+PFvJUmvfl729BSslFEJVmsk6yLHaL8tmf4C5MoDACggoqUBixsDmRsabzXTVgtm15TZYwBNOyO3TyWOTVU5LlU48Pj5nF/Q5paeLYMPHZnKJ5qgIPqcPO6p3JMjyhFwZzKSASVY6NaOff68FJad6A6jSyllXhTTzY5A8AAkPZfSTzTxLbbcfTU/usVth00wvmHgS4CnM30mD4TYNAlBfWFP5QxwZdoept/ZPc+AL02462YrI0YYTbIyHui+bChTMaHchRouHbp1k6tc+FOsoYII0RWAJ4owHfig46S78pUUhMBxHxdu7ue2TJIG9zBAi03F+ztEwM14FWzUnlefjqoCLEoZWEa4+nZfjp7nkhEr/q40r/lCa0+DNDK3BUBCHlNzFl96a7WrrNiqssLHfbGXb4ya4cho9+9htgkz/rkflWoxppNPYUZ6M+MXKBoBE5D1s+KA6kTAbZ+QSheqjQfu0rJ8aB4HftOG5bJTK8fuf6garXzdYf+zzN5/3ccj9Ex+p+2IevwynrW8l2TD1Tmy48CO5UbZSwZXi/OdPFhJgitIsndxLyf6X9J7MrLpjkFJeiCpLYL0sUixytsH2iX0tiOtSaKXjYc3DYNVofHTRfczkFnLSzzB1tXXQhTBBONeS/V1o9kUqJn0XA+QR9VEakCyhG7xYt4jciB/5qHl//dKSAefMbb1S3L24PdP8Lgd6DK2ZpbZ5c/QZ6azi7t7EtudalsRA6KzTAZyn8SmS9X9Uu83Sd8BTnnHopFUtcqCaanVQ51zsGzmFPtVaeH1AlZ5GQ08O56BHKvM6BDxUjkovBvey4Fn3HDo7LjOzOWqkpFfS3wrBPfCe8je3i+CgKfpVNCbYehhepD9bqcxDuiPnHnJjXjGhFTbVHkLGfo89OBAz6POH9v61nR/t++M/JsRHXCj+dT+0en4xBPTJg355A9gBA6kUv97YYQErObYVMUlqk3x0DEifBd6YkH7pGjhjDt/kFKPtITRSgn1OJ4GGjS6e3pkr3xhJb2GPJht7dKqwxecrJwl8Vd4QMeD9rbl+Pn3fSNN+MXfFrEnzP/jhQj2OAtcuBPpEUyagTZr6WgoxgVjAPQQiUQjb25/40IttnVdVjgJTVNFp1ES0jJDbwjrOaLEQn0I8tEjTXNhTJ4ssEINfckZNKvCxM1s82q5VehNYs0w9zY0iBYO+6B2Kvz4CHsLTMwzRmexlvjTdXh2ChXH+869NBOpFMahzz84sulvyhpeEyEjEyuw/t5uwnzk9IOXtSmEETE5El74mu/ok1CmtloqXHzZWO4kQpewxRs6SDJaALVGthIw4W9lTrYvmEm0Vrvzc/v8WA7bACE7PfqlghmUSR84kTXHGKhQXuwRpsXGBSa1nsdqnPiv6MYj2dzWCYV+VYtc94vTCjwt2XgkaCi2aSjQPSnKw5LMJIFL1dYfHWFCvlbs2M1ALxx1b2xKKV+KymgBg1mKhUsX1zaHl8hkHO0aowAHv8IF/uwMuxp0+3u3oT2+3qSmTWwnt6LYOKi+MnTWzh5vMUruMp3TjDkcErrOn0is3hNd0cK8W792h/pGvGJcWokMNP/SM2dFqK9Zz08osOFDVJYhZJxgRoCUzEvLrgR2kiRC7K7gJieRwJXxcRgr+P3SU4X4O6S3qO5vzqFx8L4M+SrosQBewgZCwb/wffp/R0p3F2w50ko8PYZk++N8vT5o6Ep0jFAIW/f7FhRpk0oEv9/EFu1pgJn4TLKERLLwKf2NBkSZ34L+sR2DJ8Xs3gkoeH16Uq01VO2UGPTo0kbHgmDHfbU39a7C8I4007dBGFIMQK+F6G2XzFw00Cof8BW1T+/wfTJyIU+qpudar/TBPqIv6CCJltH5ypE0X3klfJVT8YpSIEg+4qsKBDNZQezzHOUxWg4zyVPl/9/9udANfmyJfjCld7c9aMQ2xZ0wFmZPQ6XlYgvhLC+/pk8QgYs2GmKPZXQiWya6EVBIuJYZT4CJQR10bg0DwBr4oTqgZ+dphshICiOf8PafFBfNBczVW/n3lQtjBly0AanRlklkiXWXqtsuT2yaTNX+n4wlM5nubLDVN9UzAR9ZfaVgV8S+ChVPx7hWrJCnVEuYkLSbLeZcS+9LkaESbkZWOuZAU2aS9YRNsvLxdUoVsy7U8tgZQa51WjtG26DUfGaY547QSm4Cc9WpRHeG7Ff0D6SkY2vKuvNHsv0ExWJo6IbB5BEWyfV1dYlxysYyM/HQLEruQxxA4zo4QgJ3mtQq5W/WN8vYfv48RVDL6jZo7zTCe7QGicOK5Zkp0Gk0+X8noH9r54fG2LxxkUqAR92DRV28GM12/cBa+yzJddDncWMlfyVu/a1Sq8PIWg2ahgaArDFIKGNQuHfv/kWrJg8iLhB6N3q7bJbnAv3a9cmpzv7cRjGzXGqBhthVV6rOo7rLHhm6NxdDKo+1XLA5MxbeG4IGtKcbLxKOgXJgxblP6WiMqJ/6fy81Y0j8JSubn4PDLBD3+jJvJ66lXq4TGRiXwyrjWsffSSeHF8zJoWUahuuHEuu4A303hMldjyqeOuScBW2+9WSaz/o11jhPOSqZ3LQb6djANIAQtEy8UqLBKBi8uC8tLb5ARbrAlLW33B2tcLGfdQwBb70OIh3ZzJ/v6DNCIAWmEDsV6PTdsE6v5DZPbXKlSmfcfkO2eabuGeNjOo5zyYc3FIOdQ4Y51BWeLIvI/iqZcMEeWVfbB9hiR28+Z8OdfetqtujuGGFRsNW7QIM39bMcbr4i5fnOdv/p01hKLZe4IoeYGmALuE8tbfsAvCZDJ84nmwr21mCVjH66rczPH8kTwRJYkDXwStbHBtWOZv6cSH6nEINio4gY1gdOmY4l/6IrCmxSvTp9RTO52+P4dACxx4zMfvnt7uajVx/Uo/0tpLD/BHsN1tMAThKUIejycdY3ZU5Q4rozP0NW6Ky0nR3hoGaWvm6P9/O5Kjwbeh32dmk7dPpuTmcNCSV/bJo6DnhE3gEksV4WHYoUo0aPp1UPJU+z1nfToYRZQlgY7awSJoFE0E5hsRlOxxBgaF1R/tt3I+YuwTio52fGFOUrR6MmyyIwYy1gFqtJD0G6O6tOM6oyQ8CpKpqiqd6CUsTauxFieY82+4eHzqvII3YN0lgn8oWybYfGWQ6YXnh0p0nxvp4S2CM3qim15da2dxJQHds56BWrrpJaVG3We4ybRic54+avEA+erCLKhqV1uQbt35ftTonBlaifXDiE1nHWuV/iAkd+Dej3xBbU+w8nKKhcGPqdtgZvp6LTKMJjLYXnKtIBar8i6z1Ew2zw5g+R+os2gFiBoFKlPTlUbPYD3/UEjgELE789ayKMqgmC8IkKoNd2CMqcyk9r67CtFb8D7gAr4E1hTu061Wha+9WBGJNJ+ANMCJMFyd8pa8ukS6p0Tc/upnE2kmkX7LUN6XYTGKcl/VrhWuVvVZe56AkmqPQbwlg+J4AvAkFupDebR9S8sZjfJF+3IKOiQiJVIijYZcxzySbeL7YhUY4VlmjO0ld/NkC6I+j0BQPDrd5yJhR/gUNHtypac1MAkTCVlNU3QKjV9wYm7cPuVQId4c8ZRdOBIAbUA0bS29aenrYdd1cg6k6lbMZ2UtuPrQiO4pTrtHJXCqwdgVwYa+fC4PXza2lZG3NB0eO1qicauw+UJXXPd6eYSQ+g9ytD7wy4qO6xQjka5fKRqeebv4P3KiEqyzc6MxJclr/j2j9hQ3QcMnuvChfLz1HvifDKi+/I201nFrTU3vP1lNjzeBFvtfklyeJlS5Yjp1s18iVFWud67RCQXsX0MSGWb2b4tOCWzOzoFQp9iYxwKw2n3+vURqfunHfEZEAP+w6C40lg47lIFF22vKRsqW85xzTSIgjbTeJf93HzIHhJ9BclPiWgM75VLGoJEuZRXTqpOfOBKPzqMS/MCFKDkTTflKJOy3L8+CxoeLT++D6ZBLv0w9QGy/meM2ddqstTK7rQLymG+eB3NzmdVagg5Smbw6ypuyAmh5rxYiksjVsRemGBoC7jCyoyviYvTloF5fxutn7W5AIArqHiY/E5LR34S9btlhE0hRuLTdmi95pFV8plgOTplc6uvEp9+mXKzK/vyXvuPtKXNUnU09llcELrjFUsn8Lpr1Io3X8zSx8aZVG57Yv8Iu0lflsJX5wAW3QjcjOAIo7BOvrQjsuBTPLz29obr3Wpso1BCUlBwTNYpQ1St+MRwyA1BrDBFP0dx4Dz0NR3lfNVZ+dyfeenBgRLuJJake7aqnY0uB11xx7Aplsxsxs2PQG0tRxojxlco7ztGyBOqOJ/ulw3jzDZrSjxe/nWzabIhZgMcr9WGw8okRs1vmPK2fO/bN2SN9yPSZ+RNcttEXD709JxMyx3+c6m5JuVWTwLbwGggqh3GCsU6Axdfx/hnMORYYuEI8k9Ve6xfNPgqFqpq/gUr6Gn14vhBeLb4Dg53iNs/6kZT++ewx0r9gAXYnww8c50+9GplGHizbmrqRXs0/qfab+wZBKiu4hdL9Sy5T3AjaCJref1D8lfvACBrOzzLgJWUH0Zl7UZLk2NHZKWFiBc2lDcyS3voAyphJrs09olRYMHpDQ7q57HTnMj5TMmk/LxTNHxab1RD1QnaMGjSnf97mo46XcP1Z5MQsfq9lj7hdB0w+g1e+7K4kIi9Ea3MhgU29U1xxI6X9XBQEYZdah7xu3wECaG5DLq8OlVj6LlpSEPTbpRkERKs9qpYBAwBQE+WSxVLqo4tmPdG6x1vm3cLtXeKgeL52LjBhhFjhzgOnIrx3eEdsskf3MlabOaTMD3kYeqswhaEz/RP8T0iNw9cd10DqC5r4skYLLFSucSmL8wRV426oSKH2Q3SVR97/xOxg2ZZvbKpB4foO1yjMgGqAmBkxBBQoCHkLnJnmHSpKF/su4WakuUym9To9ImjgotTge2qcZNO2DJ4mstlz3vmNP3iyCiLwefVwdVgv6A0QKw1ygjbTM+A+Dn+T4j9FZ1USCWfVljucW4gwGl+VoeOP0OEW4K6700ifTBeaaqJCQ4c2tWXUgUhobu/S+l9K5qNUL5vpiClaoyKs2TOVKVw4rtbBs/kGgcBQr7jCMdsx7b+sXj3K5SsJWth7dkvPUjQ/gCtSaStm0CEvd+Ie1Cr0huncMwNPLodKvc6wuOgYZ2as10mi7wYNmLZgCn7Ve8e4JCBZG+zvZdIOFSMhXOO0mPtJTh0tfo+scLTxHWu2zcMO8wThydAFQPCcdtvXnsahLPkytNZrb0V9KFqqg+Zy4eG1LTpWegLnh5XX4aNbq0i9mo6+FxzQaZCGK+jWodriJe+Tl8aJxnQiiG8xpP0dfLxm48Zyd35jI9xwDC2duMdHAousgPDGhk62hQAs+rkOiitLYRejgiVonfW0gJRO64LY+gnapzjU0KIij2huSUrOeMD2C6yOGswz9JT1htkYHqEJXlrc5Z57jRJSvIs1vdHrfwpnl1FrveHp+1+bGmjJEdHsTrRd8mZrgeqY1vr/BIkthY5jdCefGS8wsUdrHnaJpiSuj1khMUN1qbC2lHcATGLvWjLMzzfCb+yQSahEEbK4XMCGIdQJt9UrgnF7LK6aTTEkhJ5sB/vSldra18tQDI30mmZf9kKAeRKRw35plSEzVX36bNJl3cSoge8I5FHLaDGT7mp4Tiorjzk1yCZakckE4OSiq/JepZCMkdhZvH+gDXfUgpy+PHpaVxFX0T0cEGr8OfnjaH/jPo4awHwsfJxBgYgUWo9aQQPFGUwt+uViQjJ6un6Gnrv0W8gvmEgl5lAphW0zQDVggBK1piFyWS+DN/am9hc3wOfuh89ocGcCvs9alog4laZrP/cN6sf/bzdbOLhdM9DLuTHjcHIY1E8/DTYmzkuT4D5WSnfHMBARQZL6DHGuCVoJXrdBlLhISVi/CJEtha1OJ5VsAeNSSwlvdB83sc1+/LbKVpu52R1FNS8XqwX4dQbGB/2SMDImcT1l6TM8IBy9oyqgZ654J5kG9BiyX7ZrW/JqCM8NM1x/HLitXroLTVwFH4RqRz2EEpmDhWxHfezEGM0c6KLL8/T81bEDgFFH9ccGI5cwJ63F7k+nXCRIshsFA/uNvB1f2YrtWUZdWNl2/ZooU9n7mzSSBXKYO523u2ZNdGYhBtFpDwV+eptg9pR8rky9+hS/rKCB6ITHaXm2vO4XU/GTyoIHJ4FSmxd2fIjw5uUC/StIiZEQ8x9YHdWXAFaG7x2UAUPBvQ09TvFaPVv4LosXaKGXCxZ8fW4C1df/it8zh59ApyixQyi/mdtkN8i+9Mua0aKj6O8/tQ7orMNAZU0w9EMjbv16uRebbdsFTdPrlnv7Xt8AWA2PMY6xYjHQ3K21LlHfaJ6139yNdPwfbnyPg739FA44dae0/7Axmhe+k++lcQAOKCyZnjatxX74NqFoirCafaTXKyhHtt8J8oiOepIoa0b7aL2H2mBR06Q4pfAYRgzh1DWj5gdTTwmtApGYFbH7TLXbdGOpg5yRQ8mmuEf1Qp5y537svzBSSZ7RR99fjSzcv7L+MKy4ohOn03r13ne8VVZ+RdvlXZSVoaq9V5HcIq5LROwlaa65kB8ma89mtl+6pjGH4DV9Z71mPdeWZzgq3BPvAXsAnOhIzbD4WqdLB4QB3R1CrEkYHIK/z5e9pxm6eJxxHc8UVijXXEL8uPWk5cfumuFYgeLdLRRJWwCKuSEvJa236UDC3t7IorVTcZQ/U1poGCgQdXdKkedAjQf452GwqayhpmncOFcDqXLLOLh6NG8GQsZoNH2WOzJH9+URLWl6qfmOXfTNjRBQX/QPRQFIHjjn7KQXrSyOUYmrdHVXuJutkgZx3YACB8Kwh/xqhCfVsZvL7A2Ag7K4Ht8c1F4wADqAn0aGeqXyEjVVTCnvPHBGqxnWTCRVMSMZlbrngKDPq2ieoXMl4gzIevMvoRS0mG/uoRVWJyhAqbaQe5/B48GEurB0Vj8FP6wv51NKTLC0tMRfGCsVLSuo93hy/FtE02aHaSVFgzlNfVP+8WLwGeQChb34Q6NXEXf/vmRTT/sTH7emp9aelu+4qImM1p71ZfVT8C06pZvXrDXuKjDC4rK9NtfkNkqnpFEXBmhtllmEGMcWZz3FUodFoEsFvefM283pmXWAPSVtVcIYY3AzmB5f7eBydURVssQk6XkFWqPchR5WTNAlW0gMEFEnXkyA2hVepKmd4v3SUwcYX5mYnMM41So6ATNy1ZeTUTZWkGTKs5FIvjEHSNM87rzL60OZvKW08g1rXJWhANTVm7j/PENvCtFhvYfpcCYcU/vgWJhtoannARIC2B7DaQXspKkulC1+hbpn3at8SxwIEkwEnWmjE57JhFUCbjrJyUhoJ2y5N+cr/M+S5OMh93b+B/G8LCVUM8xY9OWTLdhpeOfBDXEJw2KKeGZDAMr2d+Zlb/JgdXHYMGpatYAsCnEKT3le3Dw7kW9HYoaVOddid+Zqq4wJ52OfQNKdQsqzgURW+ZOmiQm3NNRHPwP9CBh1d6+ghe5t8ExcJWwU0anloPzLa5fLo8DsEihtGImBd5+ZGvjtmLz3E09oiwZcVprywuNcxGvSBytf9c7WPQNhBgIkUZ6/0Yl4Y1ykjjV2BFT7rKTR6VltOKnmjbGunnINNs8ZoFiUKdDuTnutF31ijdeJ9nN1Rv1qyKkIyKu5qqlZ6H365r63vgfLO/MOBWwp6wN3JRDOI/wIpurJAiN7Ny9cJM6Su6DLPcG+7dCQCxOVy1LHiBg4hFLXkjIm32nZCMadm5FA8RU60MBEAS5Smby2mlNuFYVj28WEQv8LCp35bqfQMi8YSTN+hfyZkGGcEgs6qldlI18h9pV6tw8HHC3mt4pi+G3WFFMV0ucWe89roq6tfQ/nvRIzqUttfZvvqNQ0gib3i4cczcLPiwvMMmLJuV57GI6IBPdU/gIIR0pjvTMbnn8ijl+CSwgJER9DP8MQWOWY0SQkNQujA5SR+31ET7TtXyloURuqu768i+HSi/wILz4GZ6E5WOm44c1659EPn++m8o38SJ7aY4twh/238zUBByy+Z7sUxcO9wgFdcGAKCckKpL/lrx+6sPcy/2l12MPR4rPzxEXSxIrLnq6UATEBdG7zq65HtxMYahcUiUpdVvN32yKBSWBESTwA+vftLp1i5i0pXvM0I+xwxpdIhYlea0r1lfFODJ/nsZBYgzHebzOGnr9rhrgb5tn6IqxF4nGDzjr0IfMF/JkqsdXtO1ZAz3FEvlP8Xk+S0m9VQI58KKYd2+I5yMn4sqkEN5MCyrXslTeql+SEMMgla7/IeufYdefmz07GhZTNo3nbd1bfXiSp4OGtYdZdtfomsKqjoWCIt4JViJ1LIpIqMvgnwXrsu/HgvzfTCK7PbsojS9zGKW5KuiZFlHAa3ZJqQPRTJc08RY+njhHOyAMJDdm4dR0vTpg6F7ZnByq39dysJ+8mMsFP2WqQ0eRhszO9Qn3gIDylcYs7nVmwt8ZEFomu7jAITIU94RxE9jAIFZPBx/ELGobt3WLDJpycTte4ociEyshLYBtu/Y7BRGms2jb9bAYKX/83HQWeOBMcMorBCZvm9rAz2jGFxDNf2seY/fBcKxy0uqER+w7wNYTjzRuqzKLv8c6hcjAXvXFvS0Yr1+s41trIPwpLHBc2OX6i+T5EqsM3mViu/D+5vIRamQ9PSe+75rmoM2pmrlKlIZjnad5wuGsHjXrMC+nzSZNS1d1GYe5f6sJv+seb6PxhCvNbWxyokNPnRHGOjFZpHtf4AkWti4VSdUbvmaam+kCPDRd6ZTS7T69ykhsXqJvp6fHJTZ68LM+pOIOGXEru/bld8l2hunJJiyS87HN547jHMJo3GumpFeNTERKWPZK20QcdDcmzg6GS1QFh4JeKkZHhQm0nsipWDGOItY5VxeSbwrycvCFdQAhw8Xy9fwQPlgdMjsgO0ah2O2a60OIvnCus15eWsul5Hdrqd7BUe1VbySd1+Ewe/c1VdAKhv+NHo6n/26S/q87NWaFahc1tHJcbSb2yGyevkYaHd+UxtdZOmgBRRBfDRtSk9KwRuhRIxpWHEUF0+u9KrQV26GY4bVbsHX3IZiuQuCekFOrYx/vyerGiLU8+q5yKCAIGOJURtG3N5ip7ez3gK8oBJkXh4pLYWC99Igk8CjzXKFuSwC/H1voTDYvBvcyJ/SH5TFeIWCV8D6AP3HEhPsCVxU1s237OYkPn2oZTz03mR65vOngESlRlNaZiwO17s9kyLGsuGo/L4zFhuKKOO/BLNDrzZf1LNf8b96G9t2XYOltaUamJ8EeBnwEmo3RyP1EdC77FFZqS7o/RcyKhgV8pPr0rCKa7Sc05eDoeKUBVpZislFOUZOOYiut5pceZYMqQL+n6ABzEURY23fh6A53285CKP2YOlyleEORwMYC9BOMvMbUoA27kkgXTalq5EOBTIV+sS6F8ThrhS/CXeVowJ7RRjRLknhxS/Yf7/goiGUf0zzD1HyMTKRvnbklZ8GoQSpVZoFuJVBsvPyTZ5OMx0WVgSbvhRaVYKonNOCGGjOeuj9I16LWsdPxkrmohqPhOcTkSwWlSWuNWDV1/onO/EFETVSL/ORwi4Vi1BFKs382/x8Uj52BXKrlYAy6UvXzWaXpUznmLj4frgrDe7pWBG8Wl8SX+S0IJt1RWudI+d+2nLm3oG8/+5yEYsLszdPUxar8PN3wFFHLtkreGOz8Au+UYRRLYwBqJ27GTjC3nRYf6NieDdx7tNmP60rzppS5jwS3VZWDkFyDkVNb4nn2W5JR+pHeIsv4y5e4eR+6odC3vLm3ifX+gOeh58SxXbKQkngYIi2JsfMTBUw2UWXmGeh4+QU1ggkN03p++fNMh+GGdSU3jlb4yit7z1tUk7Q6OKB53RaG1Y8+DJuUws245dU268Bw2RsZP8h2PWMvsU4yQQ2ebkiIbSFjDh1ohPtKm56oPVXkLznp6VaJbbNseZA9XdCT81XpK+/+zLQguU9B+4+G8meAEfwbnnMmpjyqgMsjnXsXq1xEdBK7818ROPn//oUrmK8qskzP/gtWqiSZ73wMwuGvol5VT08TEizzlh0ue1QREViZC0XuB+t4AZuo+zQjKIKDHv8IMaKD8ep4fGkzKFJNpFtLVThIc1XxBlLWDE9W1KMAj0A5JbC3eLrMZXlsUWIk9aCQeo4BwyMBgw/NhhAsvFXa8AEM4EmroeusidCjkqZ7+svD6M0VhUT4Kls3S3YDAFjFimNYgmg7VPPMbKifB2mlJMDgvEtcdrYXcg4XmEoU0lOf66b+QJ0U9CXjW6t9X6/gqCw+0nVODBPdamZklN4OHHrthqvnsbqO0noImcNb5jzodw/Ojh/NesbEu0CGs3mS1vUT/YJ8wSsu556pn0pSXuGUAbtRd0/FGU/OCdbCY5pQnd6FbCYwCJ+l+FgDsWaxdaoaFCx1t/KzAPM6dWwNJdSXQUxHkrnR3SptdHFyJWbWpH8b1SKpuKUuRdwchkw5H2eCN9bmgpYmH0KGbwZiZNfvpzPwk6uGflw6XkOWIWL7jBGqncH7sBc2PuNHLgdpBA+EmJLvRVWrEKGXRoGWNkQTQMWgGN5VNudTz29KDAjplt3NyXlWq8H8dApks0Pv/II/jykqCAPFyTdfAVD3EdVL+9VgE5jL7Fv5LZ5SA3IlEsEafO/YDVAoJOtfHer9O1ezLRHKSrSmd3kitEoHvlqa0oL7p8mAHELkLoHg1dREXw52EThzmEmi8MbhRSgNrbssTOrQAeKtVSNY2MobQwFap/9iWGTV62eXQftpjhp6r8GQsUWJP++DJdqHg4fbzALIwoU1EugAIW4lh6vVRisIBzCrjgaDoGeKm2RqCfkkuEtVpDVeK1B+K3RSiIUer6ShlmE+7DE+h44N9Cx8VThwg5lAhZuOevFUuQMi+QA8NgZJY1RUzSYyeDg+78RBKZ6P6I7a91zyNOeY79ea5jnta+kUsV5nW0Njg8zna3i8Lnzx65PK0Pf98FJqIcyhcruOe1lm1SopyK0CfOVYjFMNjXzJmPp2WxPtTv3vFdfJpGIypljaFzrpmJ7T0s5OQiDFUpzs/7X4nmA8aE3TKsk7jfLv2h53VL8XIk23mHKDGh0+70rZKONHp6p3wSHdkzc+9jUfiTOdNAp+SdOwSxBbV4iRZf/+vgcwyxgYUZK7pzoDdWQRv7jQQ9q/U2V9XQ7954kUz6sKYrvJhRZwHysRufEPYXxgQux2wZNbysKC7mfJLpIh7wG63kH+iKllUkdd2UwCz8TyF4gFQON3If7+dLkIt2Ikf/4oCO2fV5kj+vOsZBiyQntulbGl+sdmTajlCxM9k7ECjFHLRpVGC948wES3SmrT2VlMIAkyVKWRyO9Q4JeKVmKl/knolJ9Og6WEcED1c1CcLbED0w0pz5RqNMErlSC/OQTPjZGoF0mmxH6SYSCD19QPPU4E9yXWGktfeyobLP8ZnTTNQ8DoVj+KSdakjiN3MrGMeTEbmSa51aqagEPBcV1oaY6PerwMqxsEdQa0nLsU74+aRpv1+C0gTTBBFkZMx2P4PqP0aYTCCO4YwRAIUVx9dRjPSiU6B6tylDtrbJDuDOctvtrfypU6b208mNoE/ccikyR6jWdcytRaBkTQI39klBCkP+5ZqfIWHvochbU9C4dpcZhimskSdjc8AA2lly1Sm3miZzln8MxX3QnQ6ucjtqDfQSMabKw0SBCDWGzMTNNrbFyp1aTzaZY90zuOU5zPi9VTBRDMaKyiQA6gxexCmfWl1PSbOXhry+cBEH6c4Q1S2E6OCG1NIX/dDopkRKpo5gz398AJX/oRH57GGYc4bu0d7mLRpr+j3aenXvTdrvOf1+I=
`pragma protect end_data_block
`pragma protect digest_block
b626d65b772ef67a2de1b65c917dbe30ff15102963f434f1c0170f5264384e0c
`pragma protect end_digest_block
`pragma protect end_protected
