`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
7xNpdDz5fyx1clHtN9PydHos5epGFiLYii0jBTLVq69nX7zHxu2rG6MDXH9Qf6lfZrmf0oxyx0s/lEAaae+c/feZHvMGhsqbi78Ry/NijTUgSCZUj+BgDqPCcjDM3+Q9Fqb7Jbmod9oKLQa58q+8Gk+Wp5b9NXsw1LiHhbqSWNJF4sdn1LB/2H6h88aMMQtXTISAQMVHrkpZpxzxrYq38qtiuO3f50IG76nDUIC0ETioriQGeHn6TQ/+VGpoBF5Dq5V161/5Z0hti3YUnBYk9b5O81azw7i5tTsSgy0x5nzL6sxG4Iv0Cxhcqd+9P5FTsq04fvWRy0nkKlsjiNhbHala86GB8puQirpcv1y9j476L1rNe831TkkaMnGN/3pMV97SoMMObx64gAtryVVfpbizmKpXjdOlN2sOQWRylREyrhPZFeEqjNjFHocOY5sAqaU85LtDbGOp4ugWTbnrq4IzCdJkNDR7SGs5uJnOtakNkRNI0nnD3euSODLPYkTxPii/Jy0zGgGKVmw4Hf1FxJQnQ6z5tReClMGG8h/9ScsEM9AeF0IX1bGbOj3V+NxcJ320ya9aKn56rZYQuhXFJ34gqmpDa0sWLEry1IK8i+huQqvpJV9LoRjUwg7fBzHlD9f1jCDb/iZEn2Uf+GPLCSLLt9V9xXrU2/MchuU3ZFgXsJOmzOKg0+9QbCC7NBC6hLOpNEWgpiqHyFn6MjBD71mRQapcu16gx2T8ATXRqEDErZ/4inTCRU8KH2o3XqZj4XoM+7GULKYUJ5zBpR5xFbfHj3eIwNErKuYnv9ihR0u+IdSvR+fDrBqBPrHbCDasbNj7fGdl7tAmaedfF4OkRUmGt4TKplkcIO2cS01+SHYPQpufnifbs1+YPBaY7nFDQFvPthcWQE1+3QMDzjk+ZmkYLDFa4MjCMiyASi73KP5QmXUKF7ZsXo/1JD6ldw3lAWpx9WSU9SsFF//6WjLRfFQR87B/g1BAEoNW+jzgyu9dJMjZ+Cd9lQSiAGL5N4vpBP4jalM4dl+0S2vuktefYt9ZhS6FiAgFcaUcwLxOhCM+fJw2lTF0yHBl6JF+eoQvkc5SjeZ7fHs0jQZX/mox2Hchl80FvrsOcBAYTVEHN1nYD1crhb6d0dLKWtaiihb4zuJnDNGI8/syTrl1AZnD9vPQC8mGJaCxzPCWmvqZ9Ie9B90oxYflZvp25SKy+d8TXETo9V1rUhawQfe0INjTN5MIPUFF9+KcAze2/VHQzx471ZanirM9CU9/zMFE0qNu+MJzp/vzLdZIEfRoQxhqBsTHErNsSXzQlWnQRyCqKvQI8i7I9fCmZ7e+JD64KDO5f65msbXV0oNagqqKpJQdrSvDCjRmC3RIh0ahci09QXY45wYCYeREMlJKju4TRO9DNc5svFQYLLrX5+G90WDQYk/DiicpHUnAqqB+VZrX/7f4J7gGr4DIDTqSu/XvT3Fuhs7PvF8wlI8aYFmMQmZZrutdnpHh04kDguS7D0owq1Ezi7VbueDagBw+ouajUKCg2jokl1OH3xwthtW0Iq7i/QFhK5ZlWKFsYbEADAGU07QR/lLez5amAD7DwIlmruN38Io1VOwxpGOqcocS+CSDkF+UeYsXdie3dFKitR244kLKCLdrjJuFYWY9t48fChMOIXz2EOiUEz0mbubNsVd5sG8qhafWSMhGV5tNl1icx/ulvOXWsYP06pkCr8XHcpcujBQaa2MgTiG/HX20ZhBhPO1cfrIgxEpBHJNXnNhFGPVXW0PC2WRzchtGGt2PnQJAxyeEvaN3pmEbmtrUUaxSOgwaJHQ0DxbQqbFGkVydk76r3q4xY8I5nYgvfhRQF4Fpbcb6EKTVKEM9RnwpTloq+D2LTd8+I7+oZyYxkZoSkA/v0/OGFbw4x+Zu2xS3lNuHI3CEken+AFpGbdu/rTgvodxZTvK3kwmpmG7q8WaKvUXUBT3inTKRZMNbpIBt1CRTAxdvKCu7Tp1bBED1mQKT/kS6ZgWo/mu2a7bvhU9Gs5t190YJOtLtHj29Kt8vyYOOYJoq+PbkFh6o1MW87QVAlYsGddAjyt3w5NZ+mYSZO4ckJfHR8eQHbcPyqRut292mqggte9UgPUT5SZPxeOTri4Aky6+VkiyPwwcIZt7xdy9EM+vRsRVogwpwOmKhDEp4uwpx4IJsQ25R/8LHwV0nBfBF2+O2dcBGiVLQSjIQ4KK7HYoddumUaESGv6mX/ZVn+z15TWdRtIDh/E11rwyi/xhtvw1SlrWdLTcfRqGjhx9kZBAytcdmbUwpdeQkKP5LAmgN08lcvmNulln0fyAUHDnTQTm21QjVwsZ9lD6itXCapbMieX5TLqa+737luKZtMRqHDS805CTBGU2s3Njzetk0mGIOUa/avbEoS38slAZIo1q13+GhgkJ2tcelphLY93AzxBzqtWz6gKwZc81i+vuyOIDLLZGPSfIzPFNMktqxqiytD5f4kGLqJdwUR/7OCBiL1FLmhmWHB8NJGtptwjD6QLYEofmFXVHerYmyKTXOBNknsgZc9jJ+nKXhNFAUIkc7qiPkulfkbXD9OQ39Lo4M6S8mKL9Mk0rGbKtJR9EXYlsW5GMJj4qYukwOIX8O0kWh5cGBrhmKdntdZQVmB4fudj5DzM2ucQ0WGzAhmYI4QjjAcG81sXRMHwFru764FHGLkEbO0ZbCdWHYal2+FzhaL8dc8q6HaypQMLd0Z527S23Kx88tO9JUQH9zVJ6cxTbFAZ4rihk4s8ZlZWEDwpfq/uA0FSsN9LkGNYT7FIJnofIyezG6xrOYaHGe1WgyRtPIeGVDTCOocbnv6LJ3MsBdPjKUTPWHKqGEON6wWam24GFjBicXufBUG3WvfcUOf8FKHyIAa2ZAaER+Um3OHBuAEAmbLoWjyx4pEodbN7ufxSqRFJlIqczhjcRi9uEBgYJAv2fr2I4BholCAPs6EscwzrO35bzYM/6osK68Ps/hn6/UzR04JTP1ja3biWh9y8UOpuokIB1vQjij065iGvlgjGHSYn3HA62UpGnJGGb0l+E+UHx779EENmqLHAjEGEukbn+iLdsIVSsIYY+qbMGZZtFNS7DDE5ykCD4jJQK1A45Gda84RTQkptmRHf/3MJfgloOWrPHcVmBk1P7QBFIAQ/Triyg8AZEgPm4D6yNM518yhoclV+M4rwY9CtzOPm+Tv5Cm29NxK73O6AjIy6q51OrzUZDte6tkmibUes5SToN2t08XDQp2oCh0YITcjfYv97pf4RbU3QJxQm5wNq2F55l/5Evh8+UJOt0o/K3xQ/6u4GLQqMN8loaNwbZxVPsij7H/owUacmcvMS+mnVrglyUWzKYy/j5wVDrLs0TkYTJzlVaDSoafIpFCVYAyZKfS3Wim29zYx6FnRxqhSITbzJcIwhkkZcdY4mLQq9EQG3pfeqWaZ/qu2lcI6MjA+q3PwITcJmp3LT9Vu0bKhSnbXb3CUkb+2OQtNz2wOw0mTm3UdbgwjwGeoILg9LKz30+oL/Id/4lYhEjKQuzErPPgEYqBUtydMqPeG+7f8PSF5coynMPX8HoxnHNMhBz/WYCeIrEdrIuo97pKhI9NY8jlWJCAUEbaTMxsZY6hZh3yRupJLgflXZf9ni4ZPHgqQgH/SNJt8I3ioU+zirRXZLQ+cvQQS8yMPScRAYuhNSbmqhfXq4Fa5My8Mj4KVDGhGoQ3ny6WBh8Bm56c5qs/q5jmBT/E8opYp7FfAP1hPDX8MVj3CLz43CCtiwAQS3Tj0JvauC+Oqp/l5fTSVqOHjQvqI+dZNsDen/22t/VqJrZRI9rqgyiFTDaBBFhry9tSptTX30dHXno7wjRfnBuJpovKqXsUsKXqIahy3bmpERhAv7A14P62BD/V7TDilG4VblqcDbofSVa82Ww4XLzJ0TSbJ/s270orMBk3mw5w1Hya/osWJT4RLu5iXiOnnZhMF+pTCNVdfACzW5GLFdnHW5Y0rALH1hZv0DEyI7BACreogRiNHhKSGsR3rOXOGwwNqdMhDa001PKNlLmEPR5McEpJWm3IXXsuR+0Stn0AqJOLaNPacKHz42a16V4MAxnBvxJekw8ejTzAjQ7KJC5w0OEL/mW8MgJMBF7f8+DW40vmgNgK1bDYdeja7FxPx+mW0+wRI3PEdnggQA6T/KKehEs01mic4eZ94YsJv7y5mdkghACCOyNXbAChvP9tvaXl0N2no7XL2DgNTP1ig19r02xcQ/cFnqDdhO3fggYDhNql9tJEAsILn03XbF2GrdJm0WV/Cv8uc4y0DthH4LCJZGl6SmeIKhbCawv/5cjhBfy9yn1Rn0r6k0phc8EfErYoGPY2YUz+27LYeRvWGGF8Lkm/GkMMq3JrS4uHdufcKoZleU9JzCLXCxl/qappFNh7z8QUrh+mSQvzRIK+ff3Sy+nqSK7nasBlkuTQmxBDrxjonIuUZ4rTBkLv0h6ohlxhBFlXodYHh2f9gXYNYodFiZUxwSF8kHcDhJ7aJGKsaN6t9EUBo+4VvITkuZScA9UxCxNumazyzCpxntICMsdengQgA3Gy0pAFHiemraWnfSK9G9YlO1P3L6obygURTgshU04wOr+Z9abePiLmec4Bo+ECvUgED6cho6ze0L32xMZ2RwW5jJecvPL7GnkgNY6gFw60zkQBuytiYlUo774m9rWoLnbf+IeTnq94TJv2lZLMnUri5ZgKtBr9OEMUKMVGj9i3Z1XtfkNmyMURqYLNQvCuUC/dl+tZjv8xhube1Gf+YeP7Bfz1PMXPc3ednJEwQgEBNQxi7pbtCBfpB5plgECrkiZeAnWgfM9gqa/ASiWrP6w2kwMxUX5dA6AxRrGLZakQorZguXp4SXqB/RIxZAzJvaOmlgurf4M62TiC1SsOnP/W4XqK6E3hYCMTfi2vMIp7ttINQpMtuUZV5Zn1b75Xq3Ti2AsZBhreweu8A8cTfa1YUhTHurEsr1OU262BgqWmEp8cOpr2zo/1viD0dwJ9c4o/MMAITf/AAZA0bB97PpXMzBMJ3DGuGQ7RZdAOzQgKAkvHZE0HDQYnWxOvVmHLIK9AZ72JMMFk41dNFNn6LEm5mJEq8i/ZxVIOGHHfuzevf3coS9ngSvlQSAB3Zm3D/9vXhsOJwHjrnajlNI+n7t0i2Pqj3YAH1KDRmz/SZS+DuAAVJaxVlAawOHgLmm9pe9ngIgqqh+SSAVECuIoO5N7rfxfmlz74mrDxzMbPIcl1PfkFubRYhgCGoTAdammudO5LZ6H6BQc7YTfdYVmkU8SWxCdssKW6qp7d5cR05tAW1BllIjwu8W32htCzA7U1e2pAEHCNqBzcErCtnM0xdsVzG2Bu4MAt2ujstfTLgZnduX7IJrqjrVmwYwfST51JqdZJIPMxHCPIAo5DFAVa+um+/f2f8PRGJsjVRs/CgeP75SL2OrdOVw8gNt942zNuI3rNNDiqEpDt4xLTc/pfc9pVDoNz4Jl6SOfBZAVp8qq35vnSNLnemOh/BAB8RI0UlZEFKENicYCI632JC+BlcftZ580NBX3Pg5UBqiSYwazGBFwJbdFzFPw6yxTtCm/Mo5HB6Vj3UGEu7jJ3ePb7p8BhLZvakcJV3M+kw/s59Qf553KfbaeqwC1RQAfgoXj9wKEMSpvr7kngHbIlwqBD8jVlUohB4Pv+MoSeUiL+eTDAC4gPoR4hpJnXx042NXTnrlkzC2vAkMyYUUdaMoeqNIEiZKWNl3T6VCBkuhPO9Hw93YwEWIzF4m5KJ6xXFBqH5AWYheC22/q/pdoU6KsGjmICzoVcH35lAk6L2KZO/YovDFLdVD8+aVEWxvMlHxAxWQn4rX/Wu6/olZCG5KGhp4YdXqvLP60npFwALODKGofa0fFEFdYJjYdzxlHvwSAgANzp/A81JPk/dALTn0/l1/35g9z3rqlTk05lp96G+PBs/7Cpohg2bVjadvZh1NIXyNDxShaDZXUY1MV7h06YkXLfSEDLDqlVuNRKb6F8IqE6897O2TbtjNtnWKMrZyiyq5sIW1dowZFwAgSmO4ARnfnRG1+lHRVthWgu/kNPVmrVRd38adBOElmmAUU9TzzxP96Hjnw7g9Z3RO0NgQDZLr35XEsHFJsfBfuJqqZyYSfdgb1sxl2YrDaBS1eAngR+cf6pV4TmC346Ewr32ovwz7HZsJQ4lqDecBnfb9gInlKXtiRk/idwxkBPLfg1+nGqMU+mhjhryIV/+8i+vNnhhfx0mdndFQODJV0Z4p6qS5I8OytOyjSJeNgO2Q+QgULtXAqMbhVb7T7PTNsSa6u8z4sPoixEyGT10oy5tuH0VMekC4GiopxZGeF4PBwWAn+DEzhC+j8qn7QKj9qLJ1cw9QIihI08okCcrwK8aK6CzZoaTZUXcQwO78QClO4Zl1xIUSMzn/Fq2ofBhbPjIzIawmbRPZlGWuuJI1X91IV2GJT0WTCvD7O0vRjkarnKxoywkySWnLa7qw7xe5sQPSo8ob/k93KlmAy7ZHro4m5L+E6aZxGS3Wtu3wNVavXXKc3DTOLwTdCcQIay3HKW6oKkyHMm+9uT+/D6JQRNxv2feA5w9FrCtSYJ+bYEo/WMj2RHXE1WweEzovZ2Si1a7gm5G6Z1TKK2TcCwRSpOnL0BMOpDslbZzXov3pWQ1yczCP+NINDb9Uu2n1d7/Pg12JUYnqWPSkdTniYJX80+mb0oRFG+MsmjPDqEbP2I0A3zmigdNAyCDao5UwfupkmRrpfrJVM3RUT0a9yOfcudDSX2uoRDg+Yji7N09qpuq0+nkeQbPOR1nY6Ge7MVJaglk3NZmrpXcEWqY1nTWLL2APigni36zEJyieIC+/J9sIbVUrJBiL2w9kPCYUGmdu1eGsmGcLVjgTb/3203/8Td8d27fqQwQ1JrdGnQ994KxIDClLbX2SsQ4SKyRmuJAVugLRLRB96c6dMfWJ2ZMHdhqjRTBeVCcKwN0FllTlZk7i+x/uxuEM58YLF+dNXFOz8YU2A2iCL6DucfJKaSzmtGtSxA0fbvldWNEkzujb4BWTEtjWp4S9atDDtWEsMtrBiSBlUFRdO+Zq1ZJkfs+YSJ7j5BtlDdVGmbbsO/6KtVLpenNOqXk0UOp6fPLRBCn5dTFWpZuyyS5xbQvkMorqRX1dTHWdGTJE+hpz/s3UODabO4lkKwx7jLquMmpFSfgXUWFBNKaC3C965Wd9uTElgNsWlbCZ3vhTSlo+nkhv3dTBn6vsVq58YqE0nSXi7L6A/hv9v7aBIHPfZDhW+F7kQuM+fTVvKC7oo3dfpJhsRFDxFSAi/bFc3PdIJkg2Cu7y7/yCGQn0iTcjwuNHCcJ8YI6gbqUVlVAXrRrDhnJItK08x1ae90kPY1ILAAYA5YDWcZVJMeMV7cv40xKtHZzChDwja6/N0KiOI4okYqgJZKrdb4TNFRaUpZuzNHR5mlwIELtHU/kcfDILjdz/2b4EowllORu58QPSQ3Oba4nU/UVXIdbvtYgQS7etHQebjwKOU7/GLSWhWRJFm3oYQvX1QyQ4pxMfzRZx9iesdVH9ZUxgFOwCIGz9htDv0p9NFcJm7G1oPXGUVgb4e/eJ8XxnoLGSNr+7wHXWu+TaCQEnYSz5hEO1wUUXmDGIhDal1ccJkK0Uq5aGL+OdC4aYKfHgC2vj0t4/rF/qaV+fECL+uYZOAdVkbQkgSrhP6cga81EBRq7w7swr37p54r4iMTlVjPNJnlqOvdETPWCrBokf6nBBjCXpenrGCZ0BAHrggRAw5LZkEYw0U8Y8VwseH3OteGGSFFf0NJKGm7WM0wREXXtxBu1d6oH7Vb2BSwER3YlXmu3BvNfVckb4JabixZO4KK82BjcwgWCLA1T/rbZEKpQir5bu02F9/gLL/L0qM8fMbDjHrDBlNsIoh4p5/FjSaWcZcyK0XQiNdtZrI8A8e2qwCWCL8Z31uMapDH4rfmdfqiXsFtZpyhbePUQWiJXhxNMTSZ1fQ3rw/WGouREF7i6qrxc/7v2TGfhPUWstrOT2wvYhgtosbU1m0Ea8I4NhDmaHHlTBnj31WDh38RODorTkaJ6sj0FCbuu+43YWPFwBWzewKKto+p9rIXf923watW/96+hmMCHs1ii8YQ4FB/clDdGMeNTm03SIAOea5zLMAs7F3PMXPfwOHDfWtf/8djomZQbuR9N3+mBKHvo521n6SKzhd6c2uiS379Wjm/0p4e2nrcQz0rnuFqis6RVzVqYdY2+LJDd6VqXWgM6YGvn7knp0EEfMswcfl6i0gTkR+1uIU14kvb0CxU8MDxGGlxXebx/6tA71g62a9HYvOYEAsc+Tz588cH3Kv7Mc6A6/1VmW8NhXJBhsq6qS2OXamspqYMkCkXh4FXMdZrIeRddqNvsMjvQMKXlrI/fju/1obAFCu+UFHfNP4UrB0VHMny8zk3A0OcT0kwX9FkdJm8DaxKadQNitGghWffcX3x+zR6fKpsViHMJl05efZ1Aj48Yr5OZiud/Lw50/MjV/spoHj31sLDugWRaa0mtc7BHjhNq4oln/KhsJcArRZLZU4qIFGxfi5CHUTyjx2eanI1xMaWR3hjvk4elCh94egj9Wolb7Cy2AF2invsUHAMpDQiEDrF0Fd98vVgP6hRlonnlvwQSNzsemr8GgGkgz1SQuic7Z7p7IUqnOClo9JzE9XxT1ml8iWA17tLt46YgfEqdOuNCPDszHT/CSpZ27N15MoyYSZgskPMzc9KDJ6GLL6ZcR/7PAp/lsUhwAtCnFNL5eVvAwya0BtYOCqRQs/jE+8zVdtWcbX2Cv2DJj9PY8f6LDsNlB88meNlMCWwqzdsQ7qhgvdAbqh6ZvMWP/vnMPGmlGFOApJkTiyklJnXlP0yiIZXtA016ork4JRBr3IVra3+lG9yQUDJfXZbsvKvPwemzS8V0m4AMAn32PIqMKBShN6vRYeG9Ndf2GjP0ZX15sfAy/+QWjsXiCwCVURSv93wSKekkJk1BRbBMnx9fjBMOljm2tYtpEnrdzhvG2+J29TNuWidwkqj9WEVzb635FTLG2CM3cO1wAxDpEcrc37tVQv7X4Ux9ezuX20h2YOU9SYJ4QG+SqkSfIlHKIn6H34VrTxInfe5MSk+XTLo192ODIaO2/uAIn/AiP6clvTjXS5KNcRFAUafDunKdc+otOeiLQRYSV0BZdveJWAsFCyksBtf13iTDR22Sks4D9oTlICGH4UW56RgcKYTnnEYOtZ0DHIuxQ50gwukZGQYsh9SGuRhZxqof8azjpNKZLk3EEJVjE+5+2YIW/pfoXaGeMVF5jr5gK0epcNEGhAOB9Ecnoorvmcy675EQyzGNsLkW0NSDoNQ6BrNUd0xhfvZlpdEnBrACmhiqnPyjVotI+MLNm3S/NL7EdkkNs0+p2eh6r0Nn+4UHDNKy+zZo659hF6357tJvHcuvdhIYAAgMIk928taAetgNzlRLuriT0TJZSZ0CIZKPYCBHZ6fg/LzycWJmvZxZVLRv0S/9gJ93JFA2662KlYcU/d3hMX8CzVSaTbbkGL75Jqmku0iOXQWLAmvssXc4B9Kf/pAF8D0WT2AVchdOXV+7IuBpk6v7w6yQgl2T3c9n/JnzaCi2tsV67xp1ti61QRs7jRCCO87v/fRvcNYsd7lRsUN/nyWs7Rl6dfZVuSb70uSg6JT5F/EXZmiosLW2r1r5mVJJ33jjPk5z47yan3QT+yskytDjwqXHZ0LkT7BPaDycNVmBGb+CL9Q2HiHeTC7KX9QabzT/dtTU16TwFpqWZjfXWAjk3eTW2psROn3LpVu/C/arcfphjRFKxYUVdw4tv7a258tMQUFtmvHXCc9eqiyxKkRAmtHet5MLTAHLyvWXgroER706pHCfCuH+PYnzb7cwGmCybNmgsfH+VQ1SXONVq87o/jrg7UjtslKpAXVzYWZwnxLiFtOHJqrdxnx/bxs0ohkQHZQh8zH8vO1yuCGyDM6jrDUCQ0Dkj1LP0Q8P43hmsSALXEPLO1G1GFqPsMvQ/f7isrjqOhxFJ0tAaerCpOYyg6ura9e1PcU4gfsmto6NphooGyAUvC5zmrLvXx1Adhk9nqXQVJrdtui8RFrFXQf7oImfrXuRpEdD8T7fQEXhzd9cCy3Hind/W6qKfZ5yXpdloWTicllub2HvOwfcApFxGqXvcjcvcdaSY+SV3kJiUWoZyxD0PbDqlso0MLF95ilGJ50Zyk1JheNaU1KHuWr88ggxIvGClsKOdny56mTav+BQm/hInXhDT8TURwxBPAACORhnR7/JwG+fK2eyRPHGIPu+bbtYSDpqxrGlkq3/yetTfe7shKZDAN5CnQv+5zyOSwnBljcZHZaQ4DfxxMj74LW3VfZVkZ+je35NUF2GSsi9sYnjMYAztLTEmnT45ZZ6UxEfdyP3sSjvxkI29uDAM4CDlV24YUFkHetStSwxjzP8XMzAjf2t5wgoRcEJPhFIXI7EdkrdD3flMvjDehVpbqq67Az773sEk3R+a0quJkGluxN4YplR4sz+6HRMy6cxJgdl9s2ezMbwpjXvhnzyKoTRkmHQU0kFLS4+gnug8iKhv6GN6wDGrMoQPgxDMnL3JmL9HpCemlaGyR7TzUEM4crui6zqsCPAuVI5nFkIL9bWWcuvk+UFZRxg+iK8ioPx6BKPrk8UrXynji3IGNqMlPK9YXWd8Jl6zKJaxPMM0HlEUkfB+PmukiwA1cEGq3QsdW0dsljtMxuY8lgw+oQAfidW6KiKZQ0gYqKd3EJPT69RiKWiWVcxcyW0x7A1ARsGbV842bbs046fAutFbFSQajaLgIlBbe6EaWyBbE0dxSGiR99nrUcD3hgS5Ak1ja8mrt8ONq49V1h3JMInUUUAmFjNx3givZVgZ8jlvCEYcpiQa2r2DlSNOwCWkLhKg93Dp+ymLUj+CYoF8z4pRKTbi5cJnstdC8tytfeGaxTqvECSJImrPYZKanbwan2GVJH6yxTqvnaEfhhU66RI+9mPaN2KhazdGHUytnBu8L8LmSsW9fquGmPYLIrOQ3i80vBF01FufxYQCre+fPpZsfNlC5LConIRixiYwKXIos3idW8Y+Q5G1mvZYmPph5Be/AqM6a6MwsK/wbJQAqirr1jSwAoug+yi6TnQa9ecIUr9/8M1mY5DM0bxI8nUl/THQyL0A4epvdQ7S9dI1VgHOZETMAieeMA+jLKLcUcB1X18rpoM5NovBmvo5/RzdGGXPBHRlUps7OaWcSIrO4YISv0Oz9uA2yRlgfFp/co5sU00/6uKI19m42JCgUyG+lbJIQRvSQMavZSxknKCHM72tcGmpktYbk75+2EBYRgv1IjaLD5Q86AYn3YcKIvMCvGJqFikA/vy3xY440Ws56f2wPem3YKBozSpRTSDDIwnfCdAmIjTpX55IsfuIA4873YC7C+TcRwsCkbqunpIjma0v4r17vAMYNNPZC0cjJQomfElHYFetIhTfpiGxovulniQvvxGAhNs0QTqrVRZ2LeRRgXndcQT52PXwAUxP6TcW1AruY/32ZhqD4KajJ2OwpVUWjJ0bl6JGJnrpBWCHAkvWqnkrFvimzqqD8e4rrCzpC0HRdhETpkKel7aMMG0u16vXGV00sxg65ulpUw/4P5MbX6fIXrLuSzEl6kGOYP7lDXMa5p0FxmEnAFTJWNxUhLDjY1lb489U5IUM37+jydMvaGZrH6XadBUDlFRJoqchJ5kCS2Uh7LjLc5UURiKNw6PwndY8E5XTwVWeEU714r0zTW1V25LHSPc0co8Ts/SFg/0KL9E0hS0Ui4/Ppgzx3BiwPft7RMfeHIqaKbLAXpracMIlYWceBAewM6Jg5+0P+my78QTpy072YCwC+wE40keO3N8Z7mMEPhkeuMDT5/ZBXLS2dO7QSVzHqiPM5auowC5GvvHQEIHpJvJdVzBTTZnJwketnMpy6TtjO+NcIfZZqwFBAr0PelQa46ga9/pu3fd1VXASV/pZ1v0aXG/vKdf2u73qDHwIDa5b0c7HzO2c2JpAX4n6yN/+r8vgkgWWGdu5G36gP8e7GcuFGq+LqTSnB5EEx3VUFAvg6BXskYZzqeeC3QzGzArTwRkz0M8mcQph8iUjDtDWFZXY2TL8TYx8ph3hqUjWvCSfICMeLqOexwcQlpZL4sVOW0/CH+6S8UaR4o/j17wkSmIXxKA4hanpNAPnMVCckG8ac4Saxm5hWGk6UwILMbyoJwJfxh7cnA2L6Y5SqYz5C6yG1x5pZaxUEPCTelkwi5saAhb+Vd++Y3G0e+mIiBSj97sSO/3j6MBOAj/NlOQxFp+ImoNGJ+/5XxFnox27rHcw4I6uh3ARk5cwJ0QuZpL6GkDfWnNkgUPonPuM92zEXRzcFWREydirjbQj3QsGQgJuhuoflRfUTl1NFK910CK08HK7N3yE1NldnRNZb7xxF9PL5uacFCTjZWR1FyOnxcKE5U32//aR6T+DdrpytQr2MWrHNOPVs2T8NTWKguMW+BoHTb3NAaGuru9PcuoSkWkMDYLQKmaHM9FoYT3jbW5w+dP0CSVCi0iqaGiGtnmIsPHJVSncXcbOw9rymq1X4Wt8i3wXqBmolFTucA56sDj/MlMu+PAtMdkU2OgAMSzu+XXi+OVbEmCg3wPtcEBLEszrk5TRGfcZ5WCUvWnyG88DHYynr+EAMRmx3XNBilNLktSMbUW2ysqXo7QL+N7s82KH67TYku894zkqwyYYXxiLHvGrG0mqTcHpr8YdEa2ZlYKaXSGWVY6W8BSblPfMwMv4YyG5BZ/M928yjYfmdfsMspEeFe6yKVgR6N42nr4qXM/32FMAldS6zqdZ//B7HIkhJv5/kT1uQPUrJFfCrdGeEEdmD9dgd0Qk95HNlG1eXD27No3B/sgJpSV2SPUK8U46W0nMdCQAGB1cq+IHuyEAbpwkhuudoUjDxBt5Xj0NJHOuf9M52OGIm6e8DVbkoJ7+Tgr9UDv89naD0Hp2FHvHMINMLS8wEHJ8ymUtsnHOcEPD6htFNB1GdoKbJSpmDIVs4z4gBEU9aw8RBSw5XrqIYvchF9QH4/D0Lhi2EiqRorB4V0+GfXMITu5EvsRy5Uqm5FQWs59jq8weiog/DX7O6luFa7FHK1b8Ag+bZEY4WpHQzkCyoTNeT5D7qjcrHWsZBhwtCQLy9/kKxK4ip9imwGbsf3sqALb7xCVo38N8hWOZkpcxg8xPGE6jKFCvIdYK4dJtvNBLWLdAr8alAJ/M6HJjcibCT8VJkVGe+2XSKubhw0FTe6nG9sIKNEWPqlQkFHXR+wuxgY7bdb8XZ3XmD8QKOiFMys88yLB84FmZmDZIGZhpzkU7nyAHYa5QOVIXmi3JmqfZxS9KqCfA0yjBLr9QEuRisy7OciUzD7kzt60pzktgGJDGzzoH7/GptvYeish0VcThSsWasoqPCrrBfLLlLz28RmCshqySl1L7ijr788vq9AbGBIE644wK2kgsMqpOnYZ77JM6/x6CJjBsUU7lP89m8YGevtEKbbw8aOKwlgemHBcR6E/4LWHzVUpcBmcmOFrYc9/MyDV5qiOaeE3cIKSbtqtsQPLqdge9yR2kBDacJ8FxgCfMcIVDnp2+eDnY+o1NX4lzFx3FZBwLnqOJaCLKt3LzRgEwAOTmXzdr7CthtzzBiVHSlBNeLcHa8EzINbY4n/IcKRD9O6874tKEeIQZFn0eAZugCSMVr5G1UCNC/vNaocdjMvL9PJnUIMK+sIwQDpiMkbaUBgEIlpxqwsUL1RC2IdfWInH/wehlpGeWsWkkve1GKBqMc2vXikRiViuVRW88qDIbCL1tvsN9OvCbDzp3xWKyClYSvjeE7ReNrRvCg/mQum7eHKPN1xXP4+B3IK5JBniHH5lxa3lBFMNuiXMMG+F/KJ2BVcknkzy7gT/ZiJ8q+cXLrUcB432LFrU+N9STwU1myM+j4Y6T67eYNfYgdBWqkTpsF72QpxVHR5rK36A0uxYS8X0jkCyD/uuHMPFeuNi55A7VuJ7WkFEf3LyWwIq4F+mHF7cfFJEbOF1MIFjwdp7wXX+wis4XTv2f6GLEljjFBtjqeeeinlWVtdQfoQPgtvaiT8S7QNkZbuuiehXipQBWEK8Iq0EeaOsFv25AG+qdioQXXWGn3AnuhJjmjuX05PurR1IZ0E7ShpDCS2U/DRAEWnn5EyFMUMwNIPZ0XD71xtRGQtGR71J5obDeOIrsqth2WXLdF374boZpSu2PtC7r/aNjETQwLRrkABPQnomvfGFQv9u2nsbdQoaL/I/cZ1VrgbTA11SvpKliLD4EgwSkvJPU6VaTOM5L4ovVyo9KrUVAP5LpJ59/Q0ARAqimFKnou7op2RJFHdJxfa+YSW+NEUqrIdnxc5s8nXDNBNRPUfcyz450lv6ADVTiypJKDuEMSEypMaLMl7+cnFcbbBrO6a9Bsuyd7wN3qwAwwkgpuF+KOW/2tQS5PMi4NwoaUJYKf+sMlLEhQKPoZOSZsscNrWTdRB2aAhmOmKl4P7P3vK8+eSZFkHuu47Mcbtl2G/SYs35jgg6oYf7o7MhIh5iZum1yRyteQZwZTNoyqYAZLLg5lge9rkXCjLGlu0VenBKDr2pO5ZSEtyKhznf5GOGAY7/VtYqcK7LQQzh2p7swZHbaBUFALdqjbDKxDd/RPz03W9bJzwNj/jnmeUI/jS2C/xTIeEr6DUrB84FXYyWGF4+qzR2tiK0O5m7UhyyuUmG4TiccrbHpkL7Bmo0S+qSA73wAWabHi6s4pjtqrslpqpyU7drqSudG5MvvSZaE6ITuEiuvVh7FGTVaj0Q2Cavpe4DijNoEVMIdu0xnCSaZ4laRA9bO568NlKnft0W9mVi53pcNDA2JFX0ct1zAauibze2eN7jBw02Od1SoDLyAV1To/D0VymtGclnxpTP9nDrtHekIuiEaCZfi0i1K3fFIYhwsKj9T+HN5FDWN/7DxYiG5Bq841U8hevpWlOUYDAWCFhbQZXdnEucU1BcQce6GGGQx5gerKfnIVyl9h9kyZXYSLwR1W170xoquULuLjdbF+TMdXSQfiKdaFZ2pEGjw/h188tu1FZSFzVqVLCTLSLMp/eHUKLgDBUUT0G1x1lFThgJ40XyiuMF4JIXmUOBq4AVW6xZ8QOADct0JHc8W+8A9Ue5qWvUqdvyameeWpbI/iwg4PniDKdPUdz9X6baqAKJg/HrgtNuRZONKQTYg9I4QbZZAbGHLIXpYAuFWztKtjHCl+h/4/PrtCq4FLpSPYgTrCD2wIdKzq08XYcKnFD1exp0Bh00+CRsIdM6wQZyhkKclrSxIKFQEjOgP6fRxyiN0PvZFWFH/sS18pVWrYksFvjLln4MrG/Dte/HZ4D+OsdYPn+3BQ6K6kgKCvYPHAZceg3AYiyCzlX+cHj+gpv00xuShRn49bGzd0owardNuHu0Z14+qEclqxIEfgbyoOm8rzJ/z4npw1vKLIsardh1RlF24I1AsW1t7tHUZlbzf+U6pQli0raXNCHcdijPR7Q1Z6NwmNcBT+pWQ3xTj484WbA6u9hNsutFPjr3C150zM5sONOBZuf/I780/RZeJK3EyWig9CCB9oTepDxJc7ZyZdeSsYi3xm4Jc29l5SrRzcoIz1+M9o0T5W87qoVj3z2YvFnfsCcwg0JJAhMWGj3KYCwdOESgysnBX1wb9Ix7I0Ov+XKbNUeiEHtyBRRFnRow3cHZTLBE/tAsz6CvrUcOuyToGo24+JDF/W+B+jcKAH9NgUGFQT8YLNs6qZE/ZllL8skFXzFMgR48JuAQmuFMy8ZfXXJUmx1jjBksehIHw56dV5X6irrqNyzSk1nhUwP5hpfe3QRa8tJn5qBGN1RQ6nj42wTCxBQO3hy92AwsEUydyZGS8Ay3Au7Q6Om5TV5F7EVFicnih6bZjoR46mcwhWrImH5v79jpUp60F4grlAzbKpMfh3rs5AgkSQJbVFzIn+3NJTiJ8daqjMzMfhFUe3tckXeyoRJQPNoqC5wgB9jTmpNjKdbBJsnDhCtKP5eiivE6uyPKflwSRL5BuCrNsNA3jkhjX6hT2SmkkdQneZkZX2L3NAWTriflhgV/PxX18dKYkScaTT2JSCjH8O4xPQC3un2SowMhW2U2IsykgPYMlov/f81y5ugmecqJDSL/yaiHEVMtyHxOrL87T2VP2gceVl9nTgyr4qTX+0pkMNyMghiRvMUhdwuTYUal4sy3cdEnkDJYrdM3eWhoudmDTqB2KL4Pl0Ot153H/DwgJ7h8LF2DuFLD7WpDlwK9PF85HtOttcmvcT9XT41ZZ+NljYGePPMr/49vUPcNEC4ugZ9E50Siawr7bFaXiw8rRh7/6cOCUI9yaFpyyJMOGUlNmgaYeftaw/R4LNdvzmIGqspdeeEtSsfEoiKOuom0orw7bpjwiHUAlmFNbQXhd07Rk3csDJsJ+LcxRKicVC+spJf7IE75c26kMjGsBlPpAe+mf5vNl9q4vKXLgvLnNgIxVHM7k2XhsrczDb9O/fU79fhZo/uObM1YCokIK7fHfwhUpnwIgLZl9Z+O11Xz1RpN2AXUZRphwXz3EWLMHuOjx6grDdNvkqwanWgLCmHop6LmUC2oJCxsofp1yCX0XOYCZbavNWnshaolHRG6n0Pg1bVM9zC4Ts0KPifXz2hHUzhDpchy15QDZ2zH9OzzSe5ED+iDEuMyRd6wuXSX4xd1L2FEFcW+KhaJ/pNDYFw4TG835P3GZRaS4BnXWjIBV1mKj1J7v8Ka6MGE+GtvsPyQlMq6RB/HzFjkC07U3JLKw+TOFPSX8rGtzDBG7M6luJb5lGac36nTSCeVSgtoh9yFugluJ48JYIRzNEozuyWEVkWFmkxt3Fm/kyr9y6hwjzqrMkbOZMoC2l61JFcNkwz9TOltw2iw6GM1uPBN2jGvGP7M6k6ejkqnZ3IAablyXa+BjOeh7bqWbr86i0Xwqk/nQPLr0ImfDENhiKO+hh8Wdas5da4ohRmyTaRW5zGvKE+/ZN5Uynb5zL3zt2xgaBDq5quZQ4cZoS5KJVdovisFRSxtr0JByjkc2OSM1IGmc2YsulnlqcFF3H5IPDp3W586QcfBl/TOsokL9Ujk9s8jYQtaO34d2qU3tLaH1MGMnbV09u/CPUFTIIlusbTIJtnfk3pUSqJe2zFGJltflyTMWCHUEfdO6mEbmmHhz0XrBkGzF65k82ETWYjvIEJZRjbZGtmVrL0tx9XnD4ddR1NvR8MZzVk8x2QPuaYNJVvjrHRlpK9Td/cJNfIbWogNjGhDeigjeyLWPGl2j/Ku0LsuJgGgeHT2DCowMd5EXKVFmnVO1IehISfuDbqgpIkhUbw06Dh2owlBQyVBTgtCCidMalQYV9TPrmfshv2yWHx3wzdr1eGSesCXyaxBhLcVOgbXMVCTK1fgPGffD4gXTtmFMSaRZqOrnVddLho62h4kYxyatlPSn8GRBj0fQtxrmucA4aIWxLziG7g3dBYRWdSQ87FbiR4YhISIjydnEZ3qU/s51AD4ZJoLAz7rjW5kKm51GAztBfGlJEslEhDKPHnHVucgJ+V8YZKLXubELHNyD7yQHrCfYjhVIX0ATM01JdFb55oNbmMkFhkCvCDOXsVK5ANwN60A6MzRhB1URGOGK1qq47RwlJkwJj7YT64k3kUTbVqO5t0uOz4GwFxRxMIMjGBPVw5USCXZrJlJpdaS/icgPb2N3t4RZWyCv3a+ntIfxUSRx6hceK4/JoF5OpUeQTTea827wXX4VbDmo6qNEmoL0WWS1NOKr7KleZFmP32vxUwG8e9uCpxvj7rILTm5cwryh8nLs5949qJ90/Vv21JkUCNyDUuoSrm1vM/KBhXnUhSNPQuv0dS0K52ed6vjZTjnAu/7oAy0M9JwNfwoYo99PhCVLU8qZ/F4/si3Nua7QrsXhnU4ob5FyjEcCss+oYkL0l0M1W2VJQEC4cKd6Q+AzNpaK2BWYELDsC73RBTi3xpG/+M+CpU6OP+iInMqSfKuWVEPZG3jAPVVOmTgHrmkyGOzV5gpPAO21WtJ5XT6EqQ0dY28qeUKio0Lqyf78oDQPI7soR2gfeCVL/4H43gjHq2lNK8WKM9nUSi+2H12/q78rFv2HaU8SOp3X5T+XEmR2Lhkvpe6udH1SfN7LKHiTkHJUcwQFeRyPIsgh4rfWINAWi+mJJWpAQ8emKSU8FAuR/t0WurujZqeYUrpu2kOtEzhIG3F0VHVCQC6eMeM2N9cwlo+YK3EIpJ8tJXYK9h6tE4eE01lxLcH1BLQ889R0g/To62bmPn0kSuZH9ZJEA990eJePCKrf6Ul7qjzFla3YYa++zXBmWgW3JhWHW3ID2Cnu5hi//VVHiRXlRbQyiUbj+BtXdeVjJszQCgvvNzEnlE3IFOM4QLbuRC5QREmF2uW8Ts4U8+qWv4OPf81vnif6yAykV9+8muMQ076No/ZN/dAEX/NUGEnfhWYAAETWQtwx4HI/a8ulDbPiJ/2TY4adB7cRs+b9HFHyM14S9TQV5+ga6OeUHA6FP3V336FOY25y9F/d2unm9ekTaHIe2RNOFJMA9ZWfI+D0mnCfeqZbhxLqXLBWl1xuy3qnkhGAfEoI6OBeuG+UZF8oPbEVxIzomjn4vAsUMlg7lC1H2ERCU4kvYhPJbnXu6Yx+VxDv8Q1BF1cZSGr8rRYheHFNc90DVQoUvJb57kDzFzBGSeP+z4kL08YGWhoxiPHN85/S9vWdephpuhDoyarFiU8IBw0Sxh18afurs108/lhXwq3aGuCfuVMQlfMFOyBfFee1Bmc9fu6PTY4e8v94uEWEElex934fZubpjFdiO0BCnu5cgGo2bdzGQ2Iiu0AsrHwMQFd7f5lodeM/UKi53k050LTbprz+FHEg3sYBybS11a+bgrYsLLMcDeYLBxaq6waBoi7Bg7pXzCX6jVQPykoeVkSpb90sxLL8Y7UACd30uXw0L1rAzQmeS5f7FkuW5kKzs0WaFqeJLs6ZL7EMxtvcRmfOCK5y2X9T5Ur/MxIIBSPGxUnr50erXq6vA7mZgtq3eB4u9icOTB9M7NUL7/u21uBAWyYtq+ZKlbpMsruN+KSUDn96VmKFfVcwmijJPyHr+0GJb6Rvbx6xETC6FLrAUFMhT6x4wzB8rFbcwMCBEj8NQM9eGvS+KxV7FTFKhU7SMqTSTKiR92+792/RQbxIjUCc5VpnAw5l1JdqKDiSz/nJwIh94T2V5+VcFENa3oiHiQ7v11yVihzz3vK/Y2QacAh/mdAALBOhEcdgm598wtFEK6m3gHB3G7jcZQOWymBbOWBtlXANLvBgz9CKCZnjFCDqscRvOdqNEnXRhqhFwxmET/2axlcbn4pdI7yXrsFyt3/bMGFU/HvWv/hMuCyh3plYTHRjfq3AjtAbrhFa6tbHw9f4mdj9dDD9qIXg21zp7NT1kDlqjVY9I7FQ2FSNhkHO9vW9eBdGLWQb9QH/PizmxmuGAGVU//Fn5vjI4hC0r7Zkrudc7RWEGnWKs/U0uQibDjMFqJqoUklbcjw2NSz5jobpbIPwKJGAl4V+fgQAjsqokTKbAqWIw72YJBzhoRb0l1L4te/Qvu4GNzUgkhXd15n5HJvUBtCrD1x1U0TfBdPhjL0hGJoHc9ESbRBeJ1hjjnFE9B05Ve72e7zn224SLRt/Hoyk8IBLc5pUHuabeyxj69Kve6CzxU2+Wn3AQYNwEiLJyLPsgJUbYNt8LTmdwK/kCecCu/APcdWmsUOUMqS7OMNCNzyDj6FFGm4OkLEnjyKre/O80z/mFKCKiDR+QJQRDYeSCdIx7luywmNvVJKJBdQiiF26jokBCAjyjIRjRf4CN2Tf69jBgTXTR/Yi9r3ZQh1Rt6WIgBYQr8vB8FldGWIP3xGX2Nahn2zECX0ZvK6Bzo1uVLvClQ6u7QF4TbycJVKbwt/wuY+aTZTVGeKvWEq7utxdcHhAJw/cI4ddSDlmM3WV7F20fbN8QfedlhsiNPlDalN+QW3Opc0/SDjvwSqLH3h9/U5AWc4IbafaNkdhXbCzTYy3dBQkabn4y4WHh975vNcGyik0mCo6UzWUoM896RVIyGsGRdi7+SUNcUy6QeiNmCSURbGrN2VdYZgZxe2yWDCzmqMj3x6jrAEhNj2tD/blgpvfKZ9QQ61AU57EBIZwAMk4bv9wGi8Qhw/ial/9vt2OaCs/G+rEkAeFecCxK9CRptoGPVuPFufEdlfcZ+lMDliUPnnZ9f9fq0FBa/KBEi14FsDogcjDP2GGSuSqMO2hFHySiYVdJOSYEzRG0RBU48FbRJvIlk0ExEbHf45MdYNKtxcVlN/eo/SyccfVyVdSQOKsZPB+NZXdhggLfHucJSDZ19Cf+UAyZXUGlS/pEtwOm4rP2M1audhNgWKLQ/WoJzwnWUkAsGeyS7aY0tbO2leXMnyjoXIbpdHRRfXvG/LtZnrk4ZGznWeQ+BX/5+bcYcmlMbBOumQVWt2HaMjqY/zXEtciMD1f0EwbTX6ktE+MOkzyFGXEjm4XnZT+rhsAbwPT8rEYmOQMRCyxKuN6LI1noKvkYhoyWSv//NvZM3lyl7OrImvnjA6CwzT442UzDh69Got09SWA2nEoxvHd672YOzYC9fr1ZCaDs0gUlAXyhIvReM9haARkQBtIJEworzigwG0qMW1qoQoEQaA59uHrK12VG3+dTwplO2L6LI2rFuJSaY8jxAzFhOCbQwviKyMeRrYu2SU1/Its5k/Qs/p3vY9UykvjScxnr3WRUt2SJpHaNXruqVcWcW+L/GdQ1r+EZDGfqxsz9WPNWY6j9PadWZoxh1Jv4TiZBRBNOd1zEF8YEhMc85ODZ+Eop911VfjEneIFy2u0sla9tlKCYfMW79aUiXejNa0raOiTn1la1BhPe4mAP4j6fdycO6/55XTyVramRda+vAcAzGaYNy61ungRgHNxeSuIMQUt38OQx+WnD2Wv+8CdWipnUcpx/HPBn2nGZlNN643Td3vQ2r/EKwirjTilWqlqi4ulFDVO/KxCnux1RAofIvnf9K4xvfZrmPQI38HrYRze1TRfXwreIhsCBUrSy6pkJ2aO7MHlWBdogw468ZyiYHkzCIWS1qQuK0mpeHLXLpC36w3EzZN3FDjOZNx6kRqdkOJbpLBRlFChERyT5Aalpbz6VCU8CJbooT/pqvloT0Gt0Bn99QYEAbjzpDLpucZ5W3CU4/lBXgYQV3La4KXMe+XCRNPfTlC0Yu4XXLMw4gNfgoqvgc3sZ2b6mV3Gd3V07rTAdFWDPHMSDhHyCcfteoObSrPNUD08f3KNnv5WisGfWP1yt5FR024AQ50SeBVJJwapIENO0/ag7PDUtAiyS/JPm44mug4Xtj9zCW+K0B/dvv8vvudgBZt7+im6a6e2Wr9RvOjh9vjpp8DhfaQY1A/1XH0E48wjk2kV1tVZgN16GJeYruuw0KgK/CGYyjv0MBFqew4qzSA9cDoMQP9ZqFehsHPqmyaRiunJmRfC/8NMAxZeKVgdDfO89dHHaJUITvXPtIUaH3J7qQSfOMTG+agwKRYKGgi4atBFF1ji1poPq2JrofkcdUEAB6IV8fucG9KCtlqD9nSnKdwQoDmKUEHgJJuMJprAa0j3xCAx3//y5roecq5KL4jRD/bH8SHKAFA+2h1pkvw7KniVrgXpYuqPSHS8Qm+Ri5+G7dI9phGi6fpGo1/sJ1xtUhldUj19aL9V2GEZoqZqWz9QkKG486VdUMZ0gGR+YndZ3n3VSpwyvycuvW4PE3xTwrvKS9RKoHejmf06UtPlxYcysW32h3I5ZVx+gskaJ1njxAJp0QXi/6h1aYWkphCjE0KsvqIaBl3DpLvTxIrFqNP2sXkO5nCVzeY942puqREC/GGS1aqaDsAIjBGiGvn0YVoEQoGOfs1ISMBqPtZNVvEcjHTc6qeQVWDV94YEkL9DAcYrCd84+ITtTmt4ORtU58GFOGaNCHKS75STEmtOlVU5dcTKQpG0JzoCtoRUGbavbR8i3GevhN+S/Y3+cDrhjQJCbDPF9TEqV1MiGuwLhE4LGYEjEuGAwzuX1D45igqjiQAfR8Szn8A2UbFf7/c7tNEW4d4OO59oxUecJIgB/IEa5lKfQh7tLRN0enes6PY3fFOKmNa74YiTrzu9p68Q9B3G7Yy3Tih9B8xukfA/5+0dGYRIC47v+KHt1Sh+m8n5B7Ck6LibBWXG5iwNizC6dJv4sSNh05IellVk3yIMJZJt26uYtf25+7vsNDzzW46sQWqQN7UJ31qPCKExM5OP0qpgRutnbKfoPMXAgq2qU0rTyRvbhauPM177f3mq20jR0J3OwKGbv/HOWSxWFPYhCaFgxl8rbrXJXOSx616ItX8mGbi7ZsBMkAb4x+iZ2qfXBR4lwAsZjpsgtM3LYUuSXw82aX6QaG9py/j8qwwUY6VoHpvuE4DkyE0bBU6TtxNDwMH7oSeEgf9zQgnGvXxenvcili+qs58QzVOw1BSGviLxLa/i4plLjhLQhUjM2XtgFjMml0a433y1pM9k6P62iJXCnz04h8xJUVICEI6v2DEdM0CQlwfPDVa2Wha9fq9wt5PXVi5UlTsNrUTfQEw0WEa21OgRlbATy4WEacmhkWlLqrNi8YUwjRoP0BSolFB3STGV71Ehuo074ng0xYFR0f62iODs95mpmOnwxIPCu9JIO2YIOzS4yxZK2hTSQGyrgGiB0r99fosGIc6w4G/fvNpS6N5bL2+L/lawJHp9nPzhkzDsCOVGgBvFwf/WHsnX4h9PkVXLLaZjQ2D3Boq7bREaz3A6T/v2OT2CWQBj7sNv/s3vS+CNjujdWSj9+ZSp0rgpMFJPjT5/yTiJtycbAxPcDd0amkImnGlY4UedmAEGqgkFPt5qunTdrQjUPRytxEskVH5kezS42VoQbxbD8h3oCATFi2sj6g9Y6oJjnFN4JqgXWc5ruAlc3l9O0rN90sfRjXjDucCVKT6ltBydUfDe0/9OtDxfjnZf2zs+2mvPLcdFBdG/1ozWZHjPY2gjHuOFuNalN5XKovG39Gnnqs9ULMLGgj9HiU8KpAw9nSZAKUwOzV+9dCSlDNCjQ6RnwQuAe1V4XF4YGQntrSiFTu8/461cLTvT+aizSbhQK8DE2mp1aId6ltGKbnyGYlE9dcehSBZXmnwDQWWAYfv8ocyoai95Goss+YW8gNsF73ldNBbrpaLWUs11b+cYTiEhtTs+Jm9iI4kdNkRkEcMq4Cu6BAbVW3iBgndi3mp/4309j/LGYUzqL/oYHJfrFQ7yL03LJopktUGn+Jpz0I61pHqzUd7Th9qQVqvZ7ovgCpuAY/2NyR4sYe+gO2FK8hbhdlVMIOrE+4m5h4pgdYRESGgPumoZo3UP4zfVoEG6GaUPO3PyAJRqhngT4PR5EX8R4lv7oBkjcvNvYudyL2LAPE7jtPVWxErhb7EKjxZL+3FObqIvq9ReRdLWGxeXZ+dXzKmVLEV8ipyB8stR4snRK9rrtN8NsDcCL+GXo120LrNMWwPg2DEdsQMSqJSj4sn0Y+S8woOoy3GDEBSysNIwi96ecxmY5stIgU/zNValRm8YYN9dCDkbz7Yhlq66r7bVScz7ct8ciMjLMrL8ILOhYgb0Fxe+1Lj+Ba9+9H+l9OnSjAYyN9z4afQroF9CzQubNwNIBdyOemom6A2oHoL1jSr5vcLMAIR0sKEHgItkB295qujjHphbc54jN4QeJW4VGan4xm3CcdkdJE/1XwiHqmhg6MM86L3puzO5hx1VGYSYTf1ZvnbnjLOrhBH6OT5SIHIj4baPjifxUlEVkUcK1C5xK4GF/EXTZO5SVZx0a0ETy3d8HInqxzw2BXem5WD1aUk24vqc7DirM55lx0y7SvYi2RsiOOKM7A6aS2kTXmd3apvIv23kZiR0A+NdByqn21SunXNC2UNHwknYyGyOluay50vYe41VGCr7FmNChfJLyUH4VfzykIbgZBwYSolrZnPEJ3CgLhx2eb85DhBsbKd4x/eHSIt5fuO+NqXPmXqgTW1MvDpf6z7UCKCsCkahYm8hFpMu+nYuHM8JA0Pn6Er53wLKAlO0bu6fGroEVIMQR9vgetj2mUdhYzmlyOBx0zu4dZUM7CKDFSPmu+s09yLUdzh/pDOcLdB0BgB+mg4mz3av6RxWUDMbox0iuS0Y0y1lO/JntXrY7n7ulivy2wigz9TevCevf0XBIFDewPSkUh/oVPCuku6e1B/L22XxuFGuR9uLu70cxL9df5Z1M8W+gaBRmgtO/TSU/kjPBvfwXtixOs7hg/wXpPHO/HnLprgJIwCPpdc7Fu1SP1MjFRGWCmR1hEe5snm7kjTLid6MDzakFmFYmzMLjaD08ZKPUzXWzpFvKaI/FJxCe31OVpcLfIbfFjrMV3vkOWPZ6FYruadPAmwEFK1/DCZYuuQGn3qTtNlv9bjyJ4VHv+gOunW8rOneAXHcACV2pqkcGPj2ZEuoT9Ug9X6+zFynvFQQzsPwotx07C2Qu7HDNaMkXallhd48tx1By4NrU/U0Igfdo0A4fpRFJNgoCEt0a1gXVunVlSSc8nd1N0TDqXdZNwekrPtXz2quOO9lGK1KVY8fdGxiLTV8gek8lPUX3I10q8Twb5Hzm7HmVQ5yDRGwMQGoSVAV2XGXw3GHLeMNxZjR0GsDELpvB4PNsEk6dbvLnIL5qcy8mlIaWzOi0PRiAATP2sPyYa/6aTnTDzMnsFp4KQPbmKnpqmNdOHjnYbQXEAdr4ogItQ8hma7BeM5VcaGXJyDNWsMWlVFDVKXVzvVHzxFFAPJfSY600rd8bBOgAAMIDhTu8Kh+dSyaVeLNYmo73A+zPnAtt6ZNPixCNm5DAxcA0a/4xJL3IBm/1eUWj+vGHNes/SdPBZIL2iPq+x+p+uRhaf/WqUfsuqNWSU8qDNDxjj5z8bkejRogLkOoawEDQ+b6Za4B01kCJgyPzOJDLbbW9PVNkwD9WlrnR3Qk7S44uhHELK0L99DGp3VMQojkxAdpLmxgCg02OrdFqpC3tYfGxQL/OIMnvW50Xxr2XYG2onuhMoHxV8JTS+B8BmESmbyUoaQNFTh7278e6Btb6Cwd+FUrZCGjz+eFsqN6jrhU7EP5QY7aNvPl1TnmtDownAOnMvGnOOOe1aJpYPZsHCkVQhMKuqk9fJjQ50uG8OQ89Y26Hb5lO5djUMQZofNU2ChVYPX4x625ini66I016sRUrDRCRQ7uri9hpr1sfllB/YxZBp6ay2CtLmqrQbUXYy5AtOhUzReMgdG8PnZNYl2ISzZeWQuv237oCMaqfm4+5rWug3ukgLeF9Sloc4lK0/L2W3LxqbY652Xal/KBeksLDvIbqLNgPOyK5BhUmllzEyRKKXpzz+Iel47+/4GzIQ7wyRRNRDCNSO9bSjS9zQx7pyC4SkNq7EDiftfv5lKDWwXI6vlU9kg60Q3MlPN79KbkhBNVu51ZHUlOjkyKgWI/LrGhcU/isyU6DeQIOYOJIF8AWVi6nuMkOw6LehaQe2aNepBZPqgcswvFtTv/j+kISbYiLL4+85vrPisBN8CL9kP6U6lzMeZ325vmRBnui8tF8KpFYKZDUAaH1kIlquN9/LeZEcO3CyQQKiZ9tMfH5Z4nS6QPwzMqaK/yI57f5nbrGHt1F/TUeMDYVxANtpqYbDvOG2mFyzQBE9G0my3R0xBDyAdufY0Jwqvm+jA8qQrhWTj4uTy9Apg8ihyRJZVwhFS4syqoQFfSHbVEh9Kmkg4u0qt5kTGztNwSgyhiv78h53Ipu6P1axBrq1mISjYcZbHpj0vwBOIQ1sdDspBMAokkaG/8cN/X5SNe3cWE6Uld9pExGYh5lbDFIOVWlUm6K2OVj4TibVYsEzqQ+XHZYgllZr39iTmKmQSxoxbtUGtzJnuXL9bQvrHT30cE59P9mX/lywGr+ooWSQ46TZqtCPvHjSdKjsAXX7qxwnT539jLwWTCQxQI5WFBdc7jmEtwM6r5C5NlBxsE8w2fxT8kRb8bu9RlEB6LvNAIRnu2VYtVaKUQsoDtsSdGEatiT69Um9GOKpy7yQV3Bxow0ddfMNSrh7uDt7DzlztHHAgmYMDjIl+eFfqfWuVpohOFQzc+cSkzzr0E64pWTz7lqd9A1FOPkGQo+hkLoxpw6cAQR2X7NUeR9vpYKfjQd+QUbkBgh1wLLJ0x/h01aVcp/g2svR5wryeuEazAy5NybKwBaftL/qfWHeHgFHWv2D60043VENo1O+xBA3xpiYoYFvccc2EBqPLf0FKxM1yBz3v09vyVtl5EtYo6pRxiDZ3Opyyn4ijc8v4GeY7XZohg6T1TAE0BzQ+B51zkWzpzUx/In6S53XV3j0xZK5KNASI2GCBDCcBSUZGR/nsotam5tT56dExW0dFdPbaGNhABEare7W1gLnPYYWMSnuCYLwAMGSVAN5MORq5pDes+chRvSAIr1IzvCovoz7Xs1xZwmrR2awBhNU6HrKlInbKvKtjrCgEXm9WV+QtHxy6QsbsOfh98nD7QwP9VrCeZdsxtzZoHPrSSxleUx0/evNGM7HImi7/1QasAGDictRsI/Nyb67grSt3opzF4p6Lc0cClIcObCdr4IUTCdRvVojez5HOgmShSkc4Ig78iOFyo1WrIn8OloV3H5VYl8iQdNGOeDU9VGbpRi8upZVYF6uraRt/QCyh1zsRX39OCPfVBMGmWUh7bkGhulsEav5K9rE4cUC5431lQI71tlgqfoLsZCB3LsfZ+MES1RhbqF9k3M+WTMsO4LKBruiAh6gyy6WiJ3vC6cen616y+OotfhrW+zrzuswKjkL7xiOeRaPJE3eRSpjy/YOJnTzgrZelC88OpfrmJnStYShdxjZMtzc/Eu8ugZ3HiP9sS8yEtJJ0iSr6r8AE9vEtyL5FXibKh3Wg4zeTVnOJgTY5hCWL0qjE2SmXC4jFmJwubSLOD1Ytz4zrILhxZxpsT9fT9qiHbUpoq5VlS2jTiQHsI6tTH/YZioRjLx8PsUpxAOVY/oX0N+vHQPVB4s13qkRT47fEKghwzbgB+egypazk8TI60+ZQrxZ0Wt1Yga5wyOEaTbs+DJnNG1n1o6hy4NB9jSIg3KsKy4LKPrmBptxVcRRZXksvvERGxZU5R4juRwkgqyxKUevzirR/rHAwHLST4y9TYG2c/QjNUMEfb++0dfNVi3OLiR/oRiONU94X+qXLCJ5aSYbCvTuib400T8SVrz195gALS2moDujxHrgq7AX/8wZoeyCD+vsZ3vuZL8HF6omQpcgxaS9M+lCUpvkaTRoE+FeHNTdF/TFNUuH4aOjMxECWFoxVknFHrNgivQzKqcZ7pvWEASI1Q+rXkbgEFO6c6CGF/OI6FC7yosIBtbPxllo3JT/G4GuKUo3YlbN+HDUhJ1TVw+OPLpOTDpVuN+64oBXfBAKzbewW1GzSDgJh9CQwh9Eg/mlfOghsV/zfanxfO6OKGpUjtqBO9DoqxO0SjLLuTqMsTOD/RRWHrQt7AoIUXPLxtIUjJbpOHzd1S/19n6uVsS2imCERRY8/m6iomURWr1E+AXuGEYtK4zds6pcQm9aQrKlc0C44TRVMmu0k+Q8q+Nc4ZeCs+33STZLvH3wSlXzZifpsUYFn1hm8IvFU+7vlrj9c9p68q9Yk5Z09hE0BajLr/2ynQNH6vx3smj08eLCkYKi2VAarX3TDGjyGgqN9KLHFyq5VHY3iuTNUq0+BJ3kQX1w2qjiel2DMXVYRoUWvArAghHKYxPJVrhLoTwAesuOt/ez4ZG6ryeb706B6Gjo/kLU6qRo3VageJC6CB6XUfpT1LCYt64GINA8ZSTk2ls8GnF+YYeiXFpzCmpDSkRTm/jCW5Z1T6+waZ0Kdo5cMhLnM1Egp9NYaDPuBircwOOvF0KfmD6OjmfI2J+nBS3xaD423SnQk8KkCHQz//BPGuaabFWBSrvCG0QGEljHVAvL6TsPTbf9qkWB149U2fRO1A+5tsqSpdyN7Ms5NUANM7b2FnG3e1/lwBKlz2F/uaj+jKNCtSmz/9igVOAUTdqtAnW57P85dXuveeWVv0gEDpXN+feseEl7ZLrh9R3zozM/7Unt8VTOuVXkiAUvYlktX4qwZZW4qLa7zhprXtEK1eKNLTi6K+WHJfy8hvqLt8StioWYqBffZ/MNAqY7rCSE8UmmmcxWnAVnM1GUaWQkCHVlKWLHnqhSv0fNncntVd1/tNQ/8o+4DNi3Gr9XIErpfsDsJHzNLewsHMrHY8lawcJMvBx4G+Neugw3MYy7WycNlKPO7EVrU6bm37PvPkx/EpfJrm5qeokEUARe9iBjJrk9lwOFs8E7hy1OCrWOcGov6TY9W1GdbEaLWoikiN7zaQCySdD9mgrQIVHtVkj7MvZFdn6HuWMeSh29didU1XDJzvXbCS4HpcF5tgZHPwU7XRH0rDw18M3cewUYPupifGluK8BERDoJl07cYf1XbjNOjuyr77rSg1FCpjmayOSP1E+/fYA8sElEtNpnzqPVDHjXI3BlJBSJN4nwP/a2xiMVeD+Dy+/rfqFlXvvgy5YYeQIXfeYdWj1gUEZhOJxsAuvw2DpuDqlFFB8OcAz9NWmywvNoOidqjx15T6CgjG7OfEsC0WAIpXD+hFfZLNQ2kdKdbzSSZYccE8T/GHmtG3YQyXau9/X9xCEKq+RxzPe/s5CUyWqnuLTYSi3xEpPELwjA8wZC/SOLRFXVJVTZ3QPQO1nDWjZ0nW12jBf/hg7TQSQ0tSOUAuIgeHofVOJDsFy9w+e2IxAMerhHq6KY2D5WthOFCW3IglPY4goyd3oIMcc6v8RJnbBPdLcWBEx6Tu82SFqP/6APus9Q1feH3DsSkG86gU6Qcuo9jDB9Le5GS+ibDZO8Rhk6wtmv2s4yF9YDEunEK/AWbCKzjQZln5zM536CmAGfJVylawxnBZmuATb0YPMxSbS4KBHt+DJdUAlXDz1VLim5/4NrTaMk7huc7t0p97Ja4lAFK4E/8Oe5x6+C7refQXOEbx96M7qfZhL9DvF2ovebVbFSuG3M3q9crQJH+kEPx1fAquU/7pd00eAxBRzu2cDsS8amPQTNAAW4/JA3J2eppQ40E3uctHC6EmexPvcN8+bOgUzr0WVeQaKP/8qgl3SE+xQYNqNyqoPBmT3GFNE9tVeqpr3LPOjue6WAHgUNxUR/ZsgpcWHMihsH6zOb+QAgCZzpCPXH8yCcTIHVui1HkaTKoxxT3yTeuMvEldsCEPlJ5TxPEayxxBILy3UNpqcpJeIqUyNaiSAwL0Oie7vF5IOK8/TB8HVTDY0dt4lx43W4xehHxEe6QHsZY1LyV6c6HZzf50BnQqQkI9uhiZOUdxqwjxVz/mKINzTJiYRisidmL+UPi5jy7IM+204yF4z3EbXPMPOXNuk4YASyg9Hp9GaJ02IOBRPNz725VUxJokFKQyXR0BZQzsJe8Aeb4zAF304uHpBG3b4Gyq8u9l/qk8SusOeeq1B0dWGQWHLbFJbnujiThiUz5FO55QHit7p3NTugEg7b+9HgG/XQsAO6F/nj5t3hOcVsIvYHt/kLe9gnQ02Z+KK+QZ8HoX6w0TYx2BKfV5EbBMafu1T5PnC5de4Uc7weh/FyCQZrLcxd4xKv1NuLMhd3hEvWZ0zsaFF1Ihdf5KsZ/53eaMg20+PvfR3k8nnBKYcsBnJybw7h634FQVIJPBsRtLTfdcCU6BK6buPYaH6K37fDhfi+E1sa8e1Aq6PPafJvBCdhJmESeXfnR+myUhyxDBN6kxDEL8NwFYS6hM8rqx3x/t4qdzwU09IbxLkH6tnSmfZCxpbv1uk8giZF8CAmGSC85vxDopl1ZCGUlI/9cJoDGzLKr6YJV0Sz2vcOELLQ/JZDtF2+twIqpo7Drx4auK9p6zkyikYTRnBazx6mDWLtWozqkCnj3mlJ2KfUmGuFDe9e+bmTviY/5ET10j1nmS4HHi49f7Czg8BweZj7a3O+Hj6l0ZW/fJODTEdek5HtGG4m8HQv4oPgIMtNcYCuj9yAn+07mYJn6DnVdH14Y7hWlWRAF+Nw/BXfDeN3rxWjMejwSJrcLIoGfR1f0a/EVtROIQ8jAo08zwzxtTaffuasW7fLyIFZw1ar6Dj5Uv8o1a6qBWX0YreLVwhWjSCFCUXKqZWjcs/fJqr2X/b6IqfeZgPRaUv9tzhn5DOUVq3BJw1/3kY8uQEIDpQS5or/iSEiDpO6c1plDF22B1CHVhPJJZtZRyzts+GkxqCkkjPLHWhobHZ7kZyu9yqZh7Q42lKEzqvMhPpnUPDnYEDVPCqEtJ9fqk6OTJuRJEcwhir4tN9Y0uG2XTFBCONsTU7r7V6VD0uVCWvhXvvL1GBpVE9zJLIKiT5f8LNjkHnApJuCW7/zuy5ueO5SHyZ46/7HT3Ly+GECG3TVw1RglEfFIcx7U/xHneyNQOlypJuGioBfoAZzj0dc6MVuXvTDkLuQt49zf9l4j1z1i3sjDIDBF9olRjh8hepO6xCvyh/TcfwU3MpCcqVuwHrbyPeSKctRAPdu9zRTeNAVuHz3H6TH/0UJS6Ab5YI9WtmWWNGJozvWyaIf+d+nKLPwH/A1mTeZY3FFjUfDT5bHaIipy31Z/2Xoka87BMh+CKabAKLDVgSTLizczxntHOp4Lqg2GOcPcBrM2Ogq8Go85Z5+i92N3O/ZAzm7lJLWg8TdytEGhGIgOpnNAlZAp8JC9N7QOs55YE2/RXhoUR3pD762ZQSdlaA6D+RFsNMgXSJUYVrQI2rwRGwRt/lBQ+JB5nAyo4N/Tv7z/7o0C2e11PV5CmndanifRofqsstiD2aacsfjnrdkbTqdGRYm2SdKGUvc9RviTXl4NxGkYjy55XmJBpsSnfFug41OjGOM0s4CyJwgpXLtX+HiqkVQQ51hPJlsHwE9+9V24+iUc0Pp+4J9Ipfh9zhMFYPeC/dVtKJFYlohh8jiGtB9m9di03lXQOtLPnazw61s/BRZx3C7+oRbOIv/5x7893ebxTX9slNJs57Lb11OxwA4cMNVsniD7dRHgunl+inpFEp6W5GckuXbLgpi9dtII+sSCYcONoCkEsEvwS5PkT9Mw/KUQROMs1iZZGKVwnZaMQWpt00ZJ6I8moeBTb1giED6pwtukeMSoG14Hl9aMSAg2AZ4eOwZYKWhEdYiZQfBi/6q2LG5Y4gyfEa9MlY660jf/i9DM8JNjlHpgve82Vr6vG3sMvl26O6zSdOxn9FGYN8WESehIaUXX+yI4QGVB3tYs5m3QFOt3SBr9dftP4ZhF5hasW6jlrJqFj6WqYXzM1MH3alv7g/VVaE7Lb2rz+l26CWhewNa0aZfAjnmS/Sz3fZJP376NnLBENCtVlUfo1ldjhmWsmFuYYbp5l8/c3aNgI7xdC+XkFHf9bDfJC+sHrMRfHBI8S5ylwihEHx8M8YOhsQv9CkGcPmTup7JwMtGN4P/QJPjQ5kJVWWH2dCze2az0Er0CWDf7i+V/YIDWJxs3aRY3HP712txuY1BC9SRKu3D7iv5s0tquN5RYJBi1Y4Yv79gWyQfRwhZxAHbw6WCsHi9yqO8E+Z3a06V4sy4twLwcL1dctpYEt/TYI/j6sY0m/17NWcJfnr6CQ1CxPHWdqKArxNaGXMdT24gl26vASyHh5qJgkC7qwUmCiyYtQ0oaXgoUzJBAPwiq+AFkjpvCJlE2zpU4VTCWUY9HZwqj3UA0+S6HnvA9xJFS8fjKaeNqdwp4R/3vT7Vm4K2sRxexT4AoA/ca51W4f+eqTk0xzY52zxJCtGZZ5weNQ1IAr3PxvrjolmzPot2IYGZqTpMAp6eSAqg0kZEt8dYI3ZyIghmFK2Tu+Gd4ymm14y3OCoKreUS5nK37lP2YZi9gFf2dKQwPlaCl423PVQSTItyu+PWXMSmGx5dEc4eduFSXdwK7MdV5H1bx69cIN4zAFEI47KOpH6iMsCoD6B0kaId4uBfAN4H3k//jA0qD/FsgDH5nZWa8kN5XCZAMpZj24G48ziNG2EFfh6ypo+LsWsmBjBdkD9OzKHTqGuu94K7ekCV5F2RSTXWYpUO1tV6vhvd76oX6C7VDOOlMNqFul5YPOvo4TDyKA6Ns+N9YzrXtg6tFFCFJjaAoiTrD41jdXWJLk971kx0CTDZF+D1PnHLIWridzmNr+WHr79GFHaw9+8oHr6gFW9CyqXpHEQS0uhgXNMzp12Tmp0LqNnRDOb5QpYSxWA+nzfwnbFC5veE6r2AQEn2Zdmq71WObKlyliJ+T0SNvdnroX6bAwoOk424ZJUSDEyo0I7V9uetmb59HwMx9rTumCn02GXBfbt0fqiu1yFZ7HWlZ28P/+nlJcR31uO2Civ8ozaoitkLK2j4N5azmUxGb+zaD5/ogq40xg0gklDAkojwHIABcgprn8Gy97yca9VPfMuhZmwIbMOqLG5cw1UAuC7MWPc/tY4TOXlkAU1XmQMhYgyM/kyr5Q3W0er8edAhSMIVGeFY02M+YlEqvrdHt2xM3d5+xi22unsOWiVxZ0Gx8D6RB6nJvAtUvTfv1pVXpegLlZN/qDYVkOx94rTt5TZXJ51gsxB4xFQzCknpTzyss6mOey8bFXmmCBP6qXLnprHbojo/P2Uws7FAAi/hwkhd9okwZssxKJg1qCbRviGLU1975Vb0XKiqdU+HoOhZk6L+lozVxBdRx9A6tDTpGejhlSpEF94/dMgPm9rhJWwToGngnyB0jj4s4VrZVkaEng+eD12Enjy3zTmiLysSkkeyu7guSqBzDLwDDRDSwl9/fsCWV3ZsBdI6P58/ewGZhUZilBrhn/bB7gWVGyWbwQRUHpXeN21Di/Ap5ESceL15Z7aol+Pr0J7ShZ0UZDgxvRZ+4Xv5pGeXI+OKOHzVLmYRQRYy36N9LisPYzBsr9MSW6Roq1nhSbTVee1cK6834hxuOIAfjloaWqhZzH9ipC9297bREo+ynWTkTaOKSz17cybyHwsiHqRxCiczjPj5HmRnC61eS0I7Om3bqwNjCNIek1QOjBFWEgVjm5SRFQDt2P0Alnjle9hIp9C4wj8iqPc618Xu6wCFEl7LfTtU2MR8v4UUpSuSKCJRFBXi3Nb/EL0fcgwWcgEuZzQ2H3GdmBhbFkcm/HMwAWELiMCn999H8GK9IRJdaXgSbKqvR+KdjEo44S/kILahVfiL7JV6dyjQ3cIFxFBk4Vq7meGxKefk2m8oA6C/aBEly9sF1Zkhcdu1fZwHffIUzwm/vxGZWvqaaWWl6G+kACMcN8BJzKhx7cQGZoM3qG1WeSwClpWy5bUy4anRRQ1fNCStnapYmUZN0ErPl2YRc+8fNXlpTYX8u6yfKY21id6wvZPdHISAboXZlG6z/oth3y1X5vBtgEQb0cNHhshb8GMR4rXyFvT0j8tg0JIdJyEWq87CfbGtdbagfRmf9O8YYwzDfd+s8GKd7frDprLCqcOpP7soiRNzOGlyUOHS1iWbf0/mk7z+bAXD/2f45zTIFT8KBNayhvl2lMmbNtvjvwJqQXgJvRYvGdVteahkZxYLYBaDndY2I0vflF9jXOjHpFnj4XP7+2pYShCfRTAz94DdMmdQcQhR52vIXEXLJTWZfbqLSxKwbi3o65MDCXSGVN7xWJMfETLq90nLv6E4QxSIWryK4ZxwxbzQ61x8gMQb0sBypakdRK9+LJHoCoXHwfkSDby7nOTf+SF9y+6jPtMt2e5+Xq8ciX+DO4BMJ1NIVX+50WLEUYzI5oKy502/Ey4zEdSditdP575DivdymVm3weCdSOJBOya74AkgqQbcXwOsyOGgQAJNh9f+AFWVekZGS9a7qQxABhVXQDKcI0X62f+9bNGtL8jhaY0ZU4u/HrbsN0/bkt0ZVTn01zXCny8KLPaPk7LNVC31fKmvl/HcEbp/acotX4CvFD8dpllmheOJKb/K3yL/hm1c7ba3pltfvv9H1UmqXT3uIkwmQLC9rLB4LN4iX3BM/cct2rGj0LMemoieyXKsO6wX8iMO5/A+dMDgVvcTH77qjG60LXYxWAmpP6fNqvxEFiarm0Gm9V1ghCpwM6F1dt/9kAANlZWn+ikrprTjzdoQRQAJ6NEgGd+NMCnoWzRoUHfvCix32PrhIqsbUJy7SjKQndb2ODll28SVwqfl6E4YFVlugp7E29hfB69Iz+goWsc+sJlbDxgPNI5QhJjc7U/CxZVhtGnZZ/VRj48FXvY3H0XCjoOWlA1cdOdBE9FfA+iottixsGWjLjwk8k6p8kZHzAX8vKBxqy9i8jzpjLKKbLiCfVK00VNpzho+P+ZyzhRdlfV3dfOsLQvuc2k8BfM4WBAx/eLA9RmWFUoHjgUrgWinTkTWCcLRFPNfPkDqFLjCuypZI8lwxu3/0FCzEBne6kFFUdwHg68EXlZOXfCCL+NvqCOW5vUxkksAwJGJhyLLk9ibujLrN546KKfA1MahbMOrdNzx2bGw5ICzzfB8gc8mvBOxAzyHIpNzVN9rnJz2pU6fzSW+F3K6wFvgkuTPHOAvQmHPOCv/ZzVPq4CuQdp/lE+sxIjkWOzq725/yY2O7IrGOVBQWlWMjf62GVAtpIZeAMCF4xXcfjibdFRE1J4XiHs/u6yDi/SVTJxU6ouHg9ZXskQlT2zyJi4e5mg9WVqEqgGLbZBvVkRxV+XsMstg/gfdj1drVBQz+N6fuKRGx1HcXPEOdPZfLxKWvNi61u317f4iTuvBuPb9t/e92LUg8oeXe3O4+Wt5rOLHMGXUn2tZ9+1cxlFndi47TxgguYvevfPQ84jJtrMkAUUvOUWYwgyKF9ZNykpvnbrp0hKTMdbO7A4IGMKOD0BIuVBIO5xu/dLeasVViZTNgfFhYQ1XCUXMwi7xIZ8p3hSrfiAOu2WCHfQKS47x1ljEEoYBIwn5fivF2R7jM3kbTi6A33Mhe5pwHgDbRTWju1kyh7CJK4/q8JkgoH797F26/6JINvCCnIGQ70H/Y3zKRiLC/kw/jX0rqvNyWb9xKr18VXzHOG0g7onp1xiyIh+O00mMY+NYn35uTq3qCpMQQmH+A9h+Pobv982lk7nz6s4PHgGYgxWjmiUR+AqcUg72FGGGj4aE1x+px/3OOFCMO2tySQvlKJmxPk6dbIWOtMF8o6esCZQl66BxljX6KC+MDTw4ba/w9s/oUaJ9IYFqk7ARIufY8wcCULEO/qqbNb9VUuo/T/7CoIO6satm5s0qmCGkkR1Ri8aketqiBcTLXdCWr2gxuzGt0HCcnFfij9tNJdT6kQ+tzo1tKbTxNgmhbDvNMCHpEYxVvbZAnTEfY0qycvC7qRtDrnRqTCuVQ5Fc0Uq/Z15PuldW18iMcuhIuhNVt//RDR2fl6EOG73sjxOAAqiUPLCXSxNdGzKjpex9GrpBMBGxzlKkmSX2FoPzkBxRG3iOLGIqDmalO1Lj9bRocKo6nWlsE4KcxOG2MOU27DiH3oqneuhU/MOzTbxe4oS2hjydj7rXoKtx6U8Q5xX4FRnlI1TMvmeFi7MyhZvooggeRRcLX6DxmD3aisISW4zTAA1iptLNMjPwkD665+2YKlhCO/9X1oErFEJB8DZY0BAQPL+qfsGDePFbiICtktpdyE/l1lOxW9+/8QVxUWgx0S/R1wSoUrLlFjocnisEYseg2IJBilp9Y+9PAcV+YLKf+pqZ7zIpdmQHRTlAR19LbVLHWe/NiiYMRo/0+w08l9na9Ccs3xcHbq+1m+GZ26GaLDDzmVUOINWm2vVFCTRLAt4dSvSnrNTXSFg09+d/L+tQKu1+joj/9cAJACBLYr6pCeRBRmWburqKTMqLPGM93hhZR30beCL7TQPR5WduMISLHrC4j2MjcBpbuX444T06XMpb38BkYyZhCAT2zWuKtS7UHGaRW8KZod6bkSoh+u4ntOz8ODwQuDOW/cNayNHU5RLbB1/zi14HX0I3nodXQENyQIL7CFPs4ZAIErQYkEhExhV+dvNFsu3K9sAwIUkNFsUlCfiTaWg5+1gA2o4tru6CQapO65nxUEaoVRiCQ39r62F4mN1kO82CyjKFvNLw5dw9W/MODQbZ7Yj7/UysYdOK0EuaDkdmMLpBMqLLRzI9W1EdNS74wq94xYVmCzAsgiDVeU63Ezo9Cv8a4iaoNxI8r36ZNcjAfcwww9byUfz0U4U5qcPQPwA9nYYXB4os/Di4NL1NNt9v7oKLPrIVBpOvovx28brL03eWDqgoD4YzuHDx30JFjcApa40r/K7SWccm308tpcDeZgSzTPzteGMOXW6igMMWPRjXQ479O9Vx5x9ogSbnQQ5yNZJG5dngoeiwbxq2iG0TcTM4R3sw8x39Fcsj5jgMByiGzFV46uwhsQQP8UOTD/7T7mR/WcO8oiTSk0noEfwd9pmsvAfyHCF+zfIlkMXAc9eDeC4NkqdF8gLl17Pgj3JoXbmqmf5auQWIRrIWdVNKTorV4m+WPvkd3usKQRC2m2YMlSWwTCU2lXPj54CJ/3/BusoE7t8vU+V8/Fd6rFffZfXtlSG0UWBzlIFYUfPoN4dkGBY1QUwpxxwuIYaPHURuCdWvIunuDxcSzhymm1FztnatjxuLmRvF9OYN0pReDddKOFAL6D5OTN6lUGwvLi8ZR7WrbNrV4+VxOhOmjWCRrlQ4PYvKpmswoU1kPDCWRnKI4/40EdT3t7VufLJly0WZmPES1E2W1aflFHnT5B+B3V90Z9FXqHiFxwImGumBkaOisLnTjdRgdssJD/sCkAVok/m5nhi5co5IfbysfjdN7zDD2rxGBXGC0dRVs0y9sJ1q68/t/5EF0XwezQrpeyIz+JHD/noo9VzqjhtVNlJk/zSFNrtMfWV9xuHIEPRsNruS5cG3r83/ewskMCdPR+wHpkTpcg3L6PnBipt0EFrt/P4h40wnI4R98dSftFmSlb6RRhpS4sSBZ6Yywa804vAvz9A5YfihQk5H/YpeJT9KwZl41JwXx6aDtrHzGS4FNLbQLIi2so+VXuViIJeimsLXRlbelR9yCxUs0dgyeahnejEmOALwNYdQ7juQIKDwJRwW1Xxy1tSC2wgZAYswwTbzTEwxsc1LzsQ47wwQnKQ+VRksS5RytBehjcytBMDHTVULbltUMY7OVV3gsIzfxoiDG9+dEqIw4r0ZLpU95BpMJLv/Z5IX5j0n+IM69aiG9LbQNknJBYeuuJCNfnCa+doehP+ewCmSji44YBBnirqWYj6joK4pt8ItPP8UtH8K7r2Iq4yqMyxPSgfroRZr8+vd4+5xurD4MD+/AhAGzPLbtu5aDLaqJ/tYHtZSHZXj5ZThD8j8YXRg5/x6fVYDzE/4kFkr3dzeJzB+e0vUp+h1X3yUeiWy1rdWLLTSNuCl5jV8RCbovI2foqReQg3spj6zHRWbP4arTO31xqThBhsQP7tBP3NuXJoiZvniB+q4NYSQ+uckhrWA+7pcircb47p5f+y9eAuThPectuvO9MEI0yGCN1wXwJCK2215o3Jn/462J92dTv0m1z3MTTs6UK0xz1olh21QQCuUfj2YvIriSCo7jUR2JgP8GYJUgabtqmn+Q4TW2hEeKdd1gX6e/nHOqNKsKsJc+TDuvp0841HtfsovIy+BEpwCnELkxnFRa34tbzvYjUYQXp0igE/rDKHpkNHx/yunDAOXYa8dcrunVlfbhQ/ktfRMvBH+7rT6WJmLYeO6PlglNzUtZm/GqGhyPxkmcPfne/F7Cm/9aW5U/2rkrlUdxkHoxQn4ESGiuq9/eJjzNj9w3IOEis8JT8mDBU9KJmvoXhGSbEzZemDgA3f8C4DZxds+NsR6mUuutbI+7cUDiMiBExT4lXp7501m6WKDcHm3hMkFvavGjrxMPZbZxhgjIFiaS0fqe3BllwfcZxvf71KJSr7yQKMW3kEiqd55W3889Y1ar56mqWQ6eJAca9urNrHVvF9m+pmxe3+MOlW5KF0wMwy5QUUSouyMtlA5qYmmIv7nGqEFqYnbUMRp/AVwwx55B767mn8WuyILXHePwsh59mBbRuDdCI1ESz1KmnuUw0zYeDCEc/H6G4ypT9afziXQxtCeuXNvp8TXBC7bOoJVD51QRf6T8bCU9aB/Dl7CInNQxw4FWynA2OrHng0SblAPLWSd5n6t6FuFU2IGo0mX6ctUV04ZvzxG31wXfC3yaYWDoGhDomsVqL2IyitdwIJqeZrkjkBJ+Z0SH48MkDFs4UvbofQShOFAyPUFAWCa+OCzmLBwHKSgO25os4NT5aeycgF5lqAk4UV60s61P+XAdv+oQJwmnqmOGLU7QqKJL5qJILXMMCJjIubKWOy3aFrLlJ2A3Q0kLzEQxFXaihZOfaf7Ty0Y3MVTohqo2qb5XQ9Ggn0WBelRZP8ex1qmJYS+KRN1jZscXfSYlkJ89zxopi5rwakTrEF8Z4b/18tdc916aLvfOWMwWi8691KzIwVzfnHGOV16CL6tcAleA1xVRgFUuq6nfklZXa8/3+4Hojtmed/KD2bcC1ggLbd8YS4kbIAFEKesy1jsVKwXf9bfguU9rE8mRKKWsWAlZ3a7BkqoUBzh4oxOO1YyWl7PIYahVnwL4MXYwC6kH+5ui3fk1kq3Qlm5QVyH4xiZgzc/aBngzqRUdCZFm67h4ytSeeLbtLAQNUtGE2G7Rxiyr+qUuWzw7iGZQH09Vsak5exOJN4Nnr6oGI12dAix75/4w1NkUVxIzvt+UtgxoWRFWvTR4etk7GlHpHeFOoEn7nw31qDJKAdHPSmU7mrtywyoybF4ZiZa4GqiEVLXS/0KCgwUZBKJZrIipppSAIFMKSVGrmGMbe3FPbZwxYWGGdopy1Y0RaemFey+xyeACdpnzNaJsoCX0C8kURbjQG3dGtb59N3ycm6feKknkN3qf4M8630KDB4HG/nbW3VUOMFXjK74hEyh7Ibu2MRE3XQ9lHMgKIiNZAsj5c5j/RebSS3Y7bKZCBfKYe8BKiQfDcem91qE2Z2M4dFw7WOSE49L6o5BniBJttC9mBvM2CwGAiLnACk80h9bsSRWSIGHof3UWW2e7c3BQgr1SGzDIr9yBrQiaK2Y3NMHBOPuXDCEkPbZHsvbbRFCAQV0lbQ9ycfYIct2WCT11uACqLAzelfu/jL32vPxSBZMFIvB+FD/H2jtgRyK5TYCQGx28pQcuJXCTiLjiFIvIci/wQGH3m3YFGC9/GZH0ryUNScN3LiL16qmk8/6FrYsjGBf5QB2jHHYpbmRddyvAi7yiKJqQjmPIkymdJZ4Fkf/MDrpJz5rt9iC6ZnkaMrl3UTFghh/jbmopqqCwW/tbl+XKcPPqst6zU131Ifiwg2dvl6uwkSI4U02K4sSTWKfHkJY/JF1/DgtVaAwojtRRoqupoq9VQfZqYcvGz1l4bl6dFDdnqKwRTAK96vI5vs/ePU7STEU4iRB7i+ZJyRXXQ3yljbJJi88ovvRZnqOJALKI39OFR63NZ2Rasll60EblL0CNXlcRvzjuJbmxaeJQGTd8RZDmmp7EJYrrgQ/br3xSX09/DBlbdM5ME3MzMn8sASR/ErJj6HwzTMkF3z+j0I5zA3lH+EeqKTII59FqA//dQ9GhMHf3k2JQJv4/+eiABbml2Z1a7+R1SSH2HvmCE7sKvxyHbYOxH6UuNmuAlsIb0/SnCKOtkkd42VrlqbRxP+tojz/cOkNYU+x8hGE46BfQDntRtEPmQ+ejK1CWpxBBe/b/b63Z2KAtJo/vzBWu9Ic0ujPiz9sjZNNu0IwU7BiS3a90XtJ4KX17ksPFndMKszCSj8GNhpt4qwYF72AwrSZ5GjOPRMZteVcn7HTCXH71QzrpEiRz5bqXYQ6NF7CtlHfYJbVq5RfxgF8xnk5IYVCWENyW57BpQswe6Vyi0+8y+OGj75zxifFkjeo4SucmsCnac4HZ+wBfLhDg/pn/RJtWDIf/Dlwq7tt9yr+XK1Xv5F5Lak+ho3hs3DWJXSIyGEkDWved+922ED6DZbEeM/Y8GsxdbD+KUIppfFY21EhMok6ZDQ58fakPev63gtXNxrf3y6K9twmE3b5DkuSWLBiaaWU+DjcCucaZEDDxuZSrcEskLva2nu6d+WT0m402ABDfSUJmrZd1DsREboVwPM2aUXgXIzequy+e3E5KKC7+SxqzCDY21Fxt2TTk/4pa3g0K0LHgH7+RFk+ESFOqR+7w4hOQG/NH5Y33fB05javJhZEwFclPbovZz5vW57hKSCggYU7+6QnOnyaKgA8Vv1U0BZaJDcrqlDtBhKvEZXKbvLydBCpH1nj35Kjs1S9YCS6j3UhAVW7mWWlVb1tWEqzQjfnEwuF0TP9d8cDwp3vNn4TFNpdTpmG4rKCjIt8E6Yxp6Okn8jDZ27xMwSEGqM/O/Z0Tq08TfpSk5hAEScNFm3xVge2rvaasdRsWjMRI18MQz2MeTQU7MyVRFZ+cPDATa8PcFteOoDPRYCZu5SLrWmsB9Ua2rK4VsroNSuOPq/0JLT18gay+/gmQ1oAc8JFLrHjebNxbUx4uGeDbkvmNIFQ8lmPZCjl/tqMNOS//QlJd+0j3fSKefMHubVGfxPbyJcFXHl8pRWVCKbC0zqY2TKanBA=
`pragma protect end_data_block
`pragma protect digest_block
5f4beec63dbd83352e67403f9f46c593839b5b0352fe1032c2eb2f7cd7bfa522
`pragma protect end_digest_block
`pragma protect end_protected
