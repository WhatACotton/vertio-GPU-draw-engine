`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
pKvqK5JE/DeUUo9JUQF4bKutTLMfaUbC+Yw69BwA3Epiyds3AXwbUmci93webaKGd5SGeKe1CaCEUURF+H4VaTb265XdgMd9M+K66dRE0Z7KbyYpJHYigv2TE2/MRBepNKIosllM7kdsQegx0jbPDUkfXjjx9AQUcl4VlT5BB62QjmyhN9DSCoUJ/PtxKoXd6wZHU3aGd9wl855qaMCXKwe339Bu/VOU7MfUo3IH3JDqKeuqUlDFi4IhVGIkAYGVsfnIS1O2/5KueSlR+PUA+YE1SR27QVQAZ6GkSpfOft5GVOdQGwhCyqFzU3XSXYrPaGXQH5S0Do/r0BvdlEW4piVzmDtmKyrFkNG9FxY/L7oi5+hopNw7ia3XS9JLeqjgj3ZEQeBi/4ahOY6LW/NUz41lFfi72ooqFFeDJl9sp0XNs8FWhJFvwS/fQuXkEre/kqV1TYXgYc8scmwe02SXxniQKkwHTt/XzLz02U++IqVjwRbGGP6c69gpwoyt0HI+iYuT88ZAjKzjHYFhIf/6C6Gy3NXD010kiBCuo3lpfXK4ofr6OivVzPo0WKcpkzEzw2Gxco5bQnOmxIR15Rm9bKavzKfT5qn8p+KKypGImGWn4P+kUg6eGaBNHC8Zaii4Ye8/+4MzyMO6Z85YcFujesWNiFy+rsTjOp+aFYBRO2Lwq4/wlEsCUZdE8dRqbhGUjzXuAmlQCmBAVTH6LpGGTRnVZr+8JiE2PZqMHVprE5cnv6XuRR6eLLXhZbr8GnUgMVwi/FIot4oaQfzH+6VMDeZuHCzPk1wNC4lCBqzv6cgMNPsnH3CIReeLbBUKTr9vrH7ToZjW9eQKI7yo+cZe3ge9ARf6g/NEBgGhG0XlHsPhMokQT7GU29H5uL8vcIONxssUA2ikYS1wjf7vJ2Gara97Bw5HhfureF2+KTgGougW+Zdo0dGCJH/V+Pn5sgJp74ZY9PaetWRbqfFDk27qCvUWxF/xcy5hhZ6NUnAAUdHo3+4CzzAvqXwfCfnoB+gIQsUjxR5tGoJi3tfQBfN1bmcERs1LXCPg9lLublWp+H+MI3ZjKmb/6HnNrFoEq3uFAC0nG37FPm9g3UgbGxU/oF33n3Fm4IJApg0rJdgwyXmGOZ7H3iXfgij85Of39BNa1QOTogrKQoDyXHDmXOZ5FEiJFvcYS1bnkbIBDo/vtCSM0pHQ3MukHQHmwNdOwyvzWaAGRhskUmcUvr7aXxgTI+jtPDy/3KOckHE26wcd11fE+4f8zY3FWubKByG8eqpTX0n+G1BB49qudEVst6Fok4dt4wy9qG/BT51jY5xhLSC/npIRp/70Q4hcW5s8F25FS0T19o77cNdTPHEOrm4QQTUFbKh36z0rL/swHpfuGTcIDDqrXYF/QLULYDWdwF8TxumauamYJodabeYiIB+Brnfmsw6Sacs/EjivMUzCMUIyWJvQd4/kd3huixQgvo5fr+6BcdrsZ31VQjiQuA2/xkgRaaUYSp+8LwnrzJF71Y60KpPMC9mNGykQKvb8Oxz6eq6kVVtxDxEJ5IvZj/lT5/DfoYGB/EB2TA1clF6CBVcT0PUeLQxx7nKxIkstEpk41v4usrqoMHI8nqLF8es1qbJQau1BkXhi/jlk31wyfIIUXGK1Im+fcEooNS8F0sBzHtA5KjLFRW2t0ZQbjlPiXgPF/srfT1qcViCkMFGXbwizMHoQmIayAZBhKO7+zVmtsbMUjYuXjlue8Tg3ByWP6EwO62t8LrwzTVxcYfOXdZ5VqXdnefKwhr3vhFiv7S8UrXLjhY3bqJiihNpbkQR/Hvv7G17kNpT/ewDfRD08lXgZJotrAysAOJvtLJPefj+CCuiU53IitFZ5Hj4WB2nKxJpxwb2lYERq4OMCC5PvZMSe6vg0PnVyhN/7AFSgKBqtfswEhCkpE0WIKMt/zg2Fhto3okxYgyEAJMB2A6aE91Mz7w/srt9FtI05qUz3/2bNQVaPLaGS5OUHANBe8u+5lHq8rbVlTHPiw/hatjz9QpuA14N15afbLNxGgLhFn5LI2hNs+a/5SgaOfZbnwSunVmBW1tCLBS60OHtlwwEoGc8MPbX9A3Wkpr9Vu0i8rB0Odac26L05aQdCcu6wFszdVrlJSaEVfbqexOV7gmR5TCzmun/BSueoYA85a5EgKPVwzJZ3hC3aeDJ2HhSzw1Scmfg5/S3gUh9svbH8/aQ8IOxPpFJo3xAFFo+s8EohYMjmcJ1zj+SQ3mbSdY3n9Ava4BZ0KZN6mbqlvjxSPuSWNbsM1kpgrBHkliQs2ZwE9EhgM30I+qEB1Vl1GWhWKBXnylqnRZFx10IeGKIioMWsSky6vC56JiAs3o9T/tvsBHKZ41/QE/MapUzZjM+0rHM3gHdBjggxWjxLL+tAxIsf2GyIsA/jhZ+Mx+wZpcz3ZVWD4Fdxhb1jdCPajM5CPqbVi/Icu+9xqwU4eY1aJP3UmUqjb/ccGy4G1h5nb/B+CLYfUftNcx9ncdP/14w2qEHak/mdvBlCnjwAhfjve++c7ko2rRdRc7ZupvaxKDogwMHzQJS3uIf51pRfw6EifNJWiCcO3DxQPrKj+oxTOqKc8Gc8Z+rImb/ufDjBXJ9dMfdZwWPmWqHqu8iVYIK9bu6M+Ef1pLuZihmXPOMObaVUDG3b6YSWcREVhiupb4IC9McujShO8ROzBcPNaUO3xsCxRbrVtKoQBsy82kxHxyt0AjtYjQPO+8sR5x2gW8wVV7P2rl3a7/zgilLrWt7jLh3jpyYlTYvX6XJtoB4e7fz8dApxUDkt9Lmgy/EwEB9bp7xUhqHMkFrkvXATyNv9fWdQMM51MWEwYpNWjtjZ3JKnL2/FhqIF73QUQDKpY3Lu8MVJy1JwUFSdznyv9/1X2lby0dXo87PgdsojU7L9EozTofY+e13225z5o2MrznOJXxAKm6OAsK9PDJtDWQSzs7Kw30jcSbIF8kh2E0EcUjAbp+eWDUBsYDNqpe8ZaiAc1OM53ry+5DcP0QNWvdQsVSV39b2nU6CbhZTIsR6nm158QHPtRDcxg0+HoBrUyiuMXcW8hi6m6uWTTob6vSMrIsjvB9GrhVZWF93F8myW3dg4Ia2M3nPukk0QcQ9JLPKHIXO20rLljMgiII6IRQ8t8R32W/an2/jTlizeG0RqrEfrLfqc9q6ArYujx0GOCj0G7Q+6yO+ksCiL7wd2y3TekfJww1Cs9iGpf3mdnf33UqbCceRPaltAKoNwBJ5lvGnKrmEb5mXdsSPBGOdVpDBDIq+eBhJJYT7htO6s8p/KSnk7f34sECFbeCwJTUFc4lelUHbKcJe2OS8w3+wcA1CsiETdCZn4MSkbg3h/22IQcuzvxdIlBHjFxLV426oPddA6qy8sZy+99BmGxoLi2Ej60+o6HrGLIZLh7BdG7T+EuJJXBpR/SSAZnge2PAwXRjjF40p2D864PrXGxFq1GQHUdY2YWmlBbWTxU1Wv+IgR23E7E93mrK5xfgA2SYcX6r4O/Uw84ffIZkP5lKTe/PSTP1tEnwJLgx67ylgaca0E16dCdBGQZlO6iFC6ohXeYilv6G2+Zct+EsQFuAE+sq60XpKeyS/TVQwdtqHZ3zB7yGfuijbDf6ieB/IpQsZIE9gZk5VGcqxG+NeYa048j8iViMIZOGHWQppNknpixMvQo89UqsQKfAWVDH//IXlWAsz3oqmSEukL8QLmd3d2rvpXX6HTroHfdY5fSXZ2/kQw45RzNturKlxF9dPy5m51AzBaT7TJBp2PmqDVUZpZ4BIxD0vrulpUYVE6zWe5lpfgTDeNE8Vlckak0mL4EijHtj2ibfFN0VYGOLV7hjMm0Sfmu/U8AuCIWF95FhQTIuOW/p5BKwqAiAIX03GGQ7tl0pcn59v53zLcLpVKICBYXc3PFfPijpdA20TzqikKTJs3JcUpvVZt3Z2+o+l5l8ZKLvo/lLkBg+pQGBfRtRB+QxCnr7n5BZa0C6Nnz1nEAKmnMxdrBNSu6v66C5VrhBJ48i6Q8syUm0IueGzKvT+4CFkgqVWFcSczulbl4d49eJtYh8gKjI1V3bfg3K/spPivPC83k4dktKM918Xpyivo1ve3eNWcrtX9Tql+U3aL6/t7grCPp4pt09T1+Go1b3xJm1ywnoujXvPt0IEEByqqxuTuAZcLN+0VazvJr7im04eldyZIRVR82l3oiSLqyOS+X59crtacmmm6xQIwBvaLaQHKWBhbH9Aky3s3MkFOO0UMrV1o4E/7VjhvWwnwYvTDg/TFkxDDPB6BiYMnK1H4z3nf3VOhhXFEPqr3W9j8hRempeBhhYNxgwZ2QHTwmjI8Oxxqa/q1fydSQVA+CbCYtzGti5bVo3JCr7U6nsmzVaFy4c1zU90UQQ91x5RL8vvkFonekmTpjvsnDSQ4aXimQ5fknOtOcKFJcRXTp4MggCJ7VVgffFdYJSRb/D+ZTfUOLmCyksoaRcV+pI7m+BqJMaM8nIV8YKO2DIGuIqXUXTzZefCPbAIFtjoymfS/0KFjSPv0z9Awsjd1/5uAp8x7mdwyPqGLRHvIRR3bv5R/Q3a52xo931Do0MyqN4RdrZYYrKCj0A3/nJi8ElRumTrZZ8qfuI6i222ZahvtvGUvjObqf26OHjw+wi/Zf3VE7brKOm3xtQJ65ZDIScybm0SafgjGhHIg04bwjUSz/46wfR/o9gutYs18yed8xJ5OnxRt0tTM4XvwC7LWMNliPXw/72ue5AB9FAFN1NOc+h095HAMwxpMmDgN/P+/87l6F1A7HS0U3mo0pnfVq4Xh8H2VA38j8SE4kBvZEJorfVhBXFenhSr8zLMJWRyKb0QFBQUCECbAyyGyo/oHuHi3kAufSb6ZNeh74IUJ6UGUk3g2cv9ufLe32HLtWlZ+mXGxzhT/FiHbvRjWx8akzOrdh+aTosMF7wL1pdotZVemjFBqk/yN/F2ENtFjSoVQGEb9vVjAdvqM24lJyqhwSfvTc80t1evPpQ4wuZcY29Pg/qatotb6HmqO27vCEXMVT65pFkG4owKnFfXJV6+las2HVKVP6IRljLNhH2gHDUE29DVw24zBKFFrpzhEuhslYoZHahF7lF0rIKeBVbiOP7ISKTAeQx6BD6tgAIryZIpV1qH/7oeQbLfDHi3tWQjk7yulirOsUWngws4UM11eetPF9+qK66T0b9JPzlBlmkUTkr7GAXhp4hmgWp4IfgdUjmtZM5hhVWtYEDaYoQqRbebZFe7QgtuheOxDB/7EwFfdsQmzG3qvVXC+nnWZvmIjFU97PKgEaC5alcWOJvtDifJgE8ICJIxHdgvrJ+DH66Dr8J/B3LK9zUD7VK+gZoZxMsVF62tpdotdJAXZ5PWIaUcyo9C3HyLPb2fJ+xf5U2ojqUtfl0+oRIZTnuwzYap556/qjeAJ6aZS0frm/irZF1iPX+jb79AUzBPNkXZsrBItOTIfupB+94F8x8nIGAtr9KCkW7hFkk12nufJQudsBtMeAsTmSGUikmBeiLLmaz/Fu3Cc9Fazwmv6IR0j56VwxBYmQE6ApK7/Ch6/ozpkSkuMNPIUZaXwq6BpOtl95okIPla1/DJ9XVjw6oi3m/s25sbC0zu92ocZMGYR3W75EMelVYrxk+hfZbSXD8qwfYQq58cZfKQKFqVX2GaeJ0KC7MS3Sfwpu6j8uqlPO0t13/K8SzQSK/S2EP827IPAVWIsldE9KbQBMF1SKe00gdS4+HgsV22rg/IPH+qU68YcYydPhXiIfT0r5PMKcKmlYflGetKk1X1IShqetIdGwlkZkuRWwxDT0/JiielYr0jhsoCHgiNjevIOoVNfLr0XNs/tLdM7q8Dji2LmIw3PJJ4GBoZ7TQR0gFhuVehx+jqSae5ZRXPan5ObjLubDQwjbBTcVuQZEoJ9KYmfcr9iq425q9N0bYXNDIg8okX+Oky7ff50H3vjpysajB78dYgOoXzUCoqRqvv4kV4Qm7kMvWowGaRwuhT1FuxvtSz5yrhAnTjX6TnF+s1udjZLIPjerGzy4vtcpBD6tx+TllhcMcfYxWl5RQ9t5M2zB2Da4GCFdMZqbcIuQiLxdVORNVmbwuRfNLjWObeCDhlnJWfsgAlcO2QTDbvQcsB0gqcOZIvCVP8c3t5AyhTOgPCKtd4TQk82BMLFu8Qb4JTiGZmw1sujxuYEryEPwu7Ag0t0rre693nTlBsk72J07BhMBkAIma+CGz3aainDFFy02s2WEE1zSMozEyvvn6kVyFL/yba5/NHBkCAOWz0mAVpSQbRo86TSKd889VSzNdZlVKW3Ae3y1Xt8C0PPglS/q8avK9Zs1b1/ObMDYAHnWdIGTyE10CYgIOrtiD7axMjicu3+551Nw5gLzgkKdJrWIR1B5iiN1JF3JALNA4j5U1uUt9+CxRys9aR7O1y5EUJSTndXxIrAfyN+mrt1AVluZHav7XlgpmW5f9QQ3CQrzB4sPNTff6ouJamP0RsGhyEsLuW8NoBV8tpXCrT6qcgbsnNS4EGmudDkon/t173+46i7tj3p0oPftB2CcjYhX3Gq/UOYorculNLnt5AuJHHKSziK0ZRf9c7UIQO3rMB06iu8Cxwa1osNERA/dq//M6ZRtbMakEVsl/633r4MIThja+7w05vNzcdYPzB5B/gnq+jdfSHVnDJmrCe4lXeZziDRfx+NJP3kJHqQnhyjgcQ9Nr+M3IuYe3+QiZ4BJxq6yoi1jKEVJfqHn0A/xcGHD3A0kTlyxx8X9Wmj+sP4v6wCQQeXW8sX4OEI76GO2PtWUK8eF/rgIWrXTZIuJjsJn6e4S52F7V2q1/YQgS4Cm+iiE19WQmlHyqVfBNhhD4/ino3wpY9cuUiL2TGfrG5f/9PxoDnc3ZrbATZjgEWxVZlmEIQUCtFxaF+B1syXASAht+LWyrVM64vVa8OOfs+MDH9dZxsBB8a08P+Ximo38DFgfYS837SFJ4vbrRKVaywC9GvfXl9ZQ778ipSU2In2FU4kn0/VL2sbqb/XO7UPPCvVXSVeT5yqkjYtbJXtv2fNGO1b2BxUnMOCCY/K/3OSBa8TrCZFKeTR/3rf5QowbN4VSkq/4WvzkZ6f/Woaso3HIM3phr6stfSQSkl7hMvDtQjdbTxcawADtrXNK10snvmlNSSxu9YH9zLDcfyvPE6Tr0RHmw5qA+99jdBDIrnFJeYjtVkHd3LKEPjNkvZ8wHJ7MsUfkif1TFXYBR6IgwNwXLUMWTYGR6UksHNNzWIpf+xu7alKEW3e12cSfEJSfEVaTI88ZEAWPBqt8PYv9cuQ2FHM49F87Im2PB0daD+XXqQMbQeOkhdZCt6A53o04qMThap+N3ko7J8i5GVLwzlSStsJVGzXPP3YeQqvlg6aFJyhZ3hiwmSD45PMdpXPc5UmdPJ2Ye1qYhbVzWRw1jzf7VFfcxpbkllPZ2bUDDWb53A0wzl2jK1mffQiKTpT6mSuvOq4IkyLZ6Ea+dl5D84YgoQIj4k0Q0QWi30nmuOn5+IKnGXjZKku5nQ/IxWhNHRBN6s1VPu3139+zuAiW2NWCa76MP1B51cJa90zzJvD5pPbB1zzpmTYSVhU85tuCIbbWUZDCsl6JzBG0GhKMVIUgF/dSD8iKMjB6PhOj8YcJ5ukkEtvLGtaoNPP1rk2zSdwkvAAMBrBOYWtOvkcHC/Rw/g6PLGwHMzJy2W+45Uj8o3um4kMyOwTdXM/c5Hg/skbcMI1emkfgpdvvFqAM9VgyL9bAACHDHSTi3+adFe/vPIAXtfK6++xfn+XPdoXEJJrfsIgq132aQaX3CDhjjDLuJ/S3rOb8xnnbu0yBiNFuwGaQLy99Z4p6FfSzEpMIH5Bf48U4uZvlHGYxb84e9mMUyC91Zea+oloFD7LGnfecIWLkX6jw77S2wtS+U7mKecLdoO5G/p3ZXL5FpsFvKNom0xz1L68+Dy5ZbW5hfXXesbgM+8OLLpCr3TNdZ5xX2LmJDMhZQMFmZCHpJCLmznH43MNVYupW4W7Jyoumbok6/AsZPC6EEyYGLkn+orUfgGg9JLGSLJ7USMbCine9y2+TPU4tBYxyfGCxYFIC2C8Vm4AMVumMTI8jcm4qE8DCJ7nsJLAwjDUwkdUKX/SPWHsIa4T1+k45oqb8BGDbTmaCoUkuDOsEAXRgyoijJjIaU9g2dboLnkj26RasZWBexych2uJaHG7Zvt0ty0L/vlrCMXoGZQ01088JbyVaNz0Cs2dAmUhMEMXb+u7pt1HM/xN3bmpn4S4p//aZ+8eOIGEX0LCYx4eKsSBadXI+MXdeleM7UUiNaI5xbTuH0JYJQUh4pZPdc6Yr8//XfG3E3ViNatUCC46ICYA98Hnxb9hIptttoxpKsIsMLO1t1wGRM4RVQskPZCNdXdYMBpB5iE0tG7zGy6VsXCYXN//0+F3CB5ad+djvRGme55SfMEBq6SQu45y+sfyOEY0KxhmU4aFEZ5SJuosVVukx4fjI1jAK1HmYVRkdF8lCpyX/RZIGKCJLcmee9zWPYIEzeB5UE+Ne22QammkNJX/wnR/oVCfL/YFzDmAg/NItz9+wQw+cAdapDRQsuqinmG+/XOf9bS8BFCYl4ydOaEQeQbChYFzQJSVq4y2vOeKDzeyxpuCLcDuEqCvAG4OvoyO8/pgNpFhjveCLs3cIomq/Jm0bSvffmwPwyOkofDMhDVPwRrdSazuPJfZ5lUif1wOToxqS2exASs7uAZhAxJgqpxAt4IBKhBdYVpC5VE+m6vMHGpu8G2J/EcLtnSB0KnSc+pyFUGnA+iesUOV3I5015G3lJpFFoL++AAIuMZ8oIRrMNst0bMPFkN6fDGESkke0wMf/xi5Al6w0jJD79RDc9C7newCRqpyq9sKwpVfzNRtBZbcIvj4y0aQIOGyxaEqTheUDIP8wqmxBjzitgfV4H3/Nxi8r030/m6FDKKBiqMjdJnZbiUProRL4zKJulkBcdl/q0qE6rwYWk0Bj8vM+bFef0cVZ0mgxO3kC7P+eu4Y2KuIhCqQGGAXmw6p0xfACq4ySCnVwa45dm9HL6O2/uVQODlDzfsZDxyybuelg8RblmKRgqJRNXd+69vAn3otVWHAJJZZ9I/RHHGWj1bo+mfb9Mv4FCwJcIz5n+Sh2Fj+qX2d8VJnrrWFnRocgqAWASzA9vqK88nBcO9ZjCfqqieews9jagj80pSBx1doAIL3T+jMYFM99ZaAxfVWuMIOjLJqiEoBjfak/BKnsMmSnoVHTgWKmR3tZKSFZ3gu+vxKPebT14sYhRg3hH4vVneSv3BH/9K9Pm5qWQNYworbejM7SzKID0fq9nulx++qDX432jwWkXDLYVczPp3IdJA5o+LxSR6q1/3kQ/lHqS/0bV07dS7ikZ87oXDpb4/uOnNYXlgOK7ZChy8y3tQKxKtFAadnP63DVJCsh1n7tl1KkTBGvgeeTLXRqfB6ya4PFT0PYoASJeM3CRpaHFaA93gxTrCIgvp71tVoKCGX7pyrQvm3QjyYzF2AFBcLTTQJKncrf7dQx0qbD+SX1VoeF4uWxEhYSP/YdXhKulyifxNZdKajszMud5FlkbmmH9djlpJAyZxHuMvGMEr/uxdHER+lgVcC7WH6Z+gbL6n3oUinR5unXD+8y7lVWiKQRj0stYSIPa0t3lOHUFB6HdJik+DHdzImwL/eqNwdBoYI1K3e+N5OyeCtIBwBHMci1LQgJpSiCUjJiKXv3aRznEpuWGZZUL7vdc+aBSkLm2juf+8Iyenxm2lo88bnmXcuRT2aJ2TZ0I+l0ZSuCKKvGLVr6A+8CsSzR6tTcp6LXTDZlciYY8mbby3/93mU9RtwKfonZEsta1mUttBI0240xQSOlBXvdwlDvGiHWIaGC6V9dvYVIS91I5Ix0Ppxv87y9NJiuStOML369AuCDf6XnpigA8HGZoy3BpRPE2tya+YdjFA3vlJtuWgshxR/n5DJH6jNzgqVjEDfr6LtvQJvrV6EqsWUG/m+3amTPJ2sJHZb68gHbTEZWG3X9+baoJju9ap1rswYg5u3oMUJT8oDqc8WaNQwVQddiiRcQgoLDUg3CNV+XOy30K+fB9vgGHjGBG7nQwkH2ra0FpkGjazuvCP1EHUVh9d7mP+KxnL6b7IMv5yilJLgTS/unZf5PJomEK9/21ypCWigJj7WM/T3kUFwiIkqBMI6JuA33DBE8tWiGJek6MCtQJg3wPUdXzju3TtNQqLjnCOGwc9xymot/tgCFXb3Q4a8QTLJhwC0v8O4zcNRzO3aetUCyftkf1aO4ISCqxETOS2teHHc+reZU9Uy20edFu0j9RGTZlJTBGF7BCwogtF5eBSbysFAzqNsOZVGhp2gkG9GTJ429igmdNKvuGoV2IqiDoth01oJ/cYk3F3fT5Ndnrsu1UEEAAjDyy5H5P+ZBphK3UOvObFQPvbJLAG//jfhS1zu3YA/Xbn7imSoHVuLJO/r1QiynzJyMh+g8T6pQxsquG6fupYeeeSAWdPtpSZnwelcZjvdCXN9II2Uh3NCvhLI3YWKN2Pu0z/IuieHmBNXJFPF/ExSuOvp51Z7Tf+PqUi3obSarH/FBP5n+bxbftEpaDOkjMoGRrN9t+gO0bEtUbrWoyOX4d2jYiiISJbuxyGKkOt2HprCWcrZyZ5AWEgqqI4Yl/SdxIdfYAdTCdsGzIdsqKKEVam9ZkmMZpOyt/UY075LrMRg2xjTibFeVe7Sh63WBHaZV7HWk5OeLtOXdCXsd/3xzYvfnqEAKmZE9vikzauu8RwUrJHl41DiuYySkNQaTZO3Yl61z/94r/PGZADW2PU77LsmIVlhmQeJYoqsjHKNLEkjP3hmGxi0wm+etEQiYiZaR9+TpIakHJIbg0SzZrQVzB13WhNxjBxu4gugN8/cfJh5cRFjKteVwDhIEttGVzSYfbHk+kWVrUjvCfiQWkeHp0d9r3i3yT6IGJLo0MN3buvazqke6VsCI9VAlf1pXfbSfRgcFgj71APefYktDbknzWTBOyWI9pp2zIuPhiiMQXAlTK0E9d2oCjZ1US1zX79gsW8kopANkyB3HaMXj4SkCcZ7uNOPCyDzPvFUZvV542ThBqyGCGPSlm5uoPis0sfdWOiWduLkO43vrn9/tmDt2IBxQOHpttCZO64hnADZ2Z71Kqfd6X4LRPlk+h6lGlbRO77xIIGAjBOCQVbUh3BTNhw2AqP6Q8EbrNQbBorpz9/kCiejhLYH0DdQKaqEgD7SqH9SQcZ3dKFLg5mMbgBhJji7MFWUKKOn+9WppzNjHTtn+PMLYUePKNqbLdVQT47rrrnfvbYhI/1kP8AEZEabGYTx4ochxK6YHc7SvJbPADGELkt/wokvHE20d5fpv8ZzG1C4fYDn/TCW2Skx0zL4oe1Jnc9RnNA0TGmEMPal0ysRa9/k/PXH3gDFESMJGTCWt/crTUWHHaqaDv/X0UsqntMLB9ZnXmgPXz0qTbsnjYL4xOBio6z17JKURXBVK9pwIAkPvuDfR2FAW6PgK4yF+cQGT3jWpE/ajs755L3MSlLTfLihAFq9HT/UslNdnAF4rR8kWsVPyBZBVU6K0tPfQOL3Fn/2flHUDbJ66/rCmk0aL48H+4Qyr56rrvU6UfMzk9oL6h+AIGYYEmQwtx4W1yW7AxfD69uKlchKk8s8zYZ7eE7EOnJbmLFQyA8EazLUyWgffJW9RYRWkobJ65L+BCdJOkfhFmXUtj76pGva/C32XMOM6ob2iDfh4sX8sFTjsIaWE8jJQV59KteORMVK5oTDLYt7zgNTt49XnvpARf1HKXOQsSNTBG9XVcoBoVA6KXJI3tG1+lkHWhHXOSZEFr2WeinC0JxAYCFHNUOdalf7RKuB3fNj+KhxFmHeYCTdxO3ReeBgYTollAIH6C3ANjupYw5EX/eCguzxHXnWt9mx4/lMgb7ii1AOM2clFl/nKOIwFmb9EVZqFHLqJDhCpTgNE8cim4AScx0PURoLE7cIIZ7VeFSkHp7LPDTFiuvVqc20t4stbpfYU6llRNOebNfozgxHHTTLtCauoUBYKsM6D6dK4MvhVZA5+N5+oKdeIarBviJDXrdXZJO+JtVzCYijhS/YzwPajGrHx+L1Zkt+8gJfkS7WSFeq/b65gM1cbPjSArFufrky1PuKTCCi26NCVh4QzVKOb+wbC742wV/FX89+naqyd2rEykaISaR1umBZ42W9mqo2HLij2Lf/F/zfFfV6l+LJKLVJPVY+FCyqQ40EMolR4AB+d0ZlSHXIF6dCXBRyE4al7URn2JlMU0SjjfVCVBQ+BBtT4SIjo0k67UVpIQGKKGcQQ8hAxVEKM9n+Amzen2f/9gk4BBQ6NxdhGWDK0fJN64yKMepjywFCiHC64IKII+dspCIxR2b9zsYNRjqzhpZv0Hc5SJrBCfGz2++sku5gVvANu9osL3g7ONzO+TwyEjRokzSxW+iC9LE33xI4Owu+pN4ZyeYjG3a2qg1eMm/NnYHPMzWvpTzyBBoZghMNkwioflaKYkcMiislxDMqeXlw4D4Gb23JkC12tbIIofSsLaUYOq/O1rFgmxHEqaIeEnLlyuPS9lR09M1erftZZ5FePiipmSqtoa8Obq8FPbIx7lkmFkv+rieUtvx/TJKkHuScMWsZrmQK6K+qqdglizEOulICRge1pjZLgkiJqHt4kUm3xxVi4/8Ml+QJBUkRiAgg378S+zl/jp+QICrnBCezo0omAeUqeVlcUyriQwiClYG2jog0H9sAVpJcmlf3+o8Yrbhg5mrHWSJDTbDcpdC+05FP0W4ydENzJIGY3G17+TjqoVLyfg0aUVyhVWer75+MT73KxkNt8t76mxnR1Mqtgu8NIJzwBS1DJrD9U31keX8YMMwT8ubdUcgT+CRdVNcNe8WfIrGF6PqIh0737i/+1rm8bVOe1quCEqUegdR95rpKrzEKqwbEqF0f5Ld0qrC8M0IlrpN0gc4hg3sBk3BiEORKk3kxoaBLuQr9V7ZdOvC6n2GVz7mhMTI6T68jDIjpdaaNMGPpdEsYzRHVbq0qxGNqITxxhaOo64St1+XQE5l2Fstt/P4GJlM9DJfjX2dXtZkoKoaYVEFIiaLcAX931PLcDmq4jXWfT7g+Dj2Sm2WPwDrEgi8euE42kh9t+9/Qqp3jdsjfndhVidGssX1vrqT1RMT0nlYFM68zIx/GuCM3KS4pqMiK4nKhnBLwi55opdjdI7WTJPfwEVOw+XeIr09LD27MKbrSKrXQ5GuZCAKcwSQKOub/OvjdfZPMf5S48WCuPW+pRnECw2hX+nsUo0cYL+6pWdJGjtMknjYWLFV4SU9GX693W7A9KoAJ/MgkqEK0ObvDB9bNB9MNSYNvTZv/jSXSPuPTzeKzix6iEasikb6BwSCGwbMSslvtX/DJSKFiMzlD61QmJ/QOkIMmzD5X98eOE6hqamBURbLMheIcnI4gYJPh3y0J7UtoOxGXRhMFnXVviUd3B5Faeu5/vVn/xm6FEmzUZ3PSAK0/SPQJ9OJf7Y+VOQ/Wn9XtC+xHa1QHx4krn9Es9y2O9z6x4PboKAfFgceimc/p6sgtuNzARDni2pxMNzrFWdCWSobn+oG2PXcOAOd8Oj6RDmZmiCz6nVmJAQK9YYRcjD5ZWvTO1s57Sd/g75Ghb9N6MtbHh1aQdUzENdwVboRTTgiqMTG0lxITkxIFd/tW6pfFQ6jUo/HIeAvMLA9hzy8gvG+Lmlcf5rAnvXU+LdkIciZdVpW8ucKzQqlNKtyHGFy7fNjtgdAo1ZbK6DkRKdOkTp17IivASVqeJwRPMMDW/pVXmL32vZbxh/IYsbpGUZuApaxzIwtXNgSKoA+W9jwV3rh3hebeGbpKx2fH4Nuxi7jJqL8be+v2ZEOJmY3Jpw/WB+tJ7Cm2flgxW5qYZwrmcOW8zYEozH2RZI6gk1jm50ud2DvKIovsfHrZz8EWMWeOAlGtkKbqJDBMGjknx/8MDzywfBV8GNS0x3Fr+uNioFgYW1UzjcUKssjhD7E8UpGN0DUfLKK8K9xWbz1B/SL7D4vJXiLKCuyHHibaXlmjvJOvQjyDqHBHbon91BhI/d3QDon5q271V5UqltDmWHZzXEcHPLxGSYjbHujqJn4e+YT6LgMBtjqZCeIibLBBKzczHMBqutWwlWde8LRs3qpk+CgU1EKBESdQiM4JmVUvUrBIdR5+XtruIkLxKlGEE/e24l2mJZb7yC1r7iIlX75F4eX4yxcuvT6e30Gkj7wXG+PyFMW/S+UCN43ATQCGk3Agi+beNBWUG/fsyxXAKEmWdcmUzyyYz90xsjCnU2AwUZlBwRuV/YeFE0GUcmX0wwwm6eme4T3v6uWcq1D/XevRe5UHcanUjDdAonhecis1o7MhL0AggI7Kj5cDVR4W+2Kxn+MmrA0GRlVIe+DG6VEXF88aEkjzbOA02EFo1ufyynZIINntGrseFaucHYnZvyWQeYuPwkk6Ichfo5bVls0bxFiFuSOL7f3nvqHJTdwQQo5+DnY6ofUK/u4DSitALfIpWL3uYlaWInHHISJ7NMBQgc6S0P1Xe8G5O6VcFk6Y7OWvVyZoErEq+knbTBvQYHmEsFsM9LTFoJxpGt1Yj0DonF1bAWCkg6IoII9nIWFVmM/T4D+XO34btouvITCZfRSe+H9u4DN/MPp3jeWWo4CWNQfJvRrbn8ZAAI0PU+svFJLdHO5Cx3QbGenB7xOt67qiTAoLrKIujjXXXuYdR7gfuJcjvXwUPBf/UVzugBMMch9po3DlPbIGhTMTCReLL1G1b2bXjEG3GkcJRjA6MkeffHhnDUGXFNP1NNxO+QQzGMCyZf9cDLL6a0W8WuoFYmFt0bsA6NsbCEP5+U/n3JLvdquRocpFHWRcCl7ah6aBk3+fj0dPECjmdRASGxMrCqaGSpdlDDLvLeNnBGc+RvW0I3uoxVflTVghUSvxefXoQRu4YxlBSdxryYvlc/McT0EcbKuPBKiUWF/SVhZrB2q54TeYJiG7QjRDXe3IKdgiypRk+iglo2XhIMaT5XmyU1MhofazjOOX8CtukbayxmJ7q7U6FOpZjbK9t5B7Z3czwRQrFm5d8IhvQv+q6f4T9S3oV2m2nVf7auA+FqOk6NtwcD6DJlMD1/RnspNnUCPFNKPVJlO8AajneVlZtdpNhxKFzC0JSuvmJ2M7T935S6AaiflipSLR8EPPN2njXT6Fk8Q4hdAEXbrbRSAJ9fVKrEaG/XVAAg5Xz3xtpu5YgwXyTp5Ee7AQ2nNMHqNrOW2yRvtBBP6VIy0p0W54OWZNCDvQBIsXATY5lixYHSJGOMAMfJbxXvFs2qvX8WUrDt+2MeB3ItRmYVPrFZd5MQr9pvJXJHjog/RuVY2HwMRREORWL1matKyhyKiIsTGdUcfsLmyvzUkMV2v1uFl+ZQUpNW1U6AEkdm/7kOAy24Cs/il3US5AlGAiL4x9BUOrGcEXnTvAcecPoxfPIwHsi0ZdrwhrStvSG8iLVT/ahxm5rP0Xh6Kd9PQzDw+jDNKI2CbnP0Cn2naSadJz/9FR/KOXAeKzRPn0DcP54m+Z85iq+DByhpZKtPIN+0mGj+dXHJ5CdloiXM7SMgIXUNIW4Xl/f1zDqNXxVBpuTEm1XbIEln78A1A2XpUhPtAn05a7WvyDUmIlaYbcadOI9xz3LNKnJMmJ5X1K5BCG4Zw=
`pragma protect end_data_block
`pragma protect digest_block
62ef86648c29f702279cd0b05e6b3013ddc8b354731f7783a30e3b3e3063f9fd
`pragma protect end_digest_block
`pragma protect end_protected
