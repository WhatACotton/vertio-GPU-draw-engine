`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
AWGd2rdqlkIDSM2eeMmYAqAFpEXX7UCCd1UFi2sJHbPytl4rO7IrGahO5j7bIV4N+UFV8epl3WQibBY8EkBBOAZ4AnJWijkHvUfa2JNUMeGX8AQwRXfWLNaeJ1xNuI3fDuCqRWgfzsxuMBQPSkDk/LHNAErRSXSE1QW19yOQxBRsVcK/tLF0OzFpyCt6dloAGA+0NcWleCy6wiJ7tWzJz4UucQOAl6Q8IVr1jG5+C2WEcLaP1azlvh8d/FrPLxDMLVJqU1L5bW2xR+ToFy5Gv8X8oiAUQ/YQYw5itawlOF+ee9kQnSe+eOditH2s0cwlF8unZKf/6UQXUOHeLL1L2mXkNOXwcTEG7zMHLcpoz7sdUAqKGxuQWM4unEPHPym40bN6EqL6fWcFBj36KnexPkEpBNMOrCkj2ciaLvw2+9cQlcRqn7ght5c5r5xhn/7WsIBdWgxc+ic5CH9aUwQFYJONcYV17VZmOqX13AZy4X6uL0L51EXBN167nbcakRSr5/U1MRnEI942YNsGxL9qtRfKfioTatv4o+rkjvzPxPqlx1WoWvwHnZvuXnNBOIG8ukDLXnUtwcLbZ07ENCWINToy/MpIjnN+a8HVkqpyTYgpaRabdZJhBTvkg/I4tHZIFx4ZFk3ua7XAJgLGAZl8r4ptVuhs3smzD7HK66dg0XWq3PaSWYEW3HvUTceSAZJ8WsPXMwt2/7Fx4vvx/5vTWpppMRmdbQEBAqWXB3yQdakJuFvyvYSgBMSGax2xnKrhq44Lmkho3RwiOPWhvoncJrsXDeMPUionoY9nJJfS5TkJfG6jbE4GnQLT7IV3gbzifMNWhxxocsi/+UIpASxBWDjzf1gqgdJLE/Gmk/cE4kInnmR5+FQwmODNvHG+xx2TvyMNIr8/jrT6TqeI6iCLLXfu8ikT9p92aYaiLy13yP3xA4mIhluVfpQzEhdOzzMoaLGuPlTxhrgOSkR9F7omAc3mj3ERDs4Hw+GbyQbs+ayBnMTpQR2N1ytUsbC66rXtBCYvfG4ackPf7qjHdi7S/d0Lb4vsEZGovYFcD9Z8gQRnhvDZNVW2Q6dMrCSVUYdrAyWuUgrzHF0A3obIpaz/zQpPnd96pR1fcYyQMXRNZHOyqNibMzhaM3MTyovXuLuzbTcjoWR8eett/Y6jkdWVu6tu+bOXelh/OtnYtNCNHeV2Ao/sb7EMekr4kKVciKJ0/sN8mAvWPr3+sO21yNKnGn4ZDV9eQIWR6hZRvFyeWiaB+MfVajm5mFxNuacK/RCIofu90VQdCuqNHvXSR9+u/n160PbWch76LJvoxpURvdOBlEILynp+QvngMKdW3Hyol7WC5LjV8qB1QiPdwGDhk10uv7Ih4d1ECxzBN4/Hd/2kJ/Hd0IVecWwj7xkwYomx+nrg047tJXHaSDJ2EgfCioroHIFUyQW4Fz0DD0bvHJ22/uxNNLYs9InPl2NdCRVukCOcqrNgO4kjgGeAP8fx+Ay0BkG+kMxkJJMqCUzuBW7C0hUF+FUm0X9YPog10iKakw3P4oI/Q+rr2yg1xvMBLRpHGnkIkl0JZ1kaqLLQOSfcqpAv1BaZePmXCjWQ5EhxqJjjnvtHqdiFuKdE9SiVGwt2k8cOVgngGS9tdlFtVcZ8cMAwLApLLsBPLU9MjbdtCEc5FPxKBaqOjjgJ3TPe2AyPiwV7Fg1kt6UUTV2CR6Pz4KpOrLQdMJoEQwXyIAanE9NbRmzl3ZV+yQkVGMXrrKYi3H0NJLF9tguVIvPIvzh4svjVqYnYarwBtMJ9XSdfc+rJipG9BYHE7vtULB47ogI6HNvJVnEXrhJbJYoR5U6R6IBNIq1vzZ8yYXQp8EZlf8WctHPgXmPlk4wkymT3ziOzlXwDppw13kXQyF71pM8SDb/TgvFkeCeWI1XkEFf/w+h4lTax+qwM1gPp66Dc8rzZZVMccdkvcsVDFczO/oyZI2PXgbPoe8o3DiBk5QaUc1RMrl42VYzjUMiAebfT6Mo1tYW9UseI9o27Kgoa/WBMouQJpMCl0ljA/mMdNC/pH5Z7qw3dzU6eOOB7VdPVldtSm550/klpM77dTlWMCEcXljZJHazctjOvKgc8s8x5lYwmDDzWH7RwfqUK8sJ+Eji+MiYVYsOM2yOLKO21dtnwe0YJS7Y0HjUeIEaNwKJuOqFGS+mcVxZPbMjkkyRKeErtO9hxdvrgsGTNX90HO6mIZMR9DctzPx3qy09N1r46+70UinBh2belxM3BgCsKKgRwvMMqhLEpezulp1WnRK6a29Jo4y32kJQ8/IBlNAAyVFNKb2lCiIUELgMVdX/7xxTv5Dm/IAAmVwv5CwTM4+LHKzSJYi0tdjB7vWNoMAS4KJcC+VF3+miqgQrBrBSChnNci5gJELtaB9SDvDX2fEJTVkfpytVr+qM0t6UbkWjGl2JMaVrXH16aJNq+HHoi+QB3vgxIUDZnQBMQFtj6lQL2iZ/Kr3DX4nWxa7f2MbIHoLjsqED9KDcZPJ9hNdhW+NDrERrhwWkTWdPNV1H4K0mw3kSs9VZ4ot+JVuriaNdtBgvv4sUm0Yvey46N2xhWH/DMzYrhwEOVncDnTlNRD+nMoPo0c6UK/oKm/wJJ5mOwH4uV3DERRfttjKyaW0htIMvUsJdUfxw0pbsJdB26CWgCBk9sIr5rfkyR09na6zSUfKsiZzk5M0hEfOwqr0hvqmqHRTes63Ek/qy+DkmXk260T5gikQpbLpF9UYWo0uFRoCOBPn3YVc5LkMut7uMNR6sUB1iN7eoTcMB+VCZhIksEggQtlzWvPr98Rv47RjXc/Kr8480IW2HSM3WWx87aozq/qZVP99IGBdCxj+ToXvORT1/Z1TNKqtkRXxZ4GCaMkdUP4t+MVQyWZCkz+50oL8ttp2xG9EZd3rX4Pn5W4GjrDDPjVoZQX+V+XK0ea14j7bX7lUhWJmiJZlDc1BXulCl3upyexHBX+pC+zx0FHpDM6gKC1fB3aKnxz0X5opGyHd1XRafgSM/+F879fe0abCm51zp+vWWS9jtyAFu1Zp7J0sHyO/afc0zmHuLqhdbNQVwWpTXnm+MgHc1JSw+ikZlISUECH3R/3Y+Oz5x+v7xVRDE7Rht3rK00UAQkEXvLFQyTyBmX77dhz8uIo7GsZ3lE2BwPRLyQzeC75w1NV1uDWOsc9RM7ca4SoKrZXr1W0958WPfUV4zw5Fq0YobHkuuzVR9FvyFoZN7p+3ALV++MCe2WtZp4jdDxI94FILnnR+XAOtwk4k9pcfWgdPbIvSo3+9E535DmKjmDkWv9fqU2Lu9tbUGsMBRbSfEL+Hz8fXC5algIivl1oFNIUYWhO7SbYfySNH7gOJL2gSOiAxznrhOxW8eAEZZFrQ3MCpZGz1GTezsGzvEH1lv321j9vCdTgjSaf/Q2Ud95pBgQn6deauqEtQyQAJiD0nmJlpWZ9CsDTc//Uj90Q/IWPmaGc3PiAfPz2srozQVWGIMq8UEGat3lAuuR6SDuTWP/et/f9hyDhUjAPa9BKPTaCEDhWp7+Ee164AUvNKYsC10ncjG6Ht6GMK9RahgCaEkbrepHN6IuT7aPN+VobuTID3ZM955oeCxL1wOXoUr2tXv260tYrSR2kc5zNw5ryyl2+Vqy4MNXqooBArS0Xd5oKyX+bsFEZqanRlqUdO8qlpn8L2uHTe/oLyQJNKzuC8vblk9AKfASTihbBkJOrJV4dlQxJjqmCBALCpvsnkY0SzJca3FJ3p2A90tVvuwKyULHm5J0obR+GPKuvURGDlRyQP1tG39hFgihcAmyrFF2NIBps7kJ036jpwYGTn2dzQxcb+oLGRI/cd0ckHSSG721yiEsXaiIySNddTRcGw6qgWoRtCP2FAbmEugX90rartWfhWsVE432kXT7lqNhBYIjNDbsBfYJiWb2x/fJhgYJk2667zBucL1VBKqmgEWI+C530Bgk33LSwc20fdy+zUZOBSk7DEKMaJQ5TaB+DHnNSVuS/DxjM8gTCFfdXOFD0Uqb+QJ8TNT1JMk376ic9ZC/5ABN3xEEZXIN/f64GRkMxYgd9yd0K5UNhJfsiPsorwbsSh1W1epU1IoDIaPoSZmrPkYre36qTBPt+eotjI2+1THR0OF8J31PUmndJp7+y1xTB9fo+5t6QM/9D+mbCDULHGQ5alsrxWWvgT+GY9Jxg7/LJ4dWg2cW/rr7jhtaRuRYQSwFBuj1ZyBXgF4eq1mfIIvbRUsAACdB1zegSuuW1Ks3K2zihHFQ8iRzy4A0+OX4X4EPwDf15gxdmG+mG9uizowp2nS6AC3aDOZAKS0w5XenVvr13ytL676E5hmqnu2Nfgy1jdBlxX18rGaYT3gFXhrwJcEe7oIEWk9e+97+oonlS2JhpFmEZ3tGllxdMor2w2EGFSZtNisCAPbmOI0v08mMAWD3XhPSx2B8BMmi3iHpZHE+Jm5OVQmI7HADZe936MQv7kNdU76NFjXREypYZ0iJeQ5F6riekMAKDRYhN/EOgjyOlJM7VS0mRAEtwD7GVQ5jpFVrXJnTEQST4UH/Pix+oqTW6aCWysQx/JlXnaBeAuclQzV3MjhzgqQ3dh8qCvvFXm983AlhXJ7GonCajs6hMOq8IEhMrBiUDF5LR3CpxZQblNT4pfWkxJ1GlwpcNZYPCJ6NuUGdqcMtPdTOrAqNY/fMJfAPh1TDOv7pHBV3wDI/qJFVDkxFBllqybHGZqxq6xzKttnoUNqpK/dkAFqtLMHxHQBo3JhtQrbOkXR68J8pG5FkZXqCPkEG5dQLEWEtggJCyZkFtEfYQH3Px4fqKbGNCWjSrLiMEhcGBwwYOQ/gRc+tuoRJ1M4ayI2n3Kyyypzh14j72jPkAQBeFuv7cvyZYuvpHeht3zCK/+Rezk3FL7KzTY9G9bHdfhaothbPwNRtM7CNXoksPlOX/Y+1JEXyk5CAnbO3jGtJM8H1KizAtkwkdsj3vYKDhVatUtttgbAT5EwSwXr4bWGFK0DWi3wbC3M80jAaPKMw8xhIVdZzZUHeM0SveR5luLeDoH0slK4OB7UeYSXW1hBOYg9d6lRsNIwexSutXTRhO3c4m1BMUw3mpXmJOw+dKWC5oaDufUX/ukjpymYS3eH5SmYdFIDULcZevWo3EnEn+utCZu/bobzxKqxQnHdaeyWjCWblPGvoBM25qttIRoHf/2F2DlbQORbAhmGzMIYheU/HOg8ieoASzt6yamx2++Oix3oaq8d4wA5+SB0kkmGpL47866RYRJACYxofdQ+1evVu5aZh+B3DOgmbdGxNohc1nKcQqCh1Ogo6IIQy9XG58GdnywmAviwnAY4m/pV2xzBjfyPCt2NNbX1HhgI8Y4f0mdHZEeziY/s+/yGplLp3ol2Ice2zHlLXrfWMqiGRk6iwdoP2WTG9NWUdpBexfDaQ+xiiJG7l3lFrbSaHlxnbDJ9YEjMqkzJieymQYzH4nyDA/3ng0Ve++i0xC2j4GevD8kNeFUvNHvDOAgySOitBsaGzLx1mhR0lmvF+lmNuAEZDRpvfo1yB0D9FTooze08mAGjpC+L59MsKaGvR0HdFFPUjU9cNDXXANpdNCngTecY5ObO5ErStg/ZIz8CjXPXJOu05+te1XHl3EeMqxu0eFxeJd91w1eELJhlKk5LenI3lm/0hLXMeaYFCRRxrIDxxdDpy8RVMb032U6gHaz3Bn9FU4/Ly8RVWn2mqBL47XZTYSk94oxRMhlisdtVIf6IXMeaFV/x+zj1OAa9RAw6WsOPfipSXOhO4MJrChGeHSa7XVnqikk8LEEi5iWex4dqUx6Pbp8HmgeIYqkZInNYMzxHuu9C7LlYDdvSPVR1C8Igj4l3SlqTo3kCijCfSR/18nEjfV+wmugt7ZLW58dSZIohytHl8UY733wW6iSi5z7/OnGoJYCNyOzyIYZ1qZ7HQsYuw80PJ0vpx2uipZXBk10RJz33Ir6binSWSrf4ZhP5OmhA1XBSR1HiclaUess4/zsaLqtyPouMy3FmY3gXRiXvzCnsdG3dhtuUbmzXPcgSMjTEZeUDREBk/wURqAHRa0u3HQA8yyNEzS/7Co2jQxgIwWdMcviLONDMvvsYDH90ZbK674/VFEpKi7R7R2xvk81FvroK3gZhPKCSSPCXT4iSk+XHnUMgqE4X40WUhsQaQ2tFQPUj5fP3wsP5fA8wTSBRWjSRWh81pJ94fSe30rp/+SIE880EXG6wIWnj/5dzV6bdM9imTQQ8mHcpogTOH7l6YL23IXqpSPJ6qyKkkTL/EcG06qD+K4nxM9jyCuH0+4FBTs7Ax8pmYRDkxqZtyGgve3Nmh2aNdbr71oWX60tuyBoRqUxYdkM/sGmjit4SBW7T+Qbtw9kFqFPGaeJoiR1vEQYPe1i9RIGvsyYbgXZ3TKu8tg6/FYiTeCIuhtesw3gEJ4QZAz0P2hVoiEitRiAzcsRLf4VC20A9mlLVhWRiS+gIxRhZE2m2eSF8ciGCN2ei50UpyaTFGIhxj4neTe1cjeqYKF0EKmuyLZB+f3wSAJL6azQs/tAcPZa4VqfH+QAdSHGjc1MW0KFC0rZANiri2527UEYLucu5IQQmsQuvEF+WPonv/iTIRaygWLYEWq56KZq06oHqMu9R1k/3/yHymUaCiZjNAyFIxU9YlnDphzQFenc4smgekYo+ORrDeRD/q+PdNbPvWkL9Hw4vf95gk5UvRRIN4O7PT3Gu9pNr22CIjFHv/JyQ+7HH37gXJXGYhqo5mOt51DZAMB+Ecrq60bUffdbY+1L2Qyg22s6+faMDTO9LblKveBsqv7IACFg1qbtmeHZuNFuYj69bsv3+I0pfsH9/fUBq0CliW9nkVrRvq0mGXguO3dLBdoO2ll+CCrqRryAtvlJcZAH2wETqHfP6+jEoL4otDbnymY9hZnYImd4lhn5YokDPZA+1swd+XkTMm4obnoB0R5ROqpTPkdDVgdhyR8+6l6eMMJep1N+tSxw78Q9EiNG8smABuZg0Q8Qoc9A0GqOe5SSJj+P4s+1Xh2/qJZz9SFvmTDCf7CxnTbiklow7UFCm+0bEFy4q4ED3uYP7MAPqw4amfLw9Qe/UOjetfAaJtTX3RdzoMJ9Dzqk3HN7ZUUqtu+PWIkUPzyyxPTLl50EGyzvecy4+1KErTIz6hDSl6AD0mcnkg4D5g7wfMmppDTtQzT82WrFCXBrR2IxR/S8OiszaswB18KjQQaCBhewp7JZzRXzAGF/ka2QVajsSzN3dKHwDvhbotZh0mqte83d3vWyKHX34TDarl3R2aXEn6NUEqfybvswzCLsg2O8qN+yNHd5FvYNMHBce4goNNoiu/iaPb0r1c8BxabFXBjsR2JKE+ZiR9H9qqxBTEMxTGpw/ulh0goCXE1ZQaugVPYn41tSRjQGGICkpFM/rPVgrIP3ydgxzK+loKnV1Lb9BUvZ+wmrCog5RWN7tKI8Dd2NhE/nXtrYnBA4qDrnhBdczXVYF0mnFWqneB5VDFg/V+mNJaBFf6KfWnd8kGSpGLUeWK4F1shRj7USALXSoy0mQ8CrMfsyHmzNwIQ6/VASLWU07CMN+y66sfE2aKRI4u0Izz5fXoFy7pm4DgXVH1XtctCIBr4NkCHhTPvc/mOrCBts8mx1IS2Tonw9pa4z7g6vLuMVG/XheQ+DJwoEX9tQW/xfa8su5o9HpVlqq05J46B/729h7+2olGCvrVEWLNd4Y8H9ywlfiZkPHQNGtSO6dZWEKLjdJc7iww5CrhlnLZp67x1sOfkUJodS6r7UpdsqBvRqvgm98s2eDp2yWzQJVqohAiJGPNIoubvTDMuYZuy6NKgdAANQc890qCLRKkStjTEtfNPLGMLnMC/uklP8a4XRUSzOCqvU4Dg5AMUN/D+AY6FZvLQ7mXPPMdqvRJGSF4gZ5ow9xS0fYKTmLchXRDwEEA9cWrcVahBwGsDmfGtVSdtTrhq39K5v10/SXiIKPATLRQnJVk/RYR7IdJWTR65CFD6SuhQdREjDF6hCQ3Hk1rUHcgydUPBZYwE1rLvQ9dsLsvhcncFnaG6h6Oglw0ybXvh+N7KBRryM6Oge1LkY5NPNHY/UTxut9kQTxE3RywCY7IngOS/Nz1Cdksmvv0jDn/VHeFnxF5OOIOSnyd1QTfMp1VCv2cqU1/d1pL+wELoa2c4TBS10SxxWgDAVNRd2L8NwD2yn+7Cj0lGrsWSuptsuOmllt2o7p39AqBz78BeCPe2L5rJY5OqE4+poD/fjdF2hH3VrgVThI2b9JAv3ll3oKiGNqhUBkDVQxmV46UIJARZoqs3dQ0ySr1D+PbmAyqjWy09KXLazVpXkKRlNDjkDaWNU+24kZ38FhjLwB6nL7ZQxtQqAbOUsoAgLg4oJKchqJo8OhvvDjz4U0hhLlLp/iTX9HYclDhCkz8guDnCrqACxoAP4SBXygC3IDs25cWvBCXP6jBylJcN8fU6WiOX7azk1Z2rbkXFPRhWAQX+kQK5ACT3rd09gYcDeB6VosXVcL7kHucloUVO+J0kvTp40lWT6I8dYtgVra7J8ZYCVgUYaNrgrzmP2cJKPBwepLrh9O8O+3UlIl/VLd5ayWckEKqaWoSb7rkxUVm5gUIxN6DpTWwVNS5DHZ9Ktk4QfQvfk8nTsTsssi6AFhl8a0N1UEN/BXUAMG6qdrb+fFSkbZZQVzD+7uUD+I7ZsLH1k3P/mIELI5ZB0YFVolHDhi92H59uaqpRTkCPWSZDKd26XSG8YW2/RmxLfDdEaw5xKPK+Gev9ZGdcB7zFcXRj9sZk2MlfDSckP0r74GIgw5xe+m/4EpQdx5EXcOdntvb5rQ+7hbANhMnEn/XDbHmqau2Sa6lqdVUpXQg7XwP98YV/U1e8ezbfrBGAmbswMc0rc7a/StklJm2i/X3/9rYqsE6uenBRJZwswWQV5C8n8Nf5nh676djc/kNmAbIEv+MYaq1lqob5aKmqnLngKTl0Djngg283d7wlios/DKj5gjGMPALXJShwhw/lIwBIDkNB6opHZyyptEf5f9oo6kCFwaP48gomFf3jbkrc7nSVizY5UUzpayC9sD7ak9LSTR7v7XoKuKe9aL8C82sm/VN8jlUKje/Unj6tuQGmYI/MHuLaFV6qv2WxE1+UOBaK98FjZ63AnuGmKI1VMwLcfDBAGgHqkQRdjOgfFMhtCxnRb80sd1HjSNthEmyuJw5dKZbbL/dMjo3wozj4BU8yg4L44v4MXQOzwEQw59onzKsS13oTvOyUuUo4moUXkQTGRLmWaFtRbal+/tuKt5FqiJcCVFCBd5/9obFe5gH8gQrk1UAPWqdt3EuBDFIsUIZonwXJcgaoMdMEWVpSHx9pEBBrZrYOnJru8wX2Go2Apl+4bCbJSjAQZwdpayX/gIbXp/pKK+Y5CsnxU/pFHcc8u+YbOJSt0ADdA3bH2uJxIQky93RvbGFOJtSuNzjTi3ruFg7x3d8JmLIqJBNwswtfHewnoIT3f27biUf4uN/RAXCRH2GejTzPvFntmdcnIaamvMjRLlvQ3np1XAn+bFBpOSK6OAVscQjx2IAFcwhaOpemlDo6zzHIKDBwlrf9ulIlgwxrKN9hkFlz3VSrKaxz+ZzSUgf+jzRSJdI516hyffbw8Dsl7pt3nF82PYvl+M+o4sqF4kHp1HYCUTkfqXb/67X7L96qJzw96Il0/iX9AceL8nXxjXoGHsoIJ0Y5s8xAM+Z5JerZelIniaMHiz0ey5h4hYwNBPTHq+DQscve/G3d671/XvW3j11ImanBst1XwP57Tu7nV3wMLqXliHWBvhBGbK7MZgQnQdGWS4EcKHW0JaInCfL5ttWsK/edqftKjNmb1zvOax8sz9sdSt0EjA+Nvkt+XD9b9bei51NepbPrFR1/w841O5JKCHfOstOHuc2YwzGAYkVI9SLKnhipzuBSEpuwDKDMVZwBzcovNRmrtpNE+Og8BZ1hoilnZ0d9i1Xe/702CgJH6zTgmLh1iw2AqtajcGQfh0gBNnW227piZohz2EB2BtQHEciB1kfgDG2lVmkcgsyys+pvmXFHEaXn2drHCBuoMnqmZj5f76mYCgkAU5bcIcaG9W5Ju5F5ATHWnfNMSqHfvm9ntMpcR5Cp6T3xNM7PfMAuirLJVvnhtnCu6DFt7asXDnIZUOng3cCCQdWkdgKRaf780TEf+8oWSCyftzdPYwMdeoNhJuCo+ZzQcGmlNvkLifdzS2mdGhoVKE5wcdDS0uM2ZNZKI81VVzSF6EaFI92qiwyD0xYh5boMBCCiQRhZNgTlMmGW/bNN15W8gE4TFXxgych0xi6892BuQGbeXQB2ozzVzFcPwsvxq5iD+2nOhbdjYr5XJC6mCuU5w4a0nYx4gStN4he446baB1ANfy4hTv44QZ56Vv+99/WXL7rdqMmwAYkR8GVkOEoIHSxTY+zP5xZ3lq0FlYXZof/YDhT4Gxp9m78qmyvaD3QpjgOLnleROm0hEfh5G88k5q3C5/1BZruQwbMF0U1CvMMccXInnIjVA57AX8ip8lvAOgND4HSmjGQDwvYwFCKCj5BxqmhlvJHAb2yz+APu+yWLoD+jwp3CIJVabN0LcY0KBhd5KVoeGCj676InS+q6keBzTDqkgubWQ4FkCKRb3FR6O7oc6RTtqwCEBbWtn2qHff37lDsCH/2/6temHhTRg4UCpRUYR4iWx/Usaq0/BgFz+sk+TFx+cZMMaszbhDIjuYmiZiiOrQwv/IouspOj4GXlg/Jb/DXQqzlmap3/Rc3n+ctITLgxkp1C51yOqFJh0xO9jZ8jH9EuBrC9is2ZeM3z6F3/IsDrT6BzwX9eIt2jvT18U6lp9CZs3EFEHil8su6cBcsxiCtuhN2W4SAw+WTXCitjZtJYMC1o/et7ZGlSjS0oq2YNfXR6S4oQpzcIPx1q5JLt/1UK6TnUFWwoMl2S8qkbWmtjKMESaWyFCI68fGSlF+CJp0V2L2WDVqpAzhfkMSs2D8WZpYLsY3DiLLsoRrUuYQtLDp3UMHB6qPVWhWDyZNkWodMdF8Mm5gLdFXNXBHR5EQgpcR6TPeIp3ngD6uaqkvwKwY+akCF11tLlzHe9TQk8Fkv/qDQWjFJDPZO9xXlSBP3S8HvS4cdoP8d7v5gGuD3pBqKoiluPXB7u0Cwo3kPj18RH9bCj0+mQEFIeIPP/6maOXWZSvnG7rR7aLH5sasONUVC1PP8x4Meru0PjlHQI/iSv/Q94fva6nqeHkDuHxz8H4+nUrqBAodfaOiq/zZeuPTaYA8NFAHQgHxRMFzp9SBAQNDUa6KSDDjrqaT3BcVJoFbMn2QkiXVFsKCLjN/m1FqlGbyDIPMWc46Cjt5DAMlnPTwIGqB26YnrVw7PIB4PzWzMwp6BC6R/5dTgm1R4RyrVahOEzbo2VmDTRcPKxCZnJsH5QZpY4XO1xod10apFrqvUTPCC2NCIb07+doe7YBbTOB2MgGORw3idiXY1FNSHwHCPu3UZRWmGMVakDfgYn8CHk7F5eZE7aBX0CsMPqh0Hu5MriQclCug7XBQ9n34vkaG344MrnMyVnYTuvkbsnNR122DGg+LxooGQNDhjFaXRjonCMXT6h+lj+yo1lkw7OaI4vvGJM9x1ddsm7M13zTNRdGK8j4f1YWlbwywubf7NiRay1l+zbx0iIhs6Tbu9KwX5FKmOTKw0tRWyGEetVsFKPPPj+58dpEvMic/QnXvDKRVVx7e5KHLY4QplkD2sozJzHNtZb/aCytQGFdymy2puhMu2wXCOb/vOg8f0zgq4slx5riZEJu8euUBML7lR5nhQ5U2X3GDdR+c+B77sDSnVe3QNu6mak1cKaPoCnL41SlGmhktD3DuSTNDDc7kSLUc9dOwHatRyM8BNNAQMN7+lHZRJ99M9mlgTLjtQfUDDHtYEnT+deTd/aJr/y8NE7E1OqC88bHvwdvwsiNrKn4WZAjtupjA5AP72Q43J3bXWqfK/BHWilCWsfFxgUqeCIencmyap86F2BiXKoday+ay39DPfEwgX2/WMLCuFKID/ACh4A/r6lZR3kfc1+bzQQhJTrRrmN+Mq/2KEMITi6IRznfiF9DFwefkfpStdJ/O3SKi9Io6X/jPDjiJ9xGBPEBE/75GZWMvzN8ZNeHLiJgX6VEYk1ZjIirWVi1GBVionNq2g9apM6If9TARHIpPfyzctWIlPQwqcoLg74h7HEOB3eqgticUKzCxTxU0N/U5h4mv5nl06HxKJt5jaOWiT1kT1HZzYx66d866qm1SRSkicO7DXahZn988Uh/hNvo49Jnze3qIMR+qRawnGeyiBdYGzYnId3ODqc7FQjDycRuXpIX8cC7v031TqgrjWERu2qb1vP/onnIRATYeC8XwvHoJXfPOybCpeY2NHqmqmuFvJlD2aqeMSsPSMV3DhgSIUE/D3ZPRK6f6WFremGCl6u/BbqZMoFDiRrM5WWpBMwxpxC0LzmneC2iH9MdBz0Ggr/AFN52OgsvVXfIz7qrkpQ5hYYXzjRKzLHoUGG/4J1lpz96mwLlY8qFD5BJ6X8K4YMNodQyd7KA/mRZq5v/SfAtv7HEPUIgrE77vgj5Ihgj63RssljV3z6wUIjxIdqikYTPa1v9paPUAqWOLEBREmPc9HG8zdNqaqZYGLOd0m26ybfHc1nJiOS1/Msd22+e/nzp87/IQT7M3LgMyDghXiCMju0CxM/2Px3GMcmUylJnQWEG+LtWuAlyb5rI6QGFjps6px2SUkvwxn+Iwy0gIA3c1w5g2VjvQ8u8w/ZomrYi8sVR2ZZW9gCykpjvaGveO7/hXKvZxqwR7ImvQOIkYVZuyXdgACY8dQ2bxqPLdxDywSgpuy0mERwuV/L8xoxbq7cfClyGFFzNbrS67Ns/ipv2jsd8KAbqpqB/WVzF1iWktpWYYkEXRSNTccleZxjIkkgkCpz+tGJJNFbngFoteruPPjPgg7M9mnlMKby7uaCdJ0UXVutFXAsguhRd0EtskBb/QRiCiQxnu6EsKEyg/fgIPMgMBodn6FK1GJp3KwBfquSPNtCMkz/C2F7YuMIzoxPiBIetuQDMVlQyk4bY4UGYOqDQln8BCExiIiAe0U9gYoGLZhYmNdP2ZkdtpQ9uNTCUxetD0WLCQTIwQBhGo/R1XjrL7HJ1KXBC+6Iyaj8wnabCMmwiE+E4KJkrYzUSUMxM3MY9PzI03ekMDJfpQ9PzrbWcNZeWrqXVzh6Qbknn3ONzITaMcsRTcuZJZ/vtu6M0Ofi1pniiuwR3ggNMCREV4rzLx11OKXjwQZW+aDz2b30yYvmwQ7l/F0sLpx0oHMrH20tHZXv84r4ZLZWmwCqbCdwgXL4HHaZsassB+HQu+Hum6UsyHAUA1yNff7z0BbXoGndlsDdGu3DWkYOVTjzrkWSWcfN498xO58qx663hkSVfPkoXT7sWPmdERu1ej2iSXf1TXteQftpqyLdvYfLLkNHWMloQ1iKIW4FGnGq6VhlT7ys4qVSkYLCE9JmT8qsX9REZnRlY14L6aDLx/FGm8HCo+UC8jczwStMVkZTQMv7DK8vuBV4w4uikC5RLEzIDaFKC1dAW8HR7+lLsJ6KZ/fI1h5Toj9cEPRCy1oMEwRCrSd4jj8v8w7SJPkibSdTRXpG7pLHIFqzeGn0PoPXzOy7KJGoSIcxZYEFz4c8ysZV1kii57DkipvpKRql4gA8XWLsp1mDrMuo1TMbBQzLIomj9paYzXOj++oP6VUiSV3NtXwiV2UMfCd7wISg/l9JMxRnaVtg24ucnb5zR2taYjmoxZlxhpHmRSm1TZSFpNuAu6Y711Q+qM/e966hitvwJvTXKjTSwTuiVdgnTkreqzRElrBPHSowLO3xfvMyCbIC9naqXBfL5VEMpFnJlBlJ0a8kQnT+L0fFcb2aLPh5J1udjdlKVNiVOG7x66cSV3OXv2Qstp16PcKu3sF+UbbK99DJvV2Fd8L5hFD+P1Tv1ioM8X9xkAOE9aumS8iKl/YWvQXxGoCV13V8+/WcYW4JllnDO2rPCUQHPkTDjtIsiS3pgcUGBT6XDZNlRPMS5Pvamtkb8F2hosHBuAIfDTZdVOAHgJCGpM7DUBa4g+KrPxy4UKiSB1tzXDDj4mUuCl15nOtoGWNPLQJFeXB+rucLR/w4fcq5KktIFrHJQ/S1HRJro/268b/zUlhZ4VyDFvLvIOYGqDF60F0VaGnXKAodNMrSGMB0l+L6fKRZlvS0w4QtbO7zffmO2jj3GBmYC+D89lKZwD9gxTdSJx/0UmzXjXQBWh1/HmiMemy9fdZ9PXN9DWJqQQCBEBGfc2TGLFR5fhKeVH+QWf53dI/LS3pSuvrbOMv5lwszw+85t2uf2q1W6o0+DnT1Aq5MmSMRA4CK6gi7QWhvkrIlBh86wG9QoOsyE+hvbw+W0qH9edr9NRQBpoLkKUq/574j0VdfjpjFJtw/qIS7gx2fLgQiSITRwPt9MUBJXP0A/Py0WkHPi0UXkQpH3DKNvaO6E0kvuxmJwbL9dQKpLEeshgcvQYyhUIfFQSJ+vPvdtveSp+Bp2F3RVgrqdL60wwO3wT/aW7KHjFNuaGMUP6gONgCQqdjKBAb2AWF+t2xXSezApagJ7NSNZlTPbsrtmCFoJ09s5z0d5zXcH3TVOBJpFmay3YXtYM+XcAZcMpy9OehJSfCcbmuCmx3aY2O5abx+x4iAtYf2f8QWbq3rnqRVNjmZ7Nm5lXJzt11n8E6wvKYOqNFi20XjSJJraYGd/bqFkQUySYLf4YYkiG52kYbZ8eztltQCyFogMawy1bGAeNpHXsysOL/4Ic2b46NdnpXh1MnS8NjMpQmGdlqB6JzU2NcisqTjI2WCiHuU4Atktp/UgDCNxOBRi5Z+hASnVXG+KVyzf6oeY0Khc83hcgQraFS7K4XlGA81bRZQmnw9ox+sirE/rWFMYowkWgNpX3hK4EZZr1uo0fOESwfIHU7NpzPBgYM+kKwYT+dI4otlsGULKJw3NsakzJ1r0kps4f4vQksUjuKCR66r7T5ku0UTYjXGqaKDsqn4ge2m5qwLkeOz2h0KIKX2ZjuS+eTrXhcULUhQVYqlrvXe+6Gwq8/an1/ByXGQXYPsdpcM2Ei0t0FCWitNhte0vf/3IN2fvl5rjmCchm7zTlrSFrEVT84r4mgn4GMzSDiV7h+L3Mtu0130LLQFcnsuaOPug4cKPlmDsA9kLg44F36m4GIEdtfOvuqmT9RpxlFWWpTQ55v1/Bo7cfY3suATfImjyavMjjzlcsecG8q8W6ezXBW8uoDQQdOD7nJEyg/hpC8h2Jk6WbaEpgttilPkEvaYnDOQNv/aRAIjGje9d2mzD0rqoEuPK385+pKqYIYn887yK4AHi9uscxVRUCtawzEvZgq6U/mvCoPYDYyyywYeSknXS3B3PU82/FSEC3JxZJZok30E0r7yF3/Ncz0sdelyK866F4Z26zYz0S9WcFSjeR/LcbPKq9x5DeWD64ED0N0el1nxE9+yZf3gIMwDiT/7VbIRmBr3SjOx9rH8VDsxDEkzGrSW0Ns3rGbwI4xYRqzZWDnYXnbiCOEJYFWXIhexp2CTqjtyj+gW3MJI/T3VePX7Ag0k0dIHL2vF7bcTUtmTAFAekRysdHjvqGbENcmdci7TKqu0hRWFGaMRB/tuxR/WDHLIqeLFu0nxAapZc8nHe/6xpCUtw6Qa/XPjFD5t/XhyhgsfjimahzbomM3XK0US+O7FAUQXwr9hUM2JdyULfz2HnyRV6h7kyBt9uG9eI8Bo9OIIQkOr0pPKJUzJUVw8qApE/jVydJ/scBSS/r1EAz+dfw2WgyqkELJtXBwgfzR/R547EVgCfS2MIQILYdrHOBrrIoV2F9uO1GpN7nKbOfx3MNgAJJupQtDC/nrW9ACzq05Y1VveAmc32OQJH4rcxSEbuUUvCrkPDf/V0B3UXnMFqHpmhZ9u50J5yM+AAz4VIqtrC3Eiv5//ojFwOjur4JFPxhsSv/wR8qS0XxWbS23BGMlGF8s3tP9n3NcnmPjvV7LEpmeZ6B5sCVgdPPURrLMt3MKXvURnXTKX6Rv14WFa/y1a9REXe/Ij5pxMdeTMcq8FqnlpbvhN5ioy1McLGPrfWMjWgulZaHfv0M5ORu6XVjrpd43TexnjZ8oKIRC7gxJ4zsWqQYAjQYE9Rn3p1PHx86bgDDrk8gqclb1K2xOclXnKXJB59vdFFDEqEGJToM4A3LT6Iqgm5Jhvmp5sK/mEYGkD8z0FfyuN2l5BQKvaL1JvVx69QsluZuKq/L8Bs3Arp6jl3VJcUm45wf40RW6S23Sx+vnJA1nmJOau6v/P4bn8aB4NEgY0FzMePCcnnV7+e5nE7ZOC45UQ+LIX0RvdYG7QG9VSb1grKK4ASvge/O0rFzhkYYkAUW9OQS8aSuKHvXQybHn/ZpO3pdux02VkYGML252HPAnAth05Nlq0XEaas5kO/I3k1HNkXuCnNbbSn1m9EZPf6lbgJkGDavN3Q2N/gh4MNl9T3mNaDR5ttn0ERMjnBUeKdAh/9jWM6ZnfdRn1V0yCVrXKF6NeIh4PlsKIh57xp63jyGdYmmITuo+IR3tgQfCy30VEx0hlXmJaFQtXpDo47wtFzChiCvxqcQ2IUDH9afhiJlYav45xJxqUcx4CdBJOo9P+bp2voxtsITS/cH8JqHiMpkNPP9rJH61Q+vmMxYOneNHT20++eE8G/MIU43lTKehh+w3YR+enZPHa0vskr3BJ5B8WwI3UATrPtXkcH7BIlwddYeYZK4y78RYiV8QNyzwpGwOb6yHC5TrzaJI3wT0lC6YYUnJE+rPZG9B6Dy0J51ORr6/y7AJCIpM9xFR30ebROaN4MZkE+B8WxPBp7FqbkWl7Xo4UOBpcJfPCKkqoaU8sWA9EBchOrwJbVBDvx7ytEZoLiVCaH0hhsSlsw+qTyA74WRFSXY05ycZj83QynlCdWshs/pTOPXH/7yuWvKhkSDze/+cv00zXXMO0U6s6hPQGEbWq1HGRohV+sECakUioIFTg/I6f2pO27GfF1ACf4eiWrMJBP/cF2JrllsQc6v7epj+J9oKnqT6ncHpQWP2mCfV8rMk41K1CteHyeMbSnZhHYC+SrsLZIps/HhJI+wUyiNBc5YJCucQbEiF3MyWrcaeHcxYm03tItd08tfelrSFXRRXzkqNbwMMTV+1heskVO43akOA5tqddphHebCzKij+pOxwRSvNSv0tsJkn1u85aTlonlNf2y+vCF3OBWSsEId3hoWvIKeDjhWq8Df7I80oux1Bi4OJnjiksotF6KFrnfnHLM2STgsSwpE98CjB84pVa6dU9F2Gn1MO99163QduRtaMzodO4sPmEoMlNueBYJqvkeczkJdSzu+8WTjU0jaZRN6AkCJzyuU6xTK/jBX8JCNmvZbL0BQI62l5/AltasMseqXmSigJB3yO3dVXdKD234C1SmDJKqR2adj8ehBCAOR/MMNS2NXKOFN6HHa33rx0hi37rgAra6f84Z4z4StGUxcZ3RJsYpkz2gFo7ogs+cyB81JWdtvb0NpPYfbJdSyoXjrGeG9UDqvufiS1euvxSb+NogWjYQ9NO6i27aXjmn3WIf3VlvNQ4xZicpl7yMQxK8svQQgwzonjYQNCvaE6PYZT0y9b4TB2R5+NQZFPl/o041m/SsU+nXZhqgQhmH6eEJz35o1P9GERjN+62GDBKNPoYkM8kr5Cs/fVxJdNPjlC8MvfIcxZo4F0CXeaVdd64+MpOF9J3DMVFrRJrXtXhpNjJAKdULdELPLzcy98WMzv9N/crYMS7RVPSJmOWCEVUokViiATB0089H7Q9z4c8TTYU6EZy3jJIEbVLNRkoBfk9uMSqR8wzKTGnYsTaWZ/ZwNVThuD/NXgEId2ErDn0QnWRfGfyQnFxVtuD+QR4d+BuAxcSI2PAmqrE43/8QS8Q0pWjAubaivv1Fmz5bS4Kmlg3oEsVNqFxT3QofU1VjO3oGa+I1kD4DKG8dqB/SkBcdQM1h28ojANgkV4nRDRsO1QAEgSUxyk7hfVKK5D6y5O/e88HORKiubSaiwBlSSZht54PtldcIdxF9AbVosm8AXSUX8q2AkeSnYRCFykrx+0EOJ+wM61gMD9zofwLIY57FgXZWNyoiqw8FkiQbwmCI5+k/jDGGsFQWQtxcUvnXKU9q6X3dbAmSTV9jj6RxP1RNr8jfCnW9bfizpaV3AerWRLuBsMuaoOzhLcgaoAjkETiiX0yC59OgCEOFgOk7NfWVkGD2IEWcM+++qN9ND5LsgQJiq3e5S6e7hxKd8bwMcl07IOq7wKWX0XfKYXUD+UwAxL1uvbYpwDMwqGl2EGQfWUl/HFyRLVa1LW3c75gt+Mc9oYnX7euZ1nVzCafNjZD3kr11mKxiKeGxCvzqt/vPvRwEh81sjOZ0skEESKdxAg5NBBSolpa8HHOS2Kdf327HC0Mq6muZw8Q81olDcsC0yUXgDuiDx8SqseuIAX21ZHZyz8L1jGb9aUKQHp4yshJyJkGeVFyJRd5MRKDY5Od4k3V9gZsoaUQjwsDjRihaMdUdcqvdYcHmroX4byPbdJDYRgqde3wTww+AscKE0IUFYRFPmhOnSmsvqh05KFlQvqUUxOI2q/fHNU7axH+BIBEYY6Jre/PTAZ/cfIx1yWCDGBYuMo+DYshOeY2KOAcYuSMVLzl8BCk21fL9l/V0EUPNdtGJgJ7UcEFTRCmTViRZJz1ozNwWO77Mb4jgS8onIWAXleY8CAhdYkIuCXcdyPUQdmMag1BE+E74CN6WEKUhHDZMcLcnGKgqx1r8eTmInOgdA1MYqlV3sd3ekhclztPwkSHUjMKxQQoLFFK1J9KDAUg9CXYjTw47zQi8MMiuidF3un2XJ8kzWmdieiCSwYo0D5OjM6Hrj4nI4Xgn5GzGBXOq2814twMSoqccqo+SGv7aX0fyU2KqlWGsdZHYcVu8BzY4+qIREQYIIpkQ2LMDYZvgVqLTo1SOxHRRChk7bofvt1guHg/B8wd9v7E/kNTgvU+VV7WYYo6WwPpBxZic+EBsbutA5SEYpTZMvi8FxPoGw4WfGTiVXy2Kwby+jqW5rmD7lDuXUyla/DUERPkQyjhZ9AILv6dx2kwpesf0CoewiouHJmvsUEf8FaWGs172H4gf1RecOXJsbimlAkw64In9HLK+6RA/oz7mdgX1L+64u0ODxB+eIA3PeilJDZsANHiPOEswi29wCvmDBlZNm0V2q3zzQ1yJVHuoMTB/DHZRJHI9he88Skr0ZcpH5WoBlVF3a034ZpBDFsC/m+cJZz2YZM7C6mCGkse76PyzgFQCmdgJc/7wfckR9xuijLNIFi/l7VF4sNHyK/sdO557/APOpyUkPRVM3uRIBKOkYli/J7FAqQ6xVOz3wxiM7xjJSzN3Xumsn3Bz4TmEaAyYHCeggdqbQoVhnn8DrXRy1SvJCcEuC17Nk4/PeU7OUKRxXLXzQiYxtbupPjA5O2UZUM59dGwTLEDmAo1hRUp0fBmyoSzwi9FIlsT8oR2BPE9CTSE0KME1p9G5NM1IApWT2iaH592KlxwjYth83J70K6QFuIo5y7S4iAuLKNoLZQf2zihPB+Bd4ln/g0r6zJUa+O9w4MjGKg2Wss+GywTOWkb8NGyAbik9aiijUK7gtNbsBFSOpL8nwLfOzbWAevmXJ3DsAF3+/j6G+GSe4ore7+e28jQnZGRUu1Aozhb+7nquChlSOEr9dD8fhUekDoweYXItTJblsIjiF8Ds2Q6UuwLts1nzNCkqYvuScyOd0qMIEsToCJqWb/08DgCxMKQ8F+g2Bg/zkeqJIm45M8OMVn6uW8V5YqbCxGtQxA5BUm/Wfg/NBRxjOBWegc1SFTWXKRHGiBcqDv9/7vr0VJyMgSh82+eRebYE0+js8XMMhPGvgreTPkVvdokDEbnS4d8uOlb4KpEKLoo1Q/9vFkXeSnHxiALvGZF2tzIlmT4R01nFH1I+gU1GFcB7fq6E6uruChSc0RVsUb6c1d6kbFYB/NiVidEPnT3GebCIn+Os0lpkvb/EL3FBp3zVnkawUXRKe0Rf1wayWRrXhgWspNRPypJ6UXNhK3p5asP8f5j80GFBkBm0EqAkqjrmN6mB6mum0bVqoU0wyWtfgmVuoM7WQ83e37QWYyTgU+cYJ51FNIAz1ulSy5dBEGjzA8fzTtEDhOLbUv3mlad51n4BsJT1SmXiAncDriZ7reK/pTVPVpMciylUjkWHS2I1FEtnHioQ6+qLeAhcNz2ITXjm0BRCEXDOcdLmmWGe6g+O+2GRpzQrpxrmJ6aKvwEUgqExsKiM31N9oxdWt+KmzvdNngRw6KQ+Wb/RFgwzOeetpLIzqWN4+vPzEHNkL67JVv18/PID9Ybu+PPgaS+6oopZO/LFKofCQe+nWpTQWvOb+uv8FHvQmholCF//UCRgaLN89oOXZn1f6pw5WwJCwH4iUpuetoYZKdQgpOSplMMHPVK0uTOPcH9KTJnUbTCxIMdp1UxHvJuQ6sWtpZeAenQMA5rcs0/RzOITMp5rbis/mZzbRZfa2zENFOH9+Su53ctpPp6/Z7DEo5KKHqfS4ZSLnNz/xXJipt1zw4e07uAyHvJraqAVdQQUaIYKmzhfXml6mQtVXrqYsxbQx2tAncRBU7pMqHEcWNSR1MIHOvT/vq4Gxryn4lAjwmoOhQYV1bNjA79KKcCwmG3QQhyUrh1qEzvOhAq3a1mER5rVS0PGq8y0xl/aKPluTZwFSr20vVmAK27BC2Oxuv0FwhCFupOz/Zbr/ZS/Z88ezrK1p2wf4/bEOnA506kJCWVfieWpU3Axn+BYgabM4mjpflbLhNHQ68qEPUK1wWctbtL8kWJT8mk4t0q0VyFkVtQ2dEFy1aclJQAX5paTUquy+XFl6C474UT0kx0u+Vbak6fVPNcVws+DkAupRXAaqr0MzW88IYSFGatxW+jVaGRtMcgjYjoZpszT/09jfOSPBo9oW/bp87Ru9auFtGCqOxPGc9GWe4OIzB+3eE4RfQOeCGGi11HGUrWObTC4o934+hBqZf9hHH6sFWFZvQSSYtS/o3UEUL3zN3xU+4Z1OrASvDG2zowRXL+eRzSz6QXeMmK1VvjzpnoGqvkSO0lSuU0X6sp0s2woCBPw73UeJcAU/eKd0+FkQYyT1sgcaxJ5KFMJX72m6pKSHYKIvQ3Rza5Lk5KwWs9u3B3YAu4G+5Si0K0sOY+O/S2ZWwXN/sUmgspb8/uQMuDFHzO3BUYeWhsYa4+LP0XHJr2jELmXeJNhchUILcrho9YhvOz3ETLUaq1zgDz67jKsx+OyTKTEmhHTmG8TB2IYnU2au4RZ3BvoNC/D3oTRzLtWK3YG+Go31bgX/DHv8yThV/+QpOfRBSGzLTvAsdkD6xcqYqEQZFu4LaV7sNl8OIzHfaaOiUCtcPqrIWmbYGDlAOUwss6hUHMPkDzzFUE4xOhuCWukSQFg6wGK0bRCSz8iXOlUmKfMgXXA680ng2wJZfUkaB38RfC+b+PWgMUu8juLe0tdLUVhLYit3AffOKNXNezefQd/JSKXR6OJZMpCGuB0szJ+CuOqnmSoOSnM0jRc8iyELABjjdZFwcmVDYvkawUuDVLh64EPTWj8GJYlIbwp91kG/BOMxeWq0iMjZMM0QEbdA52yG5Cm6ZxaNkJkwCeTjF8eXMkZ9bpBnxBuagz82EHYuOGzKWFtVNjgsTmn9lgbEjybl8Snm5L/+D+at3dnzKe78blyHOvHBDtTghYlpA5LHpx6hVBnCre2Q27Cf9WwHCVSmayl2sEJA6wj35K3yzJMQUD3jcaA8xITODpS/0/A75x7JDLz9Tc176BEngDmG2nZWBO2zvJrL+SNOizowVrOJe/RoV9nAtJDXFSCyGkOBtJNVV9ibedZXB8s7B3kT+nJ5xPzg2LEVo68Qbo75kMs1SCyUJGckA3d5l+OgYvG8VqOe1ierZsfr0sKPG3uyRJShd0eQAKMX4zbBDf/iRlXh2EdxnSiGWrfy6LknKuqWCas6N7XXmFzl5yZ4jsPuk6JT1IfaTkLkJHuHsXqCltB+EP/sSvU9kBhipxg940kbGgM3Ltqr8vj5yJ4N0rgIeZdbR1CkOb7NRTBq1LuvOyJvaAiX+MlOwMcE/7aeLmnZ4rUxx/9Bb6xpEBREUskIf5O1+jEaqR1Xni+7r9tsl9WrWBiv8qmlu+12dv5sMvtMnOHD8GqVT5MKAjZJqPe2FpyQ7oKIpX5+Pi3PmbloGrfjiELl702UPzIy9+PFs7o2v4uOJghooqpYzUaURos7FDXruac9zROWC1IpAD74jVNuTOW8z2oRyx95f+TJ/JbNK5ZURG27usO3mVLWSg5923jQvz9H81Vrq40GF436afNcohOxpkQVU+msTA7n9B5UR09++7gU8BAANlNCj0x5z/qpDsvZGk1TbgFzVs620NjZFzIZh5d//aOYhTEoBxIeDFqRM/wFGbn5vmFlGWkOBdbMvF2lxH9POFj6yazOr13yO2DmjC6x9wCyZkl334kpq4eTNtjMAzBi7Y5Ra6ueAz7MWNjv6ys6X3nn2nn5bdFx8h8jijsoviR8Qvnp4B5++iuJcQMFyuUJbwskNJZJIPPZGwEg2v0BvQm7louYk8rmUMdIXFzzJDRmLubQcqFJk0Xf6SqYbVX428efZcbXv7bDiL01+4unXKv+Edgyrt64MLfIwss9Djk02szzyXKgRoodXeEZB4DHH+jIyMD8mFihRrNNO35A7hVqGgsbNkQB8v0D2hwO5oDnDDrblpaxy7RHgbodziRf3GIWexQLPfR1E1pbTUvzi9rQUw1r8zgPZdDhhoGYOUzV14Md9on9vz018Xo94NIeIS3UUCs4UIyCLDYVY74Wn/euaCSDIaBq7VkiWr3yv9U3ULbVXGMlK482+DmjjFcCbPxCwS3oo3LvwRx5b3gE1YxTYj4MGdY0xMUvxrO1c3EURN6zzCGDl12kz86rrW4eiMjg9bz0lRC+be5wFVv8NbeLeZFqXcvo0aQ6+yUVqYLkbYbK5MR3t3JPPNCxhmUG9vVsEve5agQlPthvSduLp/rD0vbFFb0bjSgF2APc6/g7z20Hxa/Ijn2/2+srfmafmudbiVrD4k9S+SeAuR9ZJ3JyveQc4brJFGA6yH5XuDGIAIoCV8uITg9nzQWW82EfmvS9RPk7VeP1ZB5AxhYeQzpwuyUHxKF/Wl/JtN3pBmfvs8jlgaTQc8/7rmkoVl93b3YXckLFzzs3wh80OParyrU8dmkiD3CRXR1v1awotSHGnDa5amsKOX+GaTu/PYxmaZ5IGxLVx8GVGQn+KSRF52MYa58QmEGQ/G7d6Wq2AZBIWzo3buQTPmbskfqnwfV6027m2J3ttylv2qX7ZsGRTz8CkK4BDKde/eN2hrcICvtpg73z2RBgZKnE8Mhh0wjintYk6cmsZ78hP09T1V88cQzWZh7z/4Rlekd7O9DBFp5gTVi91mW5UbTWKp+cdsfAEgnBlGjuafU1Th5liuoYnfmEYwA2mKxBaQO3TuWMyP+MhTk4a/KI1xTtd2ylJCsHxA9di523J2FdIz0+URvAVYKznrdAAEP0pwBoifCsTD8RfPgmuWfN5X779ofsjNSUo5GTOlrKgwwEQZXfTEgE=
`pragma protect end_data_block
`pragma protect digest_block
3b5728638cfef551c36fc8d6516639e5283e5b2973df2cc46e6271828e18a788
`pragma protect end_digest_block
`pragma protect end_protected
