`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
dYU41FZo4CXeao7ehcDMtY5bDddCZ5KydkDPaLpI7rbhZ9eo0s5OmxXngbOtKMiqtVfXgSQbMKasNp7256SwnFaxfLZu6bhfSYfSxBgbCsdOJ9Iv30sm/P4GcnpegS7+oqXdw034Hdv7BHN9irZxkNhk/x6ymkXd5BU46qiSylTr34jp1BJwCCYLtCoOPriUvcuf/OFERAIVsL6InCKze3Mx/2H4YyIAxR5KcRX+dta+ReTGDtv0PNPHfmdgdI6JjmzS6RKDxA7FurC3GxeNDG+VyWgWBaVKsF6J39Ru1tRpq+oHXhWUjIn36PYtHN28qMOJCPbTAFXEIHoh/lIxEAaXLrt06ehpu67r2HjiGwhkCZQOHFCE63/nYK3dxpyxJeVN6m7wu2+wrqP4jhgFcEKZ3OOwarxk+bssoMBLsbMPdjwOPNkK8KJ/lXL4DM6A1g1eqGighcs0F30lLi+hFRSiKgGaUAx0LyY/Gqoz5utgDWdXzzFjWJqrk0na+6tesvOARL2zhyDF1OByFkGEvq9OLM/+sDMGO2CfAM3yjaYlNE3zd/hEkDMKXHQkK1P7EDiK1LxnYzrWEFb7X+lhrfkr5zrQzXOmI2WCs8jfBmhk+WpJXyQS9UmMTpUeHpEKJJXZHJsCEnKcB8KUkJ6oQAr08F4qzJ8EgvFMYvlf7h9NRooZRigx3zo3kFKWhBba6AELvu3RRy64Ke0OHmypuxBNC3FDNOnqeNM3WUD8qCMCg4uSJ3dsNPjtsNUd/hhZaLzrEh+DCeAahqYGTjl5+XeODCY9AFh5Ecd4A4D+cURm9ifpbd0Wzh7LqSjnKbaCkqFPlrTOvfodKu1UmqwaT4q+iQstscywV1F2ikfdR7oGbD0OZtDdR1QYWJLfRx5Tl1sfMxP0HRshuPeHkgGhD16yM2EMuQQJInvTmonLcEx/FOncMuB4h1QFmb6i/OCmMJE+wNXzPINsW3dk37kJSjOvo3rhg/QoEow/uxeS61cm0qNFQvTTeZaWg6EteTgNF2BA+FPMM0EWNjw/eQuDesSO2ynVT9BuSh90R8TlxM2480NN6+uDszyfWLPheKI2vi6gxgaV1XSRppS+qkQmbOcQwRyEagggCCbDKrnBouqY0gbYaHIlZnDc0Ru9SjrLsJWnmXA6TmO++bIc/Xf4nKK5F3WROW1GcNLMe6XyB+MZ4gWHKMfo7Q8e3rkF1eKk0sJLSroEMbLSYcNSEAL82Wo7iiSyxcN3KC3f9njlImIgizAZeMvN8RdKb3AhOj+PdAqrasQrPUXvv0Xiv9039e+4+HLUCHSntg/dSp4cj0qEHg6CLKJIZRYe54W3gpFoifFoSpwYSBPV2I3qikm4sFct+/LWA4EWyhP97qMnWnAjQEcsK4KF4WLwhLNNjHEmd17SuQz1W8WNY+kz32Oadk2a+0s9lDqz583uzlJ+wSHros9LOu0lXss1oGNW3MlHYUlqBa/K8x4d0Dxu4J1FahfNasjDZBlJVfNUPgZUwhXicRo+b0kh8C/aXw8FJh3I5WDQDoT4gEtNqq94bHY+NTY673M/70LGKGPgOtRD6AfDTLlwzMDbXovrTeU5xIoBwD64ymcvYD9Sb6NVT1xtqDSe3QazZYgQuJJs1ETWZCYHPAuOiHWJOQGFXDaTO+4cGcJX6NXX+YtKrBLIvPxXKlHH1u3teHx/dbU6mm0/QcLmZCdzTU9jjaiC6U7kN0FqskoqU7sYPi43FKM4KGo3nDaLygEgmzTqWWry6DmejEiarVVqnfiJIQ9aQNgma1bplAi8gHIZ4yldIUSqtZVPNpnL1y8oXmRgz1I/69lrh0B7j9RZwzLVP/TtD70boThY4doeuNrYhqDTwV4guxC4y+cTUJc6xC1GJ1U6Ucz08ZIw2VV74/GaN2NI+Ct8Yp/OXdpp6YfSkh7prZdYj6/+dmNzF1uRPqrt2W9Y6qE7Cbwo1pDtnh2IiRBmq8WzKblYDmrBlFcnk/XBLqLbM8GZ1aIebgkZ4YtJIFtZveVH6t9NkUYLWA/li6ljJbAK0AxygIfhDJZxYnNznr+zTFSoeZiqosFFBzR4H6B9nRuwjV6DMWY8PSAN5RfVrKXx2eqRXCk6/VNoJS33yeTh+HMlNmNx1o6k5961u4X2W/TQH2WWvYiJpQTHffYLXdmcKV1MafuR2MqPiz7uNC3dYxanDLDMnXCGYTEHkwXpWXmtoCzJPsWzm9jn4RkSyVczGuf1MyTi+q+y/tTLKyp75kOJPtZiT/8rgR+hE2BZ5gF0X6J/tQFiDp6lZIkhNvssxQNwhblduk9MjVMsId/UWUMtwMlu3d3nLmXy5PE7PZkarsza9Eq6kBJOXNIrHDloGqZXix8cwa67esYvhffXNKE06HpPGhq113lVgriVjJY3+/SFZLL9OaRqur6ZaGAoGNS510PAS/NanNGjqvUE0EecPS1TeGLZodTwC8EntIVwcXpl03HzZIUKT/JyAhQpairD1C+wwJsu6V/hCrSca7lWfztTOwveTH3YYo4j87M5m4vdm3JG+w2weLxiyBnRKuCbd7ZCWSP3dY52cXFpdLlFIrZzC1fzEbn3ktiyW/t4Ia654YIIbVF6bwwovGIQqgyqOW4FIifTD+RpuZy+QmLerseDvwbuiNk+1txkYADKoZ+ftx4o/N4o4WALNu8sb3BDBbcaUq9TNwBU3zWF4QG+v+zV0KrO4ELdneTe5rw2bSwoawNfzFxAbeUQ2IyIwJH+K6i/3nrSlG0HcBGsMyLc9cQf1+6ua7zzHdmlYSuayN2t4NUqkDud0p8EdBwPuSHUG8L/Hn1QH91JfGZyavOIs1JbyaDqFSFa+MBQOUGjjIBW2I+GIIBrlyqWQbXsNCzG9/SKy+33vTHCtVZjFiscwqaw2eFbUpF043mlPB7xx42RJ+KfVsRqTiiEKZJH+CC4RBrfv3nZv9iSVaCDxSLrRMWc4noyqRzIOy7y/u3FV0KXovz+NDkWGriJdGogkGGSSNDutkhqcJD7K69w2VknGHuPkaFCqZintVvYgTNqddXYLGUb2jQV0C5IDmju67kuamx3948VN7Pv9USZ66JgUDj5CpFLxJke22LDFpyTKDb8FITR5bWyMPMBOHEMsyTRloPFXI2t2Q4yRBBCDpRbb3kcjHwrmk49wCgzHEHXd+NfZD5H8s+S+iw9gGK4MnvPWLvpXdiatNhW5XKfByzAbslcCre45HdgnMRp+ypfPfBnGwVB50+Ez+aYauy/MipefXGg5TEuDghMfqixTEn8K4qBz49e2fujjie1VvcyVQ4Bc1EdwwJtu0fl1h0+wraNyBS/QJd9ND0s6Hs0EQ9BXFZrwXbkIt1wU74fLt/+ts/FwBoEdnTcOyEjPGyS8af6/JKGUKuOxSc4EIYpTiirBW9nb+86Y5C49k9kvoBqrbzG/vf/D7A7N27HwnkN3UZWDKDllHRLodENQtSzDdfxlQsENK9ZR9YiptyxREpePUOSamtCuI5kK06vS9Y/3cjh5kr0ADf00Yim7lZW6PvlCQwFd+ZpM33nG7mVBeMecJn8SttPNbh9QJ4IjVkwLljvEBs+lS00XjyZ8E+62WuX0vjd9qo5XkEW8/xZvn4uJm+qq+AMIhJl32edTZmwabXVa8F79To2a4Jx1dzorfLDqRSQ0HSfzfkpitWymdbvYYh0Ix9kyGCGOJh/LbduII3kBGQwiSmNsK1GQWjM6+L/kiCcgOQUl3W4/dZGV535Zx5dLHUZoWi4adKaLPR46d3RE+ofw1/yu5nYqGgzSrgzh4VgtPs5qC8L3JakOfcxcd8xqKQKiZQpmjbnG5FV2ywGv0qlA7jEZaAB8DvgYDyJpZZJi/WlSqyiEKoHTA2kvruP0oy0SGOzNULV51twoo7i/FSwjQUrS5JjLYKzD/UZ2pXUsYnA4X4mxfi73/0x5Dlhk1XZ6nwpKfe94qjQpdC6pao3pQKintvMu0x6CtWAcYETonSUJ9VZgofbl6XpbiKfs4CnjTjMiZd5bVKNmsGFBzABKZW9HzdBrX8zcGZTzkfkoqORNf23M+boFCXTK6lZbBhvJCaBHORt6PMgTgOo4bqAilKo+tXLcDDQczUTirMboBdKGkvgS8Y7sX8U2vz66NCj2uBtJWZ9ExRwmZooV8ma0r8/3OrJ9vQqp9gqjolTFyQgzCXi6CHbihykPNAjHLPzgE4EZLEbgO0idsyhFouhH2aQ/hvlsINVEnW6S5znX6wAqL98mLAsmljF5uvj5DzJMn87RKhyQPqZ7xY6iP9RO+MO6GX9iMupvMVH0SwZlMhKa0BNpMieaUzPgDK59Gwv9TPdai4s5BN6XMyxWfyt2nEVdT7jVThXyAT3GhzOu+I1m2s45Wtj6t6yveDA4wIk9zay/KQVEFKpa3UxiFiYO4HW8EC9Knp2jANcLSiG7wXGe1pTz231M4foxcgEFKQJAhgIZJ7F+j8WMQQRLcuCkd4tYBzLACRDPJfiXxcJaMDdiHv4myCmPIS3W85vCwMqR+R+86rWAOPabmFEgGMQbNbz/KE//XmtzIaQILdig9sLQkWLSm+hMT3bbvPWn1/+bCtPiPoW86wUxCxQlD/5EByNtCnJ36PNcct/7xWko0q5ioGqIdVG1j4CEo0VCVqldu+RKo9K+SWb2l3h4u4eodJ5o0GcQFbB9zv1DbL2AeL8X6J9+iR2FYDRyJGg8F2yr3k4zY1tXIwqrq+VNfLk2iq4KLNnXYXdyDHATBvId40N/3OPzvtwBdHliRJhXyzkv5dj5zWO2JTDNs/3R3NIkVhpIyz2WEdZqUmw18dLKyISGsAV/Y2saRwbbYLZ/oz8e7p/pb2k7iEg4hcA5tkn4oW50PcySxU5cWnN6SQ4Bwa9ftf4N8Ohg/Eb670Mv+9X3qT28mQBWUWFjUySZf2OjJW1Sf6UMIxh8zzRKbXYhGecO//QRsGg+1ptuIl2KGJVADzXyagSbPTv9JTvPzxQSYhNA2S0U3h9gwrodftHjjLjOJZq8oOVvj9CSDlpfjSlhQhcvBif/s/IEN82m7c87l6isF5IXzVsAj/OdXOLhBukEeTZrJNZTHrw3GCMEnRXFutYA+9LjVpnmY4+bJYgAsOoIP3trh9iuHYXyos/c7m+57ufVWwNwoJ3p/+Wj51uQ+MTSwjWLfs5v8ptcmQdhoSIrr+YP7ZlpLoBdd+v6NkgX4o/NRbJ9S9tVLGLjBBpgot/TZlWZavdYCyAziO0BfIodt9UKK70r7hpX4nYvFXTcuyto7kCXGXs1wKjmQgbnPI47x/ocL9mlGpLTvgSPnRvjnAqi4lNnqu0U0DhiNXLuwkPVaa5v09ZdsxfzVU5P2ZaFcVETCfYffoaL1sLTYh0QCfhIO+HycN0mlLCpQ6ahGHO4IOOjd33tcRQKptlq/+1gjD3PoDsDlxH1l5hFi3/x/F0/u9KpkJPA49OcGm7A7sTYbjeMY0a5fiOX4B7KPzfho+67muf2nilBIl9i7SUxtjWNG/daCnN6aKxTMGrxX4EjYcozXLE+sAv1AYybX39iAwhMkY8TFxqpOUA3dsSXqfD9TOAwxClSlv8hUBXj0jEa/F7nUjKFYNwTALnVgNG3fJB+A1VSj+jH3g3Wy3n68x9c4ZIUcmIBwEO7bu5/b1Df0qIi0c56+blQBFtOVj00XkHDltb/aRcJu16gTF11Y1ehfxxkYEkORO90CwLvGfhKKyWcA2XMOAB/7wrHoySL/coqRMMLABYeeuenIodRgCjwdaUCI0iL1BSYJVKOe3tt2P9gwX7WipGlAmzyqEpP2TWm45Lg6EARH2KC3ltxJXaZRfASs0Zu+TLEeEbo/czxlk9sOh+QjxDXXrYIpyIhmv9Y1rFO6P8ng6GMQfy4s8D7rZpty9/Lobi/IK+0uTLV+YbpesDAb0IxtbwoZl6xOtH/yr9cd2We1eKaHJMhkSa/KuJYYudwFoeeuCY35fZLB6xTfkXtulGcM+wWQ4jE16RJwbbqw9bQ7oa8G6A+t4nNGHmGpSRt3vXXySWNr0/zHmooqoeElAusxJGB89ogh1DbqkZeuEe3lGwL4X+iqsfTly1dJg1dueJcKxJX6j8AXCZp5DHykx+pf7nhVyN69fdABAL7mihJyXgSDDOgUCYLsc/LiTpG4EhsVaJjQEiBctArY/RrPKoC/aIwJPDGnPtpleYKi3yCrv2kc7C80wW3NrlQ7rSRrzAvBV4FjvaYj9BT7+Sg1cmtyr76NOkF1t71hA+VrudzRtYtRWxWk4N4v+8iPhw8HRRf2D9b+nLxGD60DXxl9SnVD7Iu+5rBur7/1gF7X5vDw7GJ99uoxGsj+AH0uuMtjuGiZlUiPi+OF4p6UnFrwCW+mIxw+GD0wIt0xGLCoaVxFKKwe9jSzXBY8UFPq5pZYb1FU4yPAMaW9lS/Wapdn7Xdv6kBeaJSjS9FUvC60SVG+uRM+s7+I/KVoO7VdNoxKz0vmS3DOUOVd9arfFbRMSlaNLwF7wPlM57SrSTtJORYsv7g0Z4nmJm9YSDsxjLlhblCnpZru2AbOjsFJElssigTEr/OOQnvrv0cPKQdO3hDvj7yaQPJkKeLEj5oqxTwS3nqh5Mvb7hkdsr/DhpKiCpRv5Kf92yb5CwyOvfAdmaILVFVaIz1yAIbxRHxraVCQe9xwNahH3O41Nd5XLyVg6C9v6MP0VRbIDA5xmpVb0XkvsdEowFoHQwADZ/Wc0sJaEbCZcbXKPsaHhevTc0Ee6CNEVYv9wRIiJ4WgyJJxLZdV8Guk1EKqszZ7aFCmd7ClZcxC4X3ACEstHHPl2/hosWCKicEF8st1xKP+PTqE/kyWEpYh7k0PPZQecjD2n9UezEkj7c3UnX2ciAy/vjF7kMIhD0vtC/PGvz2l/LIQjFM8nqv8Gi7nv9HM+yqhyj6Y+iyZcHEu8pUUsjRycoImiAhoCYErzzpVFng5ALimwjjR3HQUN732Bh65cp/WcjdPWGoA4WYn3Jfthaa57VhAOjw4hFvduE3J39m88g2pl8611DSCShrpKbJ7EemERUApo819Cw4F94MZqFr4yPq+8KTPwDYdFFUODy0ot/x+/1Btj1PgQk1qFYn80ic1CccXeakQKJ/rqW5Nb4oWd4rFANVN2BTT9Avj5Tqdp0SLmi6WAzrdIZ35BeR7Qalndtshe1C+mWFJ+4UF8BAQFiOq5l/21X2S6WrCTJizf5U+tpl01gictwyjS9DIvnsiBgOK2BDf92L9wFYta/nvbjOGAdHLx56dTkbpN9/KiVV0qebEfOUZxaIFqbP9obfH7/aph3TiXxciclGpOCz7S/cQG/VYdAyj+sUniFb7s8HareJ2ZRTG6i0QylQvoyod6kxMnUZ/P9FOq/xjIW03rH/maW4AVOsujOdurqQp5zloTam38kZJHylzgUXYeuW9M/wR/wn8OlIb+ktaQXzbua/ur/1eEIVusu+Ekx4p4hRE1XbcXiciU9GcA5mWe8d0Dy7wrwXLn0D92evKnerPQb0b36aBPCCuj4av6Q4/22ydkz2OrIPz+SNtPmYaJGEP+qT8X0ez0m0NJ+VGNIt0ljw1i1741qJm+ZKiWSTQprU9yBOFRHBfPpKsU5njhnjNnlufrtXdP9uozYvZ4fFgyt9qbSeq0ZSBuQI5GxGRVB3Ma8gCfJhzlRi2CvuOhBJhzxJiHrYgh5StyBvUJtGnNZlY7ObNEBkgCbvNjyqBzw7/W6ffd2daOJBaJvTl2iTkNf0qDqDzkjJQkLRbx92sHiievoX6ay7EkSYtbkl6cWznxs9jAA0wQpbsQnWCC3YTFquE7DKbYADJBweahBavVTLj+iFySkETizcLHR85hQQ+IECieDuW9WNZHj/wkjptF2w6Q9s3DbksHtl6Q6TbrDOkd5eMzbxtb4ZLlZUCyp2rEpBdSD7N8tIHzdkGUN6GKgke6VC6k6ppdtd4MHZSZfAcEnrQo/9rGgmmnHCKNmDZYo3g1cLxZO+f9nj3DHQPS54hJwf1Dk1qImf4sR/L0GOKh4nnTem/R2wd1GuV2tb0xtWvFkR2Gdo6hrfWalDeppeAZ30nCXGmviaUuQ8N1mglot3dFYhk32MNvUo1grlVCt38scMoqgoXSoekIpPNeRPye/Qksf9dKts0UzMaorz27w8w6Rh5y+wBFpoqi7lLKbxjLHQOJIjUZkI03ucZaUyT4ecSMPQv38DNBUaNT2DjnYzGm48iFLS+u3/oSls4fAKaiPkFZ7AnmQbf66UUisbhmnhB7wM90ySXzrucIN+Fr93btPYSkuor+phFI59WzR4nkYHGAJr6GKHtddamPbPMT6Zy+Csk1e33+y2oahfLcgEyMO9dpYXsEhrpT8eUyd/eTVe1DlDDqr4t+ORWwIAnoqlaw4GCHmduIxt6oteWOzqv/qCbw1Z6ih9yPrtFMOSsmvFAqGuLkEMcGXTHykoleiiv3XAgMD3JF8Q5yMlKV6wT6tT4R07RQnOrHWmTmfb+591YhDjFHHD9JY3roHLZ8Qlj437vbqy+omsdzPRuZXuScb+yqqOGP1IYrvEJqLwnYXdcZE2ijRHofEPwGeVDqM8CCDzDuG7z0kUrNdzCE4OigUDQW9lKhH3MVeUV905gJWp16WYNWAVOmDLWALRzSmyW9prGlPWrJf3AnR19JO0EwyoRZbM/gZoQdfl+qeialmky/oi0tRJeOUttAQLc+FOrsRcGa3fGt7vr31Kd5jULOYxQ3nlXKDM76Ee8lNTo1g2erM44xfS5OLYKunBCBm+2Ljkv7d7BS+YzGC4w+WraK47Bdb4TnfohHtu2okZks0zc2IL9l8QP8Yhw1u+aIecjlklNkDSNsoi7w4gfsKre47trk2vYkbfFJil5qdlm/iRjH2Zah2iIgo3ndj+Mn8EGAIA8tuCNUU+rfK02liKeCWiGADBYmAYRVBvHiKnBthbp9kWWsfN6Ff1AnIC8zV7cvrpZSNmrbkrYAFZG53W3p8O2YcKUfqAczAXa9jrmZbO96LkNbf9JhyTvXNZTA5NJ4JNEBtXLqwpCw1auEZRYVSInxbrBRGqx+kZigasNSmRTMs5J67iuY+K5omV5aj1GAjdBADoZkxT5uPVdncI7wexfqU54avKrmr930zYzv1qxseSiBljEO1oF/JCIha3+XXSyG9KVQ4DbNeskQNG7g997M5EtvBTAqGiURIiBN6PDkEnPMOnar9sapUV8CClc9aqZj1QFmQTrxoZbf/LbFFetfQsyVyzkuJy65m0w4mbvzYsI7u5vlD2q7ruowdzAdd+3MaaHUNt2ZrH0FQ/Q6ybmdxrcDEAmf1OTj9RX952+SddKhsX9YsFBWMMBaHjD+dJcEpmEhlW+v9paKOnT20AWBYLKLWhqQnvvKFuRIeXJY0Tzq6JtqQtSztxO8C6E0saHjaMv82bjU9ViY7MVXbTmJ5CE8XVWRLXMK2t1sqJ1tQliUdfkH4e69tgcM2e9DFyHVGLQ1REhRfSgvXcw8P1CmuclVeUSkL9QP1ZhCXS/U/TOwxOlIATa/2LfEUVYI2+zICymcyE1w1AlccwxWaFOVM+zhkTVVdE5G1CIfy0TmN99ZViGzjAsAH7oBk3BJhBQTv5NINYM4itIFw9seMlIy1URU+bUUEWYMXwAN4i4CLP4Kxt/SyLmWwPHiZ1o2f7WkwbMHVqwjNLVKaYg8QOLxwCFsjl37KG4BqlHrmcL7kuUXraLgNK6QBsln3t7UA7CajoZ0ly7HazZdvBaPTrMHmh/OXXL6g5ap1UlZH7PBUoGKRxw5UoVUhmoHzcz8drXlzTO8yll1U7bHcJ6Cxk5L5dNQqexGi851U9d52gOs0FwnnQgPn00VpA74yMEtdr2xJ4PACb0eU949X9Xc6LZnAwn73TTACJcmuNv2Di+hA1jmVkl7B9yk6Zpb1jDi1vHxqtvGj7oiOgRDYGVBB8fbqVmqB6SJQUOqOwqn/wVYFl4UMwER9mimY6zS6lQyuf4nlUEMSV1Y0266lm4hegeV0a4M5C/9a+UkTYWBxRlS3WJ78y8Y9thXdRn+gmWC03YJ+FyCVL6SEsO7rbyIWNUTT3DJ6lh0VqJNMo7Qa7DfgYTbp7sQHPp8pX3FVyaCOWWDztaCkeCb+fAmjkAhxn3OV0EOxubYK51uyDAUmA1d/fhR23c8FjCGvMwNUEYoTlUUFRk7AcEepfzZhATvZ21ruKx32igaY7nHpOONlfQqmIwug6Oy82w8hyuwssXfcFp9KvYb/u1VN/lxl+KUqoifL8rP8rOqF+eQQQ/roVA0l8BSM9WXRb9sEvaUxEFuawjrjsVebiRHdBKPDKVhc8Xq3IwDD67RpVYHzKXgryIqwMqzsM2k9EhAyWwnarw2HUnVzxojnX4AnCOY8X6jyMQlaMMwoOGr/WtT/n9IKofE9FiG6r60aWeMKsxTixse0QELRko0oP1bLAJyEmYbIxailgazDKux4EwiDUw9SZVMzQdymTw/ZYQ+2A4h7tBNsxiCe/5vX7ds8023Ps3LKUjaRwLLGkSwRD2CRJsM7FwBQE8/vMLAcc1nVq24rZDLHbmCh1Ce0fp9rWoGlob0MmvPIhZxKp9amSaPNENhaGKn+p6+c2Kf5EuM3PDW3uWr4I8CNo5XMR4U9Y83Fr+grA4yNzCvT2ks+x5ZzC5HaHbiLI/jzBR9Cjb6eeMCcVezXI3g/YnLwCiAc9RrVHdKUvnoM+AaFBi9iLzA6CclPfD502i8plR60WsCtxIHIxldnbqOglFAhE0Bu9Hmh/wFf+VNcxIOVAGgl5+zFBJs6WoK2pQn8FdFKiu/FXiVM69CnOdZYBcQOl2Y8UvDfv5AyGXzv++OaRF2qQSKXvXyOrjR7kV7zCY7DjczCmMXHf2ZX9iiZ//MQbgUi8Ogm3SqPn50BptgERbemY1z3e9gR1DO09jAOSkjTQ29v5j76PuQ5W5D3bluDeQ52CwW3oUylNDfq5bqBV9K7oEhBJuiy/NPEib7Wohy9akVZUwj7d9gK/LhcY144VMum2JegGat35xrlv+zRJh6w9XZJ4gN5h+5vNRf9cz+lV5yJXmEUvFn2sU7jCMX9bDaaJ4Gc2/Wnb7fQVNrrihso3/tbwcIjGEObciT3wyknu8n+ohF5/q2uM0UWH/W54aStrmYexKpuxwb2Ox8yaeMq00cc9Rs7AhWbA72thJbr5UfRyGZqRYSrQvtnVcQdZlz1cvIShD3Ux0hb635Ew8H7rfbBu5QWY1NGJjxGZql8HZnUcsrc70+Zipl+Y5mH3msykF3n+Hc7dFVIW2cA5bed/hgBX9v2b0sZmMZg4uy8MSyw76qT1Dry7rZuSWGSFF8Mcf1urQAYvKuXVnFszNvprS64kRLRdY4tO4Nh7p/sG67dKrctt16LKZZyyKM9aiaB9Aq/EdkdSfF3/VKOXGFDVjSCXqNVvIXS/bjAGPCLUQouiueYcr+91XFacbyB8e+Yjo2BSfzpYDS0cS8fm1ZaJtbxEQJ5EZodKTGBvW4vuCPeyUBwzbPtpQPlkSNAFTwL58Uc4gsM7yGJcQE/Re93R+Z8pr95HNiGk2C6T/hI+gHzjdb1bhcTwAKIzw68yLT3uWB67CAW+yTcqdr4tzD56WvV8phBQXPKhL9fAsCYpTMVqjX45TuPsrUVYXHLSaUI2IXpXSRZzeSZJsoDfan3K5fgbKoBc70myCk1f6FQ7bFQFPHGprM3/BXUaEeAtH0Rz72kI8DwaNi+A7i95bb8csmM+7ZAyxcqkUJsbgoYczbLqx7s6p2QQ2haBcn/fEAIfljr2fguUrBEJ+A/5Cz0zLLF4oqxw3m+Q3ku6dd6OnmTNyIwlDrxnDdmMzdxRed7Jz0S9L4hZdcFhORVCLClhR1GAhHqq08CZQVp6c+I1sY2ZTz432MUli3loSs4TGnoSseOeLTvU0TT6gmzd3gvtL3BENP9XtCGdzatlifQQEzxvNomfrZCW1E4PWjJW4PYOI/blTe2kq0KluNjfxUrT1AxQMFQ0bcGbXlsvnJY3btpmJ1Ag2DSAvIIBLIrCmZ4N+/5sXO+hLq5n78cW6V/P6tZy7Wwf1TpTK426KhZmS42VsN+wCuc/hOx+KK60vLMqNeXOxRdixZcdzGlR0Zwha0taGnJySdDhw7cAeOFPR53tuDoHxl7r9HOeRbh0Czhjhz2ibEbkFkjFvSoWHhdzs/yuL7q1Lo/ZA+aJftIAhyCEse7R7GP35zLb0n5VK5IhTnfuVaNV2T8Azu41wlzGx4b8tBU4X0ObMvls6lhDvhloa3/Pim0vPTuo0egbr7YNYqTTAcszL+Pkzp4+rlNFOzLxY6D2qZglUis1y8m+KaKRukMPark/g6CRZu+GBcZDufMLQc3VR58n4YWycYKPrQcdPQ2OzLaflyroxJNmwtIA4VOfCPEgBh0jyuzLGpNJQ4dx8Cylg+IvCcgmCZvUWCWZLDWUh0hmTDhp8ZUzWz+VVugyndpIzsMvddFZW66k6Cngf0KzfRk5Y8vvobIxl1AchEsEYQpWKNdcqpwo/LTZsvKbERV3sjVDHfG1KxKX3cFJ05ts2u4RNURakns16qIfP+SxqN30FvVhCWpekgqJoaae5TRSMHS5U1Np138uiQymhF0KDxcaj9asj7chR8f/S04ZuU+S5RsmmjvtQlGqbC7RtWF1lwAK6TWs23vBHLL979mifXYU94uGxne0nhmge48C5HfPDoV8kPf8v+SfIRhQ4pK0NUg/3pXWsrRsw9pdjL9RHwasHuY/Q4oICZ3KSiOSFYT8pUqI/OypE8UWtrzCZFQxqDNMa7BxwTBO/dSqMe/LQfkG1Lj4x8Ozvg9D+T3tLfOPxhHhE8O5Qnw1k9mATnW5eKJ/4rTU0lt5cnhgpei/d3cCNIjj003r8p9xAAyWLSRQrmTInOF4kksiQcDZbdvEgNfBTnRB1esLDkMIpCZhyTbIzOFttQIvNFPPlcQCr3KS+qojdfWh6m4fvLrPp8qTtgoCbJo8scxHPrTjFo3Kz8vwFABaeijF48yJJBDcezUC1Qwc7532tRZiiAoonTndCOeNx0lO0ipMsVIrMCatfxeC7ehHt9bLVr1GV6c4+3KbcfdGJumcKjcRI/ZDHAbLBgjLA/w3hclwvDnjUGiJTMKxmMUatuYsR0BBHoH/BiiXMlqsVIgZFlkYnC/8gQpnqJ3FZxX/wUqLkfnsx0/XiK+LWvgKu5NWL2/KdswbJH5kGUrdNw0hSzHXGKRVkJoEzUMfWFDH0wZevwFGGHyNlKHRIkJCPA7dkqoA5eAkirHazznYeRTq0f0TVg1eIBqEkEm6WYTdcaCdxffLGo1M0iolltavHPLt1/w68hpF9eyfy53xKjxUTYNY3UOppkCRW3ecU4Nz4fdAP8BzvjyWylEww8wbL4Fq1fQV3Uxj2qPUICCv/Bcq91oPEO3dCoA8UB2AEj7WMO8InZl0HwV5NMeSLVd/InlgzTYACsbAYojX3oFuR2QySwwCwT3SUl8kTD6goWDK1Ls2TBE1ghOY0sFDodYPQzS1Nxzjm29MtXLj1ffWCr+454+vbX4b03rRaQDmxVY11PZEDcUZYlxHJhxQMT7EqO26eRg4ayiCBLpF+TbvEZnu6+k4KmVHKfvCRaPQU9JEqyQ6PLayzswk/m1ifU6MXKzZW3CU/sESOsWa0YTdmfEKXfGw9DcJ9lE/UFf/R5qkpTnShnN4pLB2OaLx3mJPoyYBXViXiBaW+D4OkzWDV+24CVilCodR3pLq5E6WsoMf4RrPRRbcMqoGdUgam6VG7aggUEZTYlkeL4YJ2G+d93aD5dYYUz22R91RLt0Xsi6kyvHXmiOCtVO21LAWQzl6JEPPIgg048nyqE35fKMqaGgNjjMKimsoWF+hXwKOjBSRq03msom4sFKH4CeQzMZrC7ushTDIH7QrzurMz2CUl6sHfnHTKTx/wzSz8USibp+oRcHZqOd6lJtQ7Y31mm8L0fIyy/sueNdrDhSQMw7CLmlDp54xoIRNKerig444k/GvYb9ThLiVjfBr2ltn/CwSrFCvmqcz6oOnH/R4pV7DjQFZPcEuGPa11a8CAeonn4qfXAZit1IMVGOz2pMsQzFfqyviIYVI9xVEZNOCFgd6/FgkaaC6y7huVpPx8splq54lOBFDOZHM5XympHtnpwGKdPoq+DzGrZD7TN+ffqWjVyQi2W2Lyw+LPIcSPBFpBb5Jn0I2OY+sqjzMyBkTYagmKoIuZe6nzb9MYlKDmP3/NOt4dWhPOtMps0zD6ehbe4XEsX8/RvdDQeG9uF66cnEewuXl0csrFEfkIZa7mrwtKoVClrfK+znRip+XyIheaeBZPWogZn4lfoJhV4I0OBenNgqS9UlBgNE65p7Egn41bjJ0Cvj3ZtNHxKvoqxYiGqAOejQApHN5eY/JOWkE/SJJs7cQZt0dD/mQAo4QRtCuGWrat8osQUx8CABn3ZNxo6uj+ZpxjMEcMVMKWTDmJ4av68JruocE2r83o5uGnyJlpksGgVELMLu0wgK3grpTXQPg/g5yorTNnn+rf0AK+OgYzAU6fLAEIYXejeStwSlH4WNSUgG9K9QFdARe3E8+YfYIOXsL9PsVuMQFtydXSBogvBlYfVuRDlYWc9ZdoY29grUKf4VoNjem9aV7pcwBKS83lTaazNB6Np7v0b3F/FhoAP77riCQguSPTAX2OrxB6mVM1oqxS+zj5tV56Yo6XfK/n4DPHVqLwfFG5IT2dSTZOs8wyhAgjP1G8We4UxTsIDJYmg80Wwqq4ivv8L5PR1WWRPQTSUC3kxeWl+v8NLBaMPwEZCyWPA+FEQYJKo8WMmwxROPkNUS8gYQR40/gmRxDJWPoBVgfbvw2yg9GvDLt49uKO7iHYMEBMVE9AWJh7/QjFONZtoHMmfUVYnXO5bMFKAHBuoRdU6gSKuzlTDYyFcm5uNeQTMp2wKNN5XFdZCl4/+AeY8npe9HB0H9l+rormX85LaIE9XtnhTA9udFZDrGvHzVVvgSMW06GrQexZubAop3VPCXEYurC5ZzJjW2nf5OgfFzAMb3p4gJdtQtFA4b7DUBEvgsy4Ssg0eyuwAbzXlFd6JwV34vgPn/oiyDcoPJjXcRD05J9F+SistOUFYJGXKPA9FxOyRiN17kqEs7ncKvrZb33FBqW18Pj8EDlxt2Sv6WB74oyhPiHF/eA+TMtR7ePdVoWxSIVPEmCuQ9vyuhDk/s1olOzcXjiIxZgQYLbVrZvCpGy0EVZhefWQIfl9jMk3ehU+qrMer6kIOMmJSqq9dj43ki4PxLdu4CZ/8j/nzXx7jh2q5rbdLqAaVyz305vyFA9PHlhILU0dZrFTUVVLOD5uYWASotW9SrPwLDBfcYtQrtF2t1Pd++icSY04m9zEeDbfG9/FkSOyQZwHBx8VJkwaxl/Rp7gKBnU6n5wRzZZHpzHfEiq+MJJJJvwuIjWRAZUwSf69u0xLrtYLueqOY3Y7ChbXAbMz0MY5ChwDFCK7XfVfG/4mnJa523vIwRxyeBjF/jsAwrYy4j/kdG/hymDv2aYq5sVZqXUl0f9sZs4ErfAKFOpDs2R5TeRLRTzgNw5+uXKJyngfQcG7H6lUlbQTXJKgaA3+bo2ec/gOsv5I6voVZMznCy+rsT/Ir0UKwjiE7O7DnR/hEhPTBEgc3Q/QnrBhYvN4XtON4IO2fAlQIzkeHXewONESTn3k/Umuj8cV0sPKbyb4RFqELBVwCll9WpXNANWsmU8linLUBFJaWGVLdQqw4hRZE1waLGrrl3YQFmvzZ9p8pm46eaBXVpQnSnfSgw92PEnmVA6sBSWlFMVzQPeVGZaTgNaSTN0SFHDIaFs9Jc7aDk2OJcp7xFmAGQrnxeAC7QC1y5K5nJxzsq8Y2C9SoumlrPWuR6kQ+13TcDBuVCrC5tDEIvaZD1dILH0YFbxPAsEpETpQVsquZObX0PjEPNpP6Tk5/kQR9lFxHYgONTz/k+682GnWEOiEceHrUcTcteNJ49r/UJx/aCjX6W4w30xSvYkMlwUAlm5DcXRFaxVQ2ARuSdX2lA/6LInANdd3VmltsB0o+FqPUhljG2gVzKl/7tZhcBit20ILBWFDoLcMlVNOAqcUgRaVUGcwSaEzu9AnZtcsl/hD4tI6MFKWQbCB6qa7kseCBfvSgUmz1ZwtPYH2Uwpc2b9njtdeHOixZR036Zuz1cZ1lZ6MdQ8pDSml7qRs6ohccRRKCHq+mK+U/E+Ww56UnrX8A458oAJIDbCIzqWdWNMZsgQ3A6sgndTwcliLVl9NuqfKaYXXRfChc2oBgNOKmBuFSa17idTQ8bwEDuOBt/3jFxnHkyXun6zDxUZ7UU+HxUNzrvgEY2dd/dtjzmLojOrLKswV8u94wgfhKdfPekqRl8IMiRNhmePqHrQ5+6gB7PSIrCWJdBSqS9cbpK/QemOMVMK5wj9kJrd9ZUG7Wo7hPGwHxbWrDrUBqXwYvqkh7Z4E6Sh90o3V6qEyAEfM2G+MXfhTnNKc2lpfleEZWgaX9xuAcF4IbGi81Hsp2Kn43dlKrJ2Lv15M1MmdQB3LSsMpdXRKDRQQXwt1BEaw/0bRFg793CP2/Zd0vvS/IbWVVlex+ngsrnJJg8qe4vsJuFMamtXEXHqtKv4evidf18sz+lo4Rze3dRj0qwnMpCQ3AzznWSE5N9Ld4+FDX2jFK9tw1L9B6O5Tq1Iqf+x6qO57MXCxtZeY7khZTZ7CbKZ0jVGlyhngTivSPHUSO9XHiX45QuaLShgj62VPcv6DbaHRGMVfJxZ9rXFNwLdxvlgUJLUpd730MfdLwVeYgKIxf1gi0welRkmSJ2DNT9BnB6zrLKtpbmZW6e01nYOT6XB3g6Y/CZwo+2LEfuxsTSyxkkxzjDaDilcw0x+uwXkHM1pb4fPb3BdcGru+ZILldmRGpUHBhGNIdlYnsTV4UTltOoo0YSt+fUxo2/urA6wRFxs5K99KJlY+tfm3GRs4oQLwcLS4lNoFPEBz8SauOp2+TUjeoE9V3yQP/x95lmD1Bs3BT1k/DvwB5krBfQuzP75AXc1AN2X9IUikOBxG2qynAOlgKEwxmJYzIKPD7M6Q6M8/GLwLNU6ujooLbEEh/Y71yFrJstO2jFEYS3XIOKPKU4CRehVVDAcMR6om5fR+ijiOUgBALOYQ3EUBO399pM15PA+yDB43ZySzZgWcdR2Jjk8y1bl9RQiLxDfPevSSa6lpw5ElI2X7xRda46CEADvccM93rLs4NrrcUP5G4WLhYqF8WN1Y2aJ+OWojT/WkVqR+lSR+TlUXPvf3rq8SUpWIf1qwdG9QPjSo+ojvYR4tW3hCLP3Zjd/P0aNEjGFFwUM4sEbi9SNemslfD5PGX5hANM9Ye+F/QvB8OkyEuIBfQG0g6RtlwQuCsJeJ3mpibRro6jC/zuopjSGCjDGWHj9p8T8eJEfOoNVd+ayLIyl5W6761+P+lC5Uf1k2moQ39aO+n3Q/w93r8Jama1GWAdZhLPam39RZ0FFL73LAaWQhkgLqB1OwaH8YgV5veMity8fNxwpJ/cjjB8Fl3FSDj0wzMn1a39mlhQEEowjWR043qdVFGNUreQSDd1xDNqfHdLMyksqDBzhzzsyZ5p/RvRxusgwj4VtldPFMgxt/QW5A7uJsnh9mAaqK1mQrfRTOkOowfoi2EYBdNIfF3YTEtKRWloAWLgPITFX3gsjDXGgd8JBoQoJ8eyNrG7s2R9bV5YmNUqnYPWHYLXolHEK08L4tBxUIdWcTDd67Wc9dY2muXplhCX93GkEnoxp/vYbxcjdKcHQaDhw3k+Oa6qMOT3lJNbuhb9Onsq++ona+1PWMhEQtO1kKGorjqjB9/ei8cu9pZKs6MSWVXyYjZO1l/mkwlxmthXSuH7eIATMJwESLiV8+ebfq51bidotrS2F4/ewWqOB2XPfsnUZeVI1qvHp3NaWnY1RU5eR2Sb/36So6dDIG4jFwVelyMm7KMdDIFwucg33b93cYxsWuNgXr2SDmAdcXyjyknoqJvNxkOBcpB4S3m8SEDfPFYcrKwP09uBIy0LAU8MBxEGN/LftevM+q6RDzkujc5aL1dPea2Adqp8bn8u24aTB7QVXhVXFabK7zJt9YBkYXjRczeONd1HFzpepBGHrB6hn4ZkV0G87U7RVovsjXROiP4Vh+WsLVzcIBorJ6NAoXPBGem6gonO5ToYskL1ZEK4hg6go0lxAwAIKVlVTAAI6we82WcqvKBB0huxM3E6mDq3wILkEpGWBMQ49W8LJRCb3OEFOVj+ynNW5dO5fAQsqIOM0DMmuL3CVE1HXwhSBpaUBzQG+CX4FNmAfnOwNOKIqMkMnDXbqwOe126eRcQeUHD2qWwV5xUoLl1KI/fVVpa9gRssU7wjmung63FfXD/fJ4vv+S9nYN8zBvWCl0C+5IDgheYswCx+SsuyEt6THcrNyrPzZjtjodoreUjRAaXonM1UinHk2uILWVudxbUQPORaDyaluanGRIIGdeVjCGkEee7h5c4ltdwirHMnI9cmYckc9s2NPqQWAVpH63SDQoPHHASb+jaRUR7ZIBtXd9c6nD5E3v3M25rUlnOz7OQr+qqroTfp1qcrP+w5NS2WchmAE8Pi0I6o10NJC42lMgh7LyKzgearoM+TCCXpUixAAg/Ad1X+fimrM4kADrkIbe+JAnJG7xiUwAZC4nnyEcU3W6gk8saTxydosfl4Dw0jvQ2+sCn7lAwPuV9LQ8Bi6v0+zdH1WOpN20h3irZWOXZu4EHH2xwr2Ka21xRlXt01vbIkYieUV5g1QCFfx+REUp2wSVkXCkwvxwBlh2OEp+xBOB6Bb5wvTdEIPioh0aFIsz2Cy+451vVqPzE+y630Cw1QZ4DxT4xl+wu3XRG8AeaL/jxDTq0gkovq0hwFNUUvQzJ+vVc7AkOyx7XTpBz7dbAOrkiVVlzJqPSesgCC9GMrtkpMQu6gfT9hDkNXZr+FcvToVY639lkinxf9QrtFVseYH+XyT1xL4SkCBDf/WABRsohLDzGk7oK7L//Pa1XYZrJSoEZLT8/ya45jnks0aXuRd2SVTVxVpkklgOU2pXkJ8niE8qIlBF3AA8qOHoFKJGmWWkc7tZunrgx5JI8/spHyJRW3tDXKP/KiFDz12/8jWylGYejqkl8xrwEhs+WhdQzhNw/wrsrsguPW7UXIyiKtYh2ZCrW4p7kPdDH3OBfDeMTvmwFyG/8a9v8LcUY7mdPbtAeIdS9O021qmc3W/KnseYiyyxnBBfAePdnNJzHqsNavzH1WUvq12D9t3aQAPvJC12rzcCybwsmq0uFKDb45BkwVxGFfcY9vD8hZwQyg4fVwZ7JNIdCbgiZ1yx+hPjgNagdjSnWpLrXSPcoUpR0DMhCO9Z78p2OkL+QJJjrdG4RPe7gdEE394+HoCv9CG7rCrgxHGZhvz1BvqWcFpWmGcmoXgiNR1JjpKiU51OIcQvSXWfZJxjgm6Kpau9k/6WOj4hytWfr5kJcxhEQCirJSaj46kgM9Xh0FsMvt/qw/yxkIke0sAPuslk4Ob6Acx8iX8TGtYhrrtJ5OX7BSF4SwvZ3JVHCUodMy/Jigo01kOhcM8ezn8gTFZNDbWVMrMvmvJKK4GjZYzsVUKwlAaB+FR1ZKaiHSspCCia9oJUUryDjN2ueUHokEoM84V4eISlzTs7dRZKOu1vseNQo0HKdPgHglIMYrRP+iheULg76POsfS5ve80UVDlPeWdMTUAOjGTphsI7FxZLNQOCJ8FMPUFf5mkqQw1YYCaIOlfBfsOud2dLwlaim3f7+qnXtoCM3LGMiRACHVlnSuQv+SLTh6VKjouIni49H5OkiEiouNYh0YAntgT5BHVrMrmcpjO/w3gKnxLBXg7jDMPKlOFX1tADXhSbT5wbDUBSjkJwdAh/mbGOQ3cnx70XqMYnv84W7UcS9r0IGdz8re309yWHVtRTjZjyTBXt2AuB7YxI5rjYPnsAD/C6Pmfb2HINEmq8UkYXGZTMk831Ia8dUX4bZS3NQSAA5drhUE170BIkeg/+7qKXJTbw1ix0iXor+TY4ihQHC7BAtK0pwbROnUVzAddIf/pIFy7AUt1oOS8tkcWKhYb2BjHAlMCRGk4wvTICpNi4Jr1JFFan4d0v5+1/hYknshS3/sUTs+oT1Ga8fLasffPLZUmdI61/klmX6cX3sUXzZLtGV1yJTi11ddNU8CG8qi+BSvloDySTC2Ik1ssjT4KTZdYLhtVuAuFROBqvs/tBocQM2Ls+t3BgHoFC/7rARlxQ53tbBdIfOrC/wPAqweYWPceT1lUJzS0GDfRDZgQiCI3j8yJ9BDnQQIkh070j1v5j0dTeisHzW4gbsG2wPP3Pn9QU42sAzos2HaCNhM6OM/kE9pl4LI3U7lwgfx4ByP4Hh2b3ZPbWnOicwfrJLCogDE7JJw+8+j9pT8XFXYmVyXqQc7UMwtGhg/6h0qzb+DW84va9JvtindPMMu0Qj3JFybZRWrzfkg2rrFds2sWySeW545Tj5ZoH1eI3X7AsW5HciIY2se5PL861v7qRoD2SuGfb5sW5qVU4QPmUXRUnuZqzyvhHLA0BATdIwM548lmh0RSN2C7/rKzHaRy6u2WmL3qeCwdul0i8kyukGPHURG0BC2kyaNnnQ6wWwZUvl6bu4JqcMLIIm57lQ4+Yps1it1eFo+eUguNanJBBgZ6z7H2WvposfcUxAmFYnpbRrXMwGILfAzu0Y4yjGxQolv6FlWLb4AySIDxfZyY1wUqA0eVvBTFKqFL/WuDu3OVXe085i2xCBkQdMCv7XsJCLQugsaH8IGFRkBJXidxRjkwV9JN7vWzNEgY8kjV0zs0H/0a/OEOHw1VPmknNsG/fwFZMKg+mVMGafz+FDnaXg4asSYkOHKg/35Nt94F4j2DK0Gp3xo03S5+zSfWcBLhESV2ttSQVSB25SWuLoIablFGaBKwyowlx/2PuvLU+3ecFlKBBNwzMKbbXEfNrO12V/WbJ8BjFgIKOMGryoLvWPxpe3UxWm+wbRDtG6emoi8eeX/CMnPJE7CYShRHbYVcnVC58T8sWGrVAg2kExDXIfYiR3ZnOCR9TVxDpMd0UtbpmjP+GsbG59LXzlJexbHwJdwoczF46Kn/gyL3lhApdBxoWf6H0HpOf6nR9bQbIempOyJEAHCAQKyExoeJlZVhZZJmyxZjair1hmRwF+x1QUzXU8X+mtuqCztf7A0nu8V8swSUVJY20DXrKGRnJQ8EZsEe2nJnpyIGHpUfcQwyz2wHB5edRda5BvLRva7NJKQgqbuwsxkOGsj1g4cvVSfh0XkwR/lrv+L9/h9SB69yH0OJ56gdr03pT2++OlXDiqKnF944xqhbcxW2BOpL9RO3cUDqOyjNgyVqdYDgjn4cv8vYKb1wCWfzSm0M+f9ZGRoQvW8LJ4RnNemdFNh6RTJtzt2L82V1d5EmwocXoIQQIMbh5++Mkfedva0JrQPA10O6MLRprk2QhA9c58g5EYB1lhWiE+5yFfzWVvh2gQR42qoYHAEvjyRC4ig/9oac3UTRTA2B5spjZBIZsTvR3mzKSRRoNtC5DZ3UcYQJXe6zRAQAkc1w/qPtOLXUNw5fjkf8U2z7fcthBXTIIJhZTLxNSmtV6VOqMbdKxwjSC/i7VnhfSoLP0iJka/rgYHKvnS2SZTc0gnMKS4Q+dA/RDkcC7wjhIWLzMI3JvwGM6ARH+wOB0M3044BmA9ZxpOtUKDLcqixWqcXFXfRbh0Y+hEUcrsojF4Z8NuYfQGlBO8mQ1UWN3rgpX7lR842GbEUlFA1rBKuhF4pXt1Sa7Z9vfP2OUTi4w+Iz9X+WYhXOBr7Z7+IXFr8KuqCKLEDiCv/oRmp3AjTPWyH6gMq8iBbVFqBI4KDunyWcKtYY9AHN9f9KbHq3uMX3IRJIKY/aMoMTkj/ewF6THFtiFrqJIpVk88L4yrmO80xgZ1T9xeBbonPjVKxFRbc4j0WZR25fafsJD9RUvzXYDr0Bkej9GpmOtpvCU9wcdbVVMlb/xoOZyEj8jI6e4yuRuhs4k1GXBWg3jtE0+GpmDg8JTWDXHhhdxH1sNn47hDWCJFtM2lbYcb1wy9cpr69tkoSQIybPQzONfORIjn6vzbQdT3QCSe1+p41idc7C3KSm5IKg/y0I7Dxt1O48+TV40KWphsX+6vijYoIQrUVojPTjif2RhHnPAMObP8ESp0ZIqoctGIvpwdjqPty6QPUHSLopDBxB2uHLCFYF2gDR4fyOF8xRqoM8hUjDNiO5V2sHcaqTEdqqQM1LrezPAnzdDIduU4sfL+P+eyf3PiAs3oHDF+WE+EruFf5WiBYV36zxXxJ+NwquTdFjnRh4UVqzTA19tZNsbes7IeqFVQubapd4G0+PkxyBZ+Priv6p7enDj6wEe12AJ+XFSZPVE9dQ8kTuEmlrB74yNEfQBYLnAK/jgNUSwIKOgmOEKiB03NcIK5UUOWSl7qBzwg8fhy5KGqlelp0j80IO67a0FNwq3HRfcQNPhrYDBKzAlHfSofs2YOhlCdZooJf0n0cYlZAqSCg38/BE9uJOfYFVK5H6S8j7KLeK7CZHX0GuOi3ukWEFc0c9ClIASY73DsE1QjfiHEnLI0pFZqA4DphFRV+jtVCyUEqabIRtN4ii1ftzW3X6czfGYX0iH0caOASxTJvEcnEye2Q5zW6zcJ2HqW86/A9Ts9kPqo0Y4RHCEzmwO2bE7Ir86zbcAAheqOdAh9OeJ1u/tOfF7xg7WBXpU37WixI63v3u+7RM8TuYm19MuCkKhinzkjapKKWgmvy7cwhOo5Kg6iEIrOo93cwnqRvnhCSgBtdNOHWALKIvvuTxnC38kEaZoZcN0xg043hcHHhMMZN8kSC/EeS/4oAW7gGEAM7pm1Kb3acn6dTXkSSbLlv5Gt4XSwS2UbeFDnAPXMRecJU1+zjaEbWvfL2rJ9e3uB73HGBHsKKtXs3n72NRCR/GHc5TBV0V9dRQDhliyfSt2KGQiRuiqi2WkeMvXn8BiHAflDc9yXBpB6meqINhbid+LKetY0lwhX+HqPPqmvdqth+3UgyC5C2Yc1ZoWeeeoQJnqcI6HpN5O2jLfMaqam0IuKp4UC+pUZOiywVoAAQX20Ne+iWSr2gCy9i72ne9tDQ2be3xEqxERJDBghjNycaLTAiXHRq2raLRl3rICnUSZrGJ/CGvdx2gCXlHBw4pNwTEWsNpmZrFuwHAwx5mkUufjQNPuhPfiBTx3JOV5993elxarg3BOItJSC3teMLjfSdIJgdBNLEPcTjCyPCxzCRg33794epabnpbMudrCNrQfZ+L8Hu9YoEryE2ug3IO8CDMRjo/McHjhM2YKr/56Kr6ApLxBEMSxphbrcYOZCISxelgwxsAHSxe6AZSFucjc6pa/QZ5F7SpPMKEhR8nyQuX5MWby5AKLK3dz5DRaiqPO8aF3Viv9VMi+hJTvnFLlfEkI26li7W8klOOgakmmsUb+LBCeajmWLRUydCYAFY4XkFGMWOfDd/UlxFpALH+eHoCR7lay4QL6lDwzyX5fPKJl2Us4m+PLnqrzCg08W6oiKMdeJMxGIV7+22HgoZWDTPmqX04yAtAzxfoZWVXmsGu8Q5zTWik4f7wQYYualcPGiPl7oDm96aB/u5g5WXrWd+sVBFp/pbr2069RIVeHAXdQvZhlmfn5N0lj5Kgv6B+BlHm8+eBtlykFq+7Mp4byh59NA+lu3JfsUGCtdZhyQxOHhUVoDOAsnEn/ybFVEKOxvmp9gobHy9WT0flXvA7Yw5dzDF5GTIKlA2hJLtAglaQccQw41ovSUVnxha2THkQZGEl08L4ieYBpM/ZzqMlKuDoXcBpTe9aeUcg76RoX3ZNOKTExB5z611EVdHy3TkmmpraKZVqBTuOq5xe6LoY+t/xDojRelzcvLjA9SYPfiMNftgl+pmwckEPONPliHj31x67fT5COk8LQjDjGpIPo4uPBJt7i99alVUat5fdLQ1ao8yW/SEFIQCwclNbyRGRMcA6TTYSqzGgvCHO9cP+zm5j8ElJ4T8XRQYkGSGqNa1Ft4It/khQ/RU9d2ryg6T7IkxVGfX7A0NUt5mipkJ/qdEi1WFu2VqTOKV9LteqRSKS4Nq1Cx18He3tWDCxzrYfnIGDwmmFeVV91wwv5zr68bSda1aWwv/sb+d9anMt0sE+GO8MrKxEFg1S+WNaNf7MamFmIfcNbLPQBAhU20AZgKGlc6TFqQo0U6XNB/oK9mzMAELX7hHDRXO1QqYKEueO+nb7rLchUho4ZXAYeYVleDaukx/5wZjxssBQQap57DzkmYqAP85by1N/KSoXpOW0hsucHOAXzqm5ecsaOKsOE+TsQXmEvMm0zr0cxpF+EXlmqDmkGa7wmfVubPUc63A2nZ/5/OdTYComqLLLh25ntM75IU9CbmB7NkImawnKuKn7k5srcrmxR178rJBlyVsxyllYpFtFH/rFkNxLtvMiDrd8FJrvyv/L5KJzXEWNa20TRzK5y+i35+QfwWthPOiJwWcmXi6eHLE9dVR7l7nl3A1odh6m/z9ly+q20JbZfZK7zde/Yx0MUWcuEz4bGVVZGR7MTFZvNx9mpLxg0IWlWSjb2ykSnDHmdKF00uD7QxN6SAfRyt6nhoryl9cbxIGEkJzJ4lMVXdYlcz7uLanNWTATIQK4/1NY0wVzTcjVqh/0ucWITvTdC/SAWDb3rfM7LiQhickmDUw350OJ3JcMzJxaK+6B2guJhdF1JWpnNgaTMpsURcDaDg29gSv2BtOZwO5STmJplwVto67bzW/orjN9vQBMtYwGmojwjEdzW1JLq4OSEUcI7dKbaYrZuB7Gd8OD3RgCjg1huud4Cm00hWibb3go0QVeAc9+2R6SxdvR4mwXjs60+LZkHEe7tzxK44C4PvJssYULNL81tvvVbOzPqi3aRorAoLmIKGUiboPb2lmsaXNsSH6kOSgKe/cBfWq3XeTVpBi9jB3A2fMLZJPs+fGBS+CGXZZxHs39kHkox9lgsdMItX8AWBIqrDcl8wRHysaCGFSlKDGuqWHMsMHl1t1lLvj4/l8nm0EcyWyxUuBmBWixnfvYAhpdocDKjEUtuUTLwssynznbYMQi8EzCOtM3mhn17N5MY6JFNqKgxUyYEv1FbqaiHrZccmZXdM0Vua4J0WraLLVFx1PaQn3rQruvZFffR9bjlsqzmJtYeXkfln3BZbNJ8SFalShVuCT+xNtT6xshBqPmvV/o48Ow5ueaeDBmaaR2IRHRCLL9OBBSLhS1ojh7Qe37jU/lPHOFvpowJ8RF4Grwovy07VQS4ThShTVZoIV+h3HJRA+Jw0A7WBCHcWGb7W7luXFtqXnLulXUL6G4KB1P7/vHDrh4egCQVWZzOxmHd3Bk8a+kKlbqQgVUGwtUCY9CRL2ZG5i3qBWByvszc6rnEh5+AOV58oXOUo9g7gjSayTl2qubhPgQ6JxAwlsmNM0gCoAnpeacH9XatX587ioh6qT/LfLMrOnAgE9U9T8OIbP6YQCobzYr3wSulnLqb1g9rbAQQM+6PFtlgp6I5LkZO+KY7wsSYYvPKiAJ3/U3DP+5dM/uQOf5YQcEmuOAQHgPRCSJFoWA/hMFYNp5RsBwBmshQUlPv9GGm0OPR8EVTj1uXqlNveEegiqivV34ytS2ExtsfQu9nSWFl2iFNmaMOw2QY/jJ4ulPj8gdW6Tjz/PKbXrXui58o/Kvsjz0Lis1ph7Id3n6SltXd9Ia3VrYTGQ4/egpA/mG47ayhBV0/Z1iXHj3CiXwLDC3rpREIjK2djnSC6TB83WomZjxfNxMeNNDbYQu+MEKDbI2l5g877thFxUCZzS6HZQIjpMlNLUNo8H5M1clYjxeAjSqeoLScd1QvZfgWg9QgnCd8MZr36FHmPrGNQIvTBFPjZmtSHFCOGiVYhresjWIJYs227KFOj+HFNhhtL+kZP7Faq/nJgix970u6M4tNFVI0ixiNtW5J4q1TmI9oXmi6cy57z7ADt5+cqz0qrG2o9ON0KIR2Nu4WKBc1o+vPSM17CS1TwvgUNFXGDHowzFvC+gj8mpsA8fWRwDx9fPc9Sw4VgQN+P8a6lBNZGO+LkeOBlVE83qP2tvlvuVM9oMh+PHmP8Dj85rSZqdMolZY8t2UESoi/OIv3ECU7l+wKfvNxn7k48k+iNjHbpftW6qgP4fi+hYA10+z/wimN9rZRZ/Uia72Hrcp7dS478VDvsiC0GjPIj//8DUQmIxUDIwFwfCgCUtqZ5zDxEPsSokEuey8MsvGIO0sy7eComDhmF4E2LZ7IIxgfGiOiy51wcYn5oisRlfvE/Tx74WedVre4yOfbmVFVTXuHI+7r3mnYhrY8tic4XO7+mntT3JlRmnoLuGzXfKgMirpX5vcurs6/iF4PQUp/D5tpJ2tHZ2C3Ub3o9vqmX12cpMQ77onVn1YuXNk1V2JNGNVGtyLXayjOsZkVcI1wbZzfA1lfGDaa25sBtW7ac6FvWdQ6gArjJKFiG5/l3A14AY2p7/YP6OgIeQ+qucdHZ6pfGYbEs6SKdtVzUbAZv1pHKDz4UVSmd5coi+SKmjlzoAUtzh5WhwUYqtfRtUqMZZLP5Ckhzxdh7AFJfKMZ0PfSpwl377CCcGP+ED/iCDKkGzapabflIKZkbLLHmyCS33JSNdViM//96pVa6fXwIOLJ5lhfkSvZsI4PUROhZTMpzQcEQZISZ3+NSe6dt6VV9M2FowWTJHGrN9p5g/tjhiZXgfdSr6UbK3VAtP34anOu7YHUK1dNO9NgYB0a7prUcyuLqFx6R+w49jY70RLJZ+JWKJ5XVzTGcqWosYoczqiXiSz/hv9D0fX+hixPrgUOzj+90EZOE9uAmm/oeF+8MbAgvVnirPhTXjeEWQOikfXII7WfGousGeHzVjU72UXYfJo1OI38br1nTQKU6ZTiQ6wZ+RPV1ZMjOW5l+TkZJOxzZbcd8EAwSxayvgwnnld1gNVMsA2bUQ782i1FWxOqlnLZnlhjzI+yVC/gFbON3qe2sLSWwleBOr9Xz2/muN1wZZ2GgyTuDIzENzglPtKJELRfbXjOtWH3xWKxYHwLAiddMHskDnJd8Gt/PDo5NqLKY/0+6v6cGe0w3syYARa3YB9A9/d/x9uBlAkr3dqtKmd/2e0r2RrUgMK47fYgQ2VaSMYPdIy8mvX12mS4Spe14zs0huiOjXk7NuO793pK8mayKgF8JjJfVTnnvT3f3Jd6rUjJr01hOws/mYMT8qx3YI1Ir7+vBBFVuAiIB9OS2ZAHPIsQraSlwlWFO7AQb+TOdI6c/6ga7WxE85pbWSc96RdCwC/8VTEQZuoYVOPUeB0Hk3r9nqQDvAyyzwknaK5MNMIiasQs9tqZwQtvTKx96qW/m96RqKqkDyZfl8umevDqOCkXA0WOr3fKTVmxO982O0Ai+CA1WrhQIYHULRV6e7BcSQ83L3kol7f4gKO0vsE1gP0mvLQ5uj72ckXVl7mA/KL4nHLXwMsZVhrlHLGfp/aKC+83z61h8wF8TGmvzn6NDuTrBNZ0PjTVmQIkKITLQ9QFgK8eGxYq1R8klYoj5x+YHBQrgAMtGPdrectBwKUEQNvF6tPA4OP78t6dHonQdDzbQqEWLCcs2SnRGqb5jwtwVDZvGwmb9Sn3D7cVs9T39J7cykqboZ65IjZyhiL8u4JfzQOkcb5i3JI4NuZ5dwn7fYOj44gUd1ux+eL8r27XmntGTWDCTrYI8KN51cKKhCulBddNCpj3ifUmX/mdmQwM+6xKlFdE+EVBsC2JyDs8LTJ0O77v1vX29/LtefI6dA73Pba0nXbmAIpLlMxEUJ/ZXCETMOdvezlCcvejFs4MLT4ZOYPz7sooIIoLYGoBmZzyD2MFjNN0cPzS+R4Vcn+LPGTikNRjUDed8wBggbJj+tsR1gAiPpx/vZApaRTKnvTK0rr/PLjTZP5iNKhGVAli8f9C3hfZSfMNYonXfqTTqQmOaicizbhVHNx2SDneMYwjNpMikmo5fpx4X8cF198DjJG81oLdz6Lvovp3K4D0IV/OttG5+pOLWlCYyMIB22H/hV84fyUEoAoHI1ZWoMnB7/lpw6xo0TtJje+cp5QImPE5w/dQireGbA4J4rxOI7odeNW1Il5JQHtQ0iY9pNQIQmnC1ZNPLes4X0MiViIEImLkYofgBJbQba24CG6JTlnhBQR8WJNsun7WbRbPqMoT/KvCL1lEEOMucSDoAeSKxEs+T7kcpa/rkAHUJzio4+DoepVwM/oK5SeaLVlAo1Z6WZ1pHbJRHHnGiLFkmz+FrBbTDr6qRdx06WEoKGT05jdtGSvUv4hfMo0mfUZa0Pt6T2WxDABPLufgw1I01KlyizTqU9wbdog7Y61f/II7gfslw9syCRnIUUatWYK1mPDi9vbOeC0OSoQRVTN8lFtVBBCT5CWD2usWp6aUbvfR3oiCY2pou8WpxIi41G1ndUx+e/orb893U8OOkZOvwv04bRwEKf2VOcQzUuXaMjpDwxUahZsET6Dw+I0KUSEJLnhbSaTGwwsbSezKR0PfixnDy0xBejMg/UYS5boM0KR3nrA4slsGfVnr6M8ywQB3qETlhI1OsTSefxNtRTFc9oH4qn+nk3B+uYUOEw/gJMxrXAs9cRfBpn4Fn2B+AaZrlp4nv1aJ3NQq/DJdcQoeHTChnSGt4lu69Fp4tXci6S3IQCX5zH5wCs31OuCvxJMmwj68Z7RszwiGl4Ez3m/gS/LtfeTksGbd/OjdtWD8purCuyMSvM8cYH4XyxbH1iOr+s03IIk8AUqta7hOYtbYY1bMrrUE8nSts07s7T5wq5VjWT4mDBpKhn5/cBJQ+0TabEnNjz1oLniamCCcKcID3XZ4+x110m0bDodxYwxbJrA9NxCgfeeDzFgeI+ZyD5JUX+laCSzDCsRwzFNTwJd1d3l/91xc3jyTKk3+yEQAm/nqiE2gAukRDl0iEfudUTYKfbEyjMymah+EXqDrwKstAg5jDiPkoXB2Ios16Na5hLBz7bTPFco0J+QeCbckkDSGFs6ohr0ZTWQFc+8Io6pw2ZLws752clNHQPhjSkkkV31FjGRvETLj5MDputKFc/6VvJ0HKQjXaeSB+ztTdrZDB9dIUEaz2l0PzAsHGp20Eim5QuBAmsWTNbDunRpV30luoYkqjrGF5goKu5qHj58WH/3FqOvsgeszn3oEjowWmW7goGTu+q2AcNZ8DzdfysNgm4wDr+z/aubcsYRgr3IIaKmuSGdzqVji6A9iLcyGahTGKa2SAJlpvLLG3os8e6DqatGrZRbGoiBb3NeY4FRFaLvg91v8nZGrfEjt0H97rKiFHvO26rOIbBvIOnMBlQ6yFEYJaPsvQGLyfAwWHcwuENNGDUuhqKFbWWGWCKpXiHXmJzYjcyhJ2YamgeSO120iD/iCslR4onxqEIo3mM1Z25f49X58N9Nh275ll3+ucJTZd94PEfwxAS6vqffUZx9fLOi+eX2pFhFoNZt4W1YMmFZnwBcx0twUxmiQagKJEEClwMmCQ9z3TfRPbyUCATR+RVDQSF0bYR+3oF14oBLI41ClJl2fRpxG60Yde43rp/naNsUyMcfBJvB48SUQohbcSk9SbmEhPlXHzMitLc9D2UjqwgSCxQudxH0MJllZkmdLq1DqLkPmZVV/4pDHaDvD4yPDQNs9oK3qmJIVc3UD0Os4ejOZMQ/i71vOglEssaPSwR2FiwKq4LwWbeYS3PdDQ2gK+4efEpKz5f0/n+Fr0P68L+6JN1YDJfP42DUUYmANlSHeGH62qaPt+X//XWaQGPtVRuj0F34xinNza+DPerX+6ztpwxJVzFj8xelJKCeF3/OTZtc9hMwBt9KKXry2yHtG/EPvLjst9W0X9B1yXMzmzLDJjtERbkt3wwA5FGZS0EFkNejtmsujsmPl1JjWl1am3DhdlUkH8fODBiOJPrdCe0z+k9TxhDqu8gNwTTNRJcdVXif3BrxOsO5/gdc4HSI0NGtK4Sv8h4fAUFfVOCzPVVMHYB9K9eYx0tEDXq0rtc3S9Y3cJwMJttlrNWXEIcdxDVBT7Mtw6XNZaF2UE3rf11dO2C07y8gUl7ejUOgH4cMNaamxmW1ChJmdfLJs3YPoS6fh9v4J6wg6OziEYcCwaYe7KVnqqCdopq36NLhOG4Ir+pFLIqxaojUxuNOb0q1OXiZITFczBNaXK52yO4njUK2v0lMWKwhBJQJmjh6dQ09lHwhLykIlIf94TIriTOJvCjoqTWq9ZMg9ICcYcSghEmdyHiO4qpiz/2B5PrzeyxdrBEOCzRey6C/eg8A7reiGmDh8W0tgtsidW/HC6J5qBPPo0KW6A3bCNCWkYOCe9fLbKfYx4nVCoATEKLQekgcwJEguZD4fPA7M0O7sr/3TT7mN0ZnQzbnpzGVsbCGLdieV9gUFxLQzxHfnr8vVL5myEmM/FdEf4cDPER7pO/p1pWBRY4c9tVvHB2iz0bJdUt2btyS0XFwYIq31qByDDVkf2qNvf/Yv5BtQY2CyhYXpBFWLPxxkOQ5AzLZ7WDDIokF9ehHLEGfvGXrDgjHzrR4j1Pcu84trdqGYXLvvHD042vaKcPp8Pg9bCVevcgAtVoI2qCdUUHV1YLu26EGV+2FP8sCCNqtpNFor0D4GZtGvhcF01QJnzfc7wLEP7d3+Lui3YQXlY9J7ewaj/Fkgete0H/TIEyz0HikGh0r3dtQC6gQGkeMmld2e0+EomKeCT09JK4XLtMaj2ZmmT9QdLv0RNe+cDj1aKJKyIP/Fs8HzJzbgYEAz5G11/7uuzVUqyE/Rf/v9K2nJt/Rilg06g2l7L89JgueNA4GDqBbNMYmKpzEGssLxpaaZr4SfON+TgnaCo9QNYVQi7HMBj+BdmwJvrbjh78m53fhLNxFD8Fao9t2dl2/YSn/WcLLlhtI2/F6sGn/AEWLpWqGwU5E3y+HiHMtiFN51vOZ04rJf6STAmEygrmWOJQdJFtfUF1/O9cO7C6BrM721/1L187je4EnzJ5SqpWau5vgMXIeRz0x3VC8MQsc1/GsJA2WQIPZOzLiJfmhA2kBMweCaRttnMOELX518vo4Oc1YJk7ZoZhMyHUD6Y962U2OyhrnQNgYjEhtvoQPLqbFm5zpCGQzuljDZQlGWtZ9/m/PPB/VjQt8syJPdQPI16zTZzwCwtP66xGJzj80uqYEPpnqq1pUITqQVtsIQnR2WG11yGXQmKvV4rtnk10R8D0cw9SiAezXtdUeY6/90S0mPvWv1BeJpT0oMNDaZ5dSAqjfS/NZF9+xjxl9In41xSW65i2zSJggMaEHhxMIvpxnUK7A3yD8L0H3VWYRpt49fD4Kf/VUdtHMUJsJhZEjxTkAImAJ/Yo0BN+ufdlvVmgtl4AwdleuK9S4U6x6H4h4aKItTsRjWQ1cY0F77lrlnwEpK9ejj7V/wz/T8B74odItm4LyHE8BTk+GcvlVeq4tq3j9ZceIUXLKyUgIr0p/sA9Cu5Pcqx8W9BrG+lAWVoKT/efyvd7/5YTv9Xx+TbCwH1F4xoCfWzT8mMRqWr13UfY34t8yvw43SAK+CeKuWo7AkWPx6IcHYUObiJKwaivEjzsOkkvz6/pq4r0kjEeM7xze9vlYOoL1cEYY6c4yLKTizV/vQQBbNxXtshamiu8e2og9PBVUtaXox31iS0TknCYOGL+W6/6qkwdVoOHo703zAAXlH7IxfbKbtATarOXSrHrUt6JA6HGPl2/144YJ68UuG0ZZQumxJqMXG3jFVFIHALrUg8BhsXKf83yK5o0o+XS0SX7IwXr34X9kKjkAgtKUuXgzrd4BCFVgK+tSrpWMbIGlTjzphk8A71gdQWfawbO/DVkRxZ9GrMtykPo4hWaCDnoK3j9xc9UOZ+NzmJKZ3sBLu29DyC0UhS3yl43agkBtwRHUJAwYK+dW82uvGbPGyhtS+L5TeBHTIko19dWcknY6CuaDx9xvf+/hkjsv0lPsQ22QafmqgGBSk22IZJyKgG7yPcgMN9dnzgPUKCGheNb6wtuNw5rQKZPd5jbhCtC4HpBfUqIzSapemkPIYbL5bmwlULPoGfLa9BAMZOFF3DDBzLmXUVjrk6d2KjPhe2otz4JiPqCJ2vk/ZP3UtuaB4LGmzY5KtG9HbkJSDNMpo0SxpEM87LvylwkHaSbGbW0DvtVYVpIKM9+zOf9OiUjMcQs5bJtIY7gs/wfaz3Rx0k62pvQhz4h/95XqKbAqPgnb/3cLv2xziJe2FWuNxZmAbeG4FXj/t3r/o0p/A3futf3LURJw/zUp4wLwNwptoNqAootllVBlg8FoeXt6/2rm8gQrM9AX1TfKQACe9/8QOu+l3i8W+0aRFbeLvDsPM45lYBWTPSL9NevvrzGm+Eg+07UoNzj92+Mia6Lp/l8uKQk7XdqJNCIpYlYfEIgwMBXibZ6z8NxAqBGSRki88mYqTu+BUjtzUrEwY6WbfIEeSYeClYGkFi58Vtmj8+M5P3RkVeVfMZojGx9d0vvOuqxcX6g1g3RixxQJypYmGbGKBFsqGP7kNDX2ySJyI6RkFVUfLnYFd6i+9nKv17WVRaziDM31bE+gu45g1pBF95hEE6XtO/CdpwNSdIFqhpn1YRAiR1z5O7t9e3TiS/OyjiiLYkjfaWccLBzhUzUe7XNivwFsCNu68kMhu5g1u9P3UMLZrejlW+w8WRkfB+nQ7Kbps96rzvAC/p5b6A/p3Y2abkjcZAGKLxPtn5wMnIiU2H5iwrEoL9eady7KK4g4DkcI5ieBojOpC6BpK5bYGWSkj1+TqdPk/u2CHpfimcNZbGDur9rWXdJrYuwTdmE1WjzrwEIApq5h2iazNk4VF/ia5bUxeidgfiDwI+iiLH6RbC3UEOSb3b+bywXpsRbBQuYU0tr0NxY2xL3lYxpebn4RRHWzL/cVQPRp4zRsMUsGSWJnqXB6cgm7KJE2dYxnODa52qL3Ta5mK5OK6yxO+ILEIt5JAkxzk3kLEA8bS1G+TW7Yt1OWRnKNCQH0Q/2ObuIQX4UEkKFasPRmR3F6YPEVhO0+v1NIsjca8fm+jaLuzMmU6xkwqM70Jc1i/FdPKhdv/JimKKvkY8BrHa72oM3MT3Vwp8YY3UTuqeUcF0VbgKEqxKznsOz1hZ0QDBQ7ziXuaHQdEP3L2S4NMjf+ClfvwfazgAk1Fq2K4lEqTc2L++ID02XEg19CIhAorjALLQhLNUZT/E5ufCP+OUk234DGWXw+5mOBJTamiLWXs+jyV6X/baDt+RgNg7ScbMNf82OQ8JvhFpZdzMg+hmlOaiLjUBanBdk62lnoiTbPSDgM5i1y94SCeFaDj1sYZIaDu8seMi6uDX7CZSIX/MvLSH9OACUH8Otmj2EmRGQyjhDPzj4ZsQJ1JwRlKMUb5bZLa0SVMIVMhg0UN8LY7UAOOwLgZM+wDIUkmhoLOO2VInEpRKFp8DmlQzPgoV3nsSJgc8FAsRKnOnb58Y1vHtG8Itw6U7VZF3J18kBf9ukUq/+AXH78nk5sP6fUGeMQgPIB/9KoUV+ASyK48/K6pyPIjlaXonlVp8vkBZxkyP3GwL0A5FKtWdx8ifxHmArTZniHxqUb9SoZWhvsc9n+DYvFN+0QFCTOb2VxbvJ5F9ejJzGCOhd42TfqqKS1CfR3eTcqNVzUgX/UWFbLHtqU2arKIIi7h0a7q8uRL1/Cu7vwIGrc4DZdQ9Vehhe8jiW3DBAum5mHBuyvLly0hrFXvps9XSQssy66rVwh/9IAR+h2c1eG+f+UvdGuiZ9ul8HaH0bgYZz+NsKFqjhGlPP2DJ3RVE/7oTKLDoBpD9QFw7+wSzWJ4Pq0uJMVDB9/cQfy1zu5dKg9jDMTH/P2QP/4oTf01uKQu2cgDURqQKDBRkUBqGYjvkDyIdta0neMGjtQnpqmE6FZI/CiYVgxmlVlWAyLTDt4dSOYn8JJR8XwmmH6Pe6WhndqHb6h1bovigj5zESaugpV8XKHw/hCpHWOkY6ps2a/ThSYkzHmnquVajB4voutr2Ktr/tF0kcsa0QwWKpKePML6qgK0EXdVm8RwhmD74/KOR249quQARWst05LFeHWJRJ0aF4nuHQzl675VPi5tzjZKyJf31+Pu1JM9SKdu4zQF0HHTI1hwlM/gm5LlsLp0LnhR9oQ2I4JNJFqMYkFH9OMxwnv9zUSfRlM9olvmSa4oWAzyDZhS1VHF7H6VnGkC2LjYLsLL1nNpNVVFud+sZA81YARunNrQk0N0fQLETMTZfsOE73MOO8aa6FW1cD+RyW4eqKZLFNXvePjT7sg+/9nzC+vXa/GD+oJG2qSuCHx/mZdhMYGRFe8aioesgJwlWoxDaNLI5xYJ+N/qvEADY3Ix9eqgSW6TbepTSYStaMFFq26Nbj8ieCQYHo5Oii8oq3XreFGJf1hxJsi1Yxso6T7NW7gQoS0SDomj/aUuGrfwyhD2Hf9Sytebny/OW4f8nYI0wBxmD0Vn1i/WDJSy7C8SbH7/PP8Nn5lGqlbuse2U6eHeVJ3yIzFAASO/pEZEG0VrZoKVA1BG5LWYWEFyC8IybpJ+3SXrkDrSkQkWJuPsDZhiFq6meq2SqQk+i6sNHb2wJJOAdvVZf4X12AGD40PhPz9Hjwkdl1d1z6W6zP01FgF9t325037q690PQw3TXkFZ0Gcmc/XbIJMFerYtrbM7U2v195cbe1C5j0uxP0iBXV+GosxOxfSXjVe3c5jDCRseyFkgxM4h7MuXd7+zA+EsKTluD1Rn/mBARoFALAwB0+sXWmFo2+SsoinLiLgqmRPL4Duamoui0geEgnFfXI31L2w++82Wt9K3VQsyZTGDhqKZR9LdlNp2hrpx4RC2lxm8dc6qJHkfpstWTr8TwTEuUrcRcVHpa9dqKTGlKXBh1RAtJycn269BpFlqtiHVJNlT+3jeC5jXqKeH6i/LY+VD9NWsL5ZFOcKLUNVM1bgusCUXPAEWydwwj0ihhCHWMwqU2QVOuW9DQW9tf337Pb8XF/kl5FBjjCy7FwAZk3DS/QKZkFqcsz4KFp7Bb4OQ3zOfROiyn0Vylyzf1VrJVE0qG96ySmwpmcqOGZmUSE5vUZlvlVnlIotqA+hrc/Mskc5YwsE8CG5gi+9jWoAxnq+EfRC/9UH6UaK7ZiQ5WQrJZepbr4i+L6TAm9Bsd5uThcLz61ls7zgGSymKe0Gvz7uLNMrmvHtI/oRIePAFC2drmaxco736xeq7Y+2G4sgulZJVl+KP/v0aR/fQzYm6xEG1ZD5u5NOIXWM037Fpq+jkyhzsrGNKg8/eTKMInAolzQrfqeoYH6RHXMNpRIORk8iMevaMqDAcIr4pA5KVd3bdPUyXZQBjhyCuqr6iHrmg2S5qE4rpdhRzx0h46wZ4xnOb+OCDWN2WrBvDFoxr0fqGZRzjqyFR6pJo+4BfttidBqSpec9q+xxe/J3/1WS3s7pCoib7m8DOXhMlGdcVxoKGi1848geVOwhsacVvXYkXp7UkY8HaeU4L7NP9c5N7RzkjmWQg5vJBCKAlxHTNgptdQn+QC9+1NB2poKJIcy9Bcb5+ppXpEU8RM2zQutLUsRfTEeHGSGB9TCgk+0FXoqJ3j9iaBQg73x8snLWH6irK22pJMtevOHWIPIkx5jBucQYudSpr4QxiCf0kbxPbe4SeE/OxqLdUgWVQegGM12A9kz41LhDH0PL6QRlCDNrjEX6fqvlEACVTK44wNgqP6T1rKGzfQil0bRTWIis1Es6ybYGnh+WivPVcPgKqxf+2V6ccmOjwEGahE2rIX6RPrC/99kLeeD3umKeexjgg4N/kzr+usU1yFNMPULmISN7hz0HqJIO2w1hxQ0P2BWdEk1nKA5qVuc7tRChqmHlAhNNYm64M3Mcd/lDcIBw7A3UYgOXjlTYHvuhzftN/N0nLXGMf48bZzAoAFSs/+Ioijzsr4eD/JmcqISMqGFHCyoICWaDW6i2QPnNbdRkt2oxGbS3RQLnX4iHsAa/v7TZ0ND2/0UZz6l4B5yr/haOdPkcMPPfpuwv25EXlfbb5HE9Tqsy/C3CiOl2ANp0bm3JmXZef49ujO1KG2ZS+/T0hV1VnfKA2lfaRqcIh18VfJ5a7n4b+BNc+xBOwQ7NQ0SBvc7R0YyY2dttAWrptFLKDIsYgVbp3YPYUk262DNn7eZdHus9Unh+X5Fj8v3t6cl54NrcxNFxlwjV7DcLEhmfq8U0F0TRFbWfDGEtmysIolHIsUBgxfctm/lOn4V6a7nrz5nKLLlftFlnvL8k7791N/OoC7uqdXiM2Fxx4LOepu6FHhPgDDExZyMes6klBc/vlhYWPh89xo5VjFOZqVRwQQe0BL6LnBoE4Ll8V0R90QTMumkUR5edQfeQ5ivCH7FwcOixUdG3J5a/Up6v9eQjjpJlRTAzp2Ay2vocvnhPZMYTeWDaVHrywjkx8XD+wkBaBaZiynPNCgKl6lbtsyphcE2fLTvzZPU7X6MdZC6pvkfxsrS4NKSTJl+Ifl7A5p6VVXR2YyGBojYP+gQjp7F2ShVzM41wJfiZ4Dp8k9MVquDboq3dSpjEAP5auwze6wGcRLRER8TiJY6sZ3Q7ymSM+lkpKid1fR3Y45JTCOX6zL3B5blumhrSCdlIlspGYAC6tP3Wt3XsFmx7H7MEjwGGkGvSzlRWHeg9vLZ0mkDjbeI7741R2g+HeP1qiW58vU4f7psYHo4b32itUX4KVIrxNKFPKq+/8K6tI+M6V7HKNm3hfRp7JeCVuEn/83aUA0R7SV1+SQNd1G0A1lP2uYsbUnJtE4zDMSdU1jVeUTtNy6+nVqQfFba8e0QYDneccnpseXXw3TL3l+AxvfB8rlXw8+d+TpO3Z675PqYVg4wlxZONfDmvUaNRJBn64pe/B5Jq0isimgmdzeAk1ycofZ7//Ka3ZbttHGjnQOuaHtIJj9vJwbPnV1Jnh4aIFtOf6OsfQ6dod82g2EY/VBAwM/1RgT6FFRif1aL4Pt5Qgf2w2nqa05JRIJy8yCgNXhHdIg0V6K6WR0s4sYzRbNVn5l/W8g5lpjpqCRX9X0d7g6SpZ7L2btWN12vOCP0U5GW4DC4HXLoH6yJBW77sib/JOLU3BdGl7ZxQNJwYbXT+xuTs9+tbSDDnTa2+V8KXd9YDV1s8P5bQOzDQ7dzJW8UZ+9X71lRA08uol9He9RZIcvmHCxbwDHk2Sv6pnn9EYzIN2WcYlAage0K/NC73ossj5gAnXs5MIEkrEXlcx1ecMcBBRMp8j/wf6gF+5Oq9G/fEDkhcloMGqR4rnTHdWq9LewN8QOHxOFe8vNfR+ABk20CRbBHOIV8et3rH85R+FFBU1UBENSGgAnJTlIn7Ss4rd3BwxSGm8vQu0PO4tbrufWSNjCbizex6f5rRAuDz49cel8au1n6mpztglPqAMidpPbfj+NdySgKh2BlzmYNU8uhHLnF8fx4i8UPaW7KWBXzTFhf39FABXF7Z4n574CZr2cVLxRVHdp4pOMYeFNbDAPw5jBfgLOzP9ZqIX/litEBcuWApcsZvQtE6WdyoOhMH5FcPTarMARsEmU8U10KRxvTm2Rj1n++fAKYmmlUrAyIEj+i44yASps8wx54HHMk4rTEHaZofRAK4sdnh/Dwl9MZ86Sas41bWjeBcrwgGKIw5pn4t9EfgbksNhlvWz2joU4VUvoI89HV1qGWKstoHhg8F7y1gtR/TL10EK3N+YwGnRdynH2iJx8BBaYax/ZhwwsjeQIZTZcUJ7xrJYY6S/SddGw9Rv6VHHxdizuHK2LQr3YXbmVokQ2N7ZPd0LhvxTWtb+QmDqH1isN9z694/EX+csFtpB5ISVs4YyNg7cjxU/TKxgvHM5xIOUYXi6kzsGBPRBB8gZkEYqQ/MSbmavMryo8sUxapaengQwkGaX/By8YlvngMKTQtsoJIyeu2KgkXC/xlhKvPqPET9yWfDezoCQXROibZp7jsfAL4j7n+BVh6fkZl21czWD0IwiPs6mu1wHoSqLNoThfcBUU0VllMArvFDYI3bzliOV9vCO3Vx6Z/BmcJRgu9YE92wDv5mh1u+EaDh6hOm+PxFx/ETucBaNSeaB/rnzEyXmACIy9kdsbpJ4KQ3SVg23ggD0nSqEGhXn+WXFClPgTdZNdgNfRHhPC18feW9UGPII/YQ7nsTr2Ef8b1ozmZX0j1TWzQwoW/DNxNGiUcqK5f0UP0ifLtNKTnfxVQZm68Pfg+2Yv/mJpbjcM0wpLWsLKMBXzEW+jS8y7TfWFCmL2q37jiUsYH8rkBlyInFjNjD2TT3Wh4vDusqR0gCfBSp14wAhXsfdrZEy/tjBstUoRgPs6wuiI/l9gHYXcxhu4JW+k79KJ1wYt5xc056VyKssSdxlEDs6yBoDL/ApNl1Ggt8t03FYZ/wFbsYE8wGs7VCAaiOJoWJapozZEAHxORlUuxSwDJrW0MIPqBUx8S07wlCEvfIWCnyQOmp9Dx4Z21LPD7MfRleCWH/gTMQvD98MAgx8LWhTFuIDZSxEr3ykk+VfoANsVLJAkXTsi1jqYRuatPP0TjZxT3MtlrAFhUUX8+D7dJJ0rmn61utJTtEofwPMB4AX5tgDkWCxkrSN8hTX24iKVjo72NoE4OJex1/UuvdI/yUxD0B5TJhB/a1yUwpuZTo9oTqpkdFcSqOl8uxnJUIOt0b6T1YtKyxiiptbRj9vNRfOl97Kw0Q2CMH0zoPL4hQwl9cRuPQ94kngkbEZVgUBpSxhUnLLFWKslckISdRQpPwIoGPitwLo4l5j8lhlVW9+RN9OnvNsLdl8PSiqKSRBqhs0nkQUTYNCwKxdg+u8ldCevd1xDr32/6s0cjaLfCEjlyTJYXRs79y531Lyz9Um3GmM2OY3SDcQd0c/ch5m5Od0r1P0fGgFRjMHEAG+VAOCqEEnJKQkuWrcfSmTGYJ7d9QYue18bZPVbzTKqCtxRSjGvWbiF53MekGcqRs06y5LPE2f2bCFqwCJ7k3KzgcLhloDuzo/5yJS1YIVw6U5ZnQZBO8XiWVlbuFXBgSOjUF9KKTMPZdBYj3HDg/ty1/FnudkhsU3SlfA5Ke8GJHjZX9Yo/mBVk/aV19x0tUMhJnFcpk+RYnvoXVLRpdlgyZO0Ld/U4fXocsVgzHiYr1zaUvU3AoWS8kIhh5imV3z6y10xt4p0eL6H5v6JzPDWeekl52GgygIHJzuhlPjMz+N1dRB/Yu668VmFMk4GngSad6bKg3QD20lSNMw50N2WXjPsStp2Iu3b4acGlJutibHlnX0sd6EFPO+0bXDWhmt40ffldbO/9gaIHVOIKQARZMb7L1YqJWVf9teoWMsSTvsvvoT1OUuW/XA5a1J5Qb2vEPBprpo3fwluOu0NGEjoI9CnG71mnIFRXoxGRh4a373Yak7dJVJ2yTjHn4FFREGMA4XE1fR3ljlQ2ZtQfE/jyBD3Qwck4Xo77bUOteaUUkSzVq4XmOYiSVd2/9tyAjPu0fO8Plmk4MibKfyPJ4zouDa2w6IBQwYPzYmE0+8KhjMCtdkMAckVrGRjwVOnZgUi64cRCNoTKLapM1EIqDjxB9Ep/iE6D3Ar1IafegAbNB5NMVVkWxdUW+norXZoqrz/TY1WrUMZYvdNeNDa0Eb6IfaCHKC7vpq+I0JZBpf126/tGfXXgoImpAD5Mo1SqGPyqP6fT5/1Hprd9KZ7rTFGp9ausi6Dk3Pll7eDbib997jig8xngAvJhzEQ/ZNyeGqB3wfypCw/ONIN6hC8KsML7ekhiGaZj1cjwhOXdGemlzdWL8PHQ7rTTDONnQtHjJ7ty9o5NzyewKUFILlub6aTTRX9MisskegN+TLLJ1vA409wo7BR1+6PEg4RqimFrML2yhNBxdXDFXdLpLgcbLiWRnG9tDAqzV7rQU95KcDOEfEr7RNBmxy1anCQzGQ4EFP5QaijDnSDYfyPbvn6vR5lwiZgGKmaQvXugc8cpSD+HFHEweHjPtiC3PNXQiX9ednrwR+5L1J8VWkEA3Z2nG0MKJRerrRn08SXNkVOrjgonHr2uW07PvhWYTwJbGJldVnGFXf/hhoU3
`pragma protect end_data_block
`pragma protect digest_block
ff21cbfaec4bbd248e67303b709e3ac1b55070d16f2c3835639802ed01557a34
`pragma protect end_digest_block
`pragma protect end_protected
