`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
eRL0GHI2519WRyPdzOnFfK+EVlW17WIk6TrA01+xh7ogrmTrjv7ULCqlyh/WpmQ0oGFLk7B3cdxR5PEF7xWIOAF0xYSRHYIaoPygexnRgpkq5hz3hnzG2MweUzM5dR4eH6PzkamSwLyj1WoUj7whqZBdcBu9VDs4DHOaIrWb2+8V6VnuHGck/HtcRNpmuh8/TG0HUyDmFieCaqoIcnOLWHlt/eC+tbKv9ynAnvbfWBWwuvmag+7ckQeesZDCTkDJUtHNHp5YNNRdKF4iiShPz39r+gKXn1QiOYhA/4QPmDUvyjhYDzVLP25Fh0DSsa6DC9z263G/EZL5uHadLqSx1NAdkK0zXvdp7ZxNQnXIYcfGNBDetn2VI19g11/aPRz5PI3dL9mp3YAEkfA65e77rgYHFaJ2CV0ywKDi+nGqT1EuXJkBsrNja6KzNN5VixrPyvgR6QmZWg28PIZVG+G2CYvt0Mpl58wO0rH4NWUJ+g9igIgLa1QaJnMRzchwPUJjPRsCO+60jHUc/z7QU3EJcgqBGflCue7XSGTZQFQnyPnUZWhAaKuiFVnQAQGfWLFm191WaOHWBee43VBNs06Y0SoEVcFwuyebGDxSWGObfyQjYXXjnc4UuWeM2YLTFV5cVr4LKfi2XazxXVFUSqPofGwkkldufYyigTA45suDG675fH+gYRK6PLZw5hHph8ZQ35t51Kl2z32JkkoIyE9alsB/ca5E1hPokyWY+S8XNiUMn63Ce5lrVMWTeAQVZRFDzl3gdt4eDhFdSJK5UhMZaCanoDgjbm+TNdMetMAbBw891tcHWKFN0PausMxwNnclPcPvwvCkoPkrFuHaQCURlICR8AN+gr45OG/iBKYbRN3OFZfZ2n8C3XApCJQSPFcj5v40dglPY17Kb4E/al22yrGmdmmUSIaxsh8xOGLy6t3UT+usZ4FPm7wZgh+k9i7TpRwpt+uXeazqf6Ud8tFzXvxOR5oLywGdXral6ObnhuPupLojd8E9i5iBdUz2FEPiNpmLCyO0/NGFmkC4A3nHLRZHloOxSgF1MRw5PlDgwkOnMt4xrTV1o8L1shRQhjvtka/UrIPjd0wo3+i6O6L+T8aIGplLP/Xd+HDB5g3lrEP0vV3TKR54VWKW3s7rPYMvSLOgys4dA2lHhujBd1wXJMhvyTWNhOhKZIlSXMagoFDxQ2Fh/S8YMF6s4th96I3FMk7zc1y8O54WUTnYsbHjQWJSu5RX/XvobdngSEXp3yZDHdB5fstZPy3sBuqILvJypMOTS2IBu6pvRy5Ngbxi9FJ15b/tCZgp/q6UToPmuI4zD/RkQo4Xl/vO469OTLs2g9pcLCcyls1CYOZ+R7KUpeJDp1JnY2HAC2K00EhXhMjk+TJzwdsOEgdmEWzdpOc3YjNVBi83JU5DlPjVNRr7IzN8fyX0KIUjDc+BQNC+FVSwJiVEMU3Ns0jGqpvy7rg7BtZUdoxHxLeoij+W+T260ItKjbJYycAs9YUnJNcB+UMqaH24hgCTt3L3urKf/TK4pXoPfQgt9dvLLO+Fay/OWCXFTF4y3IVTiz9AceN8EK+UYFrOhyoq7ozdOTf4GAMDqyMW5FuR7dhU+B5gNi2CpuFiD6LJ000SOgwmcwF+mli5MJTndC/rEQrvjWn7UHjLr2R969H2ybT4C+C34405wnbVwfQ9G5cfLm4LBCTp0O5bJC6qcKBOcJRyMH7aRUih84T6w3kcYbLf/a5mpgP/s+EGWyECHaTiOAXqHZHIWyheJLyeTRfG5vqBF1/mivpdtsiJ1eCww17dGEmYU16ZqBqxRWhAasvFErdbveoXrgOkW+dGUgyv95utgR1+KFanSwnytCW233fvqj7OHh0TN5l+2XxOS1Z5ilkCCf9ZqfwwI086We/MeZB/4S/HJtvIfsAeOV9gpcGiRXJ5uOF6eBK5wZoknJTPxO56S0dIuilMs3UvBeKXqX9lchnejstQqYvXIHnm9U62Z86hVWuHXrKWnpCAbKJ46v5akWXKlt/3wrw9CzKr12IyiPA5RkUDLSs/aAiiK8syCvJdTfwOniArKOUJzodkLiD5qY9vApr0NPSLTpKK44tnR/CwHmfOtLbBPUqiq7Gh0MOKNMiiSUsrLaTRMyeOQpgZCPSPZXJkSCPjhqVIVE8Qo+XpiZy4ABo4mDD92j3BEGYu2CwThoXYsJPEvKqEk4sTvXNfRVDTg7Sbk1YzUuyJ3DJGSDD15fhK/WZLWo4Gul/Rl1f2fIWMJdClPDzjVh9UDcBkbvQ8ClY+KZmhuhkXHKunOLmjT/d3Y2PjItXg9FEJ6g8+jRkGWP4XdxZiqUY8usL/880I5wCbToufGL39rt2WPc8DvfQGMvfQisXraTl7/mxLHQ4EzGC1ujmQaPerP/jkQyr3/h3GGikerIWR+SVzyfrrGOKO9LN8q1t8uLFHHyMH2XjPKOPadBk1EvtNUkr69fGnenEZMghIDvJXDJUOgDk3Q+0ESIAt3BO5lpw+IB8x/JXT2+wbia4X4gRzlLRMuv32WMjLQ2N1ipnaPCYrX2nW0rfUjvWcuw5pXX0BNTbeglZPVRZu0E411NtV0bxCLtpLLp6mUT+uX9Lc+8NL3mSxvSmXEWUGjgXozK8rf/X7R8qJHISkjc7/vFUmd+vRucw7b4ZpwWJ6bInSQrAvwrhJ0FkJmC2PCxl6kEWFZyHgzjAaeGxwvu2G64T3y+E6KsLoiQbQBaFFfx1hL857JCidn6qKbCcL02La99LV0h3pstneDFl9ZifMM89ntb+jVwqmv8fy/5NJICgVtSQyNFaj8FFtUXpv9Q8K3ukGeG5n5u0mS1gSpEBq9LTh7ubdO3AoMSgil0VK+iWMnqlCS8TZP9+l6JXupkDkESvE3bHTkgb8Mz2Du7pbJlq77pYf5cGa2q2xNGh9NqCNNSVE50PzvgG8kUSqca+pzwU9QSx90wXaxV93161ZO8/8N74zuiE2Wu5NRYwhsj9uoxkxZiWoD525jgFxMg8Psy2Of15kzKdnxYdIsXZ4Ux5n5dsNOrlFpL+qKkxdLKJ2mbFrM4fc4PExnRNPbEdhhv4YL30HXsaT088ohz+f4LIcdBRNxQjRJ7M4oJF0wGDeOuUioXZKwq5hGyO1oKQ4l4HJP6yU68lz0vSuFOhRQcvhkzFmoFsAYRZ7J/qgczFFXrDXqdrtnA+NoQ39NKwhjigl7JsS3cM1UtDf3Jn/B7+ewIiO+TKW0+R+OEC0YntbZzrPjiBsp5w+XpqbZoXm3m4Yf7VAXW2dCv9UPUWtZlyq+ZOz3WzgR/i4JTW9mf2L8+DDsfOLJjx/r38w6Kq4gX1cS/lfZ2NoPlRi9V4VtwG+cm1UvuXLTgMJ5b2FukFMq3GKkslACaYt7THB5M26PajecoGTHks5zgKk7uSm1GdAPYyxLRQRt1YHHFOVnWIuAJg1Qy/u8TeiZDpfMj6hux4njSnPuSZAMMqRHWcONDP3ImvIYY8YTjhrA36kcrtov5Vn/lFWvoLx1Cm4WoDAUctRmnlaMVYvSMaXhBhOAL5B7asjiLAVTmNlHCe0A5RXYheOQ1R2ST+4vXwHNchXgAD9CV16AMuYhz0Fu5j+e1HgxaboN7Ls1+5TKsyI/MzvlguoVXqWe0qSjdj/fuN5mmMshYu6uHpSTqLN8AzEwPGvYGbV2xEUR6wYUYZuHP/WDckMAAMfbMsnWfwBWqt1B7wT34PL13ajNW2+NkzLe1f6ij0h8w346+rIvxGnTilKlU4k7aO5kc9iiijo8C8islXOwCpAGynhSRc6od9/yALiz9qdd6WqAWowd7fRTtdPOaFcD7WcBFYxVuZLEKcqOe2ROgA5Rm9d/OZ4Opdc6GnJ3OVNcbQdBMtNiC5AMc3CiDQ7T5KKXQZtiV4AQGUgV4jPLcyQqSaSGhsYQeZukE5vDqQAvIQ2pYtricVdK2ku1fuCTJERwTnBjCUCC1AJSELb0uxGsPCpTjk4/Jd8+I7yX+YQeBjZYSEpaUtjuzrFHNbgpbwyMdHskOBh6XeCeK1opVnNeV/fUnb8dYc0WKj2B6lz0JsL1OFkEBVW5Fgu130PEVUaiaFQ7otoXQKxVhdgyZbdWU5RE7G0vu2nNu94k0U36pc7tUyiiN3oKcxFGpAxmoD8XRjqStYkb6SOTm1v6U0LxKgfK/dMQXF+2gQRWgzzuarGE6cMzFr2e34A3PU3kasHI/IHeJS5q8JreAgts4yEsR7nU3ipv0ohudoVH3ujctgVsmh4dsQwrGE12KmwBnKmvyplPaIp7Fy+8x2OhO1u1VMVX/ihVXFkRz6zBhN+2g5TcaO0DrwUde+EazYJByKBGxK0QYRmYiflwJVbePlL8dbTUNGXrEFDXVL1AFidu8q6216vdgPobEja4atclc3u/FfM48plm5YrV2jNyrVBcW0ZHH6eb8xtbLsAScdL1x8BhU720D0A8FXZJmvxA6JR9RVnmHFw4EkUnneqrM7E1YU0Z2mSSKXwrjwTope8JJ2rZkzg4nR+lv86Em/aCuWeZ0XyRIhsl2F3F0oewzZEoq8gRxJvstUtSxqC+d4O0BYpIDTni8HSqjBuWh2zKtfl/BDWvflaF4D1P/1jCdttJhbF7TViAWyiYCDt1zwjU+5uAvTIahdq0yy/wnpFK7gcQu3XuwHZmOlqf2QSAnGPUCX7RO3FcyO8PESOS77OUwAIW0LtSfJrMaIkOFMN9pcX0w31aeAKa3vy6TVk7LgQRjV1SlvLnI6hRYlX240gOlPRB0aWA6YjDKPYlb9zJlPNHcxK7HwLKBe5851PctSoxZSjvYuzlINSp5NmAaz9AKpwjLPIfxXuLJMz4wHMZdcKpZEZcwMeOEEvlbMKPg4m1988RZgJLYUzINQ0E9WyP4OnqogIxqJvXPPHwVRmle7JrkT4uzOqpf1+Y87uh7NdUCTv7EIuapur2fo+HZviASUdDUvbPyDkMagJaVmrmfJL6U5+jcR8ZJZ4cLdJCdQBgf9J9U4vl6gc+l3DXJVuqLkM8InLjojhJUrrYtsSqTw1GuiuhPChHpI91YE/sKLiNfjYoAbVob/EoMFU1PSteev7hl4n/uYHed9AlWqkrvHislmt2NR/PFjhBSntLIDD1UjAjy2+uZQfjjcpfNxamZEbbF4u0A4yDv7zaGK3F/bKA3V18spGoKOA9DFrrS1Zle3uKgbQcJmqW8BMW20D4GcXncKKWqmiDxODRACDtRhSJJ2gMIeFkO8LqL+r/RGC/6I06zGeTOZHtRlGiwCrKOLF4Gtu+hbhY8TrMU2CpJAehfIQ+P8BaJFVMdjJ+DSwfLWHV7wvBamTY07/U947RB1EUQbGvoW2rwM8yXoypo23VAt3wroOkk1cy05S55yDm6WKYv2B35edo8cOqjdE7kxu7YjfFf/CpPxVDmYo+l8XLQYAxAjE7roVZjE0SwPL3EIodY+gc2vIeJUZkQQleVxRWKjuuMUbGfBQL+w32ach4orfzxvFtT3bobFeqJo6DdNmcgFZTQC41q6jrcg/O9Xsg7rhXJTqvVQamA1u6HB49GIgV9ySUG8Xwd3XzXtUJrycp/XiNOudduaoUg27RjWcRGRjgaIgvC2Oww/zJONtXYDUUoSQ0kYtxnQ2BfnGWGEfQsvCzl8TIROK8aaeWNUgWE4oTbX3NwQv44657WS/yNIR3piRHvk+SQhYo3pZ9U6hh65un6CfIVk10k9MYaWm4FMoVa9yT6pJSLve7GQ4A32nzs94vC05Ln/fLlsx0uDyNFurmdaZ2lMiJUvgmtKoYTGHO97imQLPMq48aEbgUbyJSb3gtEE9oIuIB0k5Im9Xz1MoZV0q2yNFNvom1Op0naIiPMa2bH3kJ5tDoaMaspdQLfiljm8lnuJb75icA70rjDL69Y2CLaS0niN2FF33wU37X6GOQQ94tHsaGqDEXaW+O9Myr6Rd9z1md2DBGGcOE64YOIlfVtFZs+dL8m9V6BMEb7D48gGAz/UFQ7MA2PF/VmyCTBcd9x/e7Sn0kEJgaOCWwkIAwqhh82B+A/S/12FIkdObaVWTjE0QI79YoNs6cCpDch50UoZiCY14L1Jz0TIEbxfcOAFB0t4dHSxmpg8T21dTdrtcIJKaXBlXNnlzyfK+98xabtoG6Nu/nTmOzSxK7lb2Qv/3hiYNw9NUFk8+9+OC7xJ/bY7sMOjPnwFPZAZIbXn62g8XHrO+2wmdTWgdSQWNKKxEy5oZrjLn4wXKaiNe3XXzJnmGeLjUSugrxk+YNXK0tH/S7+pJOusQ/1HZ25TE1QHl+b4AKx56nPslg3jDVWHn9JEqBrsRW9R+p+xyOoVp07V317eXYQme6GlAuXdxmdQVYRTlEb0u7wv/cew7xeZZTmus8Shw+T+qo2D/HtKXO/fgOGE0szzcumv2kq7AqgtbmZLCosGB22Y38UzblcwLoG1FZNtNazEfCKIEv9cSePcAwQP30Bs8430rNLAy+3nmYVxLAfgtNtBOZjqFby0VVnDAtXCmj8moACJ/as5KyidHDnAoG8SZPPSusMGEKINhAX6+T2JKYhAVhv9ejCC+xMo2fWbEceys8ZchCfJufHt1Kcn8pqIz5QgqnWcQ9pKB2W6F3LabxDmBWmiCcTuBKtgKtk4bfJHZTDIkFiFw5Fc50uTo5dEagboHlQpKmz4uXwQHA2U6OOapCCyq2oWXtnXxgb4ypF7pwNEm0/kupwfzhFousVR3KlaI7Rz82RYETzyPp0dehtg7wgREn9FfUmV+h6vmZKzlD8GHylEY17hXN2kS1qIfglosL/DvNMlyrNzLrXb87X4nj3S2gyyY6VUNQ6BU2+b73OLvhMSFDO5DofyYMb1a0/4XFyauqI4N+R+HarDxfFxfE61jWnT82M7piLVc1J16aLnFsdjlC/0vtyDLfotCsLd/pgHQc3qsrtExPDZEUj3xM8zLXmkHQ8EK9R7W9hpDGojcwdkxlcGjnlH66xSfcO9ZnFMGvSS3k2iEywwS13oxtJvBqRR64eob2wAzZAhDfvyivBWc5UPZtCsJ3UvW3f1+Vxl0lsFxCB+dKhwu0zcKhFpnM3vTOIbsIMQ4i+w39KexpinbWuVI+5TL1vC9uISZ63MF1ScDeaWJKCFxrv5cAY/K6qugxy6A3JyhMo/lp6jingnS/57RaWOYvbSQJZnSeFrKKX20Z4be5CQ+D77S54JLHNpO/ThFRvMsmr5r5Ht+V/MJqgu0Nc94jKK8wmQC7Bxxg2aMVzxMocnCZ7rbQr+Ct3A3MdiHe5eZ6WbQOTKjucWH2k0oTHZOxwigSXWtZmZdcGMjrxfg8lMbfFfHIjAhc3a5IwMrgL1RnuliSmiOck5RUT++1Vt06TQDtrIg3uzVBi72ZN9g1VP0I35XceZ9tUzGBJp29aqu8wXeVJlp9zraVqJMIBfax46qzy2xN7iapJLIXg6zrhGupnTA7aEAqbVNbQyEr6jb5W/Hms/iCot7oRnD7uUo053lySoYD3gndP35wzQKO/NERSUdBCLW6Pp+9+Kzfow0Lmd/appwX5GRcAW8l739Tx72+JMDVfBU0B3SEE516uvLnWJZODhdO4Jh3lKa5Z1+AVtpeOWeHbHh+4htqVrGSESgkU76cCtiTBgAjFgBJpMFGUmJMJetlQ5WBpbCswLIjCX7CXsMUMcgw9i7waCxZGbAuV0HT1LUBeuEc8ql4vdcDl2Z/nsd4okdldc4KRBtaKSIdZIUmJVydGHHodz4TuB//RxOC/A3lttLFH1Rum8tRcE7Tr/GeVoBEjeIWSFnZzRjvYgNwPVXogWpC1K0twM7fbisGlcxRE/FIP4JNJqVBYRLnDj28ZLSBForzX1FSR7KMyLs8acUM18fRYinr+Bw8+evzJON/PkTBJU082db7j0HlkP8Yex2I1aTj37xRSOVVyuOUq/3pZKaS7jCNR+2sw0mEwX7zTxBucnjOExBVgVzBbzLEaiK7D1QC+9UjEJS47+1aCvIRyQYVUB6jaXbSSsnXJCtqrkPVr9BcRTEiZm0JDkOh1oJ7wGJjyksmFiv4tUOuzBwuiNlKHiQZBf6yESiLAmyYdN4+NkwkyuJxKOwhBejawOarfUDsIjyVlIT1kJhzI21Q+BGi2LailLR9aTMsB+TBvUTE/sEqtccrpQPOmNCMGE73eqL/el6c2HdnGkonQb3pkiCcPv4z0voXNAVRqW230FogyJfJnzXtgkhD9ZF1ip8qhPjChuNqlREL83TH3vqSYU3camWYGgsoYy+jteavvwq9LznaTeN5MbsKYkrCV+wJ+YGVg/Lk6lw0Xn4iCsrL57/507gP5LHAcgj/Hc9Seo/RY4IWb178vhKgqBme3heS/f4oCklAK6o4tPcIQt2Uks7IY2cuMMQP7ghhlajf0RDjAJR7dTz6XW3eZsp/o0550McLvtuNdQcjeCgLNk0X+0rNM9lXhYZf5+ZX7Y7lNLYnWAY5Otig8FehfxT73MU9CfkjD/7Wa6PAyK9E4KCzUfv22rPJdRjsYGnJ5UlrGohuulKRFYZzoeyI98JP9t2Rhac4FWQuvR6XcIZuAPVofDKlyAj5OzfjRrDVB1IWAqJxkkrya9ngvaXpPEOubSliDabDU6un7y4pixDS9CK3I85zMNVOMZiRW06khAq0cp0vqK9g7t3Y/Rb3ezk3icoV0tx+EP3sJF2aF834UO4XC+Nrt8xK3t45evmHMT3KHQ4VhZRv05TKTy9AHp12M9HsgfoBr4yToi36yt7uq4JA1rBinc5nB0KYhtU4D3+fryBTKAdMQgxZGkeT3WG0Z2lmlR65pNFT5qkT8nQvOjfAyIYFhzbm5VEXIejTmFaOZ2pCKPnhS2TMXuhgk7ErKf5iysTKaoND+hwWLhCsXj19i/MEwGc8Xpm1n2oWWtOTPAWVdgZ+scnXoIv2LEiH10y4IM+FeL3YQRprwOpT2TqpPlLosI8yKKv/d7uU/+Au9wx9YcwcZk+nfO0QQNzb5DMq0ByZisSLCV6rI16OX+Hr6Rt8Omy2pBGMKXqGNrWZ+UOp4AAeI0qJaDwLuT+E621qshv6Cqu1NsDfpgSF6xMz4qhyY6y8O+MMXBIbVm+TQfDDaAXD/4LhQnx166fW0blaK0aHI1knvxOehQppnmq0uEEYkSkFych2jpAm5Z8XjH7/hpKcSfFF+zzIBSRAxh/JkPV+1WoVw81SeyH33pLPer6uH/jbEXN7eOQkQatDh1qvs4rcSRboMEyk7dq3eVlVI7fk6sVJqfLiNT3gpSOWygKE2ZYyObZr9gWwa+VJRIRhMlg9zYxK+JO/AajSGFyp4EIiiZSzAHqlDuf9yE2M3d3aVSvpQpIWQawn56FvcNfN5uKNW9tNmSOTvQr3u1627P0VLgB14FGuruls+HvSnn20LqAs3R50PDopt4a1O9LDR80dynfUuSFfGmF2Vvvf/NdLKPGrhw66RCUFYUt9w1Jiwua+JGSt0LOn9QvfRfShiB8A2tEGmKxkkY0nP/7SYmsfo8tx8OPnt4SVeda44b5pInYNV86dDiWo6VMlc2398vSZnXg0qGf6N90Ue+Jw25hEp1bKzb9QvjSRlt+lod2XbfIp8BwhB/FwOYI0cP8ZlCE68RJJms2rlqDqeWMQBzGm3jmhFtRZajc5An4CPnBapVDUJOJbQvzkbxA1C5FVSsLl2WW8YEW9IV2ZgRYa2f3Q3zsicZLqAZAHbvrSQq6XtDMF58N+u36CQ94zGfLQWTCO6yKBfCnRZYIibV3E25LfKU2rg/Q0sUIA+y4+nBN0IS4gOwCaloqkwCMpMaqbBxH8NZ3y/rlEDIz/iXYOiL4hc9GFoNLvKqHEP9eHI8vkZQSLKfjtkNlyrqQ4XjrGCKeWWkXfut/y/OIj+ZiwYOgSiqC+4RLdvv+GQo3FOaGfMwFBewmLeaYmkAY71omQ3c9oIPuwWlUWXn6ZNG2BUCclLEC7VlpE3kdKry5uLlJx9NqhOQdG0SLkVtZIdkU0RbQxBCTcbsaBssQ3gTYq2YG8JM5k4izh1VCxhPJPFs7LdKjCex8p6JPCm/n1XlNijXCbYm7zWcyus4keAXD43lqEf65OD9adKHDfVgPQtiAodQRGNTUYOgSMqI8AAJrSAGmK1jbRyTEx5+yhodNsxqN6Jmukd/+TFElrhyCeX9eWIIv9noYMK+Ea/UaNUAXxlJE5X82Z4YpuAAKn6VyRY6MZ6mU6rTt1lpT/Py2A/ItceJIg4OoxkWCI4PmzLLJ10niD6wA3FkK0KEN7b3TIhDYaFmUS439Nu/xq+MGBHoGl8vB4O2JQpFmTMrGwUAm4cFaPogiVBXPoYE++k+O6UzXrLCmdoh/fL1ZHwsgn5U5P5UB0dqji30lImoFFdXOgPWvlV/4IzIG5zIFRBW8GeKEYOy+weHLd8sMUohRlZh8RfJQocj6KSyesvlAXsD4t6yG02nlYq7jLnD5QrsyasKazp5W2UGSlJrrMXdXuCPT9EpPckbBbIgEP9410Zp6GQ5E4l2hZMGCSG0x2bsDZ0/MGyg7HTDYJF/xg/H+FM8WpzGw9IXPTKShq76phjER7A3tjOzUSmT/znF7kLt8LBa+75tVn1iEkV/0Y87g+II2J+B6+PzDVZvHEvLsJNqqKcw3MUJ2xOFqwxIiHsIvy4oXRuAJ6SBcEjTEWogYNP48WtERPSt86ufSn8KtEKm3Nej+a1UJi13bZnnS1phgFVc1E5+3IeXZQZVD4W66ACNlUw2z85lZK5d6Xzue57xkPsdwriXnrbou6dZ6lZBQti6EFQeZTIbKO1LQsIaDOYPo6StKv6sH2MA47AKPPEC9OmXusEsvl6DxBH4kqwmdXcsmIwfa4UY6AmigFEuDvN3vyne2XwPHO5m1hKxXgmlyydAGyHNoYos9do3EkyKn22yaWzJhsRmjVuKPnez23RKSV/ump5DBtk7KnjiPYjjIK/eRXRVFTzCfuauP9Cc4Wm0oqUCsuN7nDP/TMUf/lEPenqJfGYyB/4at1kxiepagZJwfeIRT6/LA35UyjshXk8ZgCsw0v4NO9fOwJ94UmiuoiqOe8F5dkS754DziCfnDZaFdDwOHaQZXoVoyLnwVAN1yYgJ8dx7P2gD7cbMwFi2eLuPUcof2CDB7vtY+uhOpOQado269YIA+eER73ToZ99rYWet4mIGmt9aVgFPGeu3U0XF+b/Nckr8x3IyOlL3RGqFWpXFW6uaPJAd+oJq5HFI0xsWI3LrAckoDUSEEO7uOiSYga0EzCZqRaYoFjyAGwhHQqdwUYlpHXzdyIA6XxZ3MRcMsk0PzTothjBR8NL5A5uJMbbxxoXeWf4Rp5TKgyifBYz2C4RY4joeXohvfqFGL4djP1YGZY9RkRVJx5mHniqVRBQzDSF8Lh5Le+soEmXPuaqlMvwVdcUrtpyLzx32wJoFk6DZl7MPFwq6F8yyi1cim3aXa8Ba63EzcfmQkc0/2OdoGcL28DLDfYMqTC+HBP66vWza+RDa1Hpa3NEJOzXH0vrlvzKh8c2JqAvVVTsdYOpOEgCeSrFZxZt9tEzR+5TtDj6zB4lWxt5IH+TLnXZpJbK+ECwKhPfhd/jA6ax8hM45NNBIzlbb7uaYLvk975TYJTPpv8wkVaJkampW/A1oc4jPg7RSTrp9WreZBwWBZeqH1E/BBBuZdxepEB+UwW1fCx52WwvUjkeSOCiC77ot0NEhAFrhYBpKSueRmJCmGeb8QLy0fslarpkaW9CIGpffQHHVmiqtRfGw4s8EtC9q/2uyVP54ODjlhXlTXUOyPBKGmclrZGeVzx+4UlN6vZtv0w8lEK7ci/ilwDg8PtBtKUr/T+4zzU1m8yFIse0KqWETKo5xcxIKBAKlPxUi6pSyT0R967ykjVpoZKV5z0ogm7dPMoPAMYbt+W5urzBrnYuJFOtd6Yn1s9P/PxcEmEjXmqUsDev7VxUCK6xzUaDzBzzJdcixoV8fCjv183w0YaQftFKl52sbI8N0CyT9c08+DX56SvIghdxfG9djQAxVWZbbxEK+yAM8Wm1b+wJzIJzB0gtA1cimAgcrdmHQ+s2klViy+uGx6qafnFD0pRMaUwfThKplOzE5ZUkH0C7HYb2kbOdmSzc96NTJUDojdhfSEbR1wOSW45Mpp4OT8RlTYExg+C0VILxE20pyNi0D+pFpl0OvjEE5eazzEK6NmQOyhhcs7E+oQDtUPj8fM1tGan2OSFnPx7n9XWskvkYs1GLkglVrtY4EFeszlOPkK4eX0fBrZ3/KFmx2HdlIzUjWzIpaivAM8uzTF5zJr06mn0pDAlExRuOY2JotDjAl43KuJW6m1INLwYLoJWK7uMd7G5/+SmLHNYF+fHbnh0BwUnG6toUVJWK6/VGHN35SWotXMzIr2kf8RxZOI3MBbUk1gK5cPxCGNrBcd1hv+jp20IKzFFo16adR/5SOwYEkfJRY8lzNlsaYbJyehBYmynJfp8UwiI0vDedUifpi84I+qa/HkFdH1CkbUDgEJtup2lj0cd/DvSVdwr85eS9SFp8bLqJUH2xukh+/+c7zg4Khlh0VPoqtexj2gzH/1YOI4hnHdOuL+0FN8Lw6s3a05gEwbhh4HCBZqkZtBfMp+wkEMvgdpUXzPBBL5PzpRdUaWKePupdj3LSoXE+l4m+7ZiiFq3Fg1ocl2dNrs4/WzdSVqcetDm4e/4vtPqYaRHPkt544DWJZ8/OQ90ThzoCkw6WTnggeWgiFDRD0rB5GVfwI3qasA57WFatX1FoGmfY6zWthrcrHTi0fstB/khu/0L3NRYRKm7FN+nkapuADQeCfeJDtNktRkF/UiJKAiD4bczHMbsrQgzqmJCHOhxeB8yvWokVOQmbuLt1xt0adEZzgBDpRHzt/T5IRAiUe1jbwEOCgSuN03uIs9xrsW64NjQM6/qJUrDIYdE1AYqr2hYSjIgGn58nRApGKv6ta1qvA3iy6XxvmVzhn+l42FOHTyeHVgV1DT/SYpJZEPTW7YVIqi85c/ddQ3jvtPGGQL+X3EtIDhvSMAMbonyGntKLELoo7aqxQ2sgvHRPwy8ndBtD7fnYDw3Vaxskm+HpkvXwh25P5lQuEX+k+Bpe6YagWMFzZRyQJM7+gPpgIkX7R/YZO3xOh6HTHZ5iYtpBXVj+pGEC/zP6usC+O16Oj81m3vzNaqjJLBTy2R+5iJaQ96nvCQ+Mj8arrpsRyiHq1PFh3ze5ZLL/cg0TwVdoFVTE6L4NbCfKaZ54ZeyJLo+Sbq52D9UStCiMN1Z1cD7wb5aA5h8CxcxBNX9rXXdj7Sp3ZISsOC2Ve2I5CKaFMDIWqH5wgtSAIh+FpqUrRCIpn3Abp7+FyNltuAhs5RiLU7pcFQNS1IXqoOu6OCztWFd0vOKMi+4trp1NwKFRzWCi55pmalqe7ktjTW/gTl+dCTWNQseiyLR7hyHmTI44nmpZMcMpnvHkefAdXg/R6sOOvRX5upMHuMXJH8MJ+I2i92+VA2uCvx4qqYqX7GANy6u4p9gSbs1TWMnj+MQ9Bu+OUbqgeK0S7sNajcrLZ4DEYptXt6q5mSHmrJtCYiOQFi+o01sFavyaDgh5DCncIpg4mqxK+v2VHNYZ92J4a7ABJfIagNdzUQAZyg50CIE0kVSKezEj5WzAWDMxPDqw8QAU2+xyHBvNRLE0EARI3U+Km6395VlicTyAl8T2tR4bGVv7z8hhIJgYk1J9I0S0XEzPLIriMHPO2b26rwBXAsF8ZfInSWFK/SQPz28l+r9pal3CzuSimz0D0WSggt+KjKrmqtiIG1NxzbXArKiLNLtCN3uLySPGy8KvidWnFhX/t+XEwMuEg6wP+BytDh+Nh5Vj7kR2oLglr5cX/W9/+NQDg7GCXm2bEjuW+iAksmd927NQF18zuAa3jsjI8h0ySXkQa6L6PCd3gP0E/B+BTlHozTxwKkFad4Z22sn+bhe4vnomVEeS9LPQSJYSOBMuul0oRRanPiSVCCvOETAatO8s0+OkiaqaztpOfEaOUfntoHF+fEztpPhlK02SJGOKBeUgl3uEJzd/nfZJyboR4lp0jYxwEbhNkHloEaLbqhT9gZDNTDhkgGkgRsR7HkmveCSPubAhCw1fNPIgABxhapaM/EQrTsGKjMu0x7LOSr3AErgct3+8JtiGtdPDggqVZE7M43ykF04d6DaLa6c5j6U+/6DS82okr1/mslvu4WMQsEIWigWHG18obpNPCMqtvyeciYUThwomtedDVWtjk+5uiQXFyv1go4z1fr7x+Uvh2r7ltFoRDsaxAtA9npwP5Xv1agGc0ywLpOTos7Gl/F5Q96e8oPoL4OUdve3clNjhAUWct+rdl3w9mODqCApOpse7LiU4q6OXtkbcQOU5Bu1mQ4lqJi8FoTEY4QazOmfy24l00CWad1PsHyBpJGnH2wfMh4CPF3GElgAE40MlcSWBWpDDxTOsyhknDWrQENWLm8P/7mGJGxT+kjFKcA4QG+z8pALDhrvpOOi5aXcymH1r7PlU/Xk8w8Nhm3xRMWm7tKVwY7PvfofN1qg9nNYaHyEPn4AHH8LBdFtJReHyzQZ1YYvgWNF/LHuirr6sRu3R/ttppb3cw3Yny2fpMViIo9selBV1V2WPt3GOVY7RcNuXGzEv0XPevDNJ1vEsjC2ImkLkosPGnyy71X3EBiV0YE9g4nB3lp0lxn9vALpy98dX6bqEiPfyS56ksSwJw9MWSCnLbRepE2OWZETMeDFPnLJCP8vMiFKHVRA3k3K0z9Th3LrouUVj2w4h14FfWxNlKSPVI7z+6xHsu69Fnr5wykWdDijrDDcX4wWkb+TsESo0H6//dp8UmXJ/Ie7VsgZ+mmDh/OE1HyZ7EblV/OT7fST6hnpUPR1yvg5S8a4Ow1GcNLGntPtFo+LO14V8tLvmZN04/cQ08PNYEEIKpXtBEGxS32mWEmnRsFRpz195TjnUM7tR+gjS7gyfLvcG6QrlL1/LTzWjtMyyzoQNKyMcm4narK/vtN+1jLnJWS1Bi82CsiPSD0FpzHQsQzSCRPZBYMN9TqYGCqKe3D1wB8Z8EuM/DE16N+h9I6825LwDGdeqVU3PZxRazaLSAldSLXlB8VM5SfoBB1PIG5l/Qb81MtwkzLVJ+ntxb+1aeEPZ++gJ3JdrVWoacey1Pfv9e6m6R2LYR2dLIMNzymEONRVX2kEWr/axYW3NMInflhVmAZoJpPKxnNJe2L8vkuv/HNQHKEktiaqZxVmbDQykTESaxGJu01HGCoT0vyKgwH2AbZQJuQ8yqWiJDMJLoVQIgLF26RcLZIDS4Yo0V7qYsvnzlJvMiEswE+CspmFIVN8juY8sVyscclC7sLF47ZCJsB2x9ISKNfNk6RXUp6xYyBKKCqLZ5ZAN3dpkvBHaD8ucmZF2A30kW6Eitr8r1i4bbdcxgkgziH2YnKBwjwcNY78oZMCQKSgdu3+N9MLcqO1Ruw0Na2d5VXGUU8xtNF+YX+eqD5/6LIM/33tn06UPMXBxN+vFrkXz/8sgzGjSRO/SFtzh8GUoZdXx4Ros/B3j+/OVUjnncN7AiEhAPGDFRYherB5a3DBWznS0fcAzgGKXU8/SKzWFDZiGEodMpLdl/14kXCP24xa4wy6YBeTMmVt/xAKlMGORXM3Z42fQOTWl6jdIeBpDyGw5EpwiY+MN6cB6OjtshlMy758/7n4H1fcb14ECiqgAI/nWXacn3Rh7wzVEvEGlfp6pGvgOu9LzYmoxlnSs10pkQrqs9zCvSVVpNSH1MlMxWsJpZyg7sOv6s2lOrUUbZpkzVeuzoNS014IegRDiirDj8fuyTGzKLBbHrsz1bMQIteu54+UtKZupmsS05/zNz0a/Kd62127EMjJ55nqsgddEIHDtGgyV6KAfTxJMa6jEoSZAxmasdKUZLu96CqRXRkkMTF99Uz2dj7i90+fnhpBU6/0uCH5RStkmB1kt+jqkZZZcYJSOwq5bhPROPNuci8T5HC4RtLbBwnFch8MtNcp8g3kpHUMKYD85Qm92KXfgouEVbPlIMY+0K7TUv65rJei4kr8nq5fcMFXVS6h7EOmq1TWcjuI7x1dLZUrJQ+vcR9s7MNkhJjgMsLq5OWcQ4Dtka5QKaK/SDfIh653qLGyI/W0B1iBICJAZ7Wc1V1eTQCB5u8jPDu3uw9wDQ3yZHlndiZckZJQ0T4WOdCu5b7r3hXmUo+++BXDzPhAgGjPQZNorKljsntqEOwoA2nJghcmtE74em6Kpu/PjaBxASxUuwCtbkHd9phVd2D8OTGB4AzmNXaRP34evcQXcwQEaOKXQESNLG8cJ68hCOQtVnNlNRqPnoZY9X7S336jV7cjuGb89pDP+aNZYTyAYetgnUstC4TAUcytOs8lbe3MehKKxuVSZw5vAq7KD7ENNDgEwvMK/VjOq39Aekotit3yzACdhdMmDkOLzsoRKi6fLeLce6rD8bpfUA81COv/VYZPxXSmc3nK/aHtlrZYZkOT2XF5M1t4FXCl7PDG++zpFJEJqkwdf7fb3bZryMNNY5FX7XDPR8b1NhOr4zKUVTTD56DPz/CgwphXb0yZdos0AM97jgXwqAw1/DM+aH8j3zH9rcR00Bni7sny1hZ1R+9ZCYoCvY3CLdtvz5fqwTkWA56d6ehYXySa1WCaLMxPEZYgBJ0NcrW2qexmJmRx6hTIvcHL0PdfhHhau7V6d/xtGKxNEbhbMZo7knNyiqOnKZCUrO0QfOeWD4mQrkl/cucegOU/E84Yqxql3RNa3WQppbVGYhsVaWL2/9CpUYGxYQKplyaAK4D20BDO/FkHd298v80/9PJh9sPFZ18GIu6wQ5kZ7TLCN5DfAKv63Ibfp5fA4HyaLev66eRYilBcQCdyAlOQUmy7pZlPlA7GogatZEYUoU2N1DbOg9cm3lxw/5FHIuyj4fzc6m6u+5MDHeRmi1uH8gyu6Ob+W28NijTUeJSjHOXsRMOD/zjzh4uRf8lERqQv+QVESxQbatACZg4qzMLGi5LioRbY05zqAUxdbxtocpyn+GFlQ++rnvtkndHJvepVkvKEyHDnuQwPsp6So1yFS8J9OwH01PsXZ1QRdqz+JVKtxJNm8sD8mvSu2Hfm2FJLXBzTMQWc1xQ6JMKvw0a1J+vsMP5GD45VEuXyPs6eAVatLoEiScAcGJq0pasMsJxhJiyyFxvsIfoeWRN6SscshzwleYl/w4o/yB1kJEcbLl60stjiapn16d+YLqaUcvoW8eaIVfO7Ax+6wilbAXqeLHw88xBDi7IcCp8mV8vPCp60c/VDThzPh6kh3oQv8Lk8RNYi67WO2uhbTMFJt/IJ7kvEDeZxKN8Wg0Fwl/TW3HcmeBKuBksLK8V2AWgj81M5HcSAnFDoLhm3laUENFiRYHmfCa1QXSj2dGyScXA8GvB0ugeWyJsiAeZ4U7G7riVRHFHE0Fo6wUgMpdlP0f8mS6u9VUjGnughxqZ5SjkSXtpK26yJ4tB3BJXUJFvl55YafB42u3zUiIz3iEJ7OXX+H/AGtyLibECH1TCg/bhI5AN1IAU4WsN7xGTRYoQ/PvxBCWuXP70gdyTjMGYWv8rvz5cNAX4uDCIy920Z9YxZu6PNnID4HeehheFyA7NHAmbpGVGJfnIhFHKMBZU6eO0BC6AVmI/2PIwwz+0JfnKYoK5Ha0siF1SXls75dyJjPuvJH0vKT7mgTzxqwBe2JbkTFA5iZgmGSDP+5FYFQC3E63MnAeDLW0ioLTFznaHDecaPGWOOp6qzffgB9qVNXHwfAnJX43P5UctXKfEAOR4dtSYj/gf5HCh8JBQ9l1O7VZDjlkrQXXTDyIcsw0cBHe7lkzbMVg2BOTimctvG8hAKykq472U/X8/ropNSwSbbgqLi3JhGO/UTCYtm/gRIxa2bj/IOBbfBhz9z5+XzjIKOWX6zhXswM/t8r1E4fPJSV41nzcSPYfS33Sr956/TzX3Aihk2YOt1qRvqQ+P99ZkucKLScV5kD7bWMcjOAJHSdVh+BGOUyWwSIHqlyvlnmiWJGSXEN5+2Ju74pflKbR5WIR9bpcwFt19ogpTCbNx6nh7FKszGbs2f+3Rflh4rsqVZHaNw8fNwh0sFNl5N8nYz0QS/aXiIlQJuV+dFryh4POiuxHtsD+LUQB7bT4RUvGVOLsaney4cMdbWoR30fCc2hdItin/RTw3ywbICpFfZaUx5dPR30eMBPXO6ALnjQqj9aV95dHqa1fLCxhDq4+Q86BZqAL3b+r8T42hoWrVx4gztO9xK/xnpKDQp2J48cYxZZoVq42L/NZhETSr0qF15QRd8PASJ9ZbeEJIz7qn6vWDRSKAuBH/1Pqeu9m9yYYZjQ7M6BiPfiMOHChZ2+nSaXVBz9zTlc3sv6h8by2hpkBv5LDHkk2V0KMhwsz6uCeq0OOS9dkc1RaXU69dgW27QDemPnQBnjLLhnpRtHswAwtl8MNaWlIwSGVbMmkpQ5TIXJ/Cw9g2XLl9OKE1IHituaw6FcprHzSbT7VJSHDsCjsX7Oj4LBcQQhN09vww5ylCBnMQqEnGpd513flLEsZPVk51gJlvk6jGapyXdg0EPNBps+0lCcg5NSYkViUIGQ7KAs5HwpqDPCrbFpRSBu88NIWHUvXPlfI4imNq62GcIOyH28dsap6b9D8MUz4+mYwCT+/EFgMoTuyrDj8+auX2iOG5WWNRAZETvaLB0e4s5nTdjebEfljEx+Ul2uOgeJtNn9ZTFzdamx8Vz6miVG+7ba1MHjbUlc0w/O5yelBe0YZYcp8RA29n0sdB6ZslHj0wQkzQawyFP76jrMQvAHiBPMdahc4UZ4LA+RPHmna19QqJ2EfQV5+1UZeUelPBhcjX8a82Lc5DSI2MfZm4i1E5fu85BTPCPcG8WRxStHKmtq0CWrXVw8dEMUjFzgrDnfgoLuUc13794oB4L+HpQbEYl84pj36hAPxioVUMy6enZ4XvEufoRj+O0rByNrT0Sr71SyxrVjPhBn8EDk4zqohtFWnzlFkyWG5phYAgNkPgFM8J4hWnx7IJmL/kNQjWiX1DCAiXyVJLRdigwYSlI/4pLgxjNvZ9GkcJucfjnF8aDHm2TN2BPm8gxjlVVf3AT+C6hosanxDjMsc5/1XuhlGjeOy/D7qW0AkKQpPLKrUYVI87HufNGStMU7moK99xIIPoGUfe8pJSmpGl0vCMaoZ8mO8EUrpPr1yz5gt6W0aIFCyuvRNwdV8J2RfwI4CW8LDQj60PwY1Yxs8Qc02otLb318KxHqXJ2Af7ZGKK2aboi+o1uWiaR8420dxhEXKdo4Y8tvihtC5ZI+Q5SCgU7jacqcf4+7fQs3PVxSzwqOMH+3rOZQ1MGrulPwW6zsxYWOUAEyY77d1hN6vm2660Xtz83lpIGd9/4zqAv9jtk1Ys1C8zUY+Eq/R85c3k5Ypu888hfLf8O4QDvi5gJjVN7/gzPuITGIDeyICyTaC2pT0wOF1gRzVuWu0TVZnbKzx4HROJpNz7K5npV7/5/uuEma5yIMkIT4THMUzH1gZhU1bnxNOScbgXP06A9lTbZeKwjGfOQOafXGEnIPo6sq+quAtwuEg8y3Dq3NzFgLmqcKcldTDCgHkkJ+LLzPzyntFliOv/+M0n+FQfKPdCDja8ked6Ano011nVDD6IHxn0/VVj8+wlpQyTfLq1wKs0aUx0DVoDwuFpel3925+X2fcrX9SbwqVV2eWHQJaI8NLHrySQYNVrc6k933H0t7HhfTTBBgyP4nE7Sjfdk5ZqdmruYj8Rb0ZON8AcOLf2mEz4/LdJDj00J05Bi2KZEZFsxMO/dpZI2kcaHZtrSmhkE1S9wy+o+/KU876yhyXLvzS4LequC9zV0/FWADFkJBWH2S28o1xipxglXjWIIVvlwEurF/dzAZiBzqaBCLB6T2sYk3sk+Gc6zNs9dY5g9DN+wjcwlG+As7DonVdMjRVc+exM1tDsc34oF+H3dzoYxyMUa3zdrwYef2mCjLlFjhohO3HejVCzTm2J1ArGGV9dzh6TAfxoy4l7ZWSU0wt1zHGEjZtXWyCEH3yMqCkNUzXGlxhqLoO5vlZA0aHVspl5yV14kTDLwFvwrmjLTQP3DJWNEmonOabNgX07jAD71/xohqgewOdBmLKyQeM1FBBFdmKvVLtgNkb92kkDOg+9Kr5cr8V/WiHXqX7pe/Jp9vTWKdZGY7aPfhlUVDpNAOBES2BpZVcDhzZOc6BhRFhUIcpFWIZRjDXM0YsyYEaZSUEP1z72YZe1l+Otvmoko9ygn93iTEYdmQeOGL/DwH4sSfDBFAkEqoEsIJgEmvzCETupMmvDkApeOsgcRKGerpLPyd1MWIv5FPUTo2OZyAetRwMaLBI1WtJXIZOCyccm14Dc9uSwyV9X4IPbLD6jQSUqjQcLWrCxAGmmhJiqduK5uAkxEeQE3cQHvUHhpSUaUG75LkvELC6DcmmkmGepaBCx99vTt5XgOfXtzWKEEGA4KnhL81n1MgY7fmiwe5hJIk+4y94ixZEAkMOsSlBWpA+3yJDaUpw5FnQX+VjWFsFUqdAt04hZOVPevUUyKCPURx/Y5L6Po1/vwr9TXEmr8YoFbkivAJ8RdW/97x2helI9RPr4lxmUY1v83QYe3t1TegiKow731Zz6GEY3jQB10WaOEv008bTQvfYRp5yfBqn7hs+dDnpfV2hfMB/rs3crzzC1GJnHrKjgOHrybbnWVgVU4HDAm2kuzM/hsZVnaPntx9ZTrnHHlA8knta6qEKcWq4sBmMWf7Oqni7LyIoxFj4bGYYq5sbn4pJIpbKhA0wxrT8ndHZht3oxiRo2M+U69VhRlZU+ETmDXPenw2MzzlG0tOAYvQO0LVw7mnMrvh/DJUNyvNdWo58oMKXkFkZGszbJnDVnPNaKtptTGQyfthjnYRQP2s4tPkDydVhBQ9lEt8xk3vl1Fr/rWpA36U0cl/nDLY2rb5t6boz9v9xNWckyVItW5Xb+ICpkahzexgfJpTmLuly1lVF7u7NRUGlFpkrQ2RforEeq9T6eqPfPhgblBZLdaMM4NfzbaLcdxNkGkCSJ3daECSFRdX0ZijnqngmZ/f4RMRuUUb74QnYhytpwfi7E/a/CxE+ZLoCCs6hx8v7icNlAxuCp2ghH0epLN2pIlMaUr3OKZHGPwxAHx4VuObN4KK8taWtcR6Hie4zdR5j824mLbCwFhCecNnuYajQIZvz8OZu4GG5IQUCW+ZYWF43n432fRQoYp0Q7E8fwt/KRKK6CuTb5DjrQtBD7vZGKpQ+m2WC6Tq3Q6mckzTGr5QKdpEuVQFz6BHuqOrClNDNZm6AHwiQ3boga1IhuOyi1Rr7LmemidzY4bR5X8NDTlB+Mg0iUH8YyNahWm+aBkDX97ojXGUCWDUmKfO8jVI9/LLGWHcaDnjJHHTD6kU5Vv1TUrS4U+/dfJRsqj/POIX3xDdRmQptRF8CnXZOjYXoc13GdirVrDSp9aSIJ3gbG2/Bkf2/vb8/QP2sY0SdU/qWaXIM08Ts4LayzKwi/2Gc/gBnm9tP2lfjptFCL7RP9imH+4vFcHUarqu+kZvllegiffVzsHgXTdlu+ih7gD47fhgUvYvmvT/91fL4TpKHrUyd06d9dgqz4gxbvQcet9NPt/q7/WxKvVELZU2Pk+DOIi1ZOt9+Gf+SljZHfX06vxpAtdyZ2PbdXLl3uqvMSCB6T18AN8nVYMW9RAHd3PSvnp9kzPr+KuxQlc9FpmMOQBTL/Tbc/E9baqar2l72XPlR/hPLkxGBenyfRov8mTS+P5dlE99aS85Bbt8i3E/CML0f/tyMvrE4TSDp3kbfJGkdV7mQWFE8r4WayWcqzgVEyrzW+zvXylkYvARI5THicUHwXbgS5o+33zLLlpsGhMi2w21wkmn3wqkcCy/NwyXC4Jb5xJKo2qPjDSIJ8KTbQDf9PHe4Rfa2guSkCpoM9BqWkVfOLohlM4GV1V5xLE4RrOcHcib1FaoYdYQVC+edTGz7Dz8laK3onQNxUvsfttgZEcIA48bXpXf21S8UPnBV9AW/Z0n2UQyezO6MKwDFJywgs8x5e6McKa86C1svjSjQcZFOkinBbvtACt77ONT/KBExyxCbcndA6A8CNtqi1KUQUJuaibJ6dwN7szFg9/FFYeIDz08OPER5HIvklluRQkaLu0dv3C32oka0COsTmZTrandj/+RiZQhAqLgdfPjLRUDr6p+LTAMYzvwZwtcX3GdfyH0aPOVJyqkOEIWGAppMoF/jXIlMkvf31VBBTR54LSjIL12ptLLbMDEvLEFLJCnW0O+TmyZAI59ouho+3XFPIkWCNmq7n31UALBIe1K+b/Iju9bcO15931i3wt0FerR4lRBt3o6v+EKN0MpSHskXswmMUvI6nvNOtBWqKITbENGYNMbgqrkNkJv6074H6qf+Uru7UHtR4BQnOswV5ebIQHBQjW+vpjIDc5DD8agIdyGnvIi4OeGmJBQ+/NRqPOonBmrphF6FSWAhYVGqnkokWgYLcVL+p3BudECloBa6jghXqTFx3WmToCvOcyQ2PaKbKZfQvlhI9ipGDdlhGGcghvTz4qSA/i9ezLH38QJeEnvjhPlRLE1SOC2DAsdSRZOvPClrZSQHcUFFi+nuAGXrPFZeEpRkH4a3PDn0UiaMtaHXonIrR2p34v1S1gfAFmtH3MtvvqjbtArQ86x+AnXddP5J1QasPgfOQtxG356Z6yR7eY2A4bqgjTrQHE3TWxyTdHbzxu+0T/eWE8PeEcjG2LROa94Ip3gdwLzuy6yQZYjXRZFmmhEuMo82p6gIakR1KD4RjXAfA0zQr0cuSrZCj6AsKMY9gcYvql0jhhHzciCAX0q+sc4ojpOT1MeikQwc3oePxquWUCDQPDFBlwuOAK5YJ3wOOuDq5fdH3YJaojWWF0ml/vY7YeN3FuOUikXnzpN//IyYjoj2oQpZK8+jdSJBDbV3rqx+CwRuQyviVBREb/X1sc5nlZlgAnH2eHhiw3JfB+U0phCpn5Jt40PzHD+vt/bdShFXTjxQ95gckRr7qLnKMvNLdm5T2G9yUWcu/EipG/QDcfLbqQL+pF6N3+eRoI+OyfdzYDdUgId9g1d7OofoOKYVoU1BFkwyzOAL2Ha960iZ69oSLBgXcSFyBmOtnTaayLKN4fBX+GJNd+hXEH9LQp4sUWtUQx3XUQIFW6MPbIosklp5nu3kNGeeZbTTIp9kHv8CXNcSAQE+bP8hVPeag+HIXI8+e+0yyVxZsO1UVtUBhkPIA8A08rzoHGutpEAgMOBfvjdTdCl4tMiBpzsMAeov0gfGt0sSg7QNaTvagiCUIltkw6JJyLPyZaSeo4aBLn50H/5uJPscOENhYH9XKg254kP4ThsYpKwmbuXB1hUVZTRxrjH2e7Zu1/1j8iF/HiCn318m8Ii4kxFlpYRlsiYfD/FVwc+bfIF9Poa7FMmQQuFWkclTrzWK5jNS/7uQNQjlH15ZIOSxHm7jCtoC/T3T4SnZgCacWgKH8wBPnP8X4OzqS8oAyDEwdTcy7SoRAEcLG60wD9mtVlLLBDTUoNBEvyn99kiKL0/12xgdRFOQb0GOwAtcOj0tCqsqmkZEqDstAKBVlcggEvHdMEDx5QZ2irQ3HGOxRy/jZSSNCpqp+TnX+7JL1BczRmXi/5lckk5jYzW+crYJQXZPjwLjbatqiseSGtaT3Ag2ixmDoFHqQyT0PQV0ti2Ecl2W/7fcAJWqqVDS+dybV+xXPsJQR08Dg0v9tvKGlK/D/FT0XqKLGyBd1qDSLl8dg4h4Vava4EIdYF7CWjBb4DBmzdBsGFTFFFd6A4YZ/gG0dw2HUdf+aRn+CazCsAyESFEEW4MhduyfQybtgklIEK1Bd7smmzx+h1/kvgQol3e6xz2vaEaHD60QnuCTfah3N875kZzQPnvSbfjlUP93Yf3TnZESz32AjWBSkLSu7lcCIgkH13B0JWTk+VDrzC/bHWPxW/TxGsG4JPgNEpQUe0+R7TMUOZfdPZQqISgWTS8GoyWEia8uIVlfmwRj3BgByg5jDrNahN5s47oK+nPlF5jxgg+zG2xqb76rA8jaFbEPvvYa929MVwJRcj/y31Po0dcQX8io1tkSnuW3j50q0/gTlYqUuPfqDfKrr7Do2SwJfFei6qltOCE9hTaiU27sadghTb9pbJFu9ha2Tu9PSTgbjXJAsNaayI2IZN5Dv3QpkSbx9GXyXRNIgqSLQYSMTp9cyrCTq8sKZVw3ml3qFi6/EM+kDDYz5K9bk62RCj9xMN9FjN7vHwbpHXSdI0LPO0m2yonU80jEw4NAoJPt8cVPPqZ5Q/e8+vhcxrv/aTPJnHiPbc5rdGl26j6dikY03u/mjfz0qZlE4PtGB92wZwgqTCrPOtT7NhmN3X0O8StajJgSs1Xgq1su30lH7AaUtpXuB/LcPxZZIhuZYMIVTnP/yfSDdvegCmuKEkCJc6WWAWM83K0XgNBZ45Pmw5Q+Stnrrf7qSmjYqiVjPyBBK4rJbNgS1SSlWK7Ug/VntjCRPL4rLndY2UpwUcxY0HhVMOT13r1ntoUCYBVMUdT7b7+eYX4Izm/oy0y3igeXXYmNl3WSTumbH6fiweI9AJ8Qikqc+OI6+P5voSmdTKTg3bJUisPSTz8sy/qRDLDwuBilZMvYZIS4sHqf8PkFLQZPuPH0DHwbFucJOPZ5yZhYpLZs+k55TNXT9a481+GEWa3romvHyHVDyhrxs+ytjojZjQsIT0X39S94zRE8a6m7oJ6P/wVEIBSmGFEZ4//QoZsVu+mjREObXDB/KFsfZg3OfviUShIJh5e8SWRuqF+9G7Gb0Cs3Nt35foEWkjRJdPZuFrWqUx1RFiVIaBwDltUdVqcXtwkt1tZXtMKMwvuzMtBoQjo4J78q/ht7b6SBqPSuBGIbXPuGXX9JoBYUnEpRDWhrmY/nUUZJjF5u6efuYhqTLlX3MprVOM/Pf9uqYR8gUpr7/3IrFarRd1wKZ0LPzs154/YllbTq/kieh6qg/D6IYd1swZg5QaHam4fVNRGpjIERKmP5t3AaLNSIQ7hfBFXCOB94NRskl1m80QjewzTDijieqwJ9VFnJVNFkfNbITc37hx3qfILYhPoZ/dlWOCJv/lGRavAHtBZ/dKSrRC5HVJ7YZEjxAsb2pMLT5CDvn5R/ngbdW0Kley+pwu5N4xTR2Hk4kl7uiUZRo0YcNPmJktQ/lgIrgnCygDRp4iE5DIlWlImxXDPMqeo2NhIXJtKEYDFxpw1iQOYQDzeN8upE/KxSoTUpRvsZz3wuQXLNnEfWHHAOPgHG1VGPdqp/z9r711ymcJxA443fntdYybqEx2fV8GQk3naAa3JESqAddz6zyLrv8+jTjyiOjL+TVv9GjtEQTp6RtUmCRapE0qpvJisRCbnqFY8vy/LJ87mhXyaZf64B1dMwWlgfkY1sD3K9Nj9hy0zoC5/BiBVjndBzmAEsxhNxYJ7NhSAeXMkjN4xl8bIzi330Ad84D3YNdpkFHhF+IYiJUEOwIJzungKFMQ6rERjd9QCRWUkg6Kt+ZrCm0pgF0FEXvPw4ARw6H6VM1XWGJoeSR0LzlVBRxLucSAFa0Yja1OmoB2SJcfLmhB74dodx9WwtyRQWmu0dyZeajQivNggUEQu23TRhkBfIUmAyrSyJRL9Jlz/slu3PegfLSrSjp03VM+yksEGh93+gjST9B/k6Z5K51MIhZ6NwkoasKZMhu9S7VnPo0AiQmT38krusFfOlNdk5wsrHBCmzWHa7Ptm9IpgBFA5TNHRhqjZ/8GHisG2oq3w5mDaptXFsnkLNKxYIr134h6iepgten9FI067iWYBzcxQuZkKCBZqUN3U38595ikOkWyT4jYY/KRuoHXMj2PPuy4stTUpJWUHfYnAxlCIrsFwqCdUtG8HIS9mlsfHoUCUEOnEJ5LFgPYP2n78TNNZFYNnbVNaHOvLlYFaGCXst4K/3M/B5ZdxLeuFu/SlkQloznSBbDHKeb83WvrlBsbDK4MbJB/5RK3W41ySWDuwzvvakXYroia6NM4dRu40A01HVe1mdaEr7UXjgECQU1KWlO6U8H3m2V/ErjBdfOQQbuJzWsrICXWYAE5sKSuIeklEeBeb6yc/qE1rG+wrJ8JL9F+cgyamezBz/Cx5cFRuzcIUvKTnsaCEP35x2ylTHy+styP/WGblT0PO58j/bgYv590niFg9M/w9zfQUzLKlKrvSus8dDfQzK1kSQinGcpeyMcYsw9ydgfXj+X0wjvQMroagWTM2QpSPk5pw/o7pKnT4ofCh/LHLQbBDs1nfjvzTvZ547V0Hmfv6eV/Xf94BvkmvQ+9M6XpRyTXZGYnlpZQgjnK4siJG+Akt3DgW73DnD6gQ/qocxSTJtYMtJJ6oX2ZFAtXDMrt8O/Q73wLj5YzaEWgCJoP65UU3MASZX11zSkkL/exuyXIjpNuGSygeguD4o7o/QHARXtnCwT3NXl3RoGNiCUmOj23fbcPP7+jAu3yXxsr9CCFwAXYWeEkvFSkBiqebgizIkk67FbyMo8ncgqn3Fo2MXmzDoxomPzmW+lBW45g1mQeJF6+kapNaNbtCJWQVtdbuGlDzuWQvA+Im/IOAWN+Zj+E70lCTwgl1tA6P1QqIHjZyEtmBLCs3EjjsDu8MTkp/8Biv0Yv9TqdrDTGa/3cbvR6uq0SvrZEucKv4WsxnKAJztOr4XUKj3kYcWbRxj2l8oxejkZAmJii14D3yiU5C85Sd7oOaVPaNlFT+C4swN0WlPzx+/QCB4GPZY9oTYZ+2vu/6/4Fe4uQAuFXPAA1d8leWULBjgV48uFVeZz4QTGsfULx/k9nyzxYUXD4HwLMrrHrwEPQTQAwN6AAt+TUu/ZbUh0D5sgrqpmSRBOnd5IOJ89nkUNWLLqVbWyXuvBXtzlZox6dbbJ31wSSjNQ3ZFH9WlafbgZwOUPQA+9ghN0VCyIarlo4N0dz/UOzT1v/0fkSFuX+iUnsQyV055HzbFC+JDte6JRSNexEC77+ENljPIywejKBQrpNgwQAhlntdZ+RFvZIUlmxUC47j1nAUghuC4y/xjY/uZtcJNT4FPDsS3J7CmaGtIGK92VpWeWKGqtb759D9T+7dx/8SgHlsadczD+8kL468+d0/eaW/F1bvo23edUsOdE9g7DAVoNkN18rgcdnsYDXTohggSjJKj/92cJeEHLCK8rKU9+fLbafpGZxgTLV6AbeaUOq8wGDhoAE+mNrWYpZ7RakR1/YxBPyQTs6++NNKD1xd+cU1DDUOcahXB52I2mg8UKfj+oxsgZv92RzqaFYYRarlETY5GIam+9FQ4KDFZLC6L2gxhD97jed4kXMszSNBoFGF9Pcq1CWhdYmuIq4SMUd+eYMs5cUMQwpF+FViphbhr28GAgOQf0aqrSrwKlfAq7PhYM/JJPk4QNIpDSPysn8bY/2kGSaRHApYAyunxotW8jnuVILEZUJKxkBN2YRuPGRQlR7MHNtvileRBmIaZlVdHJWcjPgU5DzyaSr05e7JYbHEvvC9gDh4s752J+u1Lfw7jQpjFTR2sPFEaTigtYG7aqz2wSJAJDknE2+QztYrTD5cha8ci02aNmVBk8m5p7Q6M5Eu3J1NZH4f1FFHqCGWWcB7NOxSjdZ1DIPXwQHi4R2CPSapUIZeT4lP0Qm5SfVP+qihuLlRrtqWvMHBtyNqQqtK0u2CTs3pR1BduoUFZvmHczpc11HAqAdZ1VoCS4a+/qkgczXx45aZigTbkUnDZB9wDA6B5REMQK8/8s532axRU6sB15+ULXxgxe3o9Fa+mSrfOQv9VarQr5I3R8QeBotLVndTh2WFDDVKXx+JIRQDVFVEf9C8b2ZQ5T/PyGTfi3Od2bRM0OJ8wrGUFt6lCH7E3D6evzcpmoDrLBPqKFnTnJHpSO94l7tR/VuYFbZA0J60YTA8x1HPaO8Ik3awVmH6UIEVJ0Ximz4Z0qL4pRKqjbyXUmJZpwFy348U2GhBrXRkG81Uy/sutX7e8MbkBZ3ccqMpvFP4tK3C/CWBF3RFLWvLEOY0VzBfx7fZVdGCG1u9MCm0spcPtiBXP62nDtA2Pvp519lPvv4t18jovVEQYJKS246zRCPasIB7czLlmF1TgsJEX8Qp1Uy+H3HLYlxIuo7zMValOJWhqglUnq4VDs4aasGRBi/mbiOiQF/gZDQ0o1jxIXmOgyHqZ+qYblZcYdL2KLR42l+R+Xb5MyxobqgNLHieZhFDh9OZ+Ntc7zCFw0XISgDyyGuoTRqxnxfz9zJYIMQ1jw2/KgfHGF2VkP3k48OQrBEPK2G/x+Yzftuksx2FtYF2w6gboeF1hgHY+DIXabPvAesqQ4K3dgSfQlhvQA7H6YdYe0iDJyd/dUmIF8JbozDVkizDnNgCFmvB1beNwyJjuikVcli8UMlqjYAsu3+xwJ1CtxAwEvW+u85zkJPNjNwPVvwy4tNZ4bDH25C5g0ACu1hN0sY2N7fWwE5gvzdQ0FXyAYh7TXhyUpMOR9okCFJBKwrf4YNdworw4FbUh5mMf7AkQbfiZ2eGmSnyLnIs5RrAjJGhJjt4lIndHEDxu5liehPLse/aLiBMgXLNHDySg67wzl40U1NjflvFPthSKwUB9NqwzsG6e7ecHZrOVIDasVcyHYPb4mf3jqp8QtzTEXwlWJIgAdHSqnapuuG17aK4N8m15NBSIheUGo/ARF8zj/0wLHd13tYQf79zbwf8iBXlJXWtuxNSBFgNUv+EvApPX7ZQpV4aaHfnlt0WQwrQMviAkEVWHfVy4lVHX7OSOfqJu6dKBeHE9PoXZrgA0VtwofFv+cYxq/jucYhu17T5cWGqvMiboZ/FDjBtFK1Bwg0zGQeDLT+Ce2XLMNEDvOWbjBv6RS/d9Us5olDOM020meO51LKZgP1yyqANvR+1ZN/79Y5aczbE5ttmkmsjNWD7CxLYIZl0w2JOSgYj/CUH9uGyh0xHxE0+k82x+rjmZzK6Vo3wNG3pEmc+Vu7AGpuApIoSw3pY51c4LVjsvYQFk8rIx9JIPywU/n0kIz8lEtjt98FvRCKHJ8Du2eSCCpQ/j9lu6tpo4bww2rbi9hVVcZ5cySfib3ADPOQ/p3NYdBpJNBAJfWBI1WiQQl8BdM/47FecxI4INQJAwh03mnjK+xCQQ0pb/B9C8ZYBMFvjrUCAp1b0/E6SLNWGVeX2QIPCloCW0Nf6hss2+gcPqf0UbRGGuLG2giuMW3XEV8HQBp9R/W/F4KjrML+M6kun8WTnbAogqfYqjz+wlhEgUUVtJOh9aYunSFZSXOUZEZBwPDh3n/iMAtGDlFs5pmgHe064Xi+KWxdmkqqyan/p9nrPJmcK3XjJGMlmXWERtkgHk9QV39sZzjMadNpofUfv4dAs+mzhY9df+/J0c50/tQHxpXlgHJ3K1OsmElsHBpEo8cKe2BFNeeWCcWtuiQ9RaI6dGs4yP5uB7p7Dr2NW6bwg0oEWQKofiN5iGNTh65REsqB4xfy4BeBoKQcQAveUmRyn85co/WzwdMsQwR4XFiubgWItF8Wl7PTnp10bshAeNq8yxjeFuhnpTZ+Indj1lr4HeNH8DvI60OuozrxJoxwiiUWfWrSf6wrqY3JvfoKmzytLxY/IY4J/kO2siYpcp1CrLtBke4mF0gnyeBLa8srZvK1Ym7jfs/a55Pe+iFhSe7h7qhheqd7GjKw1rcRYI2ilV9Xrvw60TjS0wNLjxne5wot5fTv+NYryI8p5jrW9SiRjM6QOPYZ3tudInwz+1uGzPIvFlD2TDLky2m8ckWkBDJO2og8Rp7KyuGRjQdcguGSbliGw42oD7dHSlolpVo4W3My/NhXgvtdGI8SV1zsZTP2BeJDVtvIvgTQmGoAyywbrbkJyg2wrbFiphapVkVHVE6Igj8yWO3TDK0nGSTlM8M0KK5Z9StSO+lusQLpls/kodhyXnkEY4uhw0TwU2nu+7z08PCf1Q1g8kqau7fuS7Ocv4dOXXYf0R40eGCMdwUQgOkFhOShPNvRS2xr7ywO2ToI6oy23MXoHC3kR3gLJc6zvR6rNoV+/vCtUGDqirGHepmIq2fEkiPHf7elK4p0GPpeTuFpnteVyFzRLU3StscxMaS/TLbNWs+xEbeWVvIp5Kn/F53jpeURK460+Jq9oBM4cN2fC4jES9tYE6shAUv2v1vc/slNtVFdyg4tsbsgAtu8qdTisBkc6OIzy2NJMNcvBg8AmszIS3hKhWQdfXV5YjVCkq0qQVTdN7rGD034E1uaVjniLBRlzegfyToKqvel69MNTkLxpWTGePJq9h4+SUS08zM/xc6kwl/tm0S+2ydCOqmYfGWbLl0yCVxYbx5l0BkSqxTWVAHNVRghkd/BQ5c3ciDeOWb+/xw/vbaPVaSkbd1a9RG0kC6yxk9Lalr0x5IME9sj+UuEf0gc/1Y50KkhpBoskyvMnk/DCtDfZgXea3jRGfOkvnYOxq5f3yZ7Iy523iO+1emO7bBLCh8Jvk3LKea0DpWQIm0xDKrtHtyopKObAdp5BydlWwcZ0V49YgO/Pj2mOyAWoicsxPCq+wr5E7eJs3iSGNiPMtKP+pfE6KG3f56MOR0KslkLpZet/AdxwpjgFe7/HfkX5WG9W71x1b7o2idGzFoXO6Rf+adOp73KH/FOmTiauxlh59sa0j9e7rIWBMeY38fmC1zZFANWIYneewC8+prwQhb1qxZas6i60xeaDH5hXr/o9LOTIaHjYOawEtT1Wdd7YLQma0no5ADfOpuVVPPLpSArR9EswggfnAM2BgGmD9z3Hb+om+jedegxH0IVm3oZ2sDTeLaYy+UJmQPNHeN4UTBVp5tOuVdtJMkip0eFD4rSYJslbAcKPiU8nQD1TKVNzQKKXMcKz3fZ7rOzVmrMbE5i96cczuEvUXuiNAKhOgFpdLY+hI7tRQ207ARaTxxKMEMwImMMuwee2mcC7kOwRh+BEy1fDqzwmwhUrRWLenUYE1oO1JzeyhuW/o3V3HqztNtljWyNsenQaCw5JZxRC9NRttoYsNgBSPRrJHpm8nG8lwma56qz6LCkd6r5tfZeArgiU1AoCZgGgCdZQdO84YgbNVO6w9GF0rRqOeVTMEATAuDlIv9hTdGd3cPKErtOrop555wuGAOMV76iwwimETTwMgphLvjpev8J5vsx3nQjtb0Znmur6J2il1F1JAAdVajCH23kNKCP1QDkq7GDQu7dhvdxbtLehC0QvXdfE7PLb0Ru1zosWRy/w58T//rPNlnEFJqWQgBKhIKnuhhhkoYYQCuMEX+NRhYfU55AZGCXHvNDc7o9ZzexjL4ksAmnJ40oOtdaL4OB2/riEHPXaLRAuWxj+HjRu8qMQ/QiDpDx7BVQ/BFMs5yrmMwxr4Z0elQxopKee3Lsh+pGS8VZL9bbkKshOvCyuRJedHFd4So4YOXg7MDyxl/vw2O/G2lPJdVk5tp4mwpUU3AbYd0s2qsC9ASxareQ8ZBXwj4ICmgGQ3rDexUDlRgJ8OKPRDLamAWi3NpzhQx0s7orMsNtKk+jaNdTFOMYfdhB/dLa5gIbDa3Huhkm/ZNkkUaVpx731vqVg6G0TA6a7bn1SfYO11uqaDWtRAoPQ/DTdfvjod0Ro/eVnZliSReAcXhbOkmZfxoWb+rPuLtu6X6gc0pr+nfTKDmc51PhY1P1mjAFal61g+MpsXWOeeNBaNCq1/bgZfgYqmdcu5wF3LC24NNppso0G+2p5gTmG3WRaEMuk0uBWu5rlyz1OBS3b9T2qhbnzA/vv55mG6UsNvLtdCvmvXyvI3xk88lKDtEM+Mz7u9AtEtIytfKLqVxeJcvjMSZ0gaY5zQrJXgtyYejofoAmOnkZ72ZpJY9w5NYvhBWgz9ZiDTqgrgmjK0eDDD2OmgrJt50g4iDRS4Y5OVZdANS5N+aY9lUKgDl7skc0V//pTXskWcfjeGhUNbQhd7Hu6WspwEiNm+OEAGRl7buIYW23oa3b4YCTddnctm9TimetMf6nbHSTVWu7w+GU0+u7P7UP0VVQViwZJZtbAjGEBbtMsJzvsBeSzWKaiq8jUtFt3f3q6xwwcObKRB7BRUtGkbQoWd0QyiPKPt9VfljFK4ZIh2mEUnBc4Oea0n8CYW7kLZuIKrv1iQ56bcoN6Vy/7X2TqzR9LJMJ6in3razF+2M5/34bbF30pWerVR6A0/F+OLmQ9zLlHxqc1GIz4kKYvYFbMwXOTL97E0GJFg0RGk4fMdTdOGUQ/+V2Fptz3y4llnAFIr8NsnDJS7LfqvIv1suSZozp54BGhf5EYwCk/AnKKQxuKoqhLb7qdpGlVZcHMbLE42cXwlqXtVm2m3OcDQaigY6tvHkF55ZEXCJmT1XE+rA02g+xko8bRWEzC+kLWg/ws4tNFToVFmh6Sq61ZV/6EsTZsCXoK7FjEH4sZmIIqv+hJ5Z74gBSKbAKRXcem4FgQnJyIqlJ4x1Ljnsna+hVuQf3UFiXdGe5Ohvf9T8+yMUmFJfPq4dFK+B5ecI5KmZh365pE+hWh36WLPlWTvjKI4x46SsKNRxzwWpTHJafye8rrc9FA9ARNwxd31HOydXkPD/8ti+TEnm2R1fUsz8CaJWTQZHCKLZnSFx1eRIQcxiPN+ofQocon4896erout2VBg6CBRrS+FFxtCeRMjeb3rNVRfDaWeyZaw8Q/vYktXG1bBz18b2eAsGwhBJ3JaY58cl0yCGuXTHONI2iwmYY7e2odoGNpaLENGzwacpaUKFg2oi2qITeu3JX3Zdj26ajock5jxx8jdbXLnVTEAMPnbdsB4GwPdZpnUFVfWaHc6Cbxx38N4gDx//XAIC/5DTI1Y5GjHrIinb0HppoLaVF8/6ne4DQWKmsQibAQkrJJSq8Hk8nYJUc62M9VMubjtHuJOst36Wi/loZn4CoTw3hZeeg0LAcnNf8WkxZf+08DrMj8/hMQRBqgrbflG6L8Fin9iExHKOKBazzWiUUVfLMvNu1thxl6YvzSYdlt7nTykoafb7LOrho+j4AVm3Gnmpm4SjfRsvd6IEXcOJ43binQh7NHB+cGhk9Vh4pODmNYux05GjP350J5VVgR9MCQEO31HlIObLzyY1PBMsB6b0xg0lSQoW5rWOkE77xPVmWvoAJyN7UoQabNNL+N/5+hL6VFRf8IphtOh4kN74MMkWn4N+LU7LamwGv3DoukL3tXso0gbjMccNHd6UlDeLSRrgQLadlVytk60bjxfUnR3aglgVzyCzl79evBRCIvnm4EPsbAm+gEUeB7o67BJYwfuCI+lKNBBhQaOJuoZpTscpZV71DU7K32ooCM8O43vldDk/Uq0h+Pg78ghve5DMlr85tNIQhRp0iaRxjqGcaGWgBg7WAAZJMncPwNYBAwDgklll02MXT89fvzXNHNTSLLJyqsPgPAnjNRCKlMrX+NzQaZ7tuQyPHG1ixHG2EPlR1wes1339xZmiw0ydPRGaHSdA5vsd1JCftijV/GkAgnOpyC1qoJrjLe3/3Ileq0foPtcCWsbrr9tzgj+edZdHSfGU3GiUdR6Z7bUQTyuGLVL7xmw+PBYwnOSJo4I8DDJd8JWA8xW1osmvMRwuKNOTdyi3zlPllJJ0WPwpSGcbokkfVbaDCEttI0Vnt472f/N6N//j4tZ7U1OCyPHg2HoU42HmRrbqDjOnA4WNrAiaeZ0sjG6GkmX+8jpQWXE190wQucu17iGzX1zFrRNRq3M6QAXZ3b3jBQ1KPh4KbeeVw4FMUZGMKimrtNg1DniERlNrJLD+8qAagy6ILAsAifKpBGZ8xin+Nb1w+Q0MVAzYUlp4msH81MJwoxh/n/59Pg5MtGITOVvZUJaWsmCuV3rVUezGIJmhNSw7i6yxO7CouK1T9NfgvkWTPRoSrfy9+E7zYsD6yMFk0KeB7jSL77cJz4sKwq8aQYyxo06JirHAujOfD41eSml9PNt9FEdlRFw92zBbmC1JxrAsAEzaxBh2/4ZHpbSqsk34ZFdm/jIBtSx79ujf8ef4rWFt4rvQJ1AuZhxrQRnjxQv7BjG09lAL0u95M3QkzpIZQcbQQDRrZRfqFWV1jlVrO3Vg0sa/QxwPnf3EcIPML2RKHRzToflL3CIJXIxFaV/YZ6dcsF8X9ft/HrowubcZQ/HTjKUwniwH8GJN6zy3Nv+FqEgDUVW3yVN+UZZuyWhecY310OCAK7BMnhszOYbIOSFlAeelgFPMowoX7+QufpTQ5X4QD2UvnvybY9RdzFirN46Qqkl0IvNb+0zU610OkeNHOWwaOxaF4J2nq9BdUxb69oTwot8A9yEup9ZKML6Hsyf76+aom3UPCznEhE6ZcVbzA4kDUnYoOxti6DPF2VCnh1faKnx4MvvlyaD0GN3lMh0tfQHChjSPVHooVv9ze4FysSG7/6nv0L+//YpUjrQn2oIwsRDeQcIqbxMdH20eec1fGAIDjTNG+a8bxKkWG8biQYIUF1Cd2hgNzy63ZZFVxa4HHwfjnwsFGZXEVhZUm0/eBtYEh0q2TYSxAQd802ZSs+ixJ2mYI2Bh/RZu/iO6lyVJRLCjuiCYYHR23m8tbIN3nvKiJBLhCggBnRFI1up/jCH7jh9peHW/2d7yyy00GaIu0j329GZ3mMC5EDy7P7vdLyrgicsDw5OStUUgNZnmXZEbwc4NyUWzNt4o1iDQSsUwCDHWbQL846yCC17pBd5zJQC7kgnBhxOmFCO6IHwxrBh5a+3x4C0e90G2lrpqMPTsK+Fwp+ICT8OcGPb9NYG7+svH0PYZaoGkYbpfShMmrGYWLvsGTf4nEXAOmOPxb0BtwGSVfzOBddxrK5821DyuIgtLfw+z2ZHILFhclAXkTxmk7gxAb10k65qOYMdLGkkFdjjwUeK8zUtoSxXnx3QhqShJh03F00ltOseZ4h08u2WBT7yNzhmthNrZt31Ej0tq9FWp+6zVeANeyCh4rmqjbQe3G6ZaKWoI1M18b1cx8rmkz3ut1T2a73lSVkMQNWa4160/wiTLP1dQGVI5WvjZqJT7z7385pmp+y9r9XQQK2EuwPU57IIDSWPn8cQWJ3U3YPK52o/q9atqwuv+8WGGbYPrBMJPbarKTrjgOysmd4PdsDI9/k5+vIvryUVncb7dUk0r9wxQ5ik4AHWePiaerR3rkgPRxDkYcTeE1O84fiG3W/qwstL01fComKDLRnmfnCKMOn22PyfJ2qWsUz33tEBSl8TBDiDLaXL3GAe4iR0Ym9QUi4Bnw5Py/NljuXUGlwS50LInpFsMv+lxVFOguE0nPjFqCOBgmjp7bZq2bJsYNAH3mnOOndBRBTgN4nYAA+hTVZ5E8g9FLPsMotXWuzQPMZbJJUjOPtkuGm4IcwkXWDxohZ6KUlDJo6XwGCMGua1knGS3a+laBY5OprrF+pJSjPnS56vjMo+iJVBZaYc1POTkP+Zrc7ZMHv27giNtmgcwRiZzyDuMPhN41SPAMUhRLLrS9PLdEOaJ11vosDTc6YhSo3BjlvY1uujEgx+10KqgWtX/BQjTCL7BwKlUzm56iRCFHVH4u5MyqYu9q1rfbH1ufNj18fw85apH/5SvbZb5B57PlAojZw/pY3qAFS1vrvdMP8pi8ZSLbzcx+YYnVpAlJE4Z4jl5THrKC9ZMFwAP+6p48zzrVvqJ1jLqFH2haMgVAn0Uxzk8MjZvgsXPiF65vm4+aiEJJgrWB8TD6KuGiqfIX2gnko543kRWXj2TMdkHEGnfW6vu34kt1+RFOWi0Yv05+YR72ZaDt1crZstVVULTRwQ3lWG1lgm+LwfN95rPSnU4Nx4crCeSEZuusCEbRYumTlydvY+BtaMoEuFUsZVuAfjQT7zzNkS3bPbbF4em8qc/A80B/XieUFmT3yxRhJX10SfSAx6NAXmKgj8iHhZEOhk5xrVjogXVkf2UZ0ToiRSBM4G6Pog5p3lfBpI1bP+qa41j4JZ/ec+UEcJHrdJzaPnsB2r2b9DCE877BojHkwTA6TcvzpRTECuqWIyxFmbeLeDI1+r/QmrRk8eYwsXF1Rc5WPlenWlVPyRbJMaeWZIHf6QscSM5rF2zcsqg6abcfDnuftSidfe+Ln/S3Ftu2M4XXLitDkFKK/Na+I7kNYfWwgAkDPYyQAqrUrZ5OO/Lvo6EJJzm8JYW7Hv7dyXoBf2X7Chr0hKBCQSvxpbcnf8gxBbtfIlvb9k5NDnPy7L8kPsNybnfsomb7zOxjXiMo0OYjMgQbbKghubhvXlksi1egcnO0PPWrBEXcV4QzvhGAV9BVAusA94Ccc053Z4z7k8lcRbEI6pLY1MYiSVfLfy11dMplvytH8kUaPeDEyLVzeerNgVfjfTabBCeqZjnBRAx2MRNQDTQr6bHfK3+xE83Snk3X32z9Qgws1JNtc4WDHS/fEU2QQ9G+JVXYwLU8VVNL8TEz4cVYHFfS2MlsRq46VVpD5ecpMeLD8JghZNHxm1NDC4bgII5gKjCWUl4lebYCY29O6H0O53ZGZmCxniBMrop4W28I3xQ6eEH587oHCusKASboak5lw4chEv6yyc1tkI9ysULiNjeCWcrXcNuaNjnpmGvQQdSGSINMQ2LcV3OZ9Otx/UBb86LoOCiKMzWrvJHGz4OhJIUt1WaVS5CHwlxeTu4lcXqL+f1tGAeMfaLntInrw9ff2f3CxBUQmT+9VGmus4VV2JJEHnCE3kDv/CCfHoTEMAPXpe6JfjugDuDgAiPrdb2rJunCMGsdZ2hF2aI1FfD3omIqEAhJSgLRYsOqhTtaZHHw6cAQslPq14+dJvRfXtPJE1BKzw6PRprbDI8kzYjRpgpt0ahSpDhImerAN8BVG2sIMybujhl7tYZdwGcHOBchLm7m6Eog8bu5ATsNfqLxddUDCqEIOa3YJpQNYqrqT6/JlnQPlIH/TADOWDedY4X0TMYmCWIXvunnyyu7nxTqGiXClRU1CoB1yhO48MtIqhai1+hhG1rz585lkYaS6gD+R+bqfFVKs8q4VjtE6wzZ7YjZoHMb9rubUqjyaNXwTEEhJ6zXaW6S36o43fUHnHkL4T4u1HCEK/bTGa0bPwH4rrNLsLUa6sn6XaIn5Wquln5D/aXHt5UbKFc8dDlOdz2Jhp/J1R4X4ln4V3mhoUwDjKbaVgHRNhnanaqu/lEIwz19ffP67aIoSPRUsNNttXS6JIgdKFwRm/MueGAMWYeXNgaovhZOIKo4JnKGr0EbFqeWCuAo2kkyN39C8VglAlvq5phHIOXuyX38yVySKhLDlKgbL4lDZCG3bQR431/vadfSF9NEBFZCvWKzXkcDriUmm8GpSDpZyB6XEX0yckkw9/msCgkOu3oVfl746meh/jRz+WvGoXkxDpuV+A2p+nAVl5+w4JJSL9ZjQo2Dn/Wmz5llkGZvTBWZQvRUxvEi0ImN0W286eFCniday+G9sY0nxHMaqnDK18lkSD4nUDE8qi/J/A4yxO2RGQbqODOqldnDSRBeJphkaK4XJtNEONzxKuls+RcvYi+dPm/ujDzidOcDcnJVr6f8VwBLPUUOXnM1NiUW3PHtR8U0TFrHqskJlVs61dJNYepcgcGkoOgchU4OAWBv1eip6OsuoBi9gEGVuVIU/NUr4SI8tb8SIMoCrSC1BPQP/PURnIt2QZrnifuBiNRlC08DaUZpYSdpNOBX7b1wLANHg33ZFs7j+PIlXAOecpQNPcq37uA2tP5Vwg/J7y5Wo4nnPlD5p+wvy2yMk3oxJdeAaYTgFaFbPtXHQg0mu0KD72cdiQoYRQNC/QPZUrnhlsLn/1hcS5BQKJOzbelpsk2PV3+M+hsw6syxeQ4lnF3XR56lOcSXjf36PHVNs8iY7xVr4wqI2BHVFGG7z7sZPNvu6F4OKP0ScfbyyWcFdgy50yDxGsD7LpTqIyLVd00Nd3nePrZTIuQeRTaYiBIzfUDzUHpSDGlQ42jybRd981FrXOHnJ1ph+YZZCyfCycxbCnbj9EZX8rIw8sKHVnE1OkebBekaddulWwQCi/9q53SEytJFgiyEUaUhUAwJtyUw2oqK12xLdD2RcXecaNm8POsuExrvgMc3MRauq2oUDTOAjv9pLKypukU7hrgZmZPCj684OhxJpqz/w9f16GqaEe8gyxFQEo2WH+kxcpxbR5naDGkRkA2kFiR7NBP+70VqxBs2OLyhCp5CHdTjafyZZVHMX+fcM3euSS2BpoEqOg8PTj4E/FeuBK22Qw35dXhuz4u0VDfVxIo+NWyPbJpDYIsG1KrhFdZQFoh6yrNoA/+YnJ1gSBjQi43ToGn34klBQaFza6197Xw2+QpYy0/dph4m4f/PgrBImUbOg64F/PHAFAlpMvZG2lr4ryw39DYc1HX1LYOpI6XgWLZTCT1OaoAOwDJQu3+XtoKdDSr60V0ml+RaSjvDp75KFgHPyEAAjvXGkRHW7io2bC+W83q86NKqGmgbfV3cTSI6v8cO5rOdbCiK3LOGkfIHWT2m23AirdsXysain4jppz+YRX+pasDT3LF7J3Ik7hsZjmjJoGbqIR1R/PGMufmEvALNlqcLaoNqq1dNToso/49KC/WoH97Mo54RMpTx8VSzc/evY+jJtt2S05889dOIHKksP4st9WVSm/linhMfJy8g27FrxrlBGYxdheDNw/KV3SJfEMJAhbi8vsnMW8JMj7NMIkWtqOjBqURjO9M2WmdEVwjjxE0VX1Ete10w+xPLJzfKBfd7sjQM5dQ2b7kM8GZ0NOQmduwVQ6wR682wLeFz6NXgiNW09FxxYuyOiJhM/IAqrtYVRk7qkJsmJZdsdNPJ9Zk8yxXUv2Xznmwo7PV3+rPBz/Ou3puPHrK+dYf/Pncu69ilUrWrA7RJELTqkw8+Gh5doLZITAAiah/MxTQipglae7H8+3KTeSfkbd88KdBOtgGWrMlfTEY8+P78oU3rU2jjHV6proQDL9AmA2nT3pSU5Al1IKaC/8IlXtSwylACLf48/knfqbVuHx25SfsIR0nBiIHUOsJZs+iaIG522KEdvCd0L8dJyoF/N+6rfqaE4XcUXekOLnf96nAb+eyRsjXmunwWZShx8Egn+V0IqiRxp69SGH1g5F+zOQBwU5GIJORbUtU2jZ0h+uX9ynVSMyeKjbQoQZRPkQZ9DpxnFCw5Hm7ITKgpKeP9/a3/jy17VmX8xAF1eJkaMttJZNq9rn16ZrAPCtAYisfM5YuVypmx7W5gMNWHbEPv84TEkE7PNFO4dk4OOB2N+OWT0AKPmRvFrc2RYDqNZQwbAKBRR1h7K445xfkOiQlwGVEhM1DVsA+szshu+0yGies/91t/sWcFrCVXU3KmVUpG8dF3/G66NACCtgFFCC9rwrKpfOjMljFirKU4MmX95PHyYJl7c8EFUgkDLojiKr7lAChn69YmasO47aAjfnXxYJOuYj4+rCvK51wWZ9iMQUALBOAUPU+MdNiIMqVe90g87og2P8O+2dNvcvOWqmIF2k1aUpGnyrgrWRsmC3eqJhC8bflgP5T1GCupv1KJmg02Vh6YGzFNNX7iZWx4765410zHM0dPevQXLUOuqGVp7Y6B+Xa2aTTyzXlOyENCXLAPmYzJ4fzSvWF8f3aYZO3UbH5LfTdRGjqlQzZ+krT/VL8oOKV0b/VfVe2P/vcJCoNb+3Kdrv85Ly5JlPKrZPhlqO9v50t1sdB2NU/kdCEQ+9z3OAH9WRreTwyYFxP5yWDJZZNpwprh6nvrW9FaNqo7gEhUhNU9PzNFnu2dtxG/NwmoPs66yDbTIbUlMykQ4/QbFOs+7GVr4Z1aOArAs930D1IsWSxy8s3/LNZaZY1UDxF0wuzeUYTD+6301L86ozp4C6WBvSWCpffF9LUAA1tpbf7ybGQOnFRdkmehglRMriU5XhWuJO3e2JhVA+cFckfUC0XukXLMc9ehJwM1apltb5YEfMEibEHIFCzMrLNa7ozLHFMyKN+XsD2sf9yeCeoo3xXV4mvCsWiDRAuS8vgT5PPUowUsn/vBHafzx5614ihnGzzC7vuesmbmk6g1W7gEhGJsMJABPvbKxGxJhnxv5DgoklMhLXaeiHwlIDyKjOYH1A4TVDLrCLQl+Uv6yXasNoWIVGLC3A04WHdmaPwu91RTUy7L80NfQ/xT4bnCUedkchYhDRRFFxXM+N5Sme0ToJmnxsCJyqzbX4d9dR6wdk1Wi6O7Jfv5vLFqcj7B1jxoMy/RGTjgNeARVlyhs0BDX9eO26/JZdQh87075mQJK0wp5cBLeJRTIK5NE0Af5QdqutiwxW/VJ6g5afzPC41t2IJe3YvhfnYcXzQjY9kPlMQAcj1sPTzw/e/vjpg0ic6lDl4dDbXojplOKXsm0KOi4MDhRvRPhitYJIi6uGBSM/vckQ7KzpoKZxRCwZPG1IGcOszvMvGPMpkC3JPQb+RF6I+q8P8i9ZssC3ZQcLtw+sSKaRO+4xhXSQdqt5yw9hovFfjEdbhXpVwaqQ29YgUr1jVuTSQYg4qwvLazyC2B38VskXXHIqJDsE/GPU1CaQQafDsFdfnTxqQ1kTvWvN/R2H3RDZCeLhZJ0tEcTQFrymsTAXnmMK41hlZ+QTeHrmBVF0QELT/S+jK+q6HYpzEZpq/WSvqyNI3EijmVH7j5Ii9TQQbhFc5OlIkKZIvDTLgEJH1L+Zi7oj+x+5R0UMrADaOtFGb43u1husunXuE/Dm8IMxYhVBB/VbMlXVfFtnH4CZLXUwZ+YcNvXhzNfkcswEsejrdff/wLhgJUZltieVYqH19fNSewv70Zsr51tjZju9AK3vgmatBPUqWyV/FeHGeFxVf/5n7e9yAIrCnK5YzLdcVPe5cFLuNyL87OEHi8tkPDqnNZOZFDEp63rXrntQFIDAB2yvHLXz0r1mycC6SuvYsULNKOmqzbmrKu36WU5Blr4C0RX68+gi+4wt7YcaYFe7Lyrfdd4aWrWoWJDKksfO5l2+W1kykaE9AH6WUdeEVGPKkWixG+CMtI/Ne2yCv8SGNZjJTyxqHlNmNLy8HmKOOK9TzMjkykdYLh4z0ez+YBXNQUIRxKBnZ3TfqzGXHT4p0HnqL8W4EUVwlE+NLY0giz2McKnxRTFDcyEgfRJj9xZyfVvMBS3aBWtk9Y17ybApinWTE1ewTFAHozS5d8bTflGSSUZOfZvJ1/2ltVP8yf6bATQJPVGFyJRjzANKLyI587M7ic7vwQm8rBGasdRsicPtFrsRslX+ikz7HmsUnytuPo/tCSTeY1fX/4ZXK3aRzjOyDSAKddSnT+eEUAnDmdo6n0QPYqetuAiUT5Xf7XvuITKettYJuLabbOnq2TxHHIBBqL0zH6p3Oep+6WzIju3o4WufylWm7ZtpMLScAnPNj7/pfbDOfA9JQzjMdssyHcLYK1AeGq19sSsdR5lJrf+VjRew5NFaxMF7pEySSavN/JV4Ny3isq1is+Pw8Fv0lf1/GkGqoIGhk58NMLKkLsTbE8nxlXCrR8VvbwHoVZ6tOUcur7+5WqYLOFRMNanDPMyA6zrPewQWXEyOFezYHZ8GLQRBBq40Xt2cnnOoF2MhqzD1mPTeThO6vMBhHvYulEt/Ij4ColACxwOng7DrwT6EZub7B1+S4VgZfdA6cXuOswftDCZwpwDK28B2sFWeZG660TekTgRRzyH/qoV7Fy0/Ons49axtt56MCN/fkwQ1KXMF1ga3Ua8RANZvMjmUviecdCEIJj9IBhIZCxYlmpEfe8Tkcs2f/Yd7nwuT3IGd24zaszxKK/DniT6Us/7YFYLkFQLmGkqpj34mJwA9GhOnxiaY/ggINuWwYlUhao7lV6Llj3hTeMcfK8vtHDtFa7yEnTN5dcvipOXN/QBMCZmRwe+0veFqL0az34DrDX6OyawCwEr5Zs0z01ykuw+e4eXLc0Y97TfuEsPOlmTHHPDxhJOWsDp8LBSbutDj+dyAmaqv7Q9UuwOoD3F3ht9IG6JRjc32zmH4LHgmGRM+5WKGz7bHinB8WiMGt0Iiks4o4THDo9oATI4FN2gDaSdmTrHsHnhOv3rCI16xYdeFfCdreY4ETpwEssYazkyrR+ytEyD2OLc8aM4kdf4xWgW39w/3crwqac5gKs9L7j7jQjOZSChdezUOa/VIHJbcfbvVPCracFHa4TzTsWahbGX09MlGxhKgpncUd4YuYZyDzIxqNq3RVIcQB1qd5/eAREbVXRVdc/KGMrx38vUAmFJD89ET89cl2Vps7SC4UUkoYgTFBp1JcQ4TYVv6nqCvP6/Gn4ZkC+V/WLPADRIoKr7thcMZbH8RdIoOUrgLLZ/HUcbcMzfnPrLCaj0tJU0qOOBKm6pjN20twQJowQuuVfs3wQd+syDcKADbdyNwNeS5bnQ4xoRdUrHvOCZlnZEGB+KMHYL33h9HqdEYqzx0wHVockWUM3smQ0b8O9SLIpBnYhZzThH+s1t8LXafgMk0TGI09kGORc+ZHuTnoaJMzPigyJngQhZ4TJ6Th3ElD5fogTW6iY6Yxv2dDO9DcHkFUcOofTfV11CS5Eb2spDWfsP/xwSh+sz8uCBRv3C7S0b4+Jd520wWmgJmUyEfZh+GKmDwofk6tq9NKn0QoITseXP0eUQqWAZ+99v3XJI8sEbZKlnmJZdqD84993JcFoLktWxRo+Stdfxn5B0WLC9EmITTPB3hfGcKLfYDisJPRJ7oQvVQJq8oM0HYPjP5qWBQVhJ/b6EDS10NvvwZ1OYwaumIspEMt7LclG2Vkj0I48qdluQSC+ZLhXoLBzTQI6dKpgtMX6nW2+3k4QEWE7WZ1e7EyIoNlHCEUmfDvBrRBi4/cTr2Myn6JINfRpv4GedU1GrnFdoaFWml/GiaZc/r7uKy41OLq+5QGXaoVKotBx+PBaZXaKgt9ksKZT8t9EA7Pvz9stu0/M1rrxbjJitCin7YR98OI+LRXib3l8yH6SZUVxj1fhvI9meISYBl+1nfnwTefQH+iTek50ZDJmpPNwtrAMv2EOFN6QZJt2vqABSLxFJPUIC+BPlBGIdiiTmGBsG3gVRhNEEsJH4FLFIFN9l3hkocj1OBOBq2o4TcAwmEVg+mvi9iy56u4zxKfdiqlSxlIaBqwdu+wSfjCYhlCF8opRLPmb/vNw75ZxTYtGNbmhHR0JMbWz+eVHXWMSY26580tZwdpPl0Gw6SYH42ZKCbp3I8PNnGvbeZMEIugOjMgEyioB18TDw2KcmU98XNjkmiCX23fsTUT2xrD1pfKjL5VNrZh8jW2N0arCLVwWL7UuLM0gbHrY0w5ObvKEapm12OYjJ3344ZxKB+72rYVMD1/5KQfibsntwRD5+b7XwvVDKaDdXRGUp3h6Szb57ugW5WnjZ+ib8xzNdRpeEM9PAlL/hyTJiHt0b2+MxtaCAFWHzkGwTVcw7pNSIa+FOiU0wePcMOGSyq9Wl/0DrL7P+neUyp6lJMQHehnFHXlbtMV54gVL98tLJ5SGI7cXyufm633OOZIFC2p6T/HwaZBFYk31UUKSL9ujDGt26f1O0KUTAWS97mnDdruXp8bRzHawE3dsb+I5dyas4cii/gmvfRb/y3KXN4WzmzsPcZpd/qbBL6Js5p3QbiR+KkZ9S24J9zShgzoItu8tE+JoqwJGnVDoNcwU7jLBiGjYJ9W74YMRc3QQvweTCEaMlukGZKH6QOtctSxrqIWuMYn2g1o0ityzvqiPj7/sEm5ljfNMlQRSUyQgCgv/qDQLKCpVedd9R7jZs32hkTqrhBwFB0ZPR6wzibjxfbbcMQ4kccjDS3OJrL+MZ80Gzg8l23shDbXTKOAi7SxkX5a5CnfeP0fW+x8yP0dvN7a8VTPdw8QFTKg9lOSoS0Y2hoLh7LHtARi1bv+wn1trCh8IDYQiDYyDiavQRL2erXfL2b/1kK18Qz13fjefInnbYMU3zZbyWWj9fZ2lRZvjOrmtUcmpGM/iMBizm3vH1I1c8yoKsE32z1SWkcgtofsi1y+CENf4f8AX95wE3JPS9ErvvUV8rUpNAgLALLOYg1DGAzsyXy2z/TzEZ62KcJQO/7o5LQHuiyOLingWFbfnZnQjPRkFDNjLFVyLxqg69qOgFtQzEeNzj67xpDUNxz3fsNg2ZByYuwLrLIuIP6vwYFxATI2IPVNEHpSa/RRjzLrcUEfqFpOZ5jgOjwJSmuD+jDi+KTM4U5JpgURDsu3RT9DQkO/F0tXJkjRIV4H983hSmyymuoS5CVhf9qNANzAtoXH2L+qXNiQnCn1+L6QQAhIGEtkabr+Z1frNwNx3Y6K/A/GAsz3n4kSQOnAnyOoNYeWPstPZLEWAK6TbJ7CRBI9hzKlmSWo02wswZ2OvI6hIRPRa6lfIEzb6rS95/VHaZWXkl5JV+rh3FDKc+oRyLQmrTqQHCsx48LhaOGzphQYh0WcEluprqvvWDr1+8ylfneXfoikU23iKFg9INSZB5V3EY/w49maVskHyikaw3T3C/JdJMOUo5lKvlOuQKcV7n413UeqTUF01XGyp8vQyjdPKAiujapJizc4uWL4He7j1ZNMiPaXVousdkYJs2xhyx2X/hi1j9VZYVtoSr5G5gM/ln5RvJISrtBRkpXpbmTT/rEzGHlyCjdi9bmLyu+mqWs4NdJmefY3SCbF0a5Yd096gUgPllUFU2VTYY8c2C0939VBgTavy4CSRoh82E6Xc0dP0JiPwmOrtOwua0xFu7FWghRrnF+Mvg79RKZLVRgS1ctywI3AgvnCXtaiVPemO+OaNcStVChBLn0T1ekChgg6oZuoTcTO0nn8EW/GCspLfriF7SZXTgYV5aOln/p5yiFLgIq4TeCZIwvrqBK/vlCnkdMupATT19ZL7H+wQg1fTCiWRgI7B5nZm0RjcaVKzSJn7B86LnkQ88pZTW0eDch4W7wQvNswApsZLVdh8cSx6A1tAK2N2ZgkKp3HGSgQKtBlPhG6iqwCLx1f/Wc69z3mGFsAuLiclJE2hOrp/mWDR0sMokU8qa4LsNCayNNGJopqGsSZNTUn4QdvFWxnDCSsFw7Qg4zIEI84AO0Jjs0rsPtH5dsl3zn5KlOX1Zew6BJZU4tCZ4SoMX1Xu1fP3y2scPqRPSfqGYPwGeJh1r6282Av6lvXmVd/6sWEDzCHBZd3JMJ5jT9ofVQtUWG5S2JRtmatxM/mG0SUX9ECYExmvokK8dWEFharhU7O1nRqdj/vhK+Bk7YwPYVgh4X0zXax0hFJkF77DaeZ9e+GSi28+nwYkIaIhcdtGmzd+SjKuEC55ndNshrECptWo7zpa6L+vy8gvqDVoYR6sgykQTHdMjaof+mK4PBcTg9cgtl1mli9DxzJWfI8r5t5nMPC0q3CuxrV2e7Vi4fpJP1ghipDsbdC+hkSQUnN1RBO9wLNwHpFxPx4ZtN+olkWsAPsOwIB3txmP5oM6KU9Ewydl4kxzrw8yvOIIQPdel1XJQ06jLjiiHevPVd9e6MdcYcby3e+2KcMZia/dLRwkodu8PVSAmvOngl/rr94sVryz5bvBnMNnXiyNL2DD5FZOxsBLhd5a7aSauR5fOR3CVCt7bLFBf6NGw7UDV4NYT54OrAL3W50kbVUuZVcbXup+2HOcrq0BcqkW/HiZMTp+yXPGhDV1zlqjhXG06Ng2cZ2h3SNxoaR7UPtBUBkZb3hczb6d4L6xQWXmnUV9WqW5T2TmB9+64tlwgwhlMGeVXrP0CSBOtkahc3JmdIw1IeVKKgK+7eiVeLtgH3iYmt3u2EtnR3GIdlWKuoFRyraexIUztEjb1vvZ21HCxqxhsAiXAvMdjQDkbTqRYsBz7rd0lfYsMXNVe9VhQqwurfIPYA6OmzF1vMaUumv9+sepii9rZdHyZjooXVnpvpu60Zawu4Cc5nP0Z32hexDll9L1mW07dfAcw3OtBO2dxg4cizF2OYvDWv2Bit+5yik4fggJNZzqD+JcbHTPWUbEhpr76O8ZPY4poK/V5gxK72DrARP0x6OBP18yNjyE+t7nnV2p+ZVM7r1cuI7R1O/q1QoPidaYkyI0aY9zr93GsianfI7q/CfIZ3A30E5/nRd0ksxfhUUT1EETD3ectxAvwBv3RbW5t5FqKZgbsJDVbyiVthPlvAArAi4WmdhYrT17L2aNqG3D7vrqhxisVxdKSkBs2I2Y4FwdYcHk2LYiIKWtEvjX0wjCxEBsrMgkf7GvBEdZc2CF3rKq5GQiNDO7NQ8bkZwmO8lUozd8xQjd/Qg7G+sRCJvoiKLDbnZXP7xp3JwNR6N2F6sF77AMTVz4y8rqBe57pZOi3kx5kpdj/OGa5acEbKF6RDrDKkalZzk2ZhGr2slY+zUJL5UDGOaq1FVFn9UOLqF1KBJ4SjauRHeKt/Ca/yi8RGJe/ckk0AkIfMLilu3aQisxlFOTzsKfPoE6KvQ3Zu64HJN92d0TN1dfLg+i14vXpdbKGjRFRWJhsD3MrkqFsQz4Zw6V2P8whS+EFTspvQt24OrJEhcRrYKAq6QdGUySXDLWy8K6e6Fu4fkWCpBkI8aULeiLB3/6wHVvwJ0NdoTC3BYTJmOsXnkPvDfnY0PWEtczgapb4y3zKI1mgT3BmAuu3kSY7fQruIcoKUhPTj28Zoe3226TDgG9nieYgY5LTNUX0Wk0oVEZEUOZ7HfU+A1/eZNv+piue6EEc3tguIUG0z3qfE5kee0m+lxGEB/CpTJO8wJrdFkJp5OVPD+A15Msd/BDo6VxjivZwa9AFqsApAdqhX6hOvF4LghQU0TCMp/XaoAfXVzb0irBRmZdpufB1VrzwGPlwlWJWXn3jt6ROjtfy56LKhB998MfBhaI7PzJhfYHeZfW5AxJ/E5csIFWH7AI39VmgkQ91ISYARGVob48vPhqTeESqcukFUyhklZfbYZUnqvQANYvPk0GXqEQFjqVQieYcr05IhdEcB0UQxkgs3iK9UWjXiR6yqEvhF3kKX17OM/DKkQsW4wQwNSaFDJX9+IpQvFne1snTb1f/EXUU48GmZGsBPVR/khViVjY0zlRmN856EjexfcjYFw2hQAzTxRLx4rarEp2C7ZBC252WntonNpZlrl71wewiZiCAyxhB5YYbG197BPSIqmScJ5XT5a+dHDO9lPfhl3+JYMHFuen4kyKEVOQaydVopuuFRrlcX0H9CJk/uabm2VhlyiwiSLckwaOtFW/ZFoad4D3XyB5MwbDxAXfcZUtKxZdly3DW4H9cXIaeglP6MvclCoKFABRT6nFrE/S36uqpbjs1ZXIvGpCsU8nKaDScLOkePFsUkN/MBglF0KOnqG+q5FCkpA1JK/x9F4qhxMdMRaGwVPtEMayxMm8kdBosOI17Q/2L51pOFV3WK0DOUMBmI4cwSwNELnwNGayFvklaYd7I8qCmDnu4DfYXciB+YqTTqAQzeB4K53DnMXyx6QD/Gn0Dw9SVE9uxvcz3gyqHugT5wIsAMbGtnp42qUABcBC0hutddnBVj+am38WP1SJudg50sPWB1Yqqz45MvStI6gp60bflEyW3unWR5qusnzavG+ctFjdZo8EsvzpW8dghoCYZYh4RfFgOdynWMw9A3PrnLLoUczdwhlsx5SZo7q8syMDPfQfp+aIdynP1GpC+XZItkVsT9uOTOwHbJJh5BW45fGCr9mcMyd5DRlT9L9B39np+OL4f3mgddAaM4hfKNr3JRCCauN+/MAX3zmlQctN8F7Tm6UueFjPqswx20UamlVZ3M3MHIpKoXBamM3Rx9GgDhUUwI0rLNJts0tzLnxhAMoeb7Q7BxkhqHENak5ukvfbEUwkaUJ/MxHmWAsL+h8zXXKuOYzcg5ZbUxW3xUZXnFDrydnhZDBnITTWO+WN7d2Ug/uS4Q+5dHBML6y1M8bDen1gwPlq7uIWH4jzR07pgbkfg15zzFcS6vr4Xh8/Wawvi63/AvMJZ+biN4iRUu9DYXgAj2GvrrvwPRweQ9dLJpNmdJuQn13EFzpvp7gD/376hjOVDlzB+m6iV8H9V2xwg8MDfbrqFn6elJ2Gax9CZbrbB/NbfTxnrMi/dH24hPj4OOv5PSuZrtcx0C4McOVqNDnemJsUIJ7DXV06rE5g5YBFc33xDKjq4klYjFLpzG9sbsqEAhRzBBXRTEUz+w6E370Fyfn2Mdnz2xAtPWJyunMd+mXhRkmZqd3gdYocBYZQ+29CJVxzmUehyoBSWQRwgZseKsZ0NvOeZdVeaP72T9Jj6e67InY+C/FJ8xyUIaGvNWHAtEvWftHzVhofAMHJuVo5sj3JcwjlGUUph79dw+Q/WLzeEHu8zzsNa3Vt+LJWDDN6Tek8b5HKw1XWjgWH2rmCwvL88kJFVJ0F/Lp/0niwg9bubCcvl/pFqnZHNOFf2md33ol0vOF3DLDNe5nV4M1rf5dAceC286coizb8snAiuzSweL8KOQCMv+hRNsbepOCBVmzi9E0idFqnEcYqVa5nxBriZWLDiQj59FtM+coBr200RgcU6tbIGAu3QQvi6jP4TV/9mBTkN9Ey9UHkrM7DrOBKOYEfUvUXCFASPB/BlLKYTxRR+4slMKyzCmlEL3OzPX8UXywl4EMMa3kjJpOPuvM+s7qhftuzPERRP1XBjCIS/SFN4F2329a/6ffnsE+DnGyeQ5v4Wmu+sagcjJGjGRC4L4PR3/RFjOPe5lISsr5yhuCXWA9B2O57K6zsfuPUl1S1x/KI1LSkcDOfGkrpvjAuXTAO12pFMPUiICX9/MO2WDIn/LWnoKfWITkDaEjBhWEWYAii3TXtF6GQiJ4GJUALzKGRhmUyea6PiCpzG7RKfkUJtcCWViGXF44CBqn+5lNiUeCbq+7CH6L4L7CD5IDFCxZfrBjhgbFouq5jTW54PTNXChz86C92VlaVSR4gsdxMMhOzQhqToThPr/xwubegUG8NdwW2Tunl+m3LIoqEBZZ2RwzFjfvgE2bD3Jb75nPU8OhmleJCHGsbuUhu9XNdt3LX+6wox5tGUzsMlTLqvqup3CC8c/WQ4TxcPsCkB08Q9RdOahkcuWz8YYcfkkhuuzYrHvpQiamjwxrerFURKX596Z5HR/3hNm0g2SucSxRNS8zdAcdWFfVVJg/MM9KpARVXoRHhZBwtZN2a0btPy5clXQPz7xSFwGwf2XW0hycWDpnMo7I8bH7kR0okZLS8OcTx5sPLozmkS73Alkhxc/tPlaQ4vyvOdhszibUYdbiiiICtomaX7MwXNatIq6MNKA6l8BQoyXW0kaYzbCU4e7Wt7ZPs6/7y0BZk0Oe4HP1DeDQIT8qo5+d74g3Crwh/ZvngmL24m9FS4Bla5XXOYaoxEnD/B2M5e4kKKQTgt4w1jztaWHaiNbSmNdNVr5TY9gNCLSeKwDMzPZsq4iXvjrHiffL7hgVbH8kRSEBhmXgdv7fyCd4Et3cBgF6uPNBFwsAsCp8Y6cAQjnttq2b1cm651c1EyyOjJlHzEfBZtL6rIrcZstruH0EekBE/r7Ix27vxHFXYzpgDXu1NvXwXpA5WJpQUH+FgRN+ko+9e/Y4TuEfRJBJmVMder2M59DKUc/tT83TmkTxqDE5aaOAWGe0In/KliweJvOmRoO8FeliHQPfPo+GEKs63N5Gcp8nkOsh/LzlJ/v2/5Ot+43rKA4H9yhtf8Hi05SlPy4ZVGfA/9WSes45C0nJ45MPSiTGn9gNy77OJYFgjkGcXyAV6idC2XUoLXZilFKGfbkyMIOrzxNwTTSZ+9ZExef0POQVTEWwzRqCzXkiBFGnL3k06dq0CmzgFI2mc8mktpdPIakcrZLgTn24+AmvwudiS4+ECkmbvem77dSLxtQBPVZDp4EoasLJ+EzIwLVdh2J9QlLGiR9AshAemro/k/gGoebbszh4qj9EXPZQseJ1OeNT8TFkMWiV+qsjfS4IvKEnML0PvkOUuhjIL7jX0UQJSCF//VolSHI1l8bHK1xAXrUwYg0gtYXh7NFdn3V8hV/VnD0HmSE0ikpGPML6EUEG9IFQ0vdZfIcfXxJ4EW2WMkm6u1Mvp81rMKaNMxbiwQPH7lB4Vpn9Ux1pbCoITSqM/vnrMrrNNcxBeQNgc9NiMW54//AyczL96E6PN7KPXVa+HxDnjYkSsmqGHltu8XS0wK/msn78KQt6r8dfKYzq5M77Fp+Baj7gQzZ2edBQUsetrHFZCGU6pgdpdmWkh+HxJN52N1cT4Z57JsWFpKxb9YkSjkwBFYON96tRGG0nn9+qePYSPLjfNdAMU3Ty2BiUCVsIZVEstieKvRPu67Kj7yWn6aju0uJZyXvPo8UCG1rXNqZ8oLPIO/09FJHM3HTxi1TfweY/xo4WGEVTKQipYDu2ksQnIGCf5UiKwBiWdjkMAajGGx1EJZ+sg2wZOUisUwErmLTpTz06ha5f9Fa2d/WRbeH6TVg442d89Dlv7V9n4E0e1xlEJw9OC5HFYdp+7OOQFg3bZ+jzTS5liKad5M7q2npt3o/r+KEcEBwXsdjmExXL886IGp3MOTY69bBDnhl4p26O9HSFbg0z6Qrcgpn60dRASSKt/NpXg7CoYm66mYmV/fMzBtKVV8/NUQCoRnKlSJ+sgJgDl12VXv0m/UEc0hcK0qXtDTf35C5S1Dlz2Ik09uYD/FgffJliWBekll77aU8PYxY/K9zgdpj8RXguBdn3U+lW100e1LBrAwoBPNp5kZDPGfO9779aK9FvxTjq/T0fLGvcrMqqAVhu9XMGPrtsphnkTZp5CC4YD16DTbnCJNOcs8U9sgxGARoD6IZSGtu4jMfbbZxE515tML6tNRbbHtuYj0UjKGIHIGgtFVfcBWU/SJxRPqh6zfAHWWJs2fUwWo4gc0JQpd63lkcODra/t5Ophp1Ql9vxsMzuvZ5HENUEZrgI6LeSTfogog4mLm0Lm/RJz7hZd5oBzCtnhXEb9fJudZYFEsIhOqRVYpAmyuEIdmvSZIHxSLGramU2I4Fp2p+usePOJEKgDp2jGJDUGVA7qbYFH4WSHK+BDum+lVdeR4PwCOG/b9YN1INejq1e7nD7Swuf8ZcKD89qNE5J6KJ+TDi1WHzYKQWAod/iCu449xYMBX7vb9rBhqxESvsaLW67rHqVJOOMqnINElzECmTUqB+8qlubPxriDwXU0V/hyXDldxxyYseW14SM36VFEE2tfTy1SKtIVB7eVRk2UR64tEGmnEDdRTB3mw8j8sPYWcS6EgS0DOxcvsO14AY2rpVadObX2z9Zz6aJAGxBYkPOMEIs0DsFuz616yZ8koWOKHARUqkn3i/yvfBmKOy2GXYtLfcEaAm/1eR6y/6CPLeE+mt++kgw7O336Nu1JWBjsTZ/5W3OLoA2WS5oD5O6hy+CHGSnHGvi/ramUlJokSXBt1bBCQxFwDQ1bHYaIVmEn3Qv+Hlm+MBTA3xfsvkC8M73Tf9+fq0mWM0tJ4TQ/cwpXs/yR1e2jDkqwhqQMxfzUNnUU7S3D5nCpMvxL/KzGAhS0BZNHakAq/I46+2f6qAo3c6lbX3kkpQrZaOLSL7wPUkINpRnaBkmYwL8bmZNRGrXMwDtrT78p8zr27RmwyPUjeWpO5rgqib0hxAtLuD0mHZHMdGCdIyC7LZ1hmmn74L3PkVr5exbkW4FFg0s+wikUsH8ak40Zn/lsM6XxP+094iYmoszkliKnoPfk+1JYQNvS9H9KwgtCunnSl4Glc2OmDbFQ7XiKcxiGbTEpqJshg9XMQfuML8EROiTE5QAvPId5+aAnRieApWpf8CLKwjp5HpNU9YJZtBkA9SlSYZG6wQYx9c72tvcnJWzjy88VXepTuIo3fEwu5T90N2wE6rSq0CWe8tMj9GKg3lDg+xsmtfovcAPibljat+zDNLLPV7XVspNH4G5qkm4Jlr7Z/sGXS+BrvhZYSlD9tmSRWi9rJ+3PRuPMJRf9Ks+6okbsUATHRs6venW77b04LZRkdk2ASBXq+0QEBka1fy2b/bvGs35pXSBV+YZEN0MzL6B3M9fm3rf/rlg1vMjRm6sErkz77Osd/tYGwVGDRMvPJaMgUsFcwE+5b1L7GYibmImR4XvYMlY5UJ5PnopHiYXpmMVFsm2vuYWuH1a5aZtMi4lrc+/91Qam0bTq/gDz9or13mbmGK4IphojvWYa5QyOlyHlwO2r/AOMC2zMSzcJtoIIwM/d3jHH7nKMvzwAbYU7IX0clf+eiRs3BreiCcMrFF5qh4/cUnPrONGKThIQab9tuA3UF4MuaSvcZ6DFE9iWRMvmd134Sb1JBSF4XycztcALk9SehRFTqkp6Nst6gr4VQJuqkrrterIEtvLDDwDF8N1jMWnhelbqWTQTxAYaXvlbNQUL4p15qbikp8ZhFCY/Wiu3ZzPfxX4f1amtWlBwbMRyeaLODi3B2UZgM/1VInPCmF6bblz9COFzY/i1JllmLicbhSb6hT9gizGMc59NzFuKGsVPNdW0pRMHG/DRA3eTVds+udNv1oaOpOk9dEmB6jW3e2a8pCQ03m/U0SwLMx94E6neHzVsYmxMvkKG/QnaVEUsIyZXuAZ7SfeW+YEQVJriW4deUqW+rR81PWr23F409Zu0F0lyVGY/o+ZtVDNlS26/Dl6C1a+7FzCH1n1xQQsMdUPRDlU+goRQ4BcOhURiIHI70MAJEGhK2UDr+jNIASRp6dz4wU+PplDzvjk9I6QwT041yJF2JbkzBmNBRYCC0ENo50+JSORF6ZFeMcCSj3IFvYrzPLnVRud/619/jJHENYrlu8nWlPO13y2fRnyjNtC9awDCu626BzvplOpkBJR92bULBSLAdI3b1acs1E9qdvIKBLmkgqTfoqOI4Ynr4Goii0l/HqejRSzNbzCogCB7aX1s4DI/ZIB/DS/yMwG0WybyWj8P27LsJlbLmUm5r+YfKDCh0jjdmkJSzJAzBG8Nm8+A/tNy0iPRvaceXTA758mIqfjoXGuyivjxzKXxS0cn3hrs9m2lXReAtlAMw5bMYCNpLOUTSBAIaYXVwWbfl34v60bfAO2O/SqmxJXaRACy/mkJSiGR6eHYPz7BQ/2yyvBZRiUrQJBz+WZ245XK6ybmJuA+7SedB2kFPIAMu/JeiObNeU7oDN7qqreLfm9biECfa43/QPXBQeBvVYLNL8s4208pNIWwYXEktCI7CvbtY+aZ5BplAS7UEJDtlJnSlXyM6TG92iEMvzSb1KPbYFI+VpWtw33m8i7Yed4QA6Nd/uX2lA8m3wLcf/7Lju1/XJSLIlYeQaqJRFiwlqeuGNkNqVQWqGDxQ6e2L0eGhslc9dHsIjmmsgqIWQEGhIlSHHCGOUsq4MmI+fNdRje+lELRqH4rQWIAAnC1wo/ZuIrz9QSDVCJLfnXMLLlYZ8aV2pomxF+hnKm7NYIB8BFs5ANM/ehv9Yp3sdEHQGShcrxWZMQ8EDEf1yNrM/hHJKfDX5qkhDTsxd0p1VLmqTNbwynGJbD8xweKMWNXMlGrX1GzvSUiW5U/rL2sdy7aZbEZeY1YoaIj3iijHepBZc+jBc5hIugxgT8Zim7FkoGESCB2TlIZS/FDegtMMf0WC9LBdvX9BE2gjCGflAsfCDpiC0CWvYygDod4RV/QObgbWjCKNQbzi/wD9BMHbAyE8yXeI8TbXfrS1F2R9OlJpo5cCeTSK9mDMXgarAWXVJUHfjOmO1IEV6ER9OqnmQN0CK6BXi+ZbMR++l1RYsxVlO5RAxro1K+eEYgUxvUzWHWGXEnUkFW7mNdMkSri0Tx7+nsvp6ALD47yLw1q2WbUjjilR2AEp4DoBioTbcR+IVfksvud64KC++nh0Ftw663toNQQwLfFPxSl2usSxi/iOi0TmTty/mkHb6rMQbzvxYAJiOs3xANLClrrS+HISKqbOrwdSb7JpobwF7/57CYkoL2utGg/Owz02mcPuAV5Y6E+6cFciEve8WGKCncuWZOdJ+4ND0hkSQdRvybbeG7Eo7hxfFYwQoenFniSQkaTe1MSevldhWcQIPmTyOkp9f666NpUmZQPUCFORlHLYGjQ/jlTMFShEut9uz+Ycylm9O/eQrpnUYxLIcEvrSc/qcthX6MEzAZJngMqTfvbHVdJhqSUEHgBeD0KE4TpSVM5Zl6fa76upfDa2Nn2pvwRrnHmSscz23FjUdWwwgcyzgD3B4IQpeQqdEnBVIDmM7/Glp8zbswwJrmAe+qYWo=
`pragma protect end_data_block
`pragma protect digest_block
4c61b160ff1d749a39bd4e0d397f0879d16fbdc819b2b7c055cefcfbfde4b595
`pragma protect end_digest_block
`pragma protect end_protected
