`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
RDwPnVTjpv82rBurtIYz5jl+zJ8N0xJl1BwqRQh4vzZDUHaQ/cNr1vWBiMvQgpbi2sjuFEYhRU56EyccDMOohyElYffJOSY6YEuhkCPMu1yPLlIJzNV8G1FR8gPni2Hp/ThYIcChVPu785I8W0zSw6W44Ph+0hX09rEk04CX8v4GwptpA1MBfjrgsQQp/tXRX2nVArXKal2eepIqlX6Lz1p77cPr+mLd6GmWi1EdPRwh56dScF/If9ClB5NU+uhWtBKrsxUAiS798bir+grEtKxhxJZGvDWlwKrMRhHDjZa7usOvEyERJMBdvEFzki2BvdQYNDIT+V5IVergfXE/QpemIKBwrtRGMiSqehi2AQYbLHCdxDWG3OzNVNOa96G92LqloMk/63Qkpf6+3AuVkDldWiAlJidUQqmoAy8dtqsxvBhWQFOriy3Gwjw8UhXa1djroZJjkB+wD5aw6PHTY/CtEKe0i3KmCtlcfu3hVFkvr9QCgsIf+fwj6arbEfzWvFhK3zpP+s8wMQqGVXAEHlXN6wbw4LkkWj+10sq9CCSwW4adM5v6IlTOnusYUrcdV7Nmivuc0kQ+NzkNYkHlJlIrG+lnGFG2r8vdGOwFuYCuQb/njSYCqYro4eKfr7JYxrXUroY32CrMi1jaU1b6UdIOpLjftZCDNEYEWDOOt/JeLe/6ftWSPoM3T9OAGMUD6I/q2LHcOEjY1PWaFe63z1vOaQB1WTjp2xkvQS+AyZL8xu0ARXCqeWsMOVN3FGiPAEUS0fEJVEMBOoSdo/vpuA2UYwNwyAI9fK2EAUCm10C58eZ2ix+6mosRkzgpp8MJaYlR8cr6kG1OOEZH5CbR+otFnT5Gh/0SueKvJ27lqxnLKE9JX59BWubhoPPc9mAtmnFoAqsV9FX9PNv3BuBss77QHtmKImTNByg3Lv3ViRYebFpKmW3Mx0aCYtkYIWFLFd8LdkPyh3bMrls4zdsrK1fDz6ZIjfP4laCgpGzzkPCJTUru+ATHhtc9KmU5wcHcatOFN5vUrZkh03dlONUlSGNKC+nKE49HerXlnrOV8cosUt2+1fl6QeQH7PQG1BsByrUdzr3QZnM7xQGKpZ7QFiU9aAXXVSn+gYpEONQwtrryEtE4vtTo7+xAoPgwl74TeOoVmCXvjOaXpiZVkLEAS8k7KKsvnKkLREwS7avC+e1U1zes44mZwNqNitN/G7jrZ6y31dL9IX7XM+jmnB0IZ1tY3jwRGLqvx7lzo6jMTjRnLl0dz9TSBlHpVSNowCaLgNQINi8iERiaHydP8fuBgcOlqJpCXvXbrcltTYkoZgLqxBa62NYNaVKIVf4V+Qs75tzaYJnQYa5TEl1g3cToJGBweV0ZuT6qNQaaYuO6QaVtPIeffpdv2wLyN2OVK7VPre+L3vB6jgMlxe82UGmeZ8RdqXzqbyoPkvRLc7mS1A+WrBo1P+0DY6510ze4XFoTOcayGMklN+vBByKmlPZ+9yKCLLMb05fmuskyV8v/xh1PUP13QUzkUZf9uqTf6841NeW+Z/Umbi/Rji8lcW718Xqb5ol4WHRAB8LsD04lkWzwW2M9F3Q5eVW5PHL4yYNsKqOA5RvDlrB3jq52/8eqKRbn8qSpumzRCQGJnDfmefSk0DRvScZa+tVr25LUGiurtBxRnrmLJ4Y6cEeLR3xdKmxClPW9qEOPnZN/bsG58k+B1JOp3pODsoMfDoyYBwoL/nvQqk0MzK+CrgTWkZ5R/Qf8t2kgLIDh3By8NxWbrlEdmcyX+EKgbRxKRfGcg3joPdYFc624C2zN0IFltDer0+0otLN0Ti8Rbvb85M0JDWyTYZwsWnUMljj83+N/3HjZhw9CvqGgWNwjqKkSacKzhBNtXha4qplOfNCUTZBDl5kiCc0E//OtGmkRCl+4FnPZUZYMLaPq48EN5yB/nLrn8cgeveWm1HNyPTkYWJqbVapDLNga6pHdMLGaT5u4YyNad1uunSi7e5kwbrvpyo3fotGWBY5ajm7Z+wUCyPciexe1hpABPXyk4KhRUJAGq1Y1WliZ91POK6PEz3eO5eP5TJTubg3bn0WLW76HKVtD6ML7FTpv3buetUISx9K2PuKk0mvc7LXoqgusP8rvVzoDcP5zkS4qXlRjflGVphf2Ep0ot1iKUWvFUNkowaDZmMG8Pmhwb6HcxYLlHX06c32CIrFh9nF0yjxAwp+WU4COxIdAU+LowaLaqC2rG6tcJ03wHaG5VUGNYJn/tTxBSBSV7mKKXLW0/DjgRwI3JNulwhZjx6P6pqLBEuSg70pPHqZ3vOwT8miG62oP/2tjEE7beKKT0y3i0n7vIkvFUQoyzOfwtkW9cs/J1BNldhcp8qFkkgmm5Ntxvo1ezkKofD85gWfAKmnvglLqp2dqQ5cLUpiJ1CDg5yXh38OOXQabhPNIy5r4fhIXDjfIPxnAySnPoSONeZcwcUf4vqsIQvkO8hFWT0I9oIJetllBsfCnHsqBdTmlEdmt5l3bnXaYZHP9Ht7x/e1vXFJxi1p3P3MmYx6u4iRvv91uG8dqaWo3j9LF4033j9VCUaFOENrsQaeGaU8XIPr1Xib/QEzvWkCrw0ePESLMSdvMcYn1op20XNggkS42aMRBJDye7GWcJdzIyZaUR/AkdBmD0qOjljpepHu8AzFDoZ5sG03RKuhCotAJQ4QluhpQhr0p/Na6cOHt3pA8K1OCw0WiBxqtGMX8S0Lj9gsl0IKTz+PBYktBGIhyWqgkleTuFbSEklXkHH0tn5ikk/ZWSxQ3DnKsGgAxzLWoCG4C0O76mHjqPXI7ZTkk2jakPqPAAwP4yqTtQVCtuDPSoEQVa58bH9j8SV1dNkFa7K7CJWUtKnYT3X6xwiGK5bpLAfEzs89F0YyvlxZj2LQ/w8lF2lCG+J/DWgkK+2pUcMTrw0gsmDy9UUmQ9+64Tse+fGvbSVrdjhq7rowXgXxPITg7WUJZvBe6H0pKw6h4lDRPWpU8oasz0A0r5ixHA9jUs45JYPm+Pel9uyNAWdv/HyquNQvH4FDQtD9I5NnqEFqDA1Ceq0ICDGqiSQmy1+ArusZrwEQfBRdLcfW8lZd03VjjDsbmlkrUFktbg3gWZ8defHsQFJ6uUhkEorRenpgZ6uPnQj/+1b/FsnKAVtvMaUbHBwa3Dz/9xnsEp4JGSgnwWSc/IrVmfQj8XzM9DfsQqeiHUQE4UX3nj4KtJaIynVPnOuGvqlroNQjHRNQYmcKuMmFpul4tXelMOddeYv5fPOZtruEG6yq1raUEUsAUTHOCq80YQfeNjsbErJsB6wUq3BDLW/KiyXjamvt7HLs3LBgjaWFgnm/4l8CJKgpGWx2XW/tRBppctnXEr78DufM0AyG0NX3pHyH+eKYJF+z6B8vK1Rls28lpAIgYBbWuAn/SqZBYPHOVne60+mEbH/yKuEjDMgxUj/qy1LTam7HNuT3znCsQU27cIM/EEUsMjFlTmE7vrp7ROIsNy/lhrgYmdgDkrhfF+j8vPNs13U5Nu/0AVO+aSwuS/2o/ePTUgFGn5c8c8z7HuaLc/dKLN7wkoeWPia56U8hdqgBrDryjQqCyoBCkMB+64hKmeYrADfIyQ77yrqkpAnwIe483/snLfGxRmHFOcL9JxQi/uwT7h1MAIhZtYTidBuzWwJqRr5P+vnNE1UNRhyyz5mEKhP8eNNNy8W///FA3f7wjt+DyvQlS4JjRSsNpxfoGWKDaDpHUWu0Qo3PfDa8nSxpyotPo7+ylHT8JSY4KexHmQCYGy7d4pIhzdFp2aQx9zquWC7iz3nY8TvhkFKsokcp61yfRTipmRwdYU8f2wGR57OunJmgYyKZLCI50vDM5EGXNYxEjHsdJNvMvzKgMYHRasTlRqetrk3AgnTJmmCPL1itDFvOT6lNcUBOQB5UR6AqAbbah0Nnl71O4gRkV5NLSK8SHgXjW+kNgUTFpMWPwkvNYbT8H/5QAXT/JKxmoUuRf23o6B2Lap11L9umLxc1Uz1m0fqOvZbuuhE+BJMDeFWUj2uB5ZXxnVvgFZjD+smkzWFmL1YZO73hpTj7T6sbO8BLenIaALHADfFwSC6VT2J3uVc1Rxjefd5T0W8/+5UfiLjB6NgcZRLNAVQRk278imfO1sNr7iqIdb1jf9J2gPLQsyyvkUOj5ln+7piBinSo7SnMMoCYku9h+xDj63woslpYCt7CmxYrVlWf8Ode7b8zBZyooOb6RcB6vDMc4gMIpJunl6M4YEqKUlynP9AhgQVjnKtb8eAWqkmLyQRbv+LBFn73LQuKFXi6kP0rHA3W38iElFar1Q/9mWcFWY3yfyuRsVdGD8Bh+EawbMtCskGFJPzWOlWbY5LHAVQN77dVgnZG9j+GDqAl29ksRQJiEehNuUr2re2OE59o5ODmT7k/bRET5KlZfGy4D3CKgsfej5fxPpGVgVKp4t0VWj7QQAXaCiuyzan1wK4Yv10r4CfSaN+TL4/X6w7Z+mShxFbFKDgfpsHpE4nEspO5kY5E2ncC4caV8j7hWnNszCN/HJX/wkElp3VBhKB/XnZ1qnMvhAwbVr8yb4+XxQbxbPA6fwpf5gyZajH8n5zj4U1przQYZy0hNEJObh/N+UEasCJV0CFtoXOBsx3slKmMHhBLhHNoqUzKuvZLuoxWaQEUuyUxjWCI4liJNkk+cz7v4585u9gcW29aPLvRkVFN+jXqnNXBos8heq4ro9N9MaT2r9EEEBhIFh+5h+N/j0aAKj/qRCXwXNkUdRmcCPza3fmhbgn+YSvpHXKRvKf3mJ4DhOKROeAvLD9M0uvdH3hmWNzi1/dHVzh8iHF90/lcL3Plhaijr/xhuy+1nM7kPpGzOkJ3yf6sOV604xN0J2HDaEXUO6gBgvxAI8xOTmkD2ZTaPy6ysL7L6PVwCd6lhEO99jbYQmIewkYX/h1V70zSt530XiKiM7eR0tpdw0oNS0aE41BOgSiz3KFUqm4LlQ/3kvfckawvhjpaH3rAJ2tYdBh4vTLqNO+VM4JXWPr9EIFgNLcjUqt9c/48Tpsaf2jZLWYk0BHZ7euMf0nfvKPGVH4GbKFyvq2B+AJXRuWP+39xnW0NkAxczP4ZcL2ojQhP68BVusXFxsDNwIJ1PkEBobDSF3q5LSuXeLgRTWMCPmRplRmEUwkE6IkkShQ1mbsJ9Q0H9IeD0QgYOw5Hp+KWN1yVEWNl7KCQa0NuVFZWSWwJjY/Li/bxiILr6jkaoVC2KrotK4vjxkhz4r7+ccicb5KUOwiYcaoSEt1xWI/TKHnuOYfVK0ieinr4MmsOJm5TYmsyr/syEAucD6oE3sOB2lPpIiIgwxzfmKAkNZGygXaYk/lZDVlsaRe+S7tzCFUbyMyltyJSSGUg8Xkd0LyWXgtuEgG9xDJYujhfEnIdq49ataCZ7TTfY3CAVM4TSO74VBJqjw5JRWK9Bz0ljcXHWnFiyPg+epKxvHUoccbDB9IwRaSnzREJyj5OWVWbWGUB03DB40MiAOp8HURNeZoPmkaZOG+4CKzRgKcXVICJYeuthRkCqvBsnxxl/D1pUitd95SNJWh2JCuxAhFSC0O22LMvrW5TqcthsaQy9zWU2wrO1UoSZ+Lh1OLQrTmMC/SrpvIRssv7Ekq75LHm7LOlELJtZceXg6J1iOl5kkq/rEhqC+UwY0u3saQUM7mFN8Zo29vZNyY3xUERkSjV0+cQXcXYkTekq644PKiCHfPQxgNTK1EQ4QyAJ7Wy+BdIZU/5+assKDVCxYe0a+KyJDBPFeMaCknoEGVeVc1tupSV9GtMg+KOJi4zyLG5559sAOu5ATBX3umQ3eYIAWWcXnXHWe3jss91Ytmc7IPvNlK8c/kAdW1UvcDUSFqxtVIJdbNHNSYtvjGieD2FFZLuIrOF2AQ6lP8XtWX4xHwCiW+LuWBkVREULs2pFMuw/x/ysAY2YXczg46E7cbRjZiAfa4/8yfmyPv60Dk4j/+6zJ679Cj3GwFLFlU2iC+oOFGkVImbcaM1H9ibS/COfCHKWkMgL+ZyvtC+r2JOSJvNOm51TKoX5sbmywD677UFz9y+U0OL1mi5JVm5C3sYGLUkW51lzwEkBTSpvhx04emUo9kmh6AfSLWkB3kmjB2Zm2qq4rnoXfoKaDLEXQMg8tbb0JzkNudnPPbxhRHADCLXZtbAPtAHXytThoNpRi11UsGJiAsklXnqoe/Z3DojcUNFHSJv689ifr3YToWnSzWyf1dHGcZw3VAov5Wd+uaKFBDVq69r9InX0g35tnF+8i1pg92CuQJPoVTeFiFuwtVBU49clIUz7VUeN3PzWXFfzZkRkmWOhjfMjNCvYSbofHgdAEQZwW0LKk1WlPN5rcXzjsu94jdF/7WlwhE3dgBBdvNqrvwnvvnmceuXwgXsw9rcPsVucJ7pT9P/1E6tH/w4M5QeAj01hb2n+jBa2DgLS8K47da4ywIIC906zld9Haahfr5J0ktQgu7XaUXq6gjHdeDMy+gl7i3I2DFchIUFyxZ/XPsIl/OHbZyPemTsTv4fPlRxVoREGHpLQwRwLZfauxBJZs33tmvlG+xt8y3AQ6GRt1M0cZkU1stmtSxT6hxvBrnEp7xJRMy6iEjyUbajKsUVXFFKNZUjBZ+EzLhU7REXGevUcn8hsbiuGDb6IGCVeYWelbobhXHFkCoXtqarR96oZRR/8f89kAMo32sU45U5Y1Mjn3Q92sFRou4/u4Ol8wPO+kK9MtW1gK2bEVRvvcZkPjXn8Y+hzmTgrsrBHJ48pooWDVr9OJh0kcFEjBkQU520wKtKbY/qcg3W4bSCjVKhw+/h2Ad6Gx5xtlBInSs/jc9B7VMSrR+YpceB1YfO2kwNt9I8VoxBffvVbZ4ISWYg+nhQCc8vtgFLD9Q3/umX/zX7nYHbvtTWeiHXzKIYTqqBYVnsnBrHtD8zgjJr9BIejuHGnrpVDqtF+iiaQyIvEKo1mE+W9kbZn+0Skgn+uiJF4fGCi2Md+T9H5HdCRhUixxdKrXKuMOkfqR4zfVxLRQvuvPManNE96TKTd0kIKtdIVwWjoXLDMgCVmSIyWSI0NZk+R2gItQR7t5i0Pc7405giXZdxSp0p/mO6VOTeWb95V4I7Ia3N0c1aVlXPVIxQ8NbDbUMdFkrha+jm6ELL4qcrdex+7p05fW+nxzU4xN4GdSxt5QyoM/VJnr2IuUBzgXQ7OCCNIH1KeLzkGCK/RE2jr7BFcN/qG8t3pyxw6oT35D31NNOK9XCeEKFXkaPJXPa6Yc1TZ3WMFwfDC9G+7VfE2mJ9oKMEWtpwCJIxki86SG4/4b+NoVWqRqOPG1BWYAibg9EEGPATjitvPSgrdjulc1X6n9ubnarAxMRnAE3k/+o2rrVH39OFxod//JdySjUwKiGO7fSBp3+xKVwcAB/Iw6EIRxGWrJSIXn4DOO1nC+HC2PlBvsv3wkhH8I0CVhxLB8Tu0INOYIVZWeDxfj9sTZ11D5ej+kLk9/tOPTRaIp5hr4Er7BF7m9/j6sSirNm2ltlIwLYCpVkEglFRRIW1lT5WC1/I+18YMkfNZEOPqBgNRlmbOWdC5e+qkoRDNKivwxyhtJ7q3tK/rJuApFXc6lbZ9peXdMJUp7z12UMp1kZeufRFK6GhR7gZ3z0zOlgD/wpKYCK/EGF0y0SEsHqQuehd1FFoUsebE8pXft/W9cpQnZREAI/8OqQ+uabe361Z39zEgr0yg+Tp7BwL+bR8IhCQqvhL5b5uWA8FbCoKdXZAQvyAGEyLHAr9IXwNN2R5CBFt9CSWUkZQniyxlrgF9uXxcwuVtL5JEjPSL4NAEqDK7gTl+qGbLZoareHxOdBOsC73qhUDj0vyh6CZUf9EuRwjZSE+Xk4TaD2f+PfAsCcXGMKDRmeAu1ELrU7NzgG5zzrTaoBmwsSsGDv3WT9vAoTJ/D97Ey3/N/oea6A6T/wgYyN639XFVT0y5Ju+O4XA0vGo2a85BYi7kPLw8Rqc+KaUhXOs9ttl4ib+TQKUPjr49olO3wOpSfDLcSXWomJ/DesxiTZFHai/OSl+RtH8KvtTaUczxb+YEsoe/FlKbU7hyw32EeaFhu3laaMIqDqR5geF7AuOcd8xd5AvYt44LxayWXWYqUJGaEtNi3IRSJeOOufHbuu1CM+OLwGtZqNQPdikN/mRaiShKM6vgvABEVWM2+L9Dow7CYSUQ7Df4cJXE0oLgMJOGKQk88F3gFeoBQ2/bDmq4rQ6SNaoYkOwDZaf1Z57vUDXPxolR5c8UkszmhNHuIxFRUoNC6UtDzqfIA3mpqhk0bs0vFWloSGWF/kWXWC0DCfEjSPlePNT1MmeyuafyzAjTcb6122kTkeCRuaI0quo/wsWHMeepY8ZmjwWtE9F2O9ywoA2C9b8WjLT3qhlIRiD0yT4wKGhQJVFW8vFGlghhR8B6NZ2KlaRHJRuqfwXlUMmr5uakV28jt2/F1DYg0emlSKc/xRH/WaVHt1Rd0HrvADu3QonrNmJHp9eG27DVzKA1bChPi89aDCLzls93erH2kWOYEtpFS1rF8JPgT+QlsSSUF0yA3C/Xn6hdG9pI3SGJ/bGXNEF7Y+6+7ZR0fx/1L8MMZQ90wXcKoqmab/FWJo8dqK32mDWFv0QVupXVYaOFD22AgiTXYvTFPRV+cgXyIryolztp0wXul6T17/VN6cm7DNgNJrkO2o215XNsofyvx2jyFbcUGlbAVtcuNNdb2IB9lSKCLMaEorOTbbnTJQKlvsIu8d4snJ7r7Ri/6GgWeupTUH3i9c8LPcFmMGs2uS7mZkUFvEJtEcxBOFyoZdYBeAniB70dp4AQ5uSjNKS16j2YQZfuFndFwpE0YdYhOmpbUh393wCeEF+vJ1YqctEj07lmWP/aDb5iIwxCEmk7QVv9MbTh1W/qs5AwUy8cA6Ak+MCuEoUmSDa6VL24mG3a6wG1G/yH3hU2WW9GUk3OvBxPk0wtrott3QOFAhHdJlhoXY9DD3Ic3TIuUB7EGLAhLLlzKnxclhSqF+qrvb8e0YITwPz1mP2Hl/2KLXDWf6Nm/nggOIs2+isanW6JTp6OusNr4VVTZV+F31MGeTl+4YbPVupcwNyyaGM1YmQfSDAenTZd/nN1k/HBlAIpaniL8XzsLR/uTTtjn3OBK2t3WjD5QrZ3JgXDHBBAZYTXxmqDDN5O9tTNuAvtRZHyvhPg6AW6SXtVwn/Xv8cS8Bh+TrSd9WYl/MV5RdssjSXioXtdruNN4GLQGy45TfRRjAZ4hIsw2mK3NE+dLVHvI6Mq9KLZcnKKd7VkEprNOCV6+oDjFdg56lJtyrysr53zmt4rX+o8YeRj9rJD/DTiMKgLt6RF4lmmJBM8WeI3XN2AnI+1YSAbRKPUtD9lmk4AiqMmDk3NEpzPhWnC0twW+CRTNs/8CrwRFaNfrpy9IzG5b6yFNV7+h0AEiJUgrbsVnYYEBdg4WacEZJvu+d/1mkeGuAdsOZ05IkAIwKgUK1TpJcK6QxbEs17t6i3BFwYaOxjWm1Lzr2F2pD6iqan6RESGYU48pF6liheDJ01AP4OEhUD2zyiBNttV0s6JkrJNrcqgenkWjkg5w1W8YTWKq+YVP7CeORk8l9PtpFVBOvXdOofaFpp8VY8HLbXWt9AMcUhkK+RUe8Rgc9Cghp+ijPET7C15AijQ81wVqitQJRwBYp9Z+WdbxvV2sIhZIHOJ61Sxh58LcUqw8sLmAO1BtxmnvAHlHMGWi6HCfeV+0xSZ9p2ELmWaZ9lnW7Kt+JlibtItPN/MlnqEPU7/MYSFtzAjV5zFutxIg90Boc2PjxMmRdU2b5JXxDHFVxQKEW+sutR7dUaSWX2ukXrt+JItZkjfFIOjrnSjDuQCOiucYbA+rqMWYd8cHsntf4EYXqcpXoqRAk8cPPKgqCWl6Da+COEzVniE3Ry7ZXQc9k2xA0fN1UDbYQnA3NpF/MQBoHSf2LwDpBvsRoJ3dQ3yvv26WOjyj3L2rB3vXTLmAHOE+f58CMxxI5jOMqcCaTnVjNsoe/f6SERKSweyiEe4CzUVsUfYPUScDu3nq8OcK4MteJTcVTeQLBBG7CGOTdT+O8N0nxk/TLDgHjrnd7jcdCyGFUirpvM9M/YYyCdkO0V2I5fOQP6o7014Mg5yNyxh3zz6P/BbMXHanzHG19+VmXwmMIOvLziMHQ6BRAbczVYCEohPI77efj2GLwi7k2AOZgl8qaa+9uDCSS1BMSFrkgpPHxjA2gj/xCcwWQKKrHX1/5jnygLJ+OgGn5+Xs5wOTrRX01LaDPVZcsG/9aSkr5q748jlbQ7Piy5fuQ+dKkRfxnKIxTjrQsqC1PGk6hpJ5OcdDB46JB13E76E4LE92pzVUXRklZo6CxH7czMxdwoDSbtazNWT+I1NoCIEhIHEvWsudUolVxQF8qwECSDzk1Ev3Qv8QkJ2NBlxYYU+1kGFzdad3J+74DSO8WdwUBSoOiAv2XAnfFSZG71LGbsfNljO/q8JWc4ZyFWATmOZ+L0ckwvGIBOCyxdtyFpH+cXBkcIoiuotUM4nGbqO/BQQmw8CM6Lz/kfGuBdpmN6u2jRcXlzINPZsCUzIsKsqlh0lIfIFUDLc++M/A6kqQCnHWWqNrKLBHCiPqgwMlp4L/+6NpmWuhZKeLV52v4Klif7PQwg3+DWXg+G6mvhvg6cG8bgI1KJ8N24kTAzs55Y3kEaYCuJACvPT/u6XDq+Xl7JiFL37VN0k7c6VEvVzexcMg84CsAJz8fqiBnV29QIJJ486OmxNpJ+HD248+jCVPEagb8O6SPsk6DKiEoUFJTZBnMx1HvD6PE/Xd+SlwLRBQezfJvKSNnXDb6geAiXqzoxBMYtwO9qy3urpzgNKW/e8u/ArdgWkyk68hQmNh+QW77EKA4qbmEh0rX+BMDAne+9+8BfdArKMAma+x29DXc5vkeiZ4wo9fjMo33W7z3wEvJwV/lJqpyNj5tkkU9lD/Q9/ZNRkoOMeAqW1STswSBGBrn0achE/OLh093acKgFXsqEWLqT43rj8mFPEfaUl2mEsH0C52f3kI0BxobCtuI3kJjj0t+qgZvRpkwNFj/fZTJ3K7FMu2i0ANsqgdO8VgWDKwzonvSrC5W3aeLgECfrlrZTj0mqXNBybytWqqD5iyffSipFzkiiaxnGjP6EgfvcQcA1bKMNjFK6wAAuBm27MdujqtTYhjCpeV7Yoo+LE8tQQqIJTcqwLoUmj7ibbnE8OwPbLy5RgkvnP8yKPb7o5x/k/VlrjKKsmyq1F9LJgJCkzeH8+XVSLj/VIw+BiJERLGkpEqqZR+70wJTFX70Zl0TDnq2hLD1jdDbgj6DyCViPbvaNZ1CK0wLuaeYsG5Ttd8i9REoBbDqM5FEb7czj2Ntk6II6Pvk1hnh7nSvQHiM6mRClI2Esx8Pk3xBcTysd0i5XtIk1MreUXLYmAYipMgJtkrbGgUuD1T+Ba7o2K2Y3gmZnYSn+qv4vlywowy8nt33JI3kPR34giOKC18mlsCVF0wYgijWRmCArjoAF/5+zhnaXsU11WKlZc1WxNjPXApYEUjQg6H8BaMgRi+z6A/hr6HqY39+newKgHKFnC3zs1T133ryoSJaNEEqy6MArhSYzwPaQZOroFsF+ZZv3jRKc+nTq4Hlo6erzezOg8UYmrtEDw52KmXIBQdk8+UMVu9mIte4FCnp7lUAiNCg2nFkEAKBKBVMn9i28WeIY2JxN4adE/bkKdADvNSq4itKMQjk/aWKYcOp8rSi3AJLLzs17gcBprKDn4gV6yq/EeZkVoDD9rONjw1BnotvakW7zZuAgM/yXM/5tHgUKP8jKnjhMOreAeobnRrWaAI5WOE4juA+MGJyv+LPWOEUNdqVzMPfR1eHjyHeAAk+hahXQSfU/4ObrxSgGOH5/jNT6gz/hLdI8t/WtMMHknV/qutp8Tu+EOEuUz9cKiVzoeQHZbR3XGfPn0AdoK6Obn8YjHC7yUzb6miNq5uTplRyQvOFglD2zJzYr6Mwi8e/6xLMStlPJJp6S33w2ZS6nyYAlJBSZ0YW8mde3n6pm05kKWJKGK9FXWpbt+VR/nVV+2+IRvsoQJqhqUsCb/RES1vbQJx8yk+zztHkRQMVsYkCNBE141/H3anSt6K9luohByv9p6SDgxCHAgTyOawgyGX9mlJy7XKFQbP7QLY+4L+krVhbCmi6iSFVIb/mLdHHjWuyeIrlqMNVO/7bWMROMF6wPwexGxjEmP75kHB8UE1Yr+t+z7vDFRwo9slPYzOm3WIcUadRXKdYl0uSSMqeELRGh6atDJbTPTJrGyK1bea++iKLfssV/Xp4+Qxw6fjeI0IEC1N/zHxq46b9hHjyeuMWbESsNq5kaLshzY7OoRgyLRCiErVF6cs0M5kG1UfoteNGBACYdJY2JuT0BWgk8kIOUwS92iqD3TiLTmYkuYTdHnr/+r5Abap+tGbg2lRnxvonT/qulGvSs7MCIRthyqW2o9Yeyc/Fx4+w/K59YH4MEKA+epHuOlpvfYuWVJmLtcFymn6JR7bbTDlNTHrlb83b7pnqN2qVeiyzbF6fLfbrQmb1as8SoTw9aUft7+LXsoK//pVsSl+fjvEwepnp4EvwdLog1Bu4hhVK2dj71bvts82Cs/AdEb2EYDVjwhXXDd/qY5EOTw+OOIniY1ZJikqi2ynkl+0VNLOfi+UO1aQkg9/KXkXTlIyewAwl1gu90O9OTBd92m7+YXYhM3Z+V8TfSLOOIAKds5/KEBwf7AGgFQQpyIN5QOEaejikDwycHkDRrztFDm5mfooL3qF8qKPNnvNvACIo7PJqy7/YdG6xhn1S2RsMPdxaOLNa51ZMUoAOu8SnvxrCx7sUCXHUfacLbcCqzdG2c16SFnzMpDONgEFAvbOXEJffzESqH0cUas5C3TCMeyNM0iSgJhsZXl/A2jnLa1ufocEdgrOoSUUEMKrVB2/qbIBvf5UZAwVEl48sA9I3o2Kn8AHepW13iI3BcB4LyRpFdtPSCVXNNKDft32sGfF/9yMFnj0I56HBopy/PspbmVxXIUYDzFrX7hI/pIBvE9HF0ebaSugqU+aDxqIs95+gIO/s+hp4MkScYN1DYDATrhxaPVmgyRGDpIEvzyMEubotfYH/9QRTvCA4jgX+RV0Ov2OahSdhrHw2t2JbnoTmuckEu2qL39CHJ0bYK4kFueWkbouHqnpymRpZf2HhvC1PJw+q4K4KjKstukKIp6rEBMMXnqGsXgGANMKe4m/r8dG5wkyaUGZRBu0Go2tD6mcZLQrH5VJpSVN/tF4Nsa+/2bXCavUnv8mRlUwI+cx9Mo9lP+q/c31TIJi5AkuWsF2hI/XTzgr3AgvG3pdHvouynYOkpHLV6DgVvUwcZ+4Yp9y0RpA7gYtvZVAN2Rd2dyhwLG1Q5youWmohlWBT5oR92jA4m+p5Hyzd/hK698CJvzvCKTViLrXWh9Q7JxK+iARQNv39GKocERqFDiWrND/MzUDeA7U52zW47y0hh9KwL7qKhPVuxMmv9vz0rCNMS+LE1fceCCwVUbuDSQLcgQ4oBYsPXTzVdfgAnFwbbGnRPPGfH90IIQrpkoyoR33aYPai6FgzSSDMzWdQTyEVqSxAJJ6UQ3AzdsvM1HvQ2w+ZJd1e0Eu+VKdGRlCHM6csj0a5V+6F8TQBf6FM689RvlcwTgrdBZuCnVYuMZnCjUH4fcLDDJ04UuasAhzV8Z0XjdU7FQxvvRkWi4N1JVWIPj9Vxv41kiPBW9RA7Z3AT8vPPleHJuQcKxJH6LqmN3R+zc+q1tIy0MZzfxNoCHXXlbsTsthU91A2D5DzaJKxjijlGqdTG1s8W3z9N4wJDJPe2yGgSS9vx3gBAoI37fO1d1Z4pyJGe5T5FgqasHoP//rw6XzNOoUmSHR8cok6clI7Drwm67wG6/5Aoz2qr1EGu3mHIgNeNRlaX4Q3j96Rvi8c9X+9/9eKAI0oNJutdaOfrvtJrQf/bzGb/ssUTgnO1SQtAuFmTckVfmHZ2nF46p3EKMme9EV8gTWur+4Q1WYp8LT8Ie54Dq0gf7tXh8Ltbka/m3v/smQCjoDVO7xeuIO5BTtGPG/r3geypeijS411D5BCyKsXmYr6uaD4X4b2Ss/KMwGvC3WRcHS6dSaEkt9E7tBjl/F0/fOebjWrMlhCBVHO3o2od8DYGqj5XkCkP1RkUng1uDrdjlkvuiRzCs130jFt6M0YY6MaY0oN9qEA3/RQOE6bpK4vBsy+yPABps9GoTeB0sTEFBtx6RCeZOuQobajbPnWph4Q9at/TB+x+YEAc0AL7pU10AkQNsRWG9B71p739d1ZZ3JiWQ4e41e7HDFQ6fm9RZMa/MWqZhaSKUw3mfUeOUv2GF6NAB+h+8nKEJQ0SXvPc6SbVEB/o45n4ndzHlV1lGyiGPXY4mAB5m3hBmecxZgAEoRUYlbMEj6QWXRYpwKE0oPgu1j0byo89nxRIHOhiXDs2Z4IM1MXyaoyZfNkTWin6bh7OE2ZpvafzVNbmuM/I254BbdxANdkix87PNNo0IojG7NjEDyfgP/GcRCsbgu6DJlcYNTNx6EZtMAW5DLxojJBbFvAHturm2E5m9EcjwIRRLypfPjAmmQ42TAquqqIdMVWkZjYRZrtP2l9sVpdl6sMvTFb16mCfl7lsOSmN3iWhrOzPtAVcJxsMTLGVKSNXUSu2a+wtJ5OJlm7/kO55VrXJ5/nz/7XQ0VVd0ubDONm9++oj0O4gkfNM+FzLCUgRySbJnmo6XIsP4wkFmBWfNZXpkpP2S4phzjQ+ArULK4tWhiIgujyOnjiHpKq1GTiEMUE0PJIpw2o+5e4HN5Vbq2ZB7qvU/MYcfYywT/d2Hjp+Zet/LrysSk1aw2KFIQqhpdAcTvZHeyOiFdFd6NV+OyRdJ619RTh40Yhxx4QPSA+bnyFmezm+p5LOLXawLwJiJ9KG4qrvwppOCtUk0jSfARquc5DoZKxMhw1GpksF963A0cygFPhVokjDokLkjGv8Xl4rufxncMtVit7nubilcUF8HNHE1EZL6lwv1yU+6Zibp63rHf7YtKWy6qdA81s3n1a2i8ifB5lWsO9p5RWULIQc/LqFCJT95KOnUHsM9g75kHn/AMwlf1SPkKQD5c0vw4Am6cFRH2m5v9AG3gHGgOKwqw5zqx2iY4sgb78cD35QvXRlPBB/hS4edjLvf7nolHWvo3w7/GagTAys3urhwhUMkxa8U2cEDNFJ1vKfrhk5KbmySJ+0fBtaH/PgNP1XMKQtMIABmSYdcIEte22+/uT6yKSkzIsiuJBAMU2LblqiX9LjTrvjTOzQcCypgoynyGzb5PX1Cf+G+pIj4llZ30Ak/CEggtzPjGkfoVWArtcC2YTGHxu/pC0pKIBLHOn1/RNnZX2rcqRX2YatQmkNlIJFFw1RIeo+uJsNf5QEfQBZxDaCk3NirgOKsmIrkQlzXbX9fje3d3v03bNpKfbI/0gPQf47fi4mO/px62TWvnJ2OQR7jkg/GehZmCLdIolBEtnRzOXjKr2zE0/H/Rhqlc+KoE9PvJlGag0GYCnvY9jW7W1q2CwhfdCiCJxzJtIQpRLYYLeWjyKkRaD/a+a9krCsfMmHvHMqQc4h5Mj2Hvwn6P0pRvvQoECUZKCdMY+B/ObrKQ8S7Uxn4Fz/LmP+ddFPjC3WKyxSFE8Fc8MQumcSD20z7G3vq5/pxlSoJdbMTvV8t4lt5R+fDVHYO3n0OtscAND+ObUPuWY+JRG2tQmmtfDOJIyLowGfygbf0Ed6PQpdE81se6DUr2U2qIG9RE68DwY5ZGAAJWGowYNpOWyrnTHtGGKmE2FqG3TFmTaz9XaFKBqC+e2nGZa/oCFg7f25VaA40SorzG4Rm9Z0A7xRmc1FgV/EKhEEyFA2iKafAaJdStg7eE801cnrPUYjkYrQyBF3ZwwG9heR3y76jLqYEILBUZuKyEQ4S7gAisMOYRCeFKJry344ctPqX2Mr8XPIgZRO33wHzKXnHagG8P4tubH0QEW8N2DmpjPsIDAWtiFenbybWMbDFiyOKTkLm/iKx6avqan0rejy4XWXLFY7Q/xBasTx/DPm82vasKnnUDfnlhPHJ0H8G8cuRUO8kqC+oWqHG/gGchucUxloUHPHoPN82vdapZMo+n9aoUGhb8IOGD11I2v0ExAIFs06V24bFRp1lGqAacwDzGuu444FAiyudKHfE9xMDCj3wmAZLYf9KYE5G8aVXbpeE3UvL4DvZ8+SKpeNxyz0O9yoqfVtmXEL5g6g+zV8pzAa+ZK6HtI7CrWKVyrGQL2j9b3Lahj1lV/1KyuUnpXh3zfYTyilkjq+lY8S0UhpoIui3QKUG9TCeKf5VOTStDcsS2MZRPPQB6m2hn1H2MMO+dEOh01HqN4bFlUJxmofDryCqWr1Gh2ffYSlMdwiSVhaou5lO3D+Fz+aH8eTXUegexZvc+ttNRkeeXy9jkbWhUsWev+H5X7cy0fTDlBwY1q1b7xBbBXBiv65kPNtP9C0xQjT/2okY/JPjOuDND42Knful/z+t/oHZfeUco37V/IvuM734oWxucnN7MxjX9n06xD9i81SzILhIGhMEA55Q9N8T+XxuXclRF5hy5VomwgaGv/OLTTjSkLPDAqLYXEkAMqAVBWe5m3U6n9Ssuumg5+GpXOZuw9HYrEVjcGqaub/hMkg9PaJM1gvA3eS+v5qvoTYanT0khgYHEtaPHhFl6FO0h+yipjSsFKdOQSWh1WSTLXkr+sesOhvY3Cu1E47V2SgZckrif2phjX8Ki4NaJ2f4a05Xx9gtKhuxwWAWU5uTc0FB1i54SLmua5uW1XX2mGb5HxZ2voUpnNnx6wVAK5R63MfBfFh1zqaBsLXhEl7rYtkOr4ElbboFAdNt/Ep7svtAjfaonz9EZK7fAA/SDKC3puhVR6fqO1OBBtUjt54/wodkItzYoKNeoVExWnVOBFG+ex7inlTk0JpCqVQlpIloCRpfouEDDuEDnn0fex/kNma8jVWn4wwwELTpt8LAcl2xopzOME1Xw62RETCVBHGFRxcbtiKfOe+z32Y88oU+oHS8S7LSZcxT2rCZEaN/HvT6y4yUGss1zzODDY5UX7mTbMZagKphEPc/sFLGEWlpz8et0lfpbpXxIBCYgbApP1rlyXburhf0D2cAUeDWrs8ddBdVbbcFCSsW0k36VkTOVAp8/ba4rlfxFe4CdOROA+TM+pEgv+et7UGo8IxBco1t0G8uKeg+Lw8Tea7qsGWKYNU+7O+tKjnpVa/bcpRJM8ZMsCc2jXoAo8YO8TDWhNsGxJGdBXUR/Z2MFwRqMvpT0NR6XO2qrVOKg8uKHU/bUtf6C16WpY6PbjMAZatUX5ZQ95+HySk3lCUE0PASZhUE0O1E09aCW60MA2m83emyBeh3gwOZizUtdHaM68rOSI3fAEcD72CdeVaY5FcYdK7uXod5UDIjG99kJlCzmm9l60UyJIZyOAbJvX6L34bnf+s8lYI+0oOLrH3YNpgqj8rmzF3R2q7O2qz5X0oA1QG2krz6e0pLb2ckOMWNE4GztFhk6Cy0FGrzcS9l3VWquQy8Lt5eMfir5eNzt4VXdSEBlmq+6lSflCOgo0peBai1dA9+RH7uzyZeQpZCRErTCdJ97x5+F6+udVq1eT3JnmosBna8wQ4KF1u9DxnJutP03cHgDQDbZzS8P6OJk/dEjqDROMyRgWGRwad9NHrBSthbIIGsScxxUd8UAOYxAz628l7VSbdi2UwrQS4vBpxkyGbS0yCOtugjIT87icZEJR9VzWYRGMR+4qoc8uOFHrFPQl6CnbOSgu32mIRkG4D3DqGCweTcLcHhWNTWLmf+TPXFxKmcqKvr7Q43zFlEYn156RfakREtwdztn7+njyJDq4PIeFzx5C6QvQAPf4tsjCL4jVGEl8bZYEkKIODPWe83OocpLiRkmsXu5Rys6zVUoLaE2fAv0LuHem+Oi5bMUL67JTvcqFPW3+bn8ZKheitR9n4f6dZD+mfF5Y01IiG1SPnRvzCO32Tsi6rJYFqOvVlQE22K6OuUe9tSkCZKmydRJdO9hXi/09922bwgJsEBDtbaY+3y8NvgPV1Ce5JUepezyXC63/dzK6/h07PYWuYPBkSqq7otaTkmf9KmMvWyOL5ka4rZlke3iYNYaH33MeWlUnohQqiYOj3nYBF9qtAfd2E4mZQ0y3K8k1Js4z/8ik5tdQZZ4pQOcG+OSdINZ6jl03XSzSXbcSlug8SL3U9/fdnX0RpnQ5IdjjpQ7sIiaMqLWn3wYI0igDVySpao1vhS+ssV6xmRyzrt2bqQ+3z6seYQM0hIzVLetdF5KvMGuhHP0tnOgd/gXilPO6aZx3sUoC4Gx1lzgw3x4W61fj5JSRBa6KnUlbkkDG97BVSJcz5m5Z2qZBVdOqBe1BO763q3+aKYxBVfs9HQ71kjC9q0iSE6LwTNBUC4V6UYMPRrkTelgey0DuLvPTQW91msZVV5pVQyTFVkk+m2AQYWk3TB0EsVt3ZBl2cP5PqlauxGv8do9YZplCWIqyBYLbi+FWRFTEXtW50XypI0IY+fpMOb8j1/9XkUjj0x+abHqtfn5X4xHppC/ae8CrRgoN7AKowGjS8ndQWbPlxg0gc/c1O35U250zl4a4Jdjm234cyWGVTKrGgxzsZxM9y7zdq/9paJE0ULPPBQho7NDrIc+MrCbdXG4HCvpkMjBFwjS6CpD0vBYpThy9UI/a0/EFMd4jTccRiXNKw6MiKZW97hSovPWyjayUJogWGFI91bXFY0DCejT/xz41ijYg0JJ9Aw7YHhPGjCoVNOmoRGCz0OvlRwp/lr8FL3gwXAqAdCcXtF3ZW9kZFnYelcMPbOycOOIJ5XnheW+36QEzheTGetQrQUtpB4yk5XWzLz7ZoIUDDl0BR/LOBch3cWkophvv6qvHRCuVzvTPWoAcuZV4QShFVoJO6Cp1b7/sbVtBgX5REduAR9ipjhpwRvmSHwwSHNOYQVfkS0a6blxlsfzUymx0otKsho55gle5oFvcqeo/DmzbwsifFqv8N44fzQsv0IeAxTL58uZKr6oKRZgn3TRYKnmINQHXKctc1y9iszIBHs/Ev/Qg9pJcKwJx0fHXC8KTfYL+4KlWwLBBGL4/VvKsuEJ9deXRqChnJ3kmVX2ih0n6KTQvFmoGIx0lAtIPsgG5TsdAxxDPEAEmgdzKFDuWyhLc9pqm1T1l44UMOmT/DMvrEdNhyhq8HpDjRU1QWTLlfE8s5k2JXzDJDZ671If0Ifmbn2Wt4rDp/O8wIxAsiXoIMPFGJP5UfLwgnaDXU2cACcZtNB4fHG66Y+7+U7ZkGgAk/M4hcCzQgfsseSTkjx9WO+75++V/y+WNYVolRnITGDk5slEUFQpB7l7ehsh7yufLmHG1QecaygqRr8KCLSV4CBZ4aAnGMAcHdGji8kBME6IyHSKbupvW+spEbT9sQW9w1iCEhFuqWAuvEz8qLBSfetr8Ou0mixC8fd2eAOfvSAgCOOEGgE3K1E5sBXREfPXaL38V+2/27QG9+aQYNa6HCm7K04gk3fv9ucow0VINqk8Ca6B+zEu+7hqqjBl8A+0fh5Jvzbdt1eDAIF9P8cgxqjRWcrnpftKXc5QRJcYby+OQT+QBq0JE6T0Xar7HG7LP1/i8v2F8bC5aORyehT5kFbvNmDLDYxwKiMHUxegI+cZ+N42OTUEP7zJx11GIVZ9DAb9Q485BvCns6HNi6mPN/4qZD2BiWxJP/d+7UEyYxA4dwlr6G4XVsTpi0Bmk973uaZqW85ik+IhhwhHwC4PaeXsr+27htQJPt5RknZwNr2g1IHaSdMtUJsmHq2TOH+xEgINlrGbbRZGWPpmSiUui9qX8/HVveQE/0snFAUTpagftH+z/wt3w6MIqj93xUJQOeIeJno4RJcCXx3sJbq4tIIuJQF3jZRsOoD6qLmnurGRZB9etR3S+l2GpTaL2JW3Ti1K+58IOWBk5ubR7HmNXUeMr/elM4ORNxywJ7nivVWal5gvfajTGOuwdvAJ8ohIgM7WpchGMSmxlIDyXsEOen0uJ+7q/cpC71zIHuUlyt3yCvAOK7ALbiAkI8UYANXjJw6Lndd8RXT2g9CTtpelbMUoDj5wJtIpCYhasjsJxDJEnlNvwqPqVVpnygnpo9Q6b2zVKLedYhCo5NlVdBsFYbzH9922RN7K6cnw9xp61wKKFBrJGvLYpzC/OkR3YkFEcmQR/wnOJaLIvaB9Es5UM34n7d/STEbmPFpRtrSIDyiK6v46amSdYYtjslrUJvtl1jEgGHIxWfHPqE+He4Gmo2A9pceMlK22SYoksAaFUY/T4J22VMgVQbZQECBMwDk5qbXExSsHREFj73vEqOfZvgG8VMiwZPbV7xOqvY4mNhBSIBiJPNcBeL3QXupofzQxMY8AHTGlJdjmtupm0rYLdZl3x7Gzav9FNU8YEmVgp4Yp3Umnoye9SOVJz4+YR0YEp75MJnwD5Jbyf3Ses4bv8lDASGTRVGJ9GwMW4MeWM7gHhJSp7iuDRJ52Nmy1i5xogmIth0SvnnMJxALRr8RJWecB73PAhgXjo4TBAKUMEVQzx8K8SUDCzlQCCYzUm4uX2c8yayyX6s9F39q/uGg3JNjwWlWCeyoKAUYG/sqoV1nP33gxNXiUC07PyryWrrEdFFg8+wFR7+vy7VCyAAWYDf/P8Nt5pWgJ/4uohkrgV+k6q/Gy7TsJxdUfoSdqIWCxCqHvZ1FpQZBJADWhQ02Vszx9sm7odE31wpdHiDh+7qRwAAviQrDa9KlQfjoCPsXwab53gE4UuONNHZpvk9PIs3Jw2Oz7557ekHcm1qwckKvVi3jcPQqcHyENYTs3kUoseRK0dhJcf2O5lDQuw4M3fgq5JcIjVu0u/zp0ZWG8L1YDqKFWQXw9fnD0lCgAngpqK4yuFaSd4wpkkEyX6youG4Mj/dL3a6+bWcW/PlosvOffE2cnKvztkE+9rUzoIL12S5yr44YUx8rbiKEjSJxYd4sNGEoQ8zv+Dpe2Urihb6/kG9tPtSxj6sPRuhTK5T/A16MjShblU+ur9or7KHYiX3rkECQNamO8lkxE2/FjlOHq5yOjQxqggSvQdgZ2UcLCKW+8naizfyT5AZY64SMqosMCe01Ped7mqaDZhaSdADTkmlkP1SEAhP2lw11Lvqumm7Uvtj8s1jrgfBNyv4B5yfZIecEUIi72YJP2aGyE/c+nk/cM6+ynm6EPSy0sCJ+5NHRRqCH+Mo/DnpVEQJ6FVC8uhUvUlMYRMqMwwcYdgHW2V+biK6Xuu6qK5pTpC96NPxGeASh/NDimtbFh1gvc3WX2E8AbXuXB0DUFz85l508YJoMxhSlWHcyn+75pS8D6QC4IU5XhpoUnRDEXpRP0reftlz1HnZ5xLcX8BHCN4PcauNigLL6AwXpojcyr6RFsvRMPlioTBcM4ZHcm74QsLC5praJ4659QwT0FnnILDL+82+Bv7WKDdkRN1uQDpk86TPl8KIhZxv9pSVclJVvImbMzhLbBo30rt/seOmyg3CLYF7+EyELwaADyWACHLlFIOMon1mzMS1LtxONlh0NeB/O6kYS2Zjg0LqDXd2ZI+Dh2q58qpND4J/87TYPxHIZDR+/gg+00dp/g02tc77VACcXPQobvsAKGxZQU3bN1ZBwVsOTy7gahWokg2H3ZaC6y+LWhmUBO4ddpuTxY3aEduQ8a5Q23lyCg0e/dlQ/dVej7klc4eZXOvcP3ZhN25hDA/LyV5nsIUOOsTrCUXfttf56HU4o1rC0dYrxIfxbARdKrm0xoqsPu6kqHCxOhLZ8XPs1nJx6q0H/0TKEcwTg7LqweunBlaQdLoj9H6AEbc6tsvGckqOgnsaW4LQllp4UO8Lwd3CclYZQdqyIjTo1sx2bH72E0t6nylNziNvb/W01cV/jBNOvSv1vHgTaoBYrao+Kig/LhhtIQh6+MUKPOGbFytyq5ts2WVLaHRuNB5AKAcBcha0BgcLo7Uq3dvQru88DCO979BnWHZqhQ1F8DihZa5g9vdt58PCFb6mBDXU287GpGUcFKrXd8+7jXYivmLEq8f0YNuvfY9N+kfb87rS187Higps08wGcJnfmCgUG67IgWaOdrLVfUxciomDkCuU+4S/SOso6VnejIxAaGHMWbyn7O18r9ElqUk//W1Dl8Y5cG+BDvFrpReesANCmCdEfFldDqsTlcRTi+bBhLmuV9wimMRqsQ/w0mELkAonAd+qbXYlWFqVZ8k+J8+vh4LVZHlJnq29+kwKygJ7hb/mFzSxZMgLyViYg31SsiNAE3PBi+OnMvRAG3KxKAFTD7GZrIHQ690A9ix6ILNofMhe9/+ipcEjY2VP8+HKKr8hSkGH5H/fv7lx4vAcYEY0HDfNvJTPau+qGv2nlw/IFzsaaoQ0UvwNXUa8ePxFg/whSoIOMZsp6KhvWMiwAq0VyfVfa1sWx+BrjyzG7hxgOAf9h8bXz/cgpAnI2gtNqBo7wdph/4kzDpMIp9YXthWnN3r44JiSCCbVRGQl8lKvoEj40TOw6RRjPJBfYXH/2iNaJsGGtVzYoqEEO1YS0u98SHva2jcA1xAFYzgjCPkXy2EZKONoKszpr5Nm+VdPbYSeZqKaY9hWLGOae7mj3acLG8fpJPf3jL+ZSKLn6pcaSu3E5euH9jsHCJgikCSmVvww78VdG8eCN4V0SBq6wB2PgaVlasIi9R9Pd2PI5Aq4LUYMM6fD3c5eFoM6rT1wRUYoqhdmDgR4tB6nBweSbSW6kg2ryDT4g+zzAdqoCe6aVPe/tQ4rkGKvEZ/XFUEWp4G+EcB+V5YQfnPZW9cZFVQJnhDM2yXhmrbwgJeIMqdqNV5C9qIvDNsiUppCYmx0bturnqYGzAFnX8kJCsCqFMCM4uH/yZugezXSqaJNixo4sU+6za4pzdazoV9PEl6Jj2BGO6cvKJkcz+bnZUJIxjrVbU2XlikwxRYZzyuIGnRYnedevO1j1uU6RvoPkA6qn2ym41qUXnI+PlcSQQeQc1pt5vjSXBpH5pNb9JxkYJCjxCO8vU9W/nqucmM+34txHbjQA0R1F+q+RcE24pYin4V4gsqVCzblxFAsrmHcRk2evzzP2fPS4/JIvoqe8O2fViH9C2+494q9r1e/DQHuPLMqX6L1/QKpflpcak0fmcL7EmD8ddcZIp6IgkEh9auNIGAOLfDvDJd1+uI+3J+fLb/EW5fkX2/3iN1c/Dn0MDTDDAG7mhYI7r1MJCFGnFnwJ/WLj45WUKKxZTSm5Uk+6Q9Km0/QAMDrgGVzVVRdnrsrTi6yroGDQTVTjfqYIdmF+wTDrt8t1Z1zPG/5Q5OkxVUF466MAWhDa6HlILFOwiuVjPGDYXS9UbsNaXSgzZRIEIUCr+ZKa+HP0Ho1BhzP5HtekAWvWZSFjPagpekzGYf8JB7h+p+SE6HE5Lf9GvyhH6UfhN/PxpOYELL+JkoggycPXYl1V4s4K3RBOpN78QHb6FtrZv8WCfIfi7JKXWxwi35Dre9WH6k/uaBBrEqy49lYu6QMSvAD0qwiGnJUCet9lBg2uqNOgHq3kR9cAlxczRGqcWwUFVx/UmU5g/O+j/ij0cAiNaYXuPZrt8QMa3TRsJe4ekRHUDztyzP/ZpZCC9FOJrNZV8oD2jWtbkC9ruh5/3+Q5pgFIcFc2lgOdGYgyiNg2oZq348HV/gVNMbXtEsh/CNhjdF00ZF+hUVvD1oozFLuUpk+paCZjokauSQspubU1QUNNxWJmj8faY7pynoZgx1omhfQsVr82pUrJ6vvrpdJztLXZkvSCA38Vn14aBu9g5oIRto+9Gzxoy+C3eTf72Jt//ct3X47MCeKOXyE2Py4Ib7haBGmE/TW1NgZ+cIrrMpfCR0GHS9Y1YZQlQQMGl4YQofWYlRS4xATwTVdvLYdkPyNoVuRiwZ2fsz40FQuej96hVGCZtOA13o6GizJz2tRpB1pt1Mr09iNipScc1+fSJP+b16qDcD/cJJIkpjXsMCpvzopwseGAowaYE7gGznaaOoyr63NZKzUuPLW2xKcJHd/1aDeHZ1itHbUvwMAbfbIYB9ncPupfY59HUAa+it+snQ1t+a6yXfxEQAHeF74j/nSRr9G+G4ybZsW4vfXdY2IATuNc9+oUiNCgrfVV+9UBd5q6H71W7Rp7b4iMa6TfPW/Qo5cRekbUzxv+Au4MthgcwQNiX/NyuNAkR8oTWss9hhsE+T50aXUms43bgjSyt6qE/gsBWA+bgzri3hjY7Fa4+KQGwzlAaxKE3QkkXV9G6hbovc0SnuxMmCReig+womsXe3WPeMz5IxM2TRtz2nBvpGMcAHzxHMaCdfowMQIoA2xU/i3YM0l0z49ZIahSVEyjfOabPx/1hjSDTJXW6WdmZc2eZW8w9w5fazn8qvJB9MYMvCxpzAlXZOG0Xwj7LLbFRjybsLcxGk2O+QkHwDVMPqID6SQeckBMzD69L7kJUr29pFcE326nRA/UkLqUgiyUzoNXv3Pq47VCPuy4OG8V7V/aHiFb45HmBHHBu9g8UNHNNkipf6juGzyGJVEIa03ul0GGZwk3bGwdTZnhf4hApiCIxdg6D4ZP0mN3D+rXTnl41fD6fw5aR0izUMGzKdkHN8AN0v/VWrRClY0t4EBGBIDFmgEoPahuN68pyaUhhyKyQZ2Iw899ceSJjFpgKaz4avmav+0l6DZe1hOnYH0nsNNWIZ0ch01n1qcX0Hq0ijwxBmMzTjuIqrLT/kzoZxLESGFtTfgKFJ+dP7bOpTk8qsF6eoA4kQYMEp6faqAREpb9CMbfTw0zB5W7IZJ+8lV25xbtLZPsG7SYjpHNJUpQmNNhFgLfeWZ6wiVpXdJ2+dPTma+dPrjhvHOvXVYMLc9jCPtHqhQFWL+n8CaxRBUbWW0XSYPsjONrrxGJ964uszZxi6G6l1rlWxgdIpiRQngAaJTNbsz9ZMtynVRqPjyrKkfFI5Ffd1kfwF/NKPVhv/BOtKqwJpt1tpigz/xefpDOU7BHfkIybg0VDV33+aNaAgjTIVetAnOnrPqM2cfz2DN+fA+J21BTeeuQ6EXzK/KD+80DfM+o1D/BrL3qlwRqulwSn6w40gIF0rxT5eT+RfcObfu1lur6SkQIX0zuEKcDcFGn4DGpbr3D9mZzCLXVKnfolRuZ+3cPfTZ2wA/GXcwye+nYrA4R3n98JQ1MSwvSsb1HWQVvrGioL1pLE+c1p7qyzDYTNgY3wuXUqA81Q4IF9KX3ixiSfdLtqI9d5hnlucUSqWsWbeQA05RSupd6vVaF89MJdBYJxOdrzSqMA8dpZEP09noSz3oQSMcP6BiKcDQVZwUS50KlNCMDyTTABiSTcs4j4hyGe2vbjXxHEhKKE6jFhDjzU/ZsQm6EnE3Dc0bcTemMT0zVeIitPtxrsOmw8P4+zOgbc++MtS3CRUFfw3xXIX4WpmXbifH5b3nxVIugqMMHuCxXNGWQkURMEKhHhUYFl2M8unLubX1EoJwwjA7MLhhmpigYlk3AC76dPbRfW/IUb5QNg56XzjlGznhZrLR7DnGP00hnLnhr0XxhVddDPhyGSyDB1mO9ysdNHPqy1uyovkfDfVXq5aX6jQRDhVi1iVNe3DJiR9TZOZ3kzEGju2g4ZJV33tBljt9+gV1K7qVhOm1Rix8cKr72eBI32i6Xj8VDdW6RJ0T1zJZETgQ1yqdxf2enKeUFV7a7T4pCPWrfFHOqnWSWYm36mn7rq7QHQO/2FLIGlrVVDlr6tL7X/0IMCW6SAdJo5OWxwdXauD/Ea2Hcl3YePbXrd3cyR/43S9qe2zY92BFejUQGQGNV9aL9NuedcX2MCIqck8TiP29yLbaY/4pINb4/RKkTBNIQVn89UPz4uN9ym008iDVJlhbcfXfDieOtvT+A/e8dM11jLC3ZcU9bEiKXmeFjUCllQK+1zgHoKGQKYKp8MIcIkt7Fjxjv4ZTgMaoQ0DZ9R2hRzeSMDe848hpvWazZXNFf4BnRGIb/vD9LN2MqUNCY2VzDD1LzuKkmp611krdzuheCrSApBBwoz4ztUYCOO5jsGA1s8mzPMoXA7SBFE1sqkjgDgpQxylCD/oLaKtO6VtDrmF+cCMCVS05P/mFx22K5enEbZz86dTgvU+YAJLiYwDiTTrBiwhTAkrXvsPiNaHFL9vMO5RU5reu/YvrI86E71ggh2tDqwSL+Des1Or/55zPb0XBSGK2Kwb9p2K77Sb8FxXyQwfIV+xHbBrlVmQb2KgRz1HHRqVaiAx7YrIKPW/G/HuEXqY7qXDR5P1S/MBDdsGRvUZNxWx4bg/7rTAIdhd9+88/K7yPlOQrhQszeUh0kGN0AbDBqh7jp7/VoUSutWlLN0X3TxgzxOGDtzH8MHPTnVkB9RPlt92srfCUrdb1Joc1SuofbuhxhTju7ih9+dni9gOdyeb6pVOOE8VVCgFM5rrbSspmkywgfJSU3+kH2EiYyngXavV6ar9LyoDpP7MWxwjDjVRPRKVBybc42vhoye7SQA7a5wvamVzHSc4+dIS1dX8moeRY5FsMbopPfGg5YYyYCVdR8Q12DLE4GNXiHKQ26TUFA3YKy98Yjo42vqy9r+VINcwDrGEoNKMvl594JQKxb43qFQGpOX8ifw1juYPwDOcw6LHYAuzsa1W4qAtY2693s00Vurr/CDC/sHBVcVGGlza6LZbdC9tCx+bav2z07md9bxKXGf9cmbUoyp3raKHOHojew26av74l3eBjqy70E2Mpeivn8NvtsrFhBYZzTXkDVI7R+En37JmWptuU5+hVZ0E7fQstFThxWrgFJgujz3q3+5w3F8gsALzRebwtEJ/4a9i2CgNe+iJh85+1bfZ1L5n0jjf7D4oEcF14WmjJctnKOrevRpr2ln5ZKg7OH9FlP6jAzMMgm1VrHQnz6fXUPA2ZnmjuSVtXFunB9RbiXg9GiqfEfwbrWQjUQ87qK0Yur04busuTdo6Nc1E9SpXzrud+Z3b/P56LJN9fZkm2FTCRL3gH0083vG19pOzFmZUe4zQ5PUibYA6c71QvfKoLpnJbesdNqqiaUuRihSyU8yv6/+zt7JoPUVzRKeLJwwAIxBelbyeS30MzVf5GR1rGU/Bi/anUGsV2cZU9t8TwJrQOQ2QmeEF6PB0WN6RqSCfKO6BXmW92mLz+Sniwy17OGi5EHiI4qSKfZNoHkyXnWXezJWqM11uU9KvygN0TuRfdoIdI4w1OJgGXaa/BRaXCAuhmg+kVxTbUPBbW25K6JRU90+7mWMPnYzdcYe1k2TFLWyZuvsBmnT6nYJntNZ01jAUjQMJW7W2sfLHmCu81hUsUXo/pBJy/O0jewr5g/vvG1++J7Zs+sgC3vnKZVOUQ2PzQcKK9esAfT6UqCAHw+T0m6YPpRTMKgk8XeVp8Mfru9QWxha2Ffs09w9DGV2Z+aQg2tK0VdkT7Ed+SREhaWNveRA5heoIDd+jJ5vN20ZB3MKNwximxCN9HFrjZfJzrI3zht+GnSRqY5DHzhFKpsOA2gOjLZCRIwgP4WKxl9NDfIJ3PkaM+gW4DRobDxfI+iOy8wxtwvzaAQv+03wQ7MVW8Xlgv/OfGLL7AmeZ67G5zz+piNGzFAjpc6lvoMU+Q+8ZYCOJyesNX1VFnCLmpNekXgI1zZMmineAMq8f6vaARC40fZ7iSbktwwTx7YCsJPT2xpiYPMtZuLznqJ/IHfARapqEEC4w+72Xr360XZ1oap324XFUNr9yozek/JxLThndEBanV9oxAJllUalMFPcD3QCyXEAQ0CkraEEJtI+YH7n4HXe0dtUdaT/eT2CbK1UEjkhn1WoJ8pid6xgQGXKmXHUPFSVV4m4h8iMwq6i13/J5pe2wUnzQHmXrGdBRKngeotySIjAtkCFRkN8qbGz36446NBxhcNTOJjGgmreHwprS7rIm8Ea5BMs7VP/3uDiMCRqKAJHV4WiomXTyLXF5u09o7+POJNGBvbbg9c/FW5kII/i8rPatwE6Y0U2j0QbvNpmV3NUSJdjjgpIYiwGprEcNBfbqDpAtzcyxsZre5+V2XmUwHzxccVI1ae6akftNzzwmwhtYoQkmRTqjhnNsLoEZqkNdnmv9tFnaT2iA5HGnhuFyaMnNZkAEfLa/eHbqWFQthB6yOXiNDNcyby8ufdIG7PyCNVqAJCv5hygNNpHxij9Ga5Ogk4bLNSN+lOGK+lV7PcH7SsSSz1DgdKgwxixv6hfYgtnf5GxQSUO1kb5D1aTaNPFDhAjkKcUXYiOZyZSI1FZNY8Tf/1WR2oXhjMQROKOXLcs2uPjDJ37nKxO1lwgMEXRvAeSxrv0sqgaOsAu1UitNtHPcaSST+QrdluI02w62HbZsr/HvhzdmsOF5R0QuG/h2VD62EhCObykhRKsWwrxAzMQY2mvycEalqhHFlv3gQT6PGLsBnDDKE4cIgAcCHEEcJr1BxCl6j1Z8VOhUMZEwqDVL3Kiql+uur2plw+bgKEFXYNARyZV1YBqupCai278Ei260gNOP6/AIbnu7QHX67iN7xDpSfxN0DxDg/cIwexI98PNdN35KDP8bQOsGnR2EI8Ay4gSR3qHrbRBPo+JI1j2BExlc+ZgKnwZsJSLczldsTayj1NASzJSAEPoajMgr40SAShEYMMrSQJshLxu0SJGnZ+Fqx9UyFuZG6ya0jS0ah1oo/5GNcApSmylvS4sOueDlm8TJMtByzc805KwZ+LOX6/uidxegxZJeR0jr2q6SV2Mb5wTqBiwerJCdG82wstJmXkoIAYaHJQz8W0MBARuve+x6S37CqmwmAfgwZsWgX54v+OIXdwzuVZsqvabVCHoYiMs+npp7TX25VLYLX+k4BnX7vXv5QlObb9+GrRNjr2/xkMFQ1tWCjUkzDN+fmRQ+swXbiRBbw1P9udy7XUxpqwjfBErJeJTDIONOWZp3s8dGcrhYt5Pq72oCmZ4IwqHCmtWV7Yo7Epn+Z8qqePPHWu5f7llwCokNRuSDpx9z0JVjxg7w8UC9Z3wNFax4GG+11GoRsU+BjrZultJs1cMUwmci35tmvcXeDb1BViTeMOV9fcPSY70LG5BNZlzJkODy2T8jAdE3B8ktTTINpy3hVE0R6p5TLikS/JCsMi1xSiHp8IC3CWkbxh744ELqSzGNQLYC6myl8vLppb2e5DTUWiIUOmHXsZQqUSpjmHZTmMP5X2tIO3XsIwToAK4zreet+JfkBC+44XiVX5DqSczNMWkDIKDydZfIiHuaqsCPplovmuzNI3nOt5UGynrBbUxVa6qJv6CFfKCfa2zmUMCogmdYWXoaFv9p0MBR1qSk53ZrwXCjL7oxOXlvA06plRoiHqldSK3cYNlpEUl770/a0neSZQqD2BzmMLUEhGoNJqQtdlll3gmmbTo5rYXgYc8C9QpmkMh1bUwboBpShWg9Syob1fQT3Ju7tbjdpPJMrQTXujdrqViOBE+xmRAIhK4ezmWGBqT0aeiEWjB9D+3Dc4nYgpGrTQ1SELXFaBQaloJqLAJwMXIUKHrY+HsuaaaiUwzbj9bKpP4tIuLf7iXkvtF+sWJ8/hWCjJBYYXFFQ+5asvJWGQD+4RR1wGk1GlStzYz9iFXtKwkgYbE0CZZ6kQH2mfDxZkjiiFx/HSj2/sVuZtpZEwNx2vjH0aOSSooJOc7L/5+hhJKXklQQayrPfx/bKcfx/rtQXta4wp/HbnUBYQQXhYICEAozZwi7+k8fc/PC5367LQ2vpTSC+Kf0Nsjkk7aWasR9VsOVxdokYFqXnSjNqH0FHCXPax8spp/silPaPiPKXUOrzoXpHU6BTSZyB5p+ozJhvX5j1DiVbVAkAnF6V3XntioLKX/RC9+l3VbaOSD6vnEzJ8DjTIpWFQ08vjOEQqwQ3h2DGY5z7gh32LSx2nvm2DU9Jl8xkCJBNEoL457BXx2MA2NKLzRC9KjD5zxf31oaXpQZByc5bo6+YfbTelvfJC3ImDbxI+xP+6IECGI5f6Yzg7zT9zBzOAa+GAlhrzEgHKSMixxHEdrivqMcAui/WykhTJNJid99QkyjBKoZp3skxutp8307S64QzSYLjeXAq39uR6zSYzMcUGkrA6i4Az60zppcGujaxRfhR0kQBHy7dsOlJrNTr+u6FbyOyvx7Th9dWdyFXw+ejOaL718nxE1k0kxubjFPR/ja0Bk7UfXFZrwuR3o71uQxIzlLLwP+0yUQhASwitsKusKm1TMjU4Zu96nfdohhO7v2SoI3t8uD0SCm1oI/Xsog3qPbDurEVer2LCz8OM69uuHYm2ntNchqgRptbMQUstePDbPT0LbNPqZ0exxQI2SZaAw2Mq4O2afQ9lrcJYrehZdohpRxnyjteN1lnG6hVIKwA1FzxWZhDr8KVUw3WJSJFqINxv+CdfPM82D+/0ITkZlttPnCNXngpmahJ4ANAJ9EeyoWvRg8oaSZFaBbEDKA4o9iub0ps40MwSWof4OGck/Bmr+cZULQaHOBKm2Ci9F4Qviq4WhZkGdqOQFDpWYcw0pX+3Xx8SO/6XtuLQY9DqdV/zg3zelWgItoPzbSULaar/kmEVjYSuPkUG18YKSbNP4lrh2x/Gek6vv557P+sVotNvwjeoAzGS1/x7mncN/OsE3t5GDIjziYcamDXMfc6TfBvMghdqtDvUQzQVtA65up6XrHXYeloWzsIQQCysL88pYhtMYEupgJQFrAh05yqi3dz/PWhUIUbMAMLDwr2BjEZoa/plynSZjjWIKCD8D9wc9dszh9Yf24CeUj99Yzz7Z8S2ndeV78aExWUR8cMgobZu3JGkmBQZZ6q6KNmyRm0MmL/5iZkHi5/YKBccyhXyN+XusZnB7+vc6hnSHTpH7aquW2yNrY4jSMw71pB2gK2tPt0eOU5oOUJVUj3NOGc0av1LH8Td0DNCeHYLSNAw4FvjqorLcQt0NwPe4j+VkPKXu9LRoWgkUVVX1Y3SlsDDDG925ss2vNHmEU0nKv2q72dikYWYdK/Fj1QQNbBFPxmX3x8LGEp81wMo6znfwKO8HF51qrwlvY3e3qZx2SqqTcyjLxzm1NxlSCdx0uXw+6wA3iBPjMD9dcn9HEq8FLEXSdZ93RmsI2th0DNBdtMVR493rBOsVX4ekvTz6x8Ek2kvjHQMVXVOkn3qWi1TL2GlmbApL/pzsa/U2qyG9XVcpg3qOXRJU10cGqjYZlMBgEWm26gclUDiYtsWV/WKZGNkXAVpiZ2bPw2/19Tnbk8Ko12sNvbKJ+Lw+Ht0ChgPiLIytwCesVmTZDwcog1LL4NJvWz/ScMtu/GRcI/dcjeaGsz/AjTNtYGjD8keLwwhz+pPQSuFkHoS31PTeCCFaKd78n2T1DRkeljJReLN5o+kl6FogNVEyWcba+knMD/mcchPSux0Q4M9pY/0Zt5TxSLyUHBAN7+vTpIP/ToAkT0GrD/lllQv3TEl1aCOkcaJg31nCmfe9+AMryL5ekx83MKGxQ21LNg9VwV6RlmISYJbQlz5RNI7gdfegRXTLooNgJoHoAule+mFcS4pO3juBih7TU4SZsfrY4UW9UQ/jyZtrE+MMe3db/ChID+Ihy/uRMH6y8TLGlJNMi+zUmuoKIVcrBk5hrXUXTJUAge4J/kcMwuPIyQ/CCO53kZk/enHBd/aCyCruBlgJlxG82SkCt3gyClodZtW3NZ1fuEhM4JMLCJUQR5QbGPTbkmSx58Ew0nnCJxfpdymesWbteCYwya/HINB6g0XQ3KcIlWFHy7Srq6zQkJPTkrN7cg/whfVlq9WULZRudm5w2kCRnOxpFM/E0AQLeW0wSSAY9BiJa8IAzk4OmAyvp0BXy2ZZGbdcsw48gfvN4fOgU3T18csjYv1sxTkbQBlNRDDFHme1/xDVbWNlxjjXiKpDBbIF6LOAZ8GyyZptp7cypW5nukDR0J8n79meoJNWrme6Ju+RIKkR9A4nUt3sUIapNJJiTNQGEdEvchFJM2uWYwMm4Vp+VQCv5mleUQunMhxBiyhkJ+UfA/Vc4y8H07pbIKSve39jgKoXiWMaMihflX49GtmHrkTkTn/Qj6yHWBMfEV4HEQFOPp/36rKDLHs5J1IgnCddLfuto4MuTtHpQyp4Y8sos+b6G7S3FICvFniWLjtlTCMBZ8mpm1UKJXXrEZFdUpbUljDnLaL3xu5+DITsUM9SUCzWNdZn4asAxfpKOa2GFuQkxbkOlY3SmH/8lWugCtbQbxRxtGU6RLz2QSePwNW1Aw4M+b6o7Lx9sfLm5J1J5i0XsENvqIm47XDN4s7Q9buwKbrVw9vM2Xq0naiydjOAWPcWftPQmEjh/7Zwf28S+6arrEMO/7y9wC8PiZF39vDAHVpryxhVuf9vkUvze1PIb61nqiavhMyiqjypgZDGhmoE8kT10aj4r++kIzYNBP9DvbcLTXpyN6BqdresexFtNTW2BhhskgXD+Eziljiy6dcfDPktsduu5/HniOQjPMDUK3cVKYPkpHwuT/cUnsb0AihO5O69pdd/JRdLljSigt31SQgdiTi2Xzs1PkCbnvHM61PdzRmUkfO1F2xZwargLrKl+qPq03ULu0RSIZbEfqPCIoapcU2VfqmuZKWRF8/7X3SNL0JwgDJM8xYORkNhtlcefXBSPStK8/vIyNoNHSnTe0GT7DKS34lkzmELBPi6NpON0avYLQLkkFh0GHvB/BvU1dbCgxNxgnX6dwdyAsI9i5aImPRiJRAk6mY4kE1UMnW/IkxjnFq04Ksnn3liBPQ5yxoTdYwkD4yJjpBnJq0h2HlfXTH43kSnFscrjG0m25FzxgD9O+B8vpAdXAa5LfVzm2yTtuzqU04XpcgVxJQo4691bA0tCN7z2MyqiJdS6Vks5vPyQkJiQa49cizACQwtZbZuObsrzUvvTKD8Y/4UvKE0OYb5mqYZ4XhUDpAPUWGg7SErTOfEAvhH/Vg57/J+iRWKCxteJ5Tuq/ijS8i2FxKCXkpGG1kOxn/0WKNDjdUZmwQsbo9Vus2mw9OoQ8//BzXwMMuoTisHw3gFzTTZpm8prhaOlkaUC6FEu0HKGK/lzFLufQvIWiXceqcmay5MdrQuBdJZJVu5eWeHaZVHs5p7o+uokoHaZnPTv18dEHNlYrsPpF6jhs1M9NXaDWaPmLWDmUDTgrf5X1Bvybas8vtBDpVeVsHarf3Xw8xRbYNSRaut0BCxS8OttRwMW7Mzq2iVRyu880b99pAEdTKxv2T/QbL2J6QvbmC+wPVvSAW/1Pe+I+jERXHq5+9EnWvnJ4g8oAHkJ1H+FFI3gvkpstIlBmKVjk/wlsQAc2KOlHpbW3PgNspn+9f6IeUZ3iqmeEMjycxdkO4FtWIZLKRoUT4jRjwO1zP9SM3N1cerIXRoyzSkUa5JM6R82Ab45dKkq4lb3T5Zn/NfiacMC5Q3zO5UZnf8+S28JjdvfgtRna5aCO/KYsyQacQrQ6niQVGNigDTziFcaqq19ZIfqV99lwc2SRRC8YHCIziho+oE2DcLhKwM1R5DhkNkMhp9aYod6QeIWB/6gD0SZcuWCNF+4QmKxET3JMZrwc8RF/TxhxJMPDl1sTdLFisGFGtJ/gDuLKJM1Yl90mWxUKJ2RgY9/+Kqdbx/O0YSLxjd1gYAmAg2UD4IvkORTkkBCnijpsogCbiZne9KtttwXDsIk5td2k2J6SCasqNluQ4VwBdPLCHJ1TDl2Zhs0ACywPfhzsJorLnxMEzVekb4E6ScqI+plFRps3Z7U2K/UxQOTFcPZLFKESkyjG/s6B9X/lH1PboDtAowKrvoKaX+be4z+fZU4IAIsVm1Uup8ei9SzcwxMZlExhfTp6hxanB0Ztgo8pNfvQHsxLDB4hoovERu3tCOvV+xPScnYTbHbY19ffMZutw7oPWG0lWBJyIgxpzfx32XTqtp0Q6j3vqeLwhXpJCk+sjNqki+BUSyeEc54Opbljq+WXiZ50vQqrTnECj7Sy8xnXTaEZZvpmGaLC3HuelqNf2olYI9gmne/iEoHNbvsNMMyQBZdzidDVqVszY+gPjQh7SA1FhmAXpPY6BcxJL0EIHQnfPCkNp5od/9uaNuyxuWvaCgrPDtWDCsLMSIcHNHm+pYszLuKSlb58ekEWZaI8qYu9bkjVT9BiHCD2Wff5t+fk6xBLhLWUcYIUccA0omsl8oAqPLylNujihXqpcMyYnSyhFRxKdl47IsPqQJR4adVvZjLFNpzdMrHrEwy3t4nBJ1YlFltqByEyA3PoP2zBaOEfaoQFDIZT59l/mg3vHdIWars9tK/j/96jBgRknkpddQxxset6cS/Dqc2r3z3Tdoh678bYYKulvDw9kpyzCH6uuw/PakDMZM1YP0L9SW47vjPPSXU4IWz0pHH+qUF1b1j4HMwSYI1F7pD66JkXSQI90ALWafE6gb1QGc2KGsvKz+BIgiHLqLuYf2ziDDCx1An0msKkWuwcKRPKJo6TpkecwG+zZxseOrYTjhmRj8jvWB2fPPUrheTSgwEzEV3Oikcp13N+oReD8ruxw86EYMH9fy9T17TSwNgi3M5JApngc+ld+LvGkMydTPq/xM4d3StNTvyLvDpNfiLHVIArrd/wIVeb58EVz6nle+Dk6Kq8ysDh1N2yFmmGLwYiHNFG2vlg5GdNvyNvQ6SLSWB927JZIcgR39YN/0hAzSbQogNp6e/ARhzAUx5upGAShXCtu54zclkWvuEBImThMoMYW3GcYt3PpqXwamZ43v1zsBb8tbxuqWghOUekBz1ZKo2yCFYfU8hNjKFNw11Kuna+FwsbV86guoU8VLVxrmFAhJ6TYRpXesdFdJ+JJdglcVd1D0dKEEJ5CCZBBOd/qzh4fJ3AJU5euFH6UlbxitROLXZ4r7c2eLULx3wFZvKKiFJXIXNb2XlvVDvRuSpdKsz9/ghmtZ+taNvApJdTCNEjguxxpo9fol8Zmsh2boIZ8UTcw7cpPzRI4fYKHM+1HKtdI0wAIhnp3kcKedUpVn/8vWFFO9k2Tj7wcXo6nR4P/rPl1AbBhxyHzdBi8iM8XbRBbT7h8KIUi3k0VNicizAOa03SI6fvVVb+Be0WpqMo5YGa5zES85tUI4A3VZxsrPCU4a1a5c8iIWI39ko/0c/pvFzdTlKBoNNYUY2oCsh2ViUfiYfE78rP/d330eTWdEJuGAYgQV+4d+hnr24D6kBeSxQmZ8nnx6RXml6lun7n6fBH9LiK7rkwOR8eCc8JkAkKvPja3r6UQUrqAiek/163ZLPXc1mAMPZOuN0Fbxg9GNI65tvjO5k1Wa+gC4S6kG/DjTqbDWomNTMXNHJ5Q6Xkjz4GBGz1qh836yvHQnkl6s09GRx5O++TSNBtxyavBu7YHL6Owz4O8zQz4DTNE6JanQYcentm4U9UQwZeuQKOD6Cy7JQkLUYhs6sIrtEeP5Pk0ye73y5fMPZxuG3OSb/fjTa3Gj0Lni8KPen3Bn1V6FVUbomVCNbAl6WEEHMnhxvwyUZV903gPj2XeU+6exdX/yrQ9hRiWEI/IigzmxpK/I/kiireelYriPLqXIlRidqGj2WQVkxWuDE5q8wne+dVeHbNws+JAMXdapPhVoxm/ZrqcuzG7WVhg869jNTCCv13j1xmXNShKqr7jSxwAO+nsvDAob/O+idBMp9YOagWZJzNEZ/P1X2+IopU0s64rUNQvhnmbPny3cJWWM/yiESaAdS5OCWaZn9CDK41gAX7bV9LMUiLcZvH/l+ppg+6NGME9ccGMB7l2jgvn2qHZgaAOOB4Xd3JOe2gErqoVnbsc7lcuEp4LXQyF0JySjuRW5f0VFEkmtv945q9iWAKw7DRD1TqS70bGiwG83Q7++2W4u5IRdmnAF4oVzyyX+WbrhbL/ykq0K4W9B7RMQZG7qcNYDzdBZKIFh/Cs46unvBJ4cdwvhIvwG/D2L9WXb4jA6QvGrbteU7EwX9rQkf6Az4y65VKgrrZgAVB0qWL9MjP/ovCUPQ828X0C//dLeSK/QIuqLLvqAb25pztt5/+5M0sBeydjikK9otITOUJhHny/zM/eNBC+vrKcM1/BsjdmVOzlVkFgiICWJ29lCAFMAM9CfthjjcNtEktyehgN8WHLL1gqjq7efPeF13ebcLMHl4uoV8ZTHYqRlvXgjpoYtBEB8oCfsSeVIcuOoaFZ5HK2FaR73A7lGLl7/1CQlLgeEbrhipsq9Tv9JAHn6MwhGh2EbIN64zoISKYUzKJiTbjx8+uzJCLsPa29E80amDZb5G79LtQR43QgvwlEAsSN6xJF0+WOdo2SwhoUBDzqx1ZIPHHtp4lrojQIrWY4E9uvdcmQfK3oM2FT8p6p4KiFLWMmxmbFLxV9zZx8DG5kscbit6l6AloIE7fVjofR4Vp1X+KTC7V17cO/IdQXyOHfogH0Nqm1PV/Gwea+GRouuLl7RbxeR8PDu+xxz6ZzRHr3pJRnTQDqO68BrkSVSVsvqqZZcTSMvfZdSuxdj4T6vBCNxsDZrbntKzbSGHrlI/LUDMDshn3wnDe9LIYgedx9IeDZ3spSVnIbE+avUHuzg+xxnhwvYTjEWoVsFoLRdS5wSUKPZn4aqbHsYManFJVqOuWufHfqIMtgwRtpbIj1mw/m86O0P9Pan7BNgDDDpo4pttYeBxIN8bbsxOJnH2kfk0tmpqz2CDfjqI3pKFk1JokWpwg+F++zGEzmznJgGQ2N84IFLRZ/QzwgMLclWcxQp6KkSUFONVYUG1ZEzBoyEXdjSOcWoFuza7GzESN+XalPxs/U6RS/xPg1MksvpJnEkXhxXoyn1Db8mxc+NCTzyRuGOyKzF8H+qp+WBw4sdTYntRWsIeK9yJkOZ0qOXMF8F5tPPn/q6hjYGs7ywF4wvd+h6iXZ1YKbl4qsAbWzk/6RNWOvvt9Ytu1Yh0cGY2iHTpXmtZ50gJIIKkK+MnEWI6tkwK57HUeL8HRMv9ZkHQCpFL1+hHzv7mZKmG5yZS7iF9Ca+N65rJ9OLn9vmwnOefs0icHNstTRGIOlWcXol/WoBJ7cYiPLn/Gv/TAIHiqG84Bx1kBxHsR/9FCGQxKmMc523yUMoPCSm57TcSjFWQ5/QTLiFlIKMLXc99qowWhISGFmjKOLLjY+Pk+YDqyvwTr6NXgHznnTOOFi9rVGYHjfmfr/jluBEB6Qv9Xn7juNl3KYe7OhYwMWxiHsuDmzSrc8QiUSnQNIgJr6d/zp+JiL74p+hgOBv4CLsBccE6u4mcuc04tsB4GMV/C8wVSKNu0Sw1FKmoX57HhUU8B47aXTGrqd8vK85RabKteyD7dsqcv3vI0kRCI3h1gUCmlieOADqO9RNtInv7rvZrVpVcOkqKfC4uJ2+XW3qFhLDWBlboKbaATGqcH1aUJ1iq3DAo7M9mSMlWh5PPEmmjuqSANv6P/RaAoXYczuUchEuAwrubVtMUEbKBoWw1kJOzF0U+ehKJfRHTlrrRxgEr7v6+idzAe/S4fZdYfMZhXFBToKgtxS6HVHzmRNWb/7LXnjINqPRhp0Rvb9WhMgsP6JYInHSdY5fRurrwNkg59YJt8NuSTCFLhGLWDcydnNoXS57/DBylZkMG6itESbAhP1vG8NBzEm/Q4XkRQEytaG5xBcdNnvarhQQVMDtV9bWKKAf/SvikCApppL7QVk/0cZkApHJhfOWjyuJ5+kWxSruu8Eu7ikQco1JTKnJQraLJ25P60QBz5ov0N7UMUkOtRBgTltNwMezGKhfc5ZRsnR0jM8PogqT8L0wEaFXafQkYJqzBrSXtjh/pkuf4tFrMu7inIgGrDjcyAePT1qTil8nOdyraKbPBUXkHY8n490djSUEPm5BTBZ06fiOwJkHn+EDtgnR6WEr89sPUGJ771CdE3ef0yk+ptT5wZFsTmSzLH8DX4DIGd83YLqyrmo6N46AdnyrxELrLECuRap8Hb3bLlyQQHBKk2K1fCEOeXu7oqs6d9F26K+SgDpuirTNdKSjkT1Ts7Xi4smM7ACXSgiOOrN+IJ5SYcVZ3vaX6+IGNbPfhCEStINsLLubz/yfpGOVX2eLs0axFkv2bkci/HphnYJptg5u4mkJ6PzJVS9gLyUHMtfQx6+V2Nq+9XsCKPKq2NQg7DiZ4N4YTz1B5FFYNRD0OtZSjhSGiF2HS4AaLDoCLe5dFOUJRAB8e3pda1881NC+SPVkxzxuKgcauMbE82mCoWK0m0FvfVWRryfOo7igB+wtvSXFHnFs/+vP+r5PyFARxSywMT48BnrLIxOQpAwXS69eujDYK7kAnLMlf7R8tl0fqMzKaFnzNHN4yqEYa0cp7reC4gI7JvQdTCVmgA4B8guEM9O2/w8D8y4C8kjkabmxpD/7yHRAknmbieZJiYcDTQ1eLuOyy5k3HbaE6hY4htvZSYlQ20pkboIQkjfKeDCU0CGxY+Hpsa8jJUyRcOE+/Js1LgD3sKzwyC5k3x3xf1g0ZZ5qI9XX1E5jQHDXg+ph0lbQzgzYzMTj/Lk2EcilIpAY7TxHMVJQVH6Dmk+KNRY31uzb59D0hihgXaxnjwY5dvQUgqt5wBEWZckRxXRilC0GNyhLnVoDEtyqWL7ORHSZ93fvBKWTGDDY0nsLlcM9f2SLL2ZHnMncJc2f1SMk8uP7rzdyBgYShf2F8z1RyWqganKqw4KPeMaO7PYTQgOAEsheYJgr0U1jf17WYTFQnzUSoFEZYGdX0RvJyEIaCITP0TOMeLoDIGB9FKvxueKr6zPCae9jvtorjUFgh1e8zGz+7alLkyqALxHvCJAJ3iFnGF66r/0tfA4p2K5sw64C71i/yPfnUrW8CDUj8UwzCJ7TUEFOOTwrQ1U3nBdp+MEwvr482D+eJYDS7yvhNwqA5C4blqVY8FTRTI4JjO/Zqkmi3FjFB1Zg1nqQhi/s6sYr5zDPj6SgBk/jM7FttqpijLFJrLMRXkt13wMZdQU8gPnmH5ZLZOgpHTd79+ODyEfZ+e9CfEHDXPaWNsrzMgxK/4E4QIJ24NDQ2DuIjOBad3T0s+4MiPlvFUC59rKUjGsJLmp7wrBXJuTt8OllKsOmJ2rtBU8EABs9le4MaZddB84RvSRs/EJgXgiznB9gEDwssVejarfxeFl+Sfxf6fvpw4z/Y1u9fPLLskb4mTtQmlnsgvhLrAw+BPLnm/tC8LsRGCGbdionQcKomWFiQeDpechWHoGOkM8E7OgezsxhklkFTnfSftOGo67KmJSZ7Bn7KY1ZU3w/UrMbwFFXgKJlGV1r1UzNYlNd4TX8cbn9X0bmoOSn3LIUtFdpU+ceBRHrlN1GJ5SKr4VF84kAUbtwu49LE5JVDMiBRrBC9wREzRwBcxL6g0NsAbz5urS1cKvWZNKWIkz6VVfJIxdHAZF8oAhiUjqBrwcz5lfZzwI0WzZQyNjNtrGoY91bUHIopMAzI0KLyUCOnXpXesR0EQ4gtDLiTgH839IYB9C4wMO0B1lsf50ewqgr9fygJcjBfllkuKt6wbOjc7GfERN4W7x4KzO2UK6psgRF9lfdmPMn+XcW8QmhVyHEMsJhPUYDXDYduoL9rvEQZzqGuMP1xdcEABhtw5Lbn5bnN1jVICu53qrW265jWqPZdY8p76lljle8hOFjEnhyLFLln+8eAb6AA/TpIPRiqVTCOkvaBn7Vc6hsWlZz/mqrBJkRqWKCDzrzW4z2rZAKB5RsJ075SUiTkmzwZhrRYmbNiaBi38TkmoJ3zOsDKBvYpTzujIzpyBKCghpO9FWjligAIyUP/vQr5M+AUdQ9yajOU53D4i0v9s3RMLHf+pKK3VfbACdqqKkLCKQ2fqoZLqyHdy5RY/bGROMlslSqKwRACTdoTERvXLrvm09HlJpmBB+cCTsS1i3pG5mbYjaGkn13TMWKtg+573CNtin88pItWkO97Ox7zfGwleSk+4nbqwZO95ohFui4YpIIq656QXcc3oVZCHRTB/XYIDRiwluUrlOiDWwz7QI+QZPPY+EjcpeWYD3lYbqGSGpQ4js/fWsLWONh9s6ppB7b1i0ZAeeRZdhUJWVpffhX2HJ8UqGy6DLUEVJuCEgJVi8TwU9Ur3al5JCjIUcJRgJIAkt9vDwK9KIpUjWx2p14Rfkobvy9vh9vZtPoog14AWJb5mBsmlxxwaURufVkHN7CN/2SExT3pwpFgX9WqQXpjnKUnfnXN8H7eBr2/AP7Lm6TBmYS9Jn8P7L4NwMLTno6PX1BJ0+pAZGgzgZJgv9JN1o7Pjmft6NG/YJS3tXIJJAbSrz+6pmrWQGQOZcKYsT5rbvmri5jyU3/1gvDPQQYzOPweOKcioRI7T22bwqj6CfxLC/qMrdH7sSzUKlNntDE6loMwEqruhMWvMxli00yyNpVa1WvA7HpGOwLtu3wS0goo6t9Pfm9uDPr58yZwnZDkZBkbQf61A3/2pFki6FW8k69J+HN6vP+g9IZahzxeeizmuE8VnlGDeAKuCGT6utYuaILfRd+Wle/GxpEn0D/aNYP7icfL/6Ys6xZISXyhsFZ2o/kBoUVMjBYE7nUR9LBOSLwe+tmZBzuqTvBNRPyUjEeQVkanJG3CNZvU0tGKFoRCDFPJciwSQtlI0e3YJ4CwVMufk=
`pragma protect end_data_block
`pragma protect digest_block
9d40ed2fc5501cd3ee4d8fd8203c98e33f17c3281546f840fca1e54036bbc0e5
`pragma protect end_digest_block
`pragma protect end_protected
