`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
rIKohE0RUglrOnE6l1esq8bbZVRTmFbAQpba3Y/L973LF41l+qgHsTGO2NhELEB02dlyWg9AYxM7/vKzHgFigYd+3cxEhetoq8Y2sFQMNmA07fwz7WAtQy+/P/UXnZfwewmolV+V6ncKMDb19brkJXDL5uWbNknk+22kKk8MmTMjzsqh49GA/dds45eP92BxDHmq8152O50U4eUmYmSgMRg/FTNRIBKVqesGBg1GQWEnRd4+QQX8MPWd/AvgqamN/cp+Lizw7FlbxvH977N5pFqn69S1o6hYRu1OTPSOVgGwy96lpk7Sx54If/TYrJ44NVhzZe9zWyEsEGXSB4bjV2Is3l1QcqyJfKlQi3nW9BSe4CyTAOsszcJHl/WgVjzvQE8MkG1fy9Qiz1IqSVagunLA94Hoykyu9Tn8dfC+M17fBsqgOQrQfb+YZy9fhoAhY9fULiQUrC67NSDUCeCBVzxqFAyOnY9oleQ+QEgwLiv7Ch6EERmFZYcNBvFjHQMYBuXZARTFbybrR9yYS7DbL9TNsxcQiklTrQZNOAEhm0sVquX/wbg+m0MQHPw3p37iex49PTYkl43VfDXtHQf1YiuXRo7YqXZN3NN8tBnDQ+xgn3U3VOh8LkhAyWE+eeZQnKmOWA2utJ9uhl/8GudiZydvXy0xkp6ywDyuQvloO2/2mFqF41i/yUNdWMBcI82noIXz00cMdZxXEkKu5Tn3L+tkE6yzfIF0Ot0gchQ7uHl/cTFXgGA5W8aH6iYo0wEyJjKekFG8t8uF1yxLqvJs1ClrOV6TkOkG0EbWCPPQs7u6DxZ5VrNwLS7qOyjMCey1jb+ar3GwAZUGhNSqZ3uq3yTA6XhCd2tIWmePtixXw/3/O5R3M5KH++VmtMo8+AfRDlWz8tpBEMCA+rkQn9utAV9QtUWiarqFGyoq0wvuQTev3ZI9vUFTDT9w1a4tuLq04nHNKnuJcjpxM86+g5PvhyTMOaQ1NaVmKY05L7ONpW0wLFXR1KUGSDSapalPFhd3BzjpL1om7yC0QNJrYfu3IfGB7QEve5O6XbN8kX1W9JBTWOVTyB4gEs6nf4Iz8Fbm283m96xRMydSY7lIg53wu8KYdX80J2Nvxqkdjl1Ni+m0cIKhOuCZ2PKCOiy3HMbYgqTn9fUO0V9AtkmZkRZLLcLtlIkXAwquO9lv/+Y4dBfedYL1V+YtcRWjI+AkbBs7WMWLmx9MwygdS1VvShfdezUdhguncxYIBZFexSqfOlt8a0+VBt4hFvQL4OpoIx39D/d7e2XmtFF9aNrWWASXKG+5BJnz4DfHZXfplXU/giK2LsXxnB6/FSAT6Gu6OogLH1v52qW4VycC+vWHy2b5/ck9jGRKlOYIKb2TA5HtGXgC7eBXzmsI0Hwg/Hx2cyi+KIvJkZSnxom7h7iNWZOwJFoKxeqtf+9w6zd8RGiWlFcZEdIn/MJ0/tSg9Hlc/i/w3c7r3QQSvAn+io7yeLvBE8hn3tvW3Zu1+6+XVkA7VNSxFxsAfN+92lse0EUXp52Vi0ZlNmy7SQV9Jue1bSXsVjzUdsPe3KBNWYoR5REuhItTH5WIZySVVTGeQo+aoetXGnO8qXqpHhd75+e7vvKJCJdfxckkjtxCvPCsPjfgItwEnd1w1fLpmMzAa5Q4Cp7ZyrRFM06oqHwBWiyCHd9Q3fN2YjJRc1LbGreDepSh7VFwJSqqVSqCjnNPB0QQHP+DkoicIpjj9MKv6wi9INEnlT6+Jy2L+kbMMPMLNc0FxduwEVZcM/AuMImIC1Ir1jdKrPhcK65EQqiX7QqpqWG/199WNVy4ER3mPWer5MLtfBYlkM0sZNMPxnDXAXGKGY2Yh5Pud9jaMl5ql/d2UsGIpe6bQrhTHHbR8L3RL+4mBFFpA32cQyWQpapCfQBe0JAEeAYGzYcl4LE+0hVKYDUrmvsimcWLhu/cvValMniz+SaPRxFYJ+UPzOPDmA5spMjezWT9Q5FhwEQKNhSJL9Dt2elBapk6lDbF4DfVk6+AK3zMlYRermZsf+T0WSsnCbFEBznZmiyo/k3um31r4h/xe3zad2ONAqey+BcnP62cKMgEQY+mwsmj25lr+rCEdbc5fbivTK2gb3wtCC5vEYp27a9tZ+DDHF8x/SVL65ZoRbx9MHNPu+u0zN4Xy88l4FnuOBOtPZK3zwHU/9Ag6FgIa4ALDMdUuJREy1SZMBsGOfLZmrAwjvqMFJnctQ32y5bYVqwP93bLPouVtd1aSnK3+GJejycJOUi/u+1WA1yHuBAcZBL+gm4XZ231psM8pdOny8ai7fFrmt/IkpYw4v5iOTYuRb9vFeQNL6G4uhtbHvfSfv2PzfeEum0hZaw1vzSWASKnJNkKPC7lBPLJnmd8W7fDpQzMYqU7PzlRgvhN8qDPdJxgC679aGpiIBHzC4S3/1i3e3KUazyMuWr1TZASSOJgrBZA1RdxGvDNFeMZ5e0itjVjgahG5dcY4wK2L78L13TK1UWZG0aiJxdYnn+0GA03fcTHOzqhjKdkmKYgFHkViByY/PzES4mvNt3pY4xOxafNWkuh2qt/5mIakn6L0n68zB9AttciB8cjaHI7/3Nr2ilqZcE87BZ6jM1HnDudsr4L5we9pXf1mdBsuCSMRmGzVdLdqcn8LEqw2GSLh0Jyu74HOvaLbgGU5XNdww1+tge7dLEx59ETH6SroMJRRiMkNCevi/85Isa9xtf0HEXVURmkGKeUALlA1RGiLwWKov7uaC8ltXNTO1gx8RvVWirp/9MteNfEWhIkWmZTTQ9OUxKfrA6ckCAbEce5mKaPhx5L/1wmIbH/cQiS05quYlB7Hw/qRBmsL1h7GAqLqYmLJ6CtLva85P+BQBk+ZbY02nINDhNuplmiLtbryuqbobVe941lZu9k1/afh4oVqpfA4Mj4tcfExK9vQrEQaf1TaEz53PwS9eJRO1VffZmLjVdTaRY4QSrER81Mz3x/UmckTYfBNT5OHFW6zvrnAGj7jecsfHUB4V4T/KdqWVYF/98ZDLTAWpp8kmJIit2DqxqYA5rh2oQbGDmbsO04UFT7Qw/Xez/Z1ALS41dnycO8Ka6izp5X530XCh7gNzx0b1TfYU0pMjDJbO80oAQNOCeGk2puADsGOY53CTpFi8S3n9LJl8ZgLIJZOouwhX2mFdbNcft/KtTdGPxSe3Pz2qEjzyHJLcFZpSqpKzWXufc6h83moe2NnJtUbXW3RPqKM62Dknr8qHG+6poQoztgqlb4HNwbtjPj9T4s697zIMz3GayBZW/hScc9vhs2Rn4rO3NXYouLbL9c8DPq+Euh4BSarJknwh/7ORgL2b/Q2waUhhFtFgllRCy3sUD7XfziKLRH6OKOD1TpPXF3p0wpMmMS/puIbMr3UyuOEwnhwYIPzD31tq8CV3Ht82BvnBdl4nqIe1AmeXx19q8Hw4qy7R/58l64HDTsX2208SVhdP6+imZIT1udLsXZcZ8CiIqbdm3yio3h0z9Bejiedt+C65ZRpFMCdwmJaeMclj6wU2y0mJ2cRGXTzNx4SDiSe2H9acRQPmqzFb7w3jflZp8SCUsCDlyojexgPJEH7llbauxZ4vdn+d8bm8Cvk/vMqnJEshtnD3V63QvO3gw+NfGiCs5y/jHdGlyRlI3GogjggWEYzew5mogtncc4GcQL5Ymgla2rwk0Po6PXmPeO51AYta4PsR/FL24GSsDbi9xzFGwKan9ZBEcLdt+DF13octzre1R1DbktsAbMXrjO2BT1sYT7zO+rc0knEY+a7/5QRpq0vIoiEhsPNtcC7Y/uuSkteZlJlI2tmo3QaM0UI2LmzMYsqb9DIDlSpX29eJMpOSSiLtNW4FFykW80DxdHOIGQMYWgdHX26I5m5zIGHNeh9k/GQDa8H7NvOkv+gYJAH0h5v1jzr9TIaLlIwck8x6mEN/omB/t4fBO/ftyMdinYrGOtfQ7HS4kVY5+kR58fkVpzHdsL89nsW4/fiIFcBnirqDRUhQtk1X01O5xmcTUxQ9a5vZNrNdZP822nEOz6rLJW6c1VM9NKm1C1sFkhR1zUCEBaqdkgxjAm+vqdTzYFGh+vuMKCUxbk+GpztcfJuUWc1h2n91rCR/Ca3VIPQH7vlJlTbN+fT6mdhxx9SlAuPNdf/3cX84kTx1sHqbpyk+Lxc8DxMVw7pNwpg8GRkJ/To1kcyOHK1ooZLckix7NBvAjym9OAoyFufNrMuJU44/8YwFxTd7qDmosLNEtA8spXbzXP02gymzCIyD+PWdmFEXCm23iXfKIwlHGspBYsocg5GBGBvk9HerdUx+jdeMB3QuG5vZ6kg7scfEUJt907o0UQR99oGljX9j7UHA/Zd8c3EwzA6OSnTlxEWTVjaXHyA+wrjdENYiaWGi8ESyZtRWmOuvYiOHVqAas4IC7uXUV4WqkZ03Bz8ze5qVNUKVXqKD+4H+/Qi5k61i55SJy+FpNsULMPVNWE2VEjHbJ7i/QuNsoqXKGy4qJG1Op9aqb8PNlY/mlmbPdhsCK5vfg761Q3cCv0CypPq8j3qcKHQxSrnEsCCzdQt0Enn5KhLQsgADUUCv58SPNeWXM9w7Ex6vTOczadXibOWhdBfXtNs+8mwfRlnUHRzc3DRfx5N4utRufJVc96IVFBVZ//LgtDTRjlpCsA0bujNPIJmA2CnNo9+sbDBgrO04HLCwyATDL94DQlrfdcgCYDJEty4TR4voQIpwKGRxrxsdkMoAv5bkrI4skEVpW7LK8KLFTbq1ozI2Xkcza0w/7h15Cmusxm+FeGxpMhdRAvVgvQq3b/ty2RPU+Kz8XmHJfXzNgkgHcg/FE/LBYSy2MW1Q/jYdO/8ieon4iy/DcQ3OA6z13R6oIf+9eBqKL+gmP8QLTFq0ie4YjM7ml8CrvbAT2BstMIW2FSfey7X/iFgOg/wsez+zJfOY0nN2WU4w+gWBrWroZjfZ3CNQz5uXq07q/TDeKoqYRuYkV8uNjr4bCLu3Kg5KJt25ifoxciAxEVfFhnkkif6VKx0osir61N7V1r2O/5ehttZm40Nn/XGfl4KC2Yiig8twf6xG5rUKGsAjJGYXZKrgC3XSNb9dwvGa7zT9GbdrxukxSIu84mb5W1DjIzWFSdUHxw/fgOuieGCYkM4GVHcPCkvWf0GwrOGS9/cWfA5XSB2arcgnEqNmk9I/ZxJzGUbUAiFNIc2RUfb6dq7/SuxpK1o1h9yxGUSc9KK+NoRNQoC+N4/2ThPNZes8XBWulmRnPzzDC2SKdfK+41FzTO7rZgHUaWSP3fbqwfCqDGf/s+vVblLDBv/p9U+3Uk1xfex3NbjUdZyoBFDYbnuZZo2ffA67Tn2PNlf5PP3dQB0OVSAOniJ4GNoKUVBR2X/Y+0LAMHif87pk9Jy5KXx3KhlAgcH0oGOFhJXazrn5LslLaIcvmbxkz2asRK4AN/4hEbcrSR0wydusKoZbjWIiqN/dYJezItH6qqsyt/YVilBizWL+ifsDm2v8yAwDMAbsWIhtyfAHRSloY7mmJp+jM7YfXrHuzO3H8C2EvAYAMj2w8T4TMWXqlOvccohBZLwFVeDtyS6Wq1EkjkGqB2nlsNGY5Vvh6RHbXg4X6E9/FdCgDs7GYArwYwTPSGt9wIxMKDY9fhYdo6ft4yP4RbQKgAoDInuTCiM77objJOncBs0zb6VkVNWOBC2dMmZxGBq7LtvG41AbFs1WVGMlQvPrOkIeuqe1lJ4FsTlOFccfU1wROfnWrW2rx3343I8YvFUo83FPPdQeErjTlQ3dad0MrIv7FVlKcs00Yhvq6/bP6PZk6pvqku/60yGeaM3afrNrTOk5m+qU2jVcPHvGo9UtU7ohU8UY4nyQuhE8abKvtvipzTM0RMFgD9LtFkU2q8vAfjxiIiWE+gYtoT/wN85M5nzXbqwpBYmItKIELWGf7sdanZk4ZjdTmQthaY+I869SDHttLaC/09lVQT5C1WzuoRX2W9ilYUNONjFe517lO29mqi67XsTqKkUf82DVXNjkMQOuaoP1jcVQJWHGQX858rcLMlDFQIxwXy7PDSZ3bwZO83X7GkrH5dt+5HrDNGDICXouRfRjBRFNTMOCJOehMgJ7Y3knhoXQeKY59AjPpjcfl0ETNJoKd3AzA7zh0axfuZ3nJ7CI0qHZBCWjKO8fxE9FeWG6IWEcyVW5Zewidw5duUV6MSxdheHAbLb90k23F1CqqSPleY+lh7xkDeTjkSWgk692RWe2cNIe/OFIq2qhPtT8eHauJE8yWzHpfeVG5/q17jEjxEevl+xgjvO1DWydimf/wLdo880ZbPH9ClFPxix41tbF/oHLqJZf6KwhZfCeXG3INPJzEQ7frU3kCqicYBOPtaGKKOsX1NJeS2+2PB1z3arwYTYGExIzfBDjO6Tj3vP/D8XSaJ592x1Jp7HyWG5I9kxMpYjv+TY33R9JZJbdZk4ClweP9FH1bHyKM0np6L3V11UyN+5n7RyHqxbH0RL28EGWpweHleq8vVJ4kJkpyY1XouJKDVp5M7kalQN3DRXGo9scvwH0sWUOmf0/bkrFCC1K20d5ASSkzaHBambo3OHRybhY/vPdjx2HRzQ+0GeO7qJkfKfgX7eNG55gJC8JCh+z/uxwDZkQ0BDofCz2p5Xvp0BKnGvgZwombCFPCJHxgQ7NuzwaMV/SaEth+K6qxxTZqu1aRKsyr1X8xX6tG90MJfPrGPDWr/YLZNIods3TFpTbWWHrjuCbLf22LokQdFgP52Qii6xrbX1K3VyG0U6rGHGynBooJaBVc3SEkX5XVcPQKmxA6ZNYT+fv9tTtWD4e9NAmgAL9tjYLaGIw4dUMPR9W84D1H4U+27QkUSh1Lod2CJtAAvoTwBxeqD3LOMsP61v53rlDcF7XBOO6p2QUbYboZWUcfoZVC8UVZaHHG0H/dYABxAnz9kPiYIwjV9WaeZPaAUiwXGRk79+utddqhp2iKGmZO9TiJpjUSO+tCl8KWT7kqZT7PuFIk48gOdxcCqn+2BsCPy2xezv4lVyiR9y3A8qEZ8k46UZw4mx4Hv/tDEJy5pVVo2/STuqrNjXqlJM7ng+pndGN+bKoPBhz+KBchBUJPwiHuBG+EH3s2hp79PMkVzPUyzT4yVPSlAjIjUzZxQ4uDzNdS0ovu1hVOcvMMOeUlWdoCWBJGRrXFBieJYl7pU9ipCz9J+TLJyiYv53kpsMqNYUm3QQH/o8ehH48tCLV6bo2Sul+N00m3hgvc7I545m1bDqdu1mX6fj5YMv9o7QZW2YABcdkVwW/VGVcF/CW+6bZ119eY4eCysWPa1CuYc0v9vLMpA8wePNONpUMPtYcSdRdmOTnRsLkiWsZ4XwqDJ97EeWBJcA93/g31FFsIfPSbP2EpwTg8wJ72vnqQCJ2pjvtab4dnxC4P5lvQka9GNblrmKAwXVyqIVPTcM/kXHEhE7nuXVobfzv4nE+U3EgHOLvHujVroM3KzSfR6shJAC+DYZnvJpaiW9KnBM0Nrb9Z1LAEzCSUk2D4EdWwc909LBczBnxaYVZcsK4PYadBhtPJ69s5CCU9Nvto5adK0lCsW+KpFuYtK/RLJ1QK07k5Wc3a7rKrxNKMUqb+YsUTLwt/M/Lw21YLLHd0edSUfvYZ2ew99VCjZVQLhkLGo9p1McAnYN9G/dPN/gaA3LmBLa9IDCdSAxmHdU8Jbo3aN1TbhgsXW0RWdfv+x5zYbrBeorTvsQjSMfm1CB2BnvGs0Tee/ECem7Eep2pKJSDtW0KXMK85MeKupLYtKDVv2R2TI6rfXs6ZtkEvFphOFjjkcWxawNbslxfj0sOErhPPB2VhXTzPMoBwf/NtpKudBx4KvWl8HygzPj7t0wKCaDatXPiWvqdVGrHMMwnSVQeuGz0ykwzBeZP+Q8Ak5xbk4FJxWiPhQfil/5KRd+lilhiSN1pdR4hBbIfmH8zRP1wbx5jiKKfXFAdRcTEHB21MVHXLktVlPF0/BZt5lR6mKEcJzcmvR/fehnJPWJpTp3bCiM+XDacabdJDY9OZmT1/GuiZIah3l8VajOuPjJ8YzxQe3KaVW2BUSUwllqdxgRypTogZ4wDedvxmKqhY+i8qyoua24FjN+26krDhpNQ7P3NhnuoKtbM7MSFgMa6q4836+b62mwqG+hwzDtJAWYjnnDmbuM/Mcgo8+cSN8owmxbEhn2IIxFsxr0v5Yr9oV8pZi4ZJ8M3K6CM6Btn4iLVblr5u3g6ysRnn2zDlaf0NW/gUt4h1XarPbzQrLm0PRcVgu3b3TX9PnE3rVT0rmveSZ0bEPG9L+EvBgdF/s3iOHnUsCbLpx7gSClYlly5Jfs2G/MSQIjEBQVnMt5bIfmWsR4fgidKnJm8ifZ9qSmXlSu/texXCsmsrQLH9GIPtJR7fOjwwQ1W7YK3aQtbpW7m/IVZEnSkIiq4hkfW+ckiiqOXBdpBgg+f+Xm+jMnINtv8QFM1R8YTTGGaZr/e7Bl+rgOQT6noNkhEenoAcgD9ClWesvY9PbsVVkTzD1mxXPpESK9/PGRfXEFX0ZVR1xF7EBlV3TN0MfRejY1silW9o8hmB/RWF0r/4l/+eAztJ+EoaPD3BxbbKP2YDAhdRHBfcQjwNBazBlcSd8ZiT4fCwTbZbaYFpq1h1euX/JXzVLxi/FxYFmD2c1IGgkeWrUb3EXzD04Zj6cy7yej65UF6iTHNkaI3mJDTwRDqUBYB5j3BxGt46hucIGhgcH/0k3eAr6dcjuaCT5DwjeyWo+4BELCKHYK6x0ilLW7G8qLykRaJI/93Bz/WN8IQ6W1HLbUq80eQ6OFzmFUtElr5M4Zkme2UwTrR4MqlQDmfN1+52xo1gALsGXdWe53Fm8nVKMdEZBUDWI3z4WMqwCvojY3zBCYpQZgOvPF4Gu9HZNno+pND4rS8ZzNye5eUqDs1AALb8+7vcB3sIhjhR+HxC6E4Fitd9mjoJaPJtscn7SaguP6NsGb4gEJ2he7/tu2QzUaDJ2bpHAwIMxZc9/SNOe604RK3j4HTRZvdf1GlcUm5nQaswlVTpRlIfFoBLB60ZbplauUSqdTv1ATjx/zir1TABBzHP9/50vDwO6nwV+3TdKZXeLhPM3TEBW46xENY1hKzpxokL21xHNmklqVKt3EKs5nqLW7gjZhOOHLbp0Zi+JERIZqOhaDPL3BqY4SAtimtYUPkZ1i0vNyYn5Wz+kXoQ6SSsmAClACMGtkDItcKh5O39JktwK0JsfZiFmAtCC6TL0IJLhx7FpjgL0b3SK272sXN5hVpIJyNQ0TcpmMrpXqYs6VTwZvu2GwYRJN9CkQ+2BDiIp7DysGarWQi3KDzlCOFFaoHp0LJKzZrVTv9k7dv/DZWd9MfEH383Jm1OoJ2w+REO394jujbRQIFiWt3gYc0UKhQOR39YZhXHPtasjIEvUsNUb8hMSHIELs36cPfiRhFTEuhEjVe0xx6i1R4HHvkRxlIN/AEGPFhcjPmZVRFJD3gqkk90CyY1l6xbPaXn3sALtHzd3xTuAcfWaeBIwpauJtKxAG6lWlpU6KxKOdLLpUNIoBUZ8c1Y9d8DbaXZpX7vPEtE+0fY24LsR5WGoU5PyTOESOIgirCm1ABh1u9HlCaMzYclAJgiMzkUHfz2XHIRfEC7tAVQhsK8qo/p9d3sYerdZ0nfKR+CHy0obgLZ1SgLgRzxb+YedhpU44tfu2GxhTafu1zPdnoFR3u8dw5u8kUoyVlJwHB+lJ2rwkBL42OBlXtsSo3zgn/s/ZI0DfcxhWN0VMoAfxVgCLp7RWxybYK1PfqdVw4h0qDK1p3Ve2j8JVb2lmPNEK80bwjhIbGWhsytOTjdsVh6xgTC5Nu++EKp3DYv4JEfOQz+IEWYT4xYZIMZlw5jAlN1gcYrCYWwyS2muQfK0Ow4lz/jU2ZGE0ADmfsqj15ds9sGwy9O2PJMMyKqHZPm0Jc5fLs6SdRWmg2+zTijRjwrLoxgtp4t/yNglDo3lpbhA10SMwsOhYk2Cmt3LxX5/ECYsw9N2yrKpOx1GSotzj9uOfgPDluM02ln/Go1oC7zc+qZjmi/DtpIHzpXEWs3vl2ICmEsPOEM60OLKDsd5FSOQNuZ6BIuQDgXEP4Tg1A1dGOHb6WxSa5U7RYVtFPyM9xVSd9x0C70nRQbv2XKlWIkj7p+xi0EUWK4If6OOszTOrs0bzCo/NGVEybRfpmlAw5JZX26wSW++u7sjx6c3MeqpLeOwg3s9Se3fICJV3g146EcP0kSJaTTiz7Rg6GtzNfNmeCA0XDiz4VaLec7SpxqBCzw2dpVzgzR70XKZfPsF7WVFueNuYps9Xy5p1uZV9g5vvVrMcutSR5PIUpBpDLSX0A+F9PRz0ZkkaOg95buULETJ5moGesiuaVJt9ebyFdQqPZxfOUHMBl0GkFofWbElxQYWG8ln4RMPYVDQwzUdNgzHzi9pe6S0C1ILumqQuXYGOG3HLb+ZcycE/KXp4KooeL9WuGA0aWfX3W2ECdVBrb78sm1R0khsNV1gQkgXLo0ZScTNo+Rw0IoOzZ23jUHr/onVIh11bI1pb+VylTNS3KYNnfx0poZRVpX6z+Y7u1lnXnMGCVM0GyYZ5UdjQ4SHvAhJMoaSNbJ7l19FEkFZCBpabzNx5GDcmzQkYYpHAZZh4Ucd6uax1DP7lhA8lk1XgMFBRR/xRbVj2BKR1qS7QQ/j6O861i6pMfpNtjDlk3OeutBRv3HqrQkZco6r1gsymVZqK84T9EHVrA/AW+hZx1BbsKTpTV1FlRXDlu9keMRv1EX1RGdIa3v1lmaG+Mrri5c19FmK84C+zZ2ImX+f9Gy4bgrP9q/gDFGNJV6VxdABiEj0hpipIC7PgJawGRkUNx4wai7tVVf4EAbk56tHjJsDDeyVKQ/7MdNuImGLh2W1MkGD6ubpsDlFihWClyZkAPx3P6xRbBRTMXR0U3GgFk6JEXaAWeKiWLj//xcZQOH/JwrIFowDINI6xN9H9mEl6rQ22sqs481dS6eIsOQfwrSnMEGIfOdW+qcOkhLJi76bgJ/5cMATuxLU1UWD0euKsI0PVr08TdWpLIfLuXvOzJ8EOBpKLoSVkXr/wZ/kuHWEwT+pt0noWeTPixFNEr51mWx+obhY4x5Gbbnl4eWl9or87jm1jmUgPg5bMnWxlWBS+CBog6fP66v8xA7rt4x4LyRAWHx8zttxT8958ChFCiZnUEUSztZWBn566/LE4CrVHCuxl0TKuch56ySBxsybkL2UEC1oBV7xJEWP/yQyLPly/YH8YuoPByRhhEgCFgTnGAhqafyBY4i5mgLr9dgL3/fLoZgQEmKusloxxithmcLcK5g50YlZNWCxymC+aJEVWbHDKaQJZwiWjV5/tIlZuk5GoCO3xW2QUdgpIuV6T1jzmq8Zk2PJOZtY44fyQ9EuBq80Vqxkioctmlab861bvZpFC6MFucWxU9x7oD1RQwf0s70ceIvAlrCI5NUxkDKCL2KQ2cmuDgal4IDdEpmQ5BaSxm7s+kUI8inMuwYxu/BK1ZfUl+9CohXeDf6WlbjqNcS8TJO904ap1TBDicy6wrP9NTsQT9VleP8MvPA/36VsjTWJfbrkzERuc1fDtiosYUAUDfZeGvSoFaQezKRnKdauzl+SWQcLAsdtyPRespExngQtxGR1X0+2ASmQZB9VdDX51b5HHw413FY6XBL1T+YPekJTG9K7Rxjkm8r68+gZIKEIvmJb/2chfZNs0TIF6r1yN+UDs8/Ojsy99EN37LMBfjSkntdg+7P4xywxPfSbCDwiKu7Ja4U=
`pragma protect end_data_block
`pragma protect digest_block
e56fc2e1346c9d6c990422912a49ef30d92daf5262747c0ae54a3ae4d6f7ff11
`pragma protect end_digest_block
`pragma protect end_protected
