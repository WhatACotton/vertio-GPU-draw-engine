`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
8jDYxqgC1D/jzzi31bYrdmPiBNa8tcQxRwnh084v1r69ZjhsmpSNPwQKXjEU+QewRS+ho0lGsqyXsz/nLA/cqgzgCBKFJmfYwENDl+vRUC8KU2Dx1nRf+yriWgOb3Ud8MxlEqlwt+tvQdYiMQmTHmLHcOmGhZtTXDf3gaksdQRQuERdfcXENbR5LIdUCiBtCHPIrxWL6+dBbC6Jzt0m3vh1I9bcaegHoe1zJ518rxs+TTEE2DtDwOIPmkW4p3uzZVeVHI5Cx6v9auSoRHY+qhwdPtlWaVDG5RDy/+14O0LddAbGuHowhght9KxD2Il1jHb4P75Qoy1/xQdbhiMGUkfO6YNA+9vc0A7O0nkW/dV8pqqfH3nTWx54t6Zz2PM4fTmsxn6qAkxhJEZBvS2yRTcvvTQG+w45ykG7Z9ezpDn8RhS1U0YbpT3lq5TewBBIF1tybuYHcp8zZmJqiuQdZD5qTSjj6LFO0authGi8PHB4ZbmZOvTT5jlU8Y0Nz0FXlsKBc4FUqHRf3qeUC7T08Op9FRmMguWZEBO7/wDFKmKLhAvZFBKlfOu8ThIrvuDNkKOhxsEGpI09U//ki0FX4oQZypwzqXW5Z9rhz3mZzOzxHxV+mlFfoFmQXNkRBzxBfBRBpcfRJvnxm8I4rWRuNWEyoio8be3A1KEygxm1pZfTXbwo6j7K9ElvdOuo+9BYO9wyd1vchE/ZBNA7bVw8VHdWvnvwyCf4Sv0IkKtKw/YTAl5pu/yEeiPGOeMnKhTUNg7JbLBxjDja8ukXBShxBuT71pfLvvxgC/TXgmicLmHNqkXErMycOKMen86/KnGzzpC10BpTAYtymNH8L2+sUF0l8yj8cWb+HEDI8hLQMyjcCwjUeB7ZF3CDE0nEZ7hLp+ebwG0u+LyKvMRA2RbDto8JlMqvveliUuxcr55FnHDu6rlwDGLa9ManXTvy3cJkmQOdTRnycYbp3qVLwxPMJ9nRQZhe0dIk05jhRS2/7FiOGqJinfrTKYomaCfpdU9O25BFHMKGl6KK80/NCY035Ky9lHo0gykRxxqsIO2nCbtKMtyFY6dZINXVx1wlVmyQMiawntrAZNWZbFYThjUqggz8CwPpLNOVeEeRsa2+PEPhB/0/smJcQ/w2EDQraUT6sK8CIVCAHbiLUs+kfDj9mvlkarffNTiJBXrSDzl58DG4MTyDHz9CCXJQJwNMVaUVNSmrSx2Z/XFqvJ3aw+1TpHSwPbMStUHyxs7dZSfpyzq4wQ+fk0iugTlQcQNOi3eI/Pasc5YPFYYR1R3bTCmwGdPtZGUuJ4RzJ6hau40ZGAu77E+UtKEUPhnJm5uLkvI3AtMbdCwYZvw0Ei/FybTIL5Q6BeTnq4MRm7hpwFIgaP8/u0pBaNqXpA1e1SA0EMpXjoLtgjZO50xBtWwVhvyH83RjTlnYUSHwoBf/Caj/La056dU6XTUbAyz8wfD+KVgHHa1WhWBJ2G0eJ7btj4ZRncUTO1REIT4BBUTKYdXpEx7IiYnnspZfexpQaBGiIsQJ/bHV3p3tK/sao7qEZjV6y5PTvG9spUjTpX4SV0TnfE4LgimyXqwKst2KxNIyDWBll6pt+xF6gp8ibExUK+tvFjJD+uZImFYuUMMQ1hJaaVVNha3R0dyzlcaCLDZy6XGhF+5AG0eYoT8oISUVGLjBh9RqHKWDSKHgJKUdSKmoIlfIUyNVrca1Tb364YoRBAcdd/VB+HHPE0+yWNpEnK2KQG05s6/6wLbx6Egi/fDq9fbI8LfbX7u51pIA+N4l0Sc8v17JDr+MVJFpNsMPFa8J8hG13y4ftOTLKylP0U8VoSb+HfZl80Ql9RO3WqLrQ0nCz6QH3ct+PKm2hnxPisoiTO0TXGJikaQvhRkm66g5AHPg2O7xwmPUiDKUzaYkw3vBAi1Ry5uASMWy4WSvHfwBrq0+3TPJYV24oW2Q+bBfX+zbSmfDzYUCPsZeMWCvRNoeWTltc7CEp+T//w2mSAHIg3wRI6KhyLeZ8wLaNJtN3imEDX02yyXaA6L5jOqsIure/0xJVclyCLJRMstop/Fepi8c8Mwm4xVtNuIfW+W6i7BPnPx9Jx2tzfSzIfK/BWYU2JJfP3Uzn+6HTnosV0XSC/n0AtRViKNxDXDIbl6xgAh2FvFED4HAPJkwKAizCOCQgkyKj/8ywQkCczp+xfjlKv9LJNnIaKjILKzwR7BFSlZGNuSvr9IlECtOtOFL1JYU02oB8Mxz4lKVidLV5jGZBTplHYU1iS+wyllyNGOdskQZxv4JJjg0WCf/Eeb3R1iBThDYl8NEYMsHpRjvB1Vpg+qaO1N7lYZmzdjbAJUQC0hABUbIEu44rvSaUAwQ8BpG5tMQAZYQFv//1aRxMhV04jM27t3ox85lCGsOMPBybht0z1Oonh+zKY5y9RdWK8S0upGdtZuDWTp3k/jxAG0KdEDtMI9SDxeyCBO3E54VkFMb7+0PfM7USd613Udz+i9bgJLWihHl2COPVPZMtvd0HGpzcTMwQe0SX9MRft7gAUz6T5gHA1S+37fTQhPZ7n+7lTmZaVKiTHy+Hv5+bnENEwn6tnLVEsbIAmswAoHwLZ6CmtuOGD4t7BYntiG2Ke/kI1M57fsf/Ri0m03SJUYInRlPtccKtJVcdjKhCpDLam93pfiWI2fo4dcJIyqvUKWB9OtusrP7UhxLiDVExwbsxSL9TbfvG3tkagKPIPBYVqo4CefSTIgTetbFiSE3ocaM0/NnJVQh+m03PplTLYVtgUe+vzVCEvw82RjOzVWjAahYejzpwyHsFyXqxPzAiGLSyOD8YRFZNNj1CcTCoyrx+sk+dN5b9350cnNAhTpbvjR+8lxoMc86Vxj83I8dD2sgXgkoC18ZoQfNXBlFt1sjlsF5U0R4AbpZGWWNg+VK7dR2rti8Dy+jkDpIy+IyoKl51/Nkupbms4UmDS29PAaoc1B7YtlsH+mVqoYwJn56ItONBWjC1GsS3q997bksxiv/a1mQeGu+Ra04ePcCBbEpj3oqMZFdF5bMOcDuDECupM5XkPEFBfuQMZP+0n4fL70Yhe+Dc8RGFd54NFpYucXNwP1Yqq7CqHtHabGxXVikBfQ/JwnEzheu9aA6LZt4TRpN/iJgxB4mSmyChjjihIPf+sCaNnySrPC7jvb1B0aONr8lcDeNKrWyVeu7090YtRXmsSBFb3k10h475vfikULJJNx7l6wSZvnVt5bh7GgpH+5zFy1SYgl8MmvgW+xGEvkSp85HvYTflhDGzOqcTb3TVtWCzSacnQAjnW7J86iepMzUa3/O87LQnjrGcHsw1I73bJhJ378J3cQHrf5v8NCf1bQBYBsZYfRWZZZ6KU16d//z42bJ8WrPVtK5A3Y3nUaHU1iWvvot+pcXQYoZCKwFtHKcxl1DsQVLtZhUAF1uKSVceufGWTLXotf90jLmi/P28wvFyASwfsvy23gzSVNf45JtPB71S/RgjD1XbDMWjopgAxtJKBPqts9dDIAJEaTJfJtLhkNn38URHa0Oa1pBtDiRn3HfuDJAATLoTY6suKK6q8KZWeG26mk4YweP6jqcah+BHH0KhdpNP+m/40Mk/jlsPmTc+h7pkd0S4FjsXo7WMQ6EVUN/Wg3kt5G844UsE7K2Xig/EUi5VBOra+8vMMLoISVSjfBInnQXC3PH5MoRok9CJeHtjhJGEG5P5RXcpJ66G2gb38OTvgzJr0L49eTiSl92LAYYGMTooIG8ic8bgSSVZGTjod79TwaIZXD107FE1xByGvS4YOeAFjrHi3kjlBbkYMi0OQJgPJkFKu84XJQTwFrDemceEa3RG43XQGD7jHtz0GV/3O89jWLFYB0bh70/DMN5Z3zNmYI/KkehX5f2Xk/vM2CrGBTTdoLsM4iqP0Lltzah/DypEzon9G0E7kZi1ld7AE4al7iTQVZg0gVNkgT4RD5cyQKQFEm2bE30QjHxweYB2wqG9Acoa/xAU9wuhvzQjXxuiEE3onfIAeQdrFfPE7C5kg97KavfGa5iyV/nSY5fxqM67NTC7I1LlcJPw5QpX2X671JkXcxLZZ+Jt7iLzJBpgDFxKdUzx9MrFbYpY+lVHaT/N9sjMprt2WKyYSJoRn//NUbjvHypLTAQ2J2RTdTc5S3vvs7HIy+oq9W2rq7pB4rSdUUofEcNqj3ZbQGmZxqfRq7kzKV1ezwO0jw3okrXWB6PRaRG/MwkMxWHsmm4BioA2BO7TxpWQ00FZQ/TQ6Un7Dnc1jpIg6je98aZgM7tR/aNcat7eBbtdOLwxKX3V2la3s8efBqygMJi3QLx5nE7JOew10TjzhLkLtd1WFc9wfDUxhKzJVUsdUoicnJcWXoLtgDFH4bTFeWUS5IcbUDNzfWqTfoD9ls+lWYRAfFU+hFT3vXWxDzlBo6yP0hlLOwXNoSfxb7BjnA+WO15wXzH3UMnscwKoADkzR9z81SdJxws9uAcLnC1l/GSd41QLCW/PTSu5bXrawiQnFJ1BHcLPl9j+xTS+CavdJNQ5FpKzoW06p9uCec+ylmfvDtWeZc00sawUBLNghZ48QTJwadmOtVgXuIZ92FzjLpqZe/n3qg0KE4krZFmPllYUV814DgXNdRVmL0y9bzg7g2mxB5G2f4Wl+cl7rviRJqNHI+1YVBN2+d+Qn7yFbhmNwTc2iV0dEZyP0uXLXv7BZEBFt/Sjsp/CUd4t+zJ5iGNe+e5a/VPvbXjiy6H2cXO4YM6eOaHAlAHbFdhYmx94Bqz8LaCPQyMPvci2gE6JIvBsJ1EsgdVLYhSh3ZCgvj5dCETB6NmPU/TvrgRagfsufL9MjDHzRxn2wfaADSxcm2gY8S/wJSKPLXBBptdS68cUZJcCo1GFaZSwgsdiyJzmUyfQcNk3fRa8QP1Mhk0RolzJeR7ZH9qPxR1BAPfqfVf61xmP0xzVWQbvr/QhHv6r/FfZ4OFTKDRHoqDKYqNKeDai4OZdD7Yi68n6JeCXhQFgG70q3WGuwasRT3XRAML+ZW7xgv+fZNSyioAIrZoE+4aPp0LTUsFGW4EnpcAAISPgcKCSFDGSMMP/bQVzml7mbjJtTe+gyIbDopOXbxLyW1UoNnOlf7wgtL0lQ9xChUsdMaSJPxgPSrcxzUdYsiP4DAprZfhj+LBHYZuA9h6ACWsirhPB18nYBqftjBalrmA+pExyHoKgxHKAiK50CsO5oglkUHVRSWD4jpCAC8LgSZXD77FcSCLJ/UNSLOin0h+C3vVYQkjRssHMKJLITH89NmyUh7L2KgSmlopyMErKiHlXh9qaiC6f0GD77WIwJywf2qohNWT1cMd60EnQdLJChvlWt5NCncB3w/lR2DtYIi/cym2lT50zAjJIF+eJ3lMqAWKINX7OsbhNTAJ3lnwmccF+9AGeFTYWb9PG6WGWhT/ixVqxfNu6w334yDw0TxYdjpCLPBIMdejZqFvCJ3fuiv0g5xNtO8DimXnMMlemZHCH4475G4knJaK3iADPEkTNTU4EJNa//50tGeBh/OfvhSi7C73jYGHW1+dh8qPFwljodrUq/0ElUsBrzBQn3/U1xcTkbDJc/68iPqXVy3hd71RCGSDIJVb5HpPDA2VzC+ZWRO3/g5jmJ10W0urg1stckgOJThgdTGPLj3COol/PFMOtYVV7vqQXUsnIPd+X1pcqMcCzhvkkgZpFlWEE85E1B2Yl8QsS4El2j6GqYu5Atpjt0i5w/gvEoRx1tdxSHh5hzyJOpOP2fxUJReQicU9KMORTOiJhMzWGMvn+SVhERNOtF3co4hPE/s4f1f1O04GSrTVjbOS0qnIhbbMA5zA575jDw++ZkzgMlfEfGKfQblBUvbD2HXA7yECYlcV3pg0kM+U4CPFSa4USC3sOWCghg1lNOH9dCJLwAer+8p72IJjExFsPsxzXzjixGUpqOXsWAmYg1yhzdVRQQn5tb6o4rAIyrS8N3UT+gOxw6lDYVcSQTb/PwoAPpkBQyjMVGh+CpsWgJBJPQxXwC1A4YBKKnWlQa3mAqCyW7W8lTWEyoZrD2cLwdNuvNQ4kobdMSaTpreGbFahs9V7hZjkcKpV7MVMQjVq4q6CtRisDbgca7pgdr0rDNs7RtFqfAOR3oYdc8BlIWmzLBM72QQu3IRDJITRYqRBlpxBW+Ep4SIksSZCiw9YJ7vESIVF3FkItErFFuQu1LTUyNjSEKa2+HiEZgEXHeDYox10Zht+zFrB85XlWYaFeYaszsrc+jKC3REuhx80gl55a4kUINf/ZX1jd2sjFtG6pUXtcx5d0kjaFTpPJCuvBOWGsXll4dn1xyDJk/T5EvZxDKNI630sbTu4Ow4NqOts4SgEPs1XvO/gaMPBKf2mh3iV7r1K6YiPc5oNBnyk5rWKBwmGPIG+941FJihuPzZo8Ix1l9bdSO4kuqNXmPF4Dm039nMzkUZRDtGGqldKg67Ext10zALzhJfnFzbm6d3tRIbYSg2SM6XAJPTsCzEYDxUJjkHmigiUHW3Frjk21DvQlcPW6KuImwRZ+5cDuWhigaF3xaYtKLkuPWB9rCAn+XVifv39K4AoUbSPLoH3C6+PlzU761KEho3WQjH9SWdv2fk+zhQS28FQ+XShJbyW44/q02FKt/Fjdzs7FRrdbQW21JqbiAqEZDKBiMve9XgnzBfNaK/F8JoxDd+SvD5Qe37uxlaus8bb+XW8v8j3V7BA7JaqXbjfmBTcyagRrfB+GyioTRK1CGrZvtfvykyhynucdaAhSSNL/jk0kQcghkNlRL8du6Tz15HZ8aVj1lA41laaD7iIAM+pGQ6hj3NVuqYXk3LRQV1FaC1HpSyWH0kpSXLOyuOZY6pZKqxkJ4Fs4zyjhiUDiSzCdfgIjWo8MMmIvk8oTmulLgq/2Og44g6t/k37SyHgSzMkAho3W0eo0lOnqeSIN4kfCH5NLDcYRmrSc3aImF1WQ4BK3TSQ7DRalMvLAM1cl5NXpLKuLEof+jH6glvx0E8WcwcWUWji0RAzNoGmd9dIb5HXTHL9XZs23Bp+cKlznEMT1Y+Fud9LGVCsTAiOpX40oprkHJyYAfV4EUsHcS/DTlCcBG5o66JL8DbJ+lzUedTNyDksIGqZN1ApW0BwzurCiBTyCbD5qRENpSvo/8tTCz5L+UfnFzfKF6kFU/HTQBNrt8U3a3SDiWxpTraU7tZoVzXDHsva6UcUi9wnG3Z+jdikvPHkWy054X53WEgvaxdUNXz6jgzGNWEVTkPOvRQ7lP6x2fRbz4t+z1n9BKBwXDHjJCrlLLwila8x/Ow7ejAS6GTxBtMwjwOSKBs9c8eOM3/VoT5nz29eAR3BWFa5Al9/DjIbFF3BXxwHbilrtq9dQy5I5NIbhBD8FwgH949RQWNn9/dIBVsPuhnY9IEhrMnN3KvCG6zesv+0YORmHqGbDQ7ypAZBFxFCNJBX3Ep2xTkCqMjgv3XUq4wDDxYYm/L2ryagJ2I9CLx9NP77shY74WxSo9up2b8A+DPgtNKjR0UEzT1f9j9ov+Vpx6mgD44NDbe2OsfXstMFZX4fRH1iE8LyaHBP7tnvTZN0s2G2nRI/aBR5XlSCQ04eGbm7gmazi1cK8pVNwh2zL9yJlvm7Cfr6r8X9TNBZA8XJdKJRMIyUGF+C53G8Nb6qH6R3KbvFMFFxSkI9FKDgIpV50Z271lMROgQ4UmJIgIJpRrcOMe/BW8CgGCcUI9D4DjVMvnvYsqXx++3Tl+maqoVL3BIQuKk3P7QnRBkqHT4c66/Y8kC9p7CFmLgfnSAdXOyZBlMViXK40t2PKMgeWlVek8ZfLh9IBF6NHUDobJKq0aOnwkv4kfKMt4OQYCDlMcTK9iMM7lJxEChWVQkvhR2gVAwU5B/V6ao5QV/Mp4Oh3v+IkGNKuIGlT6yxPneSPQE4neZ6vuxv1T12MMW7UUMswyAey+0gqoPtG3d24auGBpJZxxh2JkawuC43rpON5+pXZpqALMJ0t/Qukw6UqAbXPMoVvK0n6PKoi8vMF0vFZT7MHdit+RS5/ELBOxx3Zh1O8s1YRUZz+ujYOYl+/Cs4eKD9mSKS01LysiNkaSghmAR3ISOroTrSNzUQV3Z8OorYHa5XzA40MBpj8dwhVZ1GebA5Nlgdpz/yuCTwq/i/s4ao0pUy0Po0YzUhSyOuCrAl+QygdBfGVqYiULV1SNu0NHDXNeh0palSZMB5RxiCKLZP9poSv/t1A8+dvuGMZ4n30hLzzi4ktMIjXe+OpzPJOfY2E03qndtvV+ZN6BU804ksYsHIuvk9uf2GFabp4uayqvx5lp3wNht6mT9P/pa0GFciz1p2Dz4jI/snm8GqORA/Wqeg4vbFuzR90XbXNHpOCn/nYWBPrJ2fyUnEsjHLUy3kaJv2JcOIbRGyBtjRcwLG1DEHbngODyTyYSc/MRgHfMr4m7qNCvOv+5cDiQHjEUgaLrSimTuUwul9WKYiTLTibKm8Db9S5O1bL9CrYpkzacgHhQX3DvAD/PNJMmi6SYCE3y78EL77uszLFdXkt82DzdKpFXSW99ZANEblSntmutIisXcRbqC61G8PYHB5MGKT+b3wD/Vn+bN5yx5LO5Oqah1MuiaTeeKgRLZREtxdf2IOEQXeulmRzShdxMILCSyWimrc6OnnhLwwOotnKErwN1VDLiiZfiWOZCvI6ah7VxTJ9tTrA8FIMQbokd77Z6SNpmtxERvosgFnrwjgCx4ruX6pCbB4G+Av98oYX5mMXcuFo300pATSFkutGpf/BqiAqsem//LWS30cf59aLDxABWP4P/o3NsJ1x4fb4FHxSxrNKk7W3Wy6+a5grpZcu7vtOBlxR/LKKENTsaylJ8AgQHkpClUW3dqgk6q969W+64Gbq96GVwC0qU768NHEIqkQMm/jnpLJc2p7mtgpTJ8I024uytwi0abD/Vg8UlerbaWLYQytoNW6Aa1s9WSK2UN0jXBcJOLkB3qhABTIDPgBLhUz/gVkLVq+FY3xyMx3Mc6qkF3BDAvEe/9xW4ypZcg5aUc6UlLhGg/kRrbmh7yzFF+8ovopdyiap1q4kvR0M26MZA0HCnn9D51nc8S0mS9nZHNxW2p1ULeozhJD/7IeS44gxsK81v4fDc3dyPkx3gyDNxSYXFaGk47yXI7DWglqmFTktRiaYDZDkol7UTmeIqGXzv7eLiaG+JiwKq5jG/MD0xZdDY4BvVC3dwKdLRILZKtOnr+8R79S9UKgZjIPylFBR2zPqKg9tlwFwgW+AQbV+uikY24/qnTZ6gjD4yP1u9aSkf5a/3TgsHtQyNqVIxLtfczHuThIxhCttITOUH2GH8nKOzSgC65FAm3LZqSdzdIiCuaYVdyKGQlYeuT/mRYvGNaPgSCi39j25x4pYM+qTUvvYST2MIUXMKZm6BmpldfX+qpdKZlHFyM8C8wBfTOZ5cGZcVkJ2U7GOSsOcFsnf02Gdxh+RYDwp5F/zRKWh9vZtVof2shnFKpcSQzaoJzk2BBp7Gxs7ecUTpBmGeSQQZMJoJoCDRLB9C1/ivhGx11dfBR9brjIInMXy+mHa5GbDkG2uLmTNIL+Dk2sgWru0+Eim26Hl6idODxn3lrqQfgHvCjIk5n3Ex3ZN3dypl/20lsM5i8/WnjyVqYIFwMziTUOAv6Nzl8+eFT4mhUbjev5YJuxRLrjAauthX7fLPDj4RwFJ13MiMHtQZB7JRQT7jxVOyFWPD9VyNIMt9IslFDtMZoQAItqHKwsJAr8TsrH4CgsLN8w8rEBGPtVK9E2TeZ6ENCGgcIo3PiqNIccf10q544kezMe+0zwHV9ka5VSK7irBER96CRy+EFbdeoMG0Nho3i0kjThDc3LOwpHA6W6C18QxaC0yevCffOsrNy/jQl2xjT6DPF2tytZTyjpDgCkvRPkP/WPtJnLwg1fNLVc6fh9/h91pJA+2Wrn4hC49cjbHCD4YymihwyXfUx6zW50ClzuelgUEpQLHW48JDtG0CjEt8ZsLTfXln8D1jhxCjto34g3Eu3/osOXdPxPxovQlXbSsgzJAnnnOizeCVIgigkyaxt4rHzMokFE2BY839S8MXQZTTeqi76K+xBF+piPB5g1aDEHkJBsq+sJhsZVakQp2TeHVuJHLsLJ8OS4BtqTQaAESISFXc4Y1pPZ7EB+LA6od6Wzc2wWGGAcDuYXWczMdhqDHcd5MC77IZr73nUR1LpYWFzevSh/YX1hfh8UK/vgsfWMpff8RUEF7CTwG8LcPT2Qeob76FLl0XRIUPb/enPkoE8leGfZtgTVUdbqtAeSDv0EyrBNQMJvZc4IRXys4QkG0olCwzfoNlGIIS6k8CD5KZdq+ANnav+hFIBuB7g7wfEyALf/T4sBNzv5KYfEnqKS+DZQwcLEq5IVpkOcI3skXoNRBdOS1z1yGMtRA1mSrf01REHDLghP4nD+Sw60OF2dsm5kBvCiboOMk626RiSgWBEtbeLeDMpCPqgKdpUAOdKjtL9OeWUDEcQk/hddOUFBiVdNcD6hekqDNSniF9Hp3eDrY0i/EqhqIHh7/QIiuHff7iZ0uiJE6Oz+VcM4HPIMX8GqOi+RbJAG2xyqU+4lF9Tfy/bNX8FtIs1yy0zRCK/RvxMrSMR4nNkW4cyrbTd8wVIulPDoUbOY0Epx0AM5YG1eWbdMzuThdCmFh6B5BxE5j9D/zBzotFM2VYAYTBhfM3toInUYcvxgYvTd7nWeSHnIOA8hxfxJyhh7eTzfckGyp2U7HtIzex9bR9oBY47EqLRdCrUDE1qnHIqitsRRCAr0Ji55oveWo2aI4EVMXyxcdv3np1quY4bpKC2FfowTrNOprMpvJw+fxonvJYmeSPr2DuFVDtUj8jg3p7lA9UBfh3r2qHY8/Rp0qYbAZRwW+Uaqt8KuLmsF4//JShGA3CF8nvsZqjOFzQ0iZRFTvxpj0IDfInVQY2bXDKqHzDdaSJjAEPBcvFLjaeMsbYCnQzUcSXQyDZ91Qjjmz7UJdHu63nimuqRSUEe8slnIvyty99aufaH1rqZFQtWboo11chmHlZxSSVyfhoxlyFjuaiCiUZyq2npTkqC/q7kQZurNvUbR4FBsjW5uQrHIcrUE+edefZSghRSY0Zpo7i2ASqCrwImd0+woejJ80FRtZDtg8vhNJOuwjWUF0y2tw0oxYivazPenGD6QokpP5QUfR/WWenW6SWKAkPjCQ9InWBsfQhy1lEb1+cNEy+PwRLAapqAdfNP6y6xGO2xusmk6xFtyebaTO/rSb1hScvPNCLRqNd/UQVl5tMjuj7vthWDlG6oz0Mypi6ObOfbYYXEhuJGoeLh57+jnu3CJYBPsWaXjJ5ac9G4giET9Tl4FDzoEazjQlCJNO1eaV2FOSO6jUZXfe1fqq/1ptjdg45A9nQN0fT6gFqHONgBjxxuK/474zrm5NgHiHdis6He40KBQduTGVy0LZ2F93+jpga+WvVsQmbKjLBS4S0u+T6i8GZ8dolXrVX14k2mtqF44yLYn6b+La4tzcDr7Mb5OmaIpSJVNNajJdk2P6KFETcXOZ/VJK/lpQKnfxQt6R/4N1adJvMD5qb3QNUuHLaeIJGgmH01rBTUn4+5kikp3MKPYrYvstunlpDPK3HJ28IBcx8hJlCwjkA6pr8P9aO5ilunw0/NUlfYL6SQDYE7gMBtiP7f54XPw1t0OoqUmUgD33jS5S5zGWDThJZIhDHQS3S8wLmhZvtbqsxIzuzm2JkQ9FN49dza8bYvZRZ8d4vNoK4UU/fVZUX7eIHv32yxd7OEvfnXvcdtqWwmiBkqg0V1pVQsFTHSXy88F0z5jOnwAGgFsEEKP3LDudHIcLlCpboJ0nfkNe3A8a3CzOnmyjjje4MdhXEujmyAH/mBhrPA3Mn7Y8ifSatrkPEuJ/ri/chQs3nsAKcEQSl885md39G9+WosGlEOSo+INVfqM/QxuKIEvcPmCryil7KLnoKsC59VE7vPOXLtcYCWOKBZTIcQCUbBZk3dde8zlMrvFeRxNdBL/rZo60Sylb9Hg13uaG+svm3aWQNmwzTdOeTAhDlks2EXQX3RGOFO2Rc/aLJTh9f7eKbdFENmut3Lcy6sJ6ErUvrmdI9dv5rWnW8Feq4l2/cAlHOt8zeQplBvmBX56ieb6pWZGh9maJOKbB9keYKN7CRLBBxzcmLr59eDOtYU72wlRUnA58jMC83t0X/sGveBhpCTunHyKtZBzFndxSWWrRgznzfHNfpwhYdm+Tu6Y9e0XJF6LhbB2r0nAKW+TgAftKNSZjFWfoh3YnhMleVgqRirv+QWb3YD42ZXigldTji6VPVSwRYOpqK+0Px8T/vD76iuWTV1XwdwvmRe6wMHiK5IVFcJOXq7L5yKom4qVdcpzeLfTLKel2Kn35TiYZ5qcDuZ7WZ1DECVAh7RkyvkTZ8BE1ORDkGRhiufHGCMjLWPQjpYbkWKXS7OGbqPFldQQ7IcHucZxSPdUwocR6XnSAJw6MdlThghi5DRZHgzTPgS7g8O/7ZQ/mlzoNLi3JgCvrnFFY2k/rqoSVxXojozujPgIqet5IJOwSYVZEYjNAigxK86n7YSpw4LWu+30q7xmS1dmts5O+KJ3hsGF+ZS3PQ697UM01A89qAi5UrIhWK1IAqed2SjikO1bvgAfXtbMo+GD7peRd0ehHes4LAieUJEXES499I+/AjeK5ReQF2JSm4f/H1We1Wpt0B3piocsHnCFsMb+/57mCoJe+HCvNCA29ADnH1zEC+fEThzB/MuA5Aj1oavskv7UG2BilsQ3dNzPstUIiLs52tCUWKnFzAAD5R87XJmfB/kUvk6w+r4MU1OB6xB7hSzpvYBVjsJu8T6M9W3/4CH/Vbun8xT/2kBmJpPQpFDb07SQu2KQZp7YJFUwUmcDy0Ar3jtzaKZoef1r8fK9T/FO0hakxxL1jlTlkdGlYow122uy7l9oxFHdpZo4XPK2Q9E0c1lx+K7/gP3KgYyQcAGBmwBVvffo6sZJkBgogmhdqyoBWvbI+XFlffyFxlbhdZru2EE9qlIfObdzjYB29xBVrW5MDtGTGmuE013RsxeAoRdGYSXSlhyuJqyeBQQNvhcLrusGcAMTQBdw+arZE8eUX8djcOQ4JV0lSrXYH9cJghD6YZRpCkX4E5NJ/TDe+kRMG/A1pU4CNwqW4r3udOfltl90Pi85B67Jj9AosXbAoLQHIjwhJJsiCeTv4+8k8712jIdCJ0L6C8RyFGxsM20kh6smu3rkKBz9m4ks10rrK/qg61JM2kX91vVeJvU3a8dmAvdWCGASNPaULiSAMcwRxkafNwjKs/BnmUGr0BGmGGtHLxZzWyzef168nCTnzpSKTKEcCkM5L1FPBD1IJ4zKMiPpDcFO48hHFJ0Vds2PBWP2ZkmAlzg/lUhnWRzgoW4AkRRknEolC2G+LF9CcmGo4v6ricOv5YVBhZokVkdci5A2Pjpriyy8JzsD+pwEwz8gNec5kPoBqR16p4QtJ2W26No93BQ8NBCIy7nlgUENCvxo3mMeahY59ImSVB6WFDkCt+im+G4RvWJNcSzpdqWiVUxmrHobS6VHfm8GrP9XA8F+cGVRFCgNq/74X44KRpvso6qbtEKwJMQKLE/XnGfXUX+hSQ78QmughrdQS0Lu6GX6CPE3G70TH11rFAMzEvcJpn4f9RTqtwIEVOksyW9pynsgmbUvbEbQbET9m2c0J2TQXqSAU5qlYCQ9VCBjBL4mFMmwgf3zI7YcErTOTGcD0s2/FoIZqdlK3aR2cztP2r19e/5isvs+A+v8mduZe7ooog+G/qp56uLSIiNibFgzr86oyxLqC1GrWEoCI3gwmgXkRsaymyTp7hkl3TjXH6MY3TUkKz8+ec2g3tRkNBtOjdOVorbMa6qcbAN17k/b5UCRhy+Grtw0Cmme4ZiN9RgG+SEILolae0sL5Xm+SrDf60A+naRGvp2Tm9d/C2njITEfpr86s8z/ecF5Vktxyjod4+l9pPA4BXhJOJxclrWDvBTF84PiDkdf8cVewLk/SyU5hUOEE8AG2Clqhjoxb0T5Q2T0jaY9igxo9CLG+dKlEpWEVPBNCyhnM11aNQR1MGOrmG1MoIM5VNFJdEzG5tM3AxKctsW9O8+pVL5hzzK8+DfBT8Xx1sj3XGgvJ/palgMRRC/AZkKbFAq+QjzlPv5IDOG5iqC6niCODs5PBsWfKUdyz+x16lanVkgbVHhX1zRIvsihdem+iToP2k/RjFovAk7+x1nAD5/xFpH1L4W4E1cdEA40uCyxxDXIyt2G1AG9vuE6wj1QVQXjHDTmJaT1zBOATMhgkdbsIJ/lrUQ3L9HKIJhvV8ezC1pJioIx4y1ZwlJIuMeHbi0m5Fgkt6g3+Jhe9TrWo7VSlUTdhIsit+nJS/x+9hrk0qObvswFy4ukJ+AvAVyIG6aGRgbaFNYKVI6pECbwlvFIFLTQDX5scqc/hM5bVyv/drtNS6TW+5Jd7p6nyltId/91MO594zDCmzQ6poCF7q4d0ubVmtI52YoB5hOQpoUOP4pC7qdgpFJ4FUlFfzXbnOW/14EPKx6ogs46/kTbmi6YFVFfle9tsGmlV7MnNyrm6XdQp31KaU5qXUz7reZVuv+D9cMj4zl6PNSAcP0BvfGV6TLeHDvH1/F5vn4+EOEi5k4YOuqa/ZOJs15vCePSMktdT9pxsPUnKT2zGVjcrgvzLUdG507ihvXSTFtn5N34llB1egblsDXo1l421I19HJd7dOQUcY/XPNElPfymVDA2zpRbi4xJdIyN9cZOx30b/Som9YuyY/FAlVSU288MEL2NDSkTQAzwAjqC1ZUKCbO3YgxoNU3ZVQ9BnYOKa1kyn+KzfX/LUWxf+VCN2ISTJ+J35xAW0Eo0E6/cqlZYbfJRBeI+koV7LDyEs5KNgsMmC0OEc4Bst7OwDegVtDgkoo6YLfBFwQ4tHSUz60I9U0+5QuyJYEXSF/xkCX8B2OXsmHuayqlbh7ViLluuft9Ii4KgHFXbzfMUy/xSI2R6pKrM66trW1yYDXtNGC78hbSWGVfQU7B2dIgcwufX/MqbiPIH/lV4vSLqSHQX5+ssHxiBe9iNhrL+jefdKZhZU2QEzE/sKhzXNXmF1Nr0hjAQSHwhSqncEsIqAnFMFTJtFFwE+8isd9g7A/RWl5v5S4TUiUtW+YMN2dA8QVNhb7FgH/9+WGbcAV/agec2GNR2sqfLlcb/wEClGHvDFgL0jI1ObOLoxY2zAO/5wiUsvnpwF3Tm8HkPhYSsFvVfPVVpjHGgm
`pragma protect end_data_block
`pragma protect digest_block
5f157034633aed897f753696c4ffd629162a9330a83057b457f7f4155ab147dd
`pragma protect end_digest_block
`pragma protect end_protected
