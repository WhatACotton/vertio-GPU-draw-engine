`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
Ve8RFBZBGG7+s1th03wSn4Ergn99TfllJVQ6YembtTi7wAVTFs0r0b9QJse8fWYOgZpgZcWsks3eV5Da0sTi1xQ7CxA3lZ/w+86jFARLCf7yhO+abjuNprF53AsgGtCX7UqqGciSPA1jKaGDWx5uCoD/LkjiRYbeYE4W6vHXFE2FYR19X9uKRFEjg9nY25gzYfYdGcbL8eURso/zJcR2yM+JLdTXGKIYJG7lHzowE4MU9f4iRtcA2WEZE5huBMCBGXPveUxFXtkhvw2bhkdp4ul9kS3GcuWOEBHrT6s1FHiatYNIUQ1MVjLu/mkhYM9/7LDdLbh5C5EY3dJRMsuJrjI9GGxirMfhiMFNS/3T6KDsO7mTYMaULlDr+tLt/JpOF+PXAc8MQWn1IZBCDfLyid7NdeTpIBFvEWQxTjxeJqrWqmwREhxgmiG8mN8Z05aEyv912sYYO5YdYA+op60f2AqMKand8I6I7GB1yfyC1iEpN6xCQAeVieNH6ozLHi+1EyvtTBQbFGTFAtfDe444V2WCywpkfNwRFpgV/qYiM+yipk5FDd86dSl82gNXpccwj4sRiFsAvTKbHcrZ2U6eDAGFFputRk6w41aHDQ7lZBHBUUJG3i6aY0qWzOIu/ZnkNdT2I5QXLYBc2piRBSXryzhAKcy+Mdcz2Xw2HfErwW5YL0AQYkO3qq3k0CYkZH8v8KXmdR3d/FN6+AdtyWNfA2w3KjPlUExQIUMNWGv/1h3EaBtNI5GU0yNp1muVse4KYYLZ1mblUb0bBHO1y/UZxaTx2p7htTD3Q18Rs8ItMoGRjdpH9ve3CPdXBrW4/3rRB7ykUKh5evxqHDcDaO/PVcphzbRrQ47ZJG3xHxwbVm5mUHDffyRpZ3CEswKv/EFLuNAD5qxoH3Ey14OIT+AIie6inxmDS0C2Qkn0BKLTezBU1ZBMgn7I3iexar26/H4QVhlDK026FXQu+ASRH6kAMjXQsziHBMwJ65W5azK+uwnpI7ZadeD7jFYNEw9zmDGRtBW6v5FfESEEX7RRYerYDAPtBsfRvmB9P67Mvb/TzP8Rb5mVaMZQTElwDJzfBc7nyu5K+gUzV9etODlY7Fsp+2RKcbxUG+WrchjWsWy1cu4q/OrAgHAyKOUm5saCfC5GqFbABdpaKXCww2rY/PsMu5Qw/hz5+jWh3hvunp8pYqz9mIMRIN8IqjUxPysmaDHPM0LEtapB131x72I/Fq3LTyCpCTabtt9UAKF3syPSHWKViZQkJW1ZCMznjsJModrrpZ2vck/eLWLaMK7wRoZ4QZbgiBI5mzVMP4+qIKHqR1MTIhe8ElU+HvP3w/QTlJ8hgYfU9Vw7Mewoo4+fRALaRKHRtBFvRhIx/XjSZCKM7zxxno0rBqOySj+kOQ8nbFw3FjQZbI2hJldGiTyL5R0zOdtjkUZFY7FWT+cd/ebXWizAb3CcMLsMA6P3JO5HA0vbRU97Gj6bmPEKXyqVpzOw+Y7wUqHsKmrJAM6Ah6HYzcoIb5uotqtD6lCKJES7JaOTEyrSIFZJKH8bSuTu/L8GkYx6u+VSupW8L9XX8xb9UNNPHEYr4Wzo93uHokA13XMBoWiuAIUM7jKo1vlmQ9bsUPM8M1oH15hvZjgwI+Y2YrDAag1JXsaJRltk/lSY+fFOOapAny4P6Yl8rhS/LQziDpixOdRcVO1PU6Im5/MmoJhrjkIlvijlEOotRGL3RjfaRT1DGZexT04OFarzwjuC3ddsUXfc+M1iGnshavBdAVD/jXMahVuA4gbZRwb26ilEBa1ZSGSQbyak+km6Wb5+L/9PctNqZ8rApkZfZEYAg5kM/G2mmbaCujwphb9Z7pZxrO8PN6rBB3OLjNqidBoAAGxldLz4a6olbUmbPxHxBmvStbzkR891DF66roHCtgDG89D9Yn0A3LQl/omSpVSNACeHJRqaOIgNsC/IA1OoyDSbHTEO0KHuqjOwnYCcg5cMR3YLtCv5XuGNJGzZm6+CWduuwaBx03xUxO45n7sh5YhMTskfMmsPFTCMfXP+8kM+458JshCFRSZ3pTGd8rApYilGUAdFauxKlCaGKCk3vIb40jdOz0tvv89f3+2QoVrBRT+iMmHZcDoG5DzwpHxXmpOFZ8IR/1ZLzSgexNEnBeDuDaR+GQGF3LHKfbtY2BYi3A9SQxSKv/CmiFOQtIVLy6ITLCakUGsZFmkLhp4iJR7lrPYz9m3l1ab/EztwI17gU1iEkfo1hpJwqman7p970hfAiWxilp2NiTGgMry9K/Mnzc1tb+MOcIAGlsjsYIyHyCps3mxYUPp8YxBnVDyYzKkV6PbKvtIn2rNT/Kmyh+3nEESz9BLVutIZVtp8/2dpSWc9pHJuzdJoIjh9sUKvHawyrGeHufRgotLgeBkpKQm4DQqS0p3U9Od1ik4fJQ9Odj8KUOfH2kHBl3E8nv30qPRTk9BddJSE98gBztH+c/2pDmW14t+TVmA1JQ82wyCvZBQE74gMA6RsKO8dCtZ3H+86BXVU25m3fJwIW6bNzZYazvK+UXlnadaxOujWavalP1bz+7iEDQ2DFrgPnewHL1DNPq2DwLet+vug/JlSUnPmQXyoFWVxQuzCeze31oOgaRVrl1ve/hZvgl+erPUYBVqrITg/s5vikojR1cJGGK6ppeCJ85q+szn+Ekztd8KM7kQVXNB7fZDk1EKVXmv4hMFRss6zQITM7BQr3OmiI9YnmH2Ue+3HwBJkk5iZB7Vyy1skO2CMc+KXUj51WnDCSaRfC4OYTl8fzSMnolrfWGPSOFComPZ1qX034zFh1IHZzP+T+3mHeW2LjAIE1jjLKtEOxebVIAgVxqv2cc8KCvP7fMlxev4uKGxs4r7atGwjsx7ERYKP+KF/WbKdQgkLaGVcYgM43ZSk34MCcGDUFQMGlaHYsd2LPTkqoUyrncSMoG/bzX7ZjtSaCylN7wdxwX2aSodgugzyk469TTW1LLPsQhUq7rTN3fhTAMcZFasEdcfm636eywbHKriUzMZVvaIi797Jbp18tAPIzNBJ+KoOunyFVICnEVfFbI7hImsa3/x9n7itQlr7IE+DDARAtL0Z0y2n/p0dCjM3h6gyed1HC+2gbwlULiUdxxaZCFlM1sYG2dqLTcZrurLOcxl7xsrm7ZDtgNtddMK0y79Bdffm6AMLr0Hyn5CaVHpBu1t2GgwnOCDSQOk1W+VJtvv68T59t+rtkBrza+aPcNU+NzFVv2CNZqzd9hGab5NYX9yZ79od4X4QvGUNoBhsg5G6aqK6qHvvos0dw3oCS+hdj0d4iKYm7a/Y08361PqmjlAWb6ihdrjuyOkHtUY6VPD0EKzxlOjNi7lC3awQy6re67aS/XwLxpujH6jtJtAhFXifX5qETjKakEDHagzgaDfdhMrSrMTygot99pAT+oPlUXMv6uzNsmfXTRKpX8WMBAG0frMHjm61MgDLLYxVAHTwoS7sOGJ+G5KMxRvvO1sJGAk=
`pragma protect end_data_block
`pragma protect digest_block
63b68bc38b9c1a71aa2a783bf8eb204208a3485ee2c645d4a765dc57402e7834
`pragma protect end_digest_block
`pragma protect end_protected
