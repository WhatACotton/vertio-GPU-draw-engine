`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
T92hqEZhnOUDG3I2EFEkmKFYp8Ndcokn4/zhclIkU5Ih0JF+BDe/BsVoAtdbjrN7tKdLC9MmjsY6CunHbTtJVHbqUuuASpvcQCWPAVQKl0EOl/jGBk4ICuxQASVjuVlXmw43A9DUZNk4IseZeAXBFkU6cJFSnxafqYvNySlLLP8HzPxsU1exs5slp8zGPf++7kmK9wom12p6G5kleahvC+suZilKX7vR2tLBETpyXaTv0mTx7X4ok2rX4r6ub0IIc1al0Lw1t27qIsBhWSDRnqBGRK5ZeQAJtWhETVWwUJnEftBoq7e3g0g/rnAgRbqQ6iJNj8oFhbYBKmkk4hPstuxOnDcgbXFejF31JbDzAJfVOI9FD+9yMaEXGLOw8gJo7cy9+Rgr3lGJwVGpdbWDIW5RmnMH6LMn4RDhN+nUS3D2+NmQEPATGxF5+BDItzn7fUDZC97sjsJM9fkulcksapAWEGrjG0G6PsS7xpNmeVPY9kA0sOYecynly2SjLNjpF5A1YoNKUty9Mymn4FPeOMigHfEVP5V2yEjdaiDr3YwT8S7AH7UHqwXtqefY+/HXzo+6YcsKn4yZStO9f9A+QLzxsgWHJPu2IxI9lXbAZ/0cSvWmmkHfkyToRGvcAJxBb3N5vy3/sFXn9DoII9smemZGQEiYTVbNPsO6TuoTPIw7PSYz2gxXiF5Vz7g/73Vy0lGIbiX6iWRrQzYyDqiUUMh1xE9C7QbjRvbLrlrlkXLJx3q5CBqq3ySogTMuBl7omNtjpce3g3ywt0A+liQTamjsl9K7VWqFnS/CQwTjPuDN3SVSMeAs0LAnarg3D8eT2u1BfYJ6H+i3FA3QwPZ04ZsOtZ0ONcGQle9rKQQSnUNgmEA+L4yCRm6sEajVYYKCBK8F/CZbO+9WIhC0wrDTqBea8wWYvnkvFRTuBqLO8q8cWu4XoJiavvowzunwAOxrIN2Oasf4BqBeFQEjfQfYzZNA1Sk27mb1whHREJfemUppeuVZVy1pyx218IckywRDF1cReGVeCWQuU1XZ+tQKa4ET84XrNQpB0cezuBrhUDTxm7TBIQC2TJeVPe/p/JWVVLzcmOm2aeCWv9D8iuFCb6SZpGX1W2w3DEnVWoMoGWZAidWCSZEhZHFIJkoNZPfPOK5lxMFZSgFByJ2HzFVFlA4YzHo5pC3fVtbCvVsgtHQiXoD/BjS2wy9vT2S5O21u68QV3guwSOjyjPy3zLHvvu5CCeIWZ0RkbxUVqULE0yw3a5eS8W4gL+AfX7HpC7fK9wxJ+wdzJ7nhk50L04taavEKG/qdaNdKXHSAwQ1jNw1hQ5hacBOL0ono9Z9BeQ9OIJaNylRUxuZJR10BSEhuVYXdkiek+nP1KsYUSYZyByCZtOCfEAVzmQNaAH+314UBnS0lCq2DofROfm3CzQh8qj53/9iJgkci006sKhcgcsixfrn3TRyeGbYk78h6kiGMSxwn1yhkEXCtHmWag/wzywTCHlqWWuvOCoCvhUSx3vrVB/Bz2YRSbAOysN3pMVspnJ3YsSdyW8EuJ0RMgVnW/0ibH8/903I1QlV67bzsty1PdH1wz70gFgGWnA0H0YeYd+Jq/3DBLtVdK+jZSptI7MeWMU/6rkRa1ECDYlOO+K0Z1Z4H6HCYxj+b1BHVobvw6J1uRhaPzKTPU0xwTZoCjBgSRSXAJX8MQz7uTaaLs0ZjYGR0RwEO46cPeZnGa+ICyofleLWOpYhkGr0AfhhqdIS05dC8aUABvnPZ+cHXnqW9AiI2AtShQrQ5/g0zN3yL3u6V4ckJtOQDKZmzJ05BQmHWTmJYoAYog8WlUOxIx1YXf+Stcr08BAx3wAuVM7KLmv/cUuBZ2Gd3wQSCcNKKcb1XmyBf/Q8Q91DxbyRY3S+9wBa+wjLK9sY/aqQ8FruoY97YldIicVrkPIYNQaqaDOo3LT3QI87FROpOJbDx8NRn4Y2sz1+iGiL4H7nrFfooURYnQLPH5brWjC8n4LCLYWSlgZ3trfnmzCfYU7wblqYrn+pw1eXHTonWKNpY0p+AkDdBxEc///vuMzWYEXkxxqTcjI4scjJMlOSvGbtZvqIjrb3rhBA+Uaf/OeUE8CWtZRlbRKPvfK+W6RMCSr1NC/6lOfi+Myrh9NH0D0Wgi5Q5Fuvb+nnf3j4gIWGQK+KQutfOHt3Ure1hDcUjqZNMWOTClmdrsQsxve0QR48KzYjxLsvLbpEC7NzUk4WIqpBGzVqD6uSk2AbVZ3GEDriN6VNzPBeL0OMpj3qCa2W5WoM8zFmarpyj2b1slUiTIl84mq8iALY6CsutH4j86YOxH/woH4/BInUIDVevqjQnFoj4c6TFSkmH8z/DX5RAL0BuTCgOVCd5brw+8A+cLF8WUJz6OCxT9z5R1Sjcz6b3xxsDmbV2wxMaYtxb+rXUQL9SrGmcQFBKBUv5CufF0G+yQNj4sYyh/RO15okdMHak8+ZpCf0uQO5NCeZfoKByhxxVMyxGq4JDNqhecmxvlcvI7TA1rivZ496Cv119aP4kxEMW6/3UtbOQY443KvZmfwww2Y1SawaO6TtINXN6yS5bhStMML8nBDa4Eeg8pRvJ7vQUybtHuRwzaLYH/J0tqpNwpWADpnw1zqIeCKvL+uSMUL7bLNuIwU/e5D1MqkrxwOjbw2bBzlAwDGulu8/71CUbYbYh+IlEP2CzdZiQ9gntserJbEQyIpRIFI6LebIhLBJrU/J8qoMiCBu+iL+aP9CMXLFU06e4HTBe9j1naqLfevfud2CrRUKL003cGX0UTlbT5gOVy7qN1BfQQT6b5qpqY5NarvyiokMHKgk4K9wSj0naW0zS1IIk6G4Swvpm50VXfaQPTOHl6BsjCTkex+XG/3liWGeULEKxxt1WBS18nkFG5yLzI+Jja++tdl7S+i7G2JMaar2/oP9eR9gCTbBbTslWPA11rkgyWXVdpmzmubgaUjRJRN77ZNFCNl38XZ8YLjQMbj3K8E/MsfB8LLRrZorwu6hQrs9wRf8sYm2ZGwt/h/IZuGAzRIdc3U1MK15CbVrOJvLTBYD6LhpJGPHyA6WmfbMRVZ2krmgxK7uoALxGaqtRerVTxEDqoQhTy9lTeLccdEO9ndR/Y8rOWJQjbs44FZ4hMDbcwcj/zlglYWofDx1xn39lZ7w0ztsgEz3foL58+6JQtcQ+2qvB3kqnDG4nfACsfKbMEE/RpDDxRGzVSZ40rFyWZTmAkaovq/C2H/d/I+Y9ZxjXIK4TI3vQ/Mn/dE6Qkfp5NOye5hrEuv2AbM9bgKivYvilzfmH2Z3pe7AyauO6F0IcK7mX/XnflDWAeGhCCK6QFR0DVK0vFtXENdftWlC8zkjxv5uuw7CNz+jlnXg1Ztrhrd9JKUYV/CPwtzLNCLEMrfaox1KaBBcFmWWASod+be8AE9gsaa4KgbTAiBZ22zUpFH9KB5VlxLMEGiwrMfaV7oXLOAKvUi3OczD+Og1dipVSWH2RmkgxvSMuq3DAJ3LUi26TFafUlktnZz3actBFHh/asSMwkuqKfE32qUB5rwvDDB3wquPd0eJ54EvquCbzIR3ml9PXk4KCHmAnzYjK9lNPVy7/LRqQ7SMFYMB02AOu9gR11scIfZXn99nXkLVBNMU0Hu+0t+11kw5WKWd5zGx0dZpSJA+H0dMDFQ0SxkRbPDhhqSnb4ykjiLO4ihAaquUf+6O8CcrETdDUKH5f4eZwGWhQJFnDU/Vpd/M9sgRgxWIJtOgg8NziELkxaFqaJwa9lUdrVlU0/BjY/4RsIPCA1Y3bj4yxVPL+ovJow/ElscBt8ijm+QGRzFd2RLX9AQYJqnW8E4rXiGdCo3fIgfI/iYSeiQIsbCn3R5wciCQ3aevInCqhPVpng3Xc6H+kfFN3cd42aSczOWFE9w45rsT3PT13C1Z3mIWixiLJ4vU0cQTEWd+HjyPOCcZoeTIhBQIpIyVJB8ZJAhEKqQOKrTNdvEmX4z/CuubYCY6xgyhl2L0R3SY7cUY7Xn+Th6vENyH8ineLMKrY1x55cP/mwEkpEx8vCyJWS5Gy3p9XeAlmh/hCA+dlXJgyK2UgpCWNM7uZykWQbOaxTBwMADZhE+i1tluwfhm6ZhgHJ78ONgp2CD2MYoVhmHRXxCC4GSIGkprVEJU2+xAzQZpNcRjOaquZ8LATxcFShHxZVNFyIh2k5YApDS0++lPLDYAVxykIK3W85ojZUkBQsSQA652vO9lq/59B4wBO150bQAyEVUbebcwEh2BWFPu3E3SkxTogfOw1jY0pW0r0FnWnc36EjaTktUJnXyGxghsi17DZV2WyMI6Z7OHr6drs0+hU3kKMUY6lLXQK5ZUAmt6iuQvyzfg6/U4/UjTRgHHVEwbBdaxAE7mcbYZmjtmavgtDCgmJF1TCHJmqo54XUs1sLswCZY/TtArt9gW1eSO/z+HWd9x7ZMBgD8k+ZbHySprxr0AIJyzKgdtT6BhTe1fHjpbtfxfV6s9ZSk/9gzV0rfHTDQMzRdYgekrJnm5Qm0DvUXCFozLqLqx+zkkSPAqoTldG9cUg4hjLsgIL4ljAboMQAmOlP5I2IFaSbNItC4TJeXCDdzkZkb4UBW+WT8az6uNnt4e+ay7SL6JKWZXafSpzJ2sUOA9CrFYsw8trH95/+MJKpfk0vEPqB+SiZlZ6MRMgtjHDtKFZ+gyEj4jxlYX8tTRCSopoU07+Y+6/8qy8qet0wUUceQI77/iC4KpUQnUpNcGjKozek5TRD0FNkpFe8tLIQ+iFC4zlfrOKE5TTUWAx+a/t81jA1CO5HLJhJRx+mhNMfYroz5PuAlk/mk2Itj0Z9RO6c4VdnY0nA6ZDJt2xAEnEEXXMOd7jk9anGEoENHK3KdvGYEW+Jb9ibITNvOMtmuC3n8g3n6sgP0xvkOR8cVDpAiL+6fCO9fvJDwFI8J9SWmj5qz718n0tDI6fs+fJRb+d7v4bpu6MFtbik0fGzXGapaotlA/kjWJNC7g+hocWo/IXy3cpVfOVguv1/kjioVS5alR4jtgXX2ksI3S1IZaZ6jhNfLtemCQ5APKCL1Z33qeBxxIjKt32WmMadS+K0qsZECQJ2CaE1kGPhileVSVgMzK4p3vC9YFd78G1muTRpvJBVbhjqHCHhrrC3DPSg1m+GZ09PwXvuXp2gIje9GuKrcp/ilpe+9zmYra7i2y81MTE9IC1SW6GkAQd8EbZmKxVREhWCpVkc+MskT2V1OkSKmK5UyushOoOHtoTG6Qm5T9vt39U190VYi5lTYz/qIPvzkVFjjKgi52XVOfInB4pbRRrXq1YhatDvTR+CGSj3Tsmgh+G7E+3jMkNBlmdzYYtCmQQlKNUn3QhaobWCYU1OcbxnHxvWixC2R4XUMz/O3kqPqmVPg0jtAmEeYJJFOB0zXKJDmJlBX6sGiJU97cD9w0aGf2zEtia2UovaDviWdahD+VSwb9bgvMgQNpR1He84ZdI3V/sz7OGUPd8L0b7FRkGI5LktyZH/pJ4J7sWFRcUFT+KBOIilTKxVbqwOGGl/EfTF+a5WdC51f/vbQd3enxlYs8M3iLwBPcGwRy6zmcEI9rrwe1AZ6p8PUa/YRyrZ8hWm7umlOPmoN+E+35I7FrWa0AR3fw+FAY2vakkiuJ14kpgbQVcXKHdYLrdE4JpWZhdcKg6SI34tHzYpcZ9nTym0nPUwu94dRuo64v4ncU5CJDxTjVD4aJ7O9rM4xkV3J6REAGXP+GLLgi1PLSGzYfvGItSI3rFif7/7ldoVUU1hmeTNyG5+h41f+iTfzQlylYQVKsn/Q8jdePSHhW34u1SBVcjPbnLwcxdPtNNtM8AKwHwZmGfujK6+jgImZPOgdD4DxNipl4TerCovEOZj9fiPntbdVPywqyF0woWyDm5mSWTaXWGZPqtkOS1N56TdEItwUz6DJsvSkAm9hfJM/b/Q63IF4T4Aw5BXGosed5D4wJKhxnXn/lHW8H6ebfqJuY9tlRB6+qW3CmuoUtRzbni88Ous7ocRQcAe31njZkPfTwtmrOrqaVkd5fEbDWp6uKmsOoMaxNNscTvPdhkXcb9ArX4pliFzD7QfWp+a3h6KGxEHjl/6zC+6pA9WzOi2TznK6IFcuQpNsr8lerwA32WXIgnDT32wmfhLEtQdYq4G+gNFO2gmxAtfWjuWBB2dYFRbHDh11Rnu+sStV9KyyYriUg8Pffrpeba/R33RNWKc4I3mkBDYn2pwNzfXAe1j/5nxE8fRIBKq/9hiTxZC/j6kC/z8Edy9Dwpq3KBdhul0feDzdeIzaiYF+YwKylyc+npkA1oQcKwCgysBjCNz5i4PtOLxi34tsjEAXy+V774R/8c8ViQywyDXY5iCzHc8h0wygL5Q/RGjn7n2/6yLtJHXyKJD+taWN+M7HTf7Zgh94gYsFeMKX18MkgWMh654dfMPogNQ67w3kZMPfhkRYLdBnehJflDCqghlLPuRWt4+MuaoB+1CeCM3CdHBzfIwqZH37F0O+S/rUOJP9zOwtXpvkoKD0bqcY7KnCyKKYn3EAF7DEGMGB7agCFtUlzmtqQcOL0Qz/wgX+7yvezIN2aYPAhhemYEikJHmYY/I5Z2AvWsqEPu7CrJdnLh2wxHXjzCK4jGWaeTfWL8GLjjdEMGR4SprfkkWYg/oToxYDcGrAc0Gkk5rZshdrHKxaxKS6wYRMopVhfIeatZ1cfsxDADvXavN989pdhjXIG7tYhsZwf48UPqS5ioclyA26DqXeiy1B1GlFuv17PVBuTLes4fNoz/fxIElbOMpr+nnJL4ckoaLPu5VvhxU2hsF62yATtOsZCcLtDgO3aE+2xxKxWch/ij0InoPtaLTTWHMr5bL9br271lF/IjAjTo2WJchNbmGrcrXSIyTpanHipkjxR8EYgJ+sSGL+OCV5plMCxhf6jOmlA0plPs3yb8QBjCJt1AjHSIz4iV2m4RgeV91R6ly/O3KWfC86Fnm4MTlMNU+pDidiAWn2kpUQeDSTupCzW/q+6kf4qUShQXFUG5W66gluOxZL5h2CkEvgocfR1ALNIR+ob1vB+XQOHkJ4eflzi6TwzxhjRP7NFYyvvzW3yj1+KPB7BfZFQYoVIBZfZjOPdiufsOd0nreWlws2Wbg6/RQcqn8hI97dHHeemzfa8vB1VQ6XdlNIWxmdvWEshkZTGLUxTXDLf+3UM4T8lR9ZV3LlOgyREbJ8ajw4n6kEwgCVdF9fjaR1ut+HgQIRWhK+8Z+2uOixjefq5uKRrMwXaFw2QkiKHZWSSXyOfRpLGWzJEIuIv/YtxeytJ5zT01w9anNxxMzmZPOT/gZ+oprb3PiAXN6c4FvVZhjR3j/DUSacLmFfNn5PIn21TCyS3LTYy8to4Iab8m2J/YINfI6MQrbxn3w/poD6UdRsem+/qUuduNudKWfR2FxfSeyBLkXOJYd//EBDwWp6tGIu+Wu5es9v1PlFm+5/PM/N8VJ9qrBu9lXCCZv2t49gpKh1afthd/wPDhYXK2B7dz+R1Bofpzb07S2MGZgwrdNQ/mX5ZdT7i0ckgRivTMi+FKWXuuGmt/6abvYT27WGsnpanFzcVF4XTK4ui8zDDilMQQgROItcdKuwHJuepSIcWThEvRnVX4wWqFh/MSWEq5B8vrr0UzkferZ4Jiwo0XAVodoguHkrNtSRdwCgxJ4GnOQzAyNV4wiMVVv34k85zY+/2lgB4i11l9U9HejbP/BNFcvqKfE96gOgNyhGi/58FQ7hD1n3dZVC7l9qLTmZZ5EMTWHWwaegfOqTsouRzLUPUyjLJQOSuCBmuQY09MkkDINV8wQ2fO6IYCAhFF613WozAVEbUl1xJoxdq3yACQwDszrhTCPqXpkl+j+Hk6/dLO5+67FNQ1hP28GFElsGJsWlRix4hNWMkajmGfGT6pIqNLkYhbKe7LvVdzOQWwlMQHmzmm56ee4VuYUWe+/51m8xLKAvuKfYMziOcZL4jYjLPFt6oGi06lRwMDErOFFWtdAVlG6zTWi81UhI0euV4iGck3JYiJ+EkP2fFbpAv2q4Y8ECrZ3hZVrQmqCAG0/jATBNDaVDttSKLX/tE8w+pSX1WchE4BEA+mBggQJKb1R4el6m/x7myn+5twYMNELawtjl0btRv9n7A6D6s0kOFL/9myPu39HzqNeLHoioJgcAS41oS3zKrnExAooJN3INWbPhBIdJUXbiRIcxZyUEWnfzAGevCwVJPCmPzEcbJ7WKTpi5OvplJ4J2WCJCJz4xCXtnQaO0gKu4RQxwtaJRXOh0cF3QVZR1iA9Y/gKL1zm5dWwBSf5NNfeNZKJnaJHARoXidp3GKyxLRPXoxdJXAqYzOOuWZfk11gqD/IlEdvXDFdoochkzNsQkQEGmiTFaTNhN+TbLOeSEPsN91QN8H7CFfevGZGAdctEr+kJkm+9/y/Y2gp3ElMlFl7PEamZ1dZUjuJhdU4tvxWl7vESFsfIvWStNKQQA8EMJXS/F8DD0u2COZZ6b6HPmYMSptRnNN8dYArcDCLzcmc2ltQ2133ZPrshg0GzoB9t/2WlscTOx3anqVEF4T6yUWkbCy5oQBFUlajx8pfEC9I6c8I+28ffGkeppKTa49TAFHtdYpBuloH8jBtx2CTESUgaD/QAJZsLKrmesSckHSZiV6K1POtE6Ov0XEoRS67EJUAzxRw02nvNaxxVXjCJR9sDtd2LsUbW7AW4jpo4uf+SXk5hqcxt6K8++vATzcmuhMMiWGfaz/dG8PHH6yJNnqzLF3VTxsRoPs+MokcQ6xR9LR3pmuI8uQgMwargh4pN72+9GB4YeHdaoFEvIhJWhx52ZkLVeHyk92Ivb9SftQJL4NA1+jOsrWfGKD03YGmHz08RMvFM6q7scpDmwq5OpMZ9v+BQACHfkKvnBfxoLYNIF6m8sqwdRNWstsOsMKY9orYDbV2aoIZGkyhH6rWBkkK1lzTWj7Y//dsF55c7W+Zg2P1ltb/6NUOWeYrpcpghnNObf5T9XP9+KQT4RFSlhI08EOmn/b+7u7X2Q1oM+bKca169KzhlZCsEpb/G41tpFqo7BispiYxY6gOfnXOG7l/6kFDe9ZtwU9IIdeIqfDtXHLiMtm43B1NmpLljVS9CtaQfgLICBDnoL+GXgZm3GaKpmo8q/aHL+pf9bs4+2SVODgrbYDBNUnBSYIrRm8E/5/zLOPd3k9THQVFE3fQambGuQRCUhXHO1ZNvta7vhZlx8UPXYz11OeRg4yU7UESkJvEXfpQBsO+YNkKjzCSeBlBZygpffZjR1IkTwyMj5K4jJy6tZIKDzD/qsYTU6qsRZblx6dywb415aiP4m+B7peGRGz4wzTR9IA1y1hQgSjTNxys/Qzj3SY58cL3BTOGK4oF5A+fqnwA7MF5M3TsVjPTMFd2rU4XlVsp8lskVqNCfaYWQ01G+3ElDcz1K3qWujeKB86ZwQy0xrojOZtkUV+1zQBVAu3/aFJqjYfLsGFXK2VnAZzb3b3o26Dw4QuhhLbfownzoTx+kT5fJ1VvCD9xUvQhcmDCSxxDlh6hrOpMm3sJWxk9jHXDC5keEKN91q++psSa6uJJbeaXtESX+7cPU20rxWz3Z/lLiBBES2Mb0LAUOTRKYKzfqTWL8JuXW4FHo1+pl0M2/fvw7NCdPXE6vFmuR3HGh4LZ7hAuhzBu92AEhp2JR4rFCIn6lgsV9fNs1FqBYPUNZSce0R5U5+WgojXjgDXqkK3XBnYWOOa/ZScY0BlgnB8mmwi4n/Lirx2XrsL9qNmZ0JZNbQdHzckg3tJY0Vk6RMBPZ9Lh9hxhYuey4bZd+ozYMe+hraZcleNZJZTEBewmYXoZjelu0GME/DT6DwVky5BLsTpi90jTGURJXso74kVlDhcfbWdMLlbqlGKg40zp4/VORG78L9K40mxHNYXsmaKQmIhdTRyRdYjmqR7NNVA6FGmTCi0UUqn+I68hmUZfedwJIPaUMx4mizULYfH9iannmBFOnp036NyJqbj+5dOYkim9kMLtTJazd1CS5+gDKLzsMG6Buf4u2aO808XqM4PgtKXGLWM2AzvwKGUmrNalkIPKhAX6gpRLqVQUlDGv4W+1ioqu83aEpX5FVRaMIzQz7T2DqobZmV0u1iZA/q6Lr5+QtJVRkNtiKdik6WnoiQdE6TttLPjFBJ8tDXER2Mm0i7Pcq18bhbSE5kKnes5RqFipjKJqT6xiZVQkeFYPff7EZ9Gf2E4QPg8RqcCsFcP2XkV7wkvByGm6HSciim2a6COpwF7hGKbFYhZeqgVmJxljHr86yOGrwv3OfV6UuuQHruu85Z1oWm10XDS3/u7fEu4owFaeHH6MXc1EURVWzIlYvr+zP2rNLrJ6RbIj7Uq8nlWfya/fzoNksL8IluiPzMMMTqFrFW+3xjhqt2ROZEKwDhnTdOAhu2xR3JRzbY8jv2DNb7UrSYO3VxNr0zYM5DY2DUjNr1CojaOkGiBxEvTtiu6TC7VuoI+j/2iGsNFjjpw8hftvVkh2bzvZhr0yRuxSp1AYsXHQwt+UXXewChA5bMxmSGxiC35oyUSLZOUVi1uTZuZE+cB6CdtztmjyampJ0jYMVnM8toos6jZp26+bNi5rZH5vhCFSXiIOAmhab3GILd9SgIxHe0j9W0liMpuPkxqBA5IDLGDjHa3WguoRRdO+eUyVzVjnZgxjRX6CVu5lp9+U4i6EKG+NPkMqNPI9NE5tdCRlEbsxRB+i3SOIbOeKMHCLHVk/fBj5iYZkADpHYw2LFTycilpr9LJvIWITKFGAYmALEsNFb5RJ0te3bXwD9zW51Obbrl6oNKeOQMt4XzkrMhKRoPQLwUr+bkOXLaFLCeqFQ0afGrkdXkiuD4dsAGiT552cnyfQghO2MyeE25cfrozPMeYvXZXMb9jHk0RYfK5HtYnnITNRKeqbGSklGeUAQ+Wy0tkd/2GOnmab+fbzcGCCr6g2s09G72mKDorTc9l9+TLNvFcq45pKq3lVd8t4zDM7BwS8wuVgdvjyaKqZ0E+fvjVR/WY9E/XPcXVCyTklsevXXlO0vv4q/5gXK/hEQCh93BFZ0MPiZoDW+OJ+27CbnkYUOTB2tlfoq79W0cHRBFVViC7BIsOTasHoGeWDSlF2WYqSwc4CVga7kELczAGW2OtHVn75sKsEvbyJLchEPrkO0Hg5o1pfxIbkVsKlkDS/lo2tp2WZWn6BzjT9vE/LpgHbgmFcc1C723H2Gb/UOh8v0sHQxSeo24I1YE+RvwMHnBanNPx+wo07cBLFZeyYj6w47eruPu9z0xNDPVa9YnNT2IRRIPkOGEv9IefwdLhI+2LLP6O1Sr0lfl4WHPMR6JNXV45hfc6Prn9a960pyln7lTXQP81IJLpp4MVg0D64FvkIrR+xdDA+85D7ZvsllrzMCeuoL3VBFrLJ/Bcg2DbpUrRuDz2EJOgsQa49vs8+8tQ2pFyf42EB9vb+dm/2yGw+pEMzkxxO/JA/56T8eCcxUkdRBvWHcPA3R7+Zp0s/3jDdJ5ykW8apwCJVoV0RQyGipmeaJkzqselwrPkXJmyxGvU3lSekKtIXWYrUokzH9WiOBc7gqFV6v7wCh5a8zjOnl2A74PjgIpFYgCoGhDstYsrFZ2MrXunqflgjfIbm74JAfVfNkZEmn5AcezxLkbSqdc6Zc69nZ7ObV/I5SvSgKgkuiqpaOaXE9mVeVBSMxR+mqd+eGcEcFNW2DfkpbkMBOpZ2yTYesrZez4EyLBT0L4JJ00XTM51dH0OhvdD4e6fgpSc4p1HOicT4ADC1U8Jnp7dG6+Xz1VjHQqO5dsndpuLVpuORZ2HrdW0EJRfM2/6UI7EwDtsLD1pvs/i2z7+6WYNJQdLx5SpfNm/HXuSyML/mKeK0YPZdsfd3m7/hKF3MkDkb/piQjkm65Q5u2EAmtmv2PmmOBvYDtXBMWZgWS4uC2uV4+ZHKeFyXhQcCmo9aQKVvSvYKnMXmzOtPRWc+iXORFQAuSfz/jj0IAjvFYpnDOtp6znuV33L6aDYfSQ4ddLoC6nrrCwP7ns59kC2bRefg1Y7miqqSdlyEr3/Cl7Tzwk2uBIqpFez4I3cvrCccsxMBmHJUlXCYupSdsfytGkB3AlQWmB+7xyk/qIF8FaX5KSEEabz5qvxnMTq9/6omVFtVrXS0S5NYtnsjOp+WHoEBn8PWf5Yh52KbKPjWBDRusCJVVk+tdxbxPxsaWEIm+LzLUIDVDOZjaBHM1PbUnwlokxzQGpztHDyJqvLa35+G9qVrMDXvr1H4sz3cV2rrMRC59fPMf7bcJUWjgppLBrqwThZQTV/i/PfATaOMwrHmNOMUS8b8ZYQBt8PGFjzszb1aQ6nOn+ehu/jV+C+e1VOP11UNEqKJF0LRjL9c7QKIPEKphuZ5ayT2Y6BnBeOy80cKdkbzQCwzrc+dszPa+RR5G4TlP2usEc0rXYAjP0Q5mpOvR5NUmivmKdrxX01nDoQMejwtgh5tZvgGPLgfhYQuglC8gUe2WR5CsS2kPv0FHnQOUwLwCKVzYXe8l44yPOySbGa5fveFrMFIwH5ZID3byvESI9GaRn9rwDiL09XiWaYOX4VccB4aT2xgW1BFaBGcHQRxUzVWfauBbS9wWmJYM3bWIuTao2GUNl6dzwM73uPJpeLf8bHeS70pGVh1uEYJdvfjsE77U2fczxj3EtA0xECK2bD+/xecAJ7uXfSz6TOLDqrEZhi9NHHkIQ8psEcEY79FugyLpbotdht1VSW6lXji7D7T03pNcKWKGDje9d8X5t4Paf08bKbcVTO1/71rDMBzUNz5gVIkfs+gOw+k7145YUcbgWrBSHVgl9uXKrRxHzZh7CXJpYj9/SJIDaJNoTdQde3uoAKu2Ifdqss7oROtPvaCoUWVEvOV0aSy309F25CWItom9qM608dMMP2ufVxeYcCiw8t3mlVthm8m5zCq41Wrxul86yE7uRnDPUoNEJfb+Zunob0cylQH4hP90vzoghrgUrt+8/0owkpBFnKDEEAesyzPOdzSVCZX27dMBTgXrxrZ+b26WK+WelLRyBE2H4lv2xd9vH1aZQuOnqWZAsL1SshXKn6rYLJyto7tUWw6eUyKzthjnOjbz5K9PtGTi2GSZJmaO06Y4JrUI8vkkjdSc9jofZw4jUcEQPagMst942ktPg6XjkG82gZCeH+eIEVSKab2D4qv9EtcJ8YXzVaGvJiHkhQT9lUUD7P1VtdqMBUwjmnk0Fh/dic7D5TR/ioIua6OUp7dteQUL/RoPS5h0nIkJwLi8xwTHghADBAoS6KTW1daqE162V6mhH4ceMT0o/8E7FHtEjjpeKXofImstHFcBqGhmjM600mFCLc3dBW740BhodDIQDkXNbg2KhoABv7ZbcRHPFlEp6OMFqNIQ+ZINdAX1Q/SvXozS50J6P8fo/E04NUckWoXybWeR14PLq0oeOZu9iKIPN6oGodyqfdYAt737MHnQPHbheCx4KHl1NtgWnvnNY20VYv81uYgGXamwJqtNStCtOZWJCfCVk0Z5xNaX69vu46JLLwyUQD72k8ijwkczXLixNsVUNeTnX8hSQkLJU5O/81o/xHIAbOhmzfqr97Why3yxNG0bP8JRYo2c+AL+v1o+2gAqaT/1WCZ9Ltj5yDfJb5+XwRXRMZlLvKLq+J/ajGrf/g6gAChqnFsJR9XuBvZWCd0TLflAjpvqtSYNw8fEUr1GGe87uYcDlIE1Zfk2GkbpW5Q80YMdyf4eBbhKW5Cr41J1gqzvJz0ZGvdb8L5P8T4+jmi9SZNIUYsqKfOsDhxABfMF3auzG1Cett/TDhPm43XEp7OeY84Nv/GF1JGlsukTr5MHynH0LPoYxygi26GE7xt+2MoeacOlFZtwQcARol6LVaHckZh9+b/Fp7dMQYyjE6ZSZpayNcEE+YLtZRv2uPgylP9BgeIwT/DSJbiv4ELMLXruY4Hlm262TUljvJVH4M5G3B58NpWTY/Qj57kKG4zuBkpj7ENj8rTFmk2aQeO7dJzHWsZjV2ykhklHwKGcs/4G9aHstrzSU0hDKmGK7Vdeh9I1MoiFFb8t2wiu7k2BJOmLznW/pjPICpoo5E+J3pn1YBKWhQ1eLyqOgO8V03qfxHPpPa40ncdKnMqMTCSP6dgcrRLtSC+HPz8eTLqIe9izpI6McTi90fp0sEtRB6eqcYiX/PidABMRlIBwmv3sk+MpZNpWqcW7tUEgWzT9K4Z+DN0y7pXrpNOtuNg0xVakdA9QaG46SmJ+Mxwy81HOL6Qa2ve0tJAloC1pNJCV/kGgivf+5SguiEytsdgv3JvE9jd7RBHY6PAGvpbLbl58fm9E4RhRBOdZ/RviEfXUvRsPWFgVcyextSoiRllMaOFpaLjzVTrdM5qvxRoydz5GQM9nh7znYDECY6sxyrEE/pWxsuaZJP9YgsSt5LlKPuHoC7HXAZB6vRmcypNzWP1SgC4c16LlQeiUUjSIlWFSC6jzcG+BvA6QOPx0A0k+lU81X4TNDU8HMKTJT7LcHGwfgSXcoFPNv/XoL3veOjBBfZxQvjI+lEd00b8hWHLQtrMxqH/GHVp90te1O2W6eSwZLABYqapAkOrZYJUjT37xURAOuXM2d9xBcfjPlKkSdWN57vD0ZZhONje9dYBU6QwKcx64WiOiRFyyk+z/hmQ9elsIFDmgsGBKxjBxLnCB0fBhw57U/x1RbDfDP2GGOAN/LprmemeANF3OwCjFeaCB29DPYCUOS4TiUY+3fM1LZlwLHM4MWRF7vkm8whfgxjkJtZYYfNxTcQztwvE3L4fmUwOCDFS3lxjLqeBG5cLNaV2LHIeAZK0LJzC3tuYzF+pQ/OqPKq7F8Xnvm5nGFLf7NReFOU3JtlgHkXUYtoiXI5CTwfMgRZsD5OVR8v2SI2/QMAiqSnB2sNHqQyM/43kZXjnbU22lOC/+F4szwfVhoBVVSdP4B4VW85tbNwxCPB24XbUYxF5Y1s5VvOaWKClv88kabnm2AFVmc//ggNKI46vviCYOi9vxLKfHRvMj9gf+jbw17W8FKJWDmoaQAcDVqauY+WXFbSBTCMQGJzdmWRBCaLdzPKzWuc2tJclrop/8TbqfR3xR88cWCrs+RGaapDerFnniWqEN8IKxOHxhXplndHD5MNJX+zCSRPPrrcPcbk/Z8NNG6qyl0MKIaNAw1keGMHVbno79o0SyUS4jFIg04o9jFJkmo0AN8QP8xLUqM6UHiMCoAKiIZBaX8Pn3i2r4Zp82hnG0oaMqjjni/ha1L7JX2vRTW1FfqqUiry2R/dwBfVaKB6ou9II2HlVK3QLyG7PBLNLHbdRdF+dKBnxzUfhLf2Ui7PP5bWIyCtp31PfCrrVWThpad2Sh67t2eaPP69dmlJpDmlJ0uBWmO24YMQi1yrxA1bSTR8vOZC3yrQVmJZHdIcn8BAiYlBxoCVP8vSmF4zR+DizA6aheOUxw8kcQCxkq7GVEn8Oci4uMEkFfxdmGWSWLhU6OWXBK3pjV7o1KKoUcCqxPJYZWzQn5vk5Z4vDNPsgDIA4z5fWZZwRelsz27j+pW26GhO2xnlkgswagMBSuCNjl37HW0DHOD+6JVpmUmdiNRg2EvPenrS/aglpMlhJfOwjT8V4z50UegSzyjWPLLdPb7ee+WM4NrvPlOVY3fk1iMMWW5J0FFFPr0DA3/XUI4kHkSE=
`pragma protect end_data_block
`pragma protect digest_block
23dafb0840e65c0ab543349e04cd796c7dbe28cf520f1bda8b9459a782594e33
`pragma protect end_digest_block
`pragma protect end_protected
