`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
XqWL7FYb2bdGUfHkgjRCjRF/1OMeSBwSfKs4Mck6h+O/uPyM7i8pJhy9l8uqA/STvdSYNeWOYTnOxBUUBW7Ve8Es8qr5t7DAILv/b6pZ9Fapfw06e2TFDULJ458lAM4vnQIz+BImjo3ss3sXYp+7dBiJI0F3S1ua/ulBschwfz3BtXBrmddb5HwsnNfybs6RIkhImgnvgrqmRqcheSImQo/EmqwFPkveywitOjkai0gfTn/htpajCn97tX6qsLUgUjyfd9a2z9MIQKmEQIzIY50km1VcWMOkh93VWwb/LJxNhzuikpLleBdHN5OjcO/GmHIwvmmdos0fiOBoztIG3IAmiic0+hkVISkGEBP3uchx7njdVyiM6qKnc//NkWV84pV5uD/eOfcMgG4CjLmDb/mgCDRachnS/zDLQhRK8Ikx4pEQHYls0gJA5ss+qs3i8ckbDvrMwOUlueinawEkPscWVbbVKMo902dk0h8kfMLMUUsXl9ftXcv1xNnxeApo9jt8JxZOVR+pDs3MnGPzzgniypuFQlQh8z1mAkzT1/gsI6sHuo64e/sfnysv/tJ7Dla8x3taLMyfGEvJPOxrqzZOoHViW5M4DF3yEGNfOHqcLEFH7wFPZfN8n0fjknI0KwTqJdPVKHdvn+yExxNGkDvd3sp6kGi2bHt8SFMrli+9eKxe8fDybupYSBV6c9XYgi0jgjTSHq9V1ievg0syA30gQycz1TYHh2+NKkKzHZZexuk4hLS7YOEQe1hTGbdww+d2fbktOSHGVIl9cTYip83cDg6G4VF39JXRhTEcYCmaufawNf+wLrOj6GYkTOgOEot7O1Gvsyy8PlMSN3SRXik8RZt/5CNC93rVVGWGYpsFAm52URl7anMLu+KQQ1rYfqvioHwznUQNjeyoRzE/M/Ou837pp2NNjxsaNvop3UI8MzHkSNBekEcx4IHymW/vL1SJXS+4a+VvFKRO+KmENk053dOn8LhIxGhO75HI1l0LD6Bve8AhQcmJ8g9Bt+IaiMQpuOdalDNuufYrbnpS3nOyANZ0fdghRdtc1ezgttWRkLb+cJRMIPrvf926V/9brjPVH+nLX414pGT5v9ZTb3u3A4PeG4um252b/8QGuoaZI1jA10uTiEzplTpEnNZGKrgfZ0+OR2TYYGR/WBzQJ5JWr6uNwqnA1BtxJAXw8mSIONu+YsTDwBAWXqUWwl4n0ix+43XGZAiz5aeuA3HJ1Cz3+xtZP6P689syRm4vcxl2y4Erdl4GTi9TElMhpEk9PLrjKZ6F4dwrqCPiB2mZ5TZnaCrx5cMqH40cCAx1f1h/Qa5/nd3etcDpF4QAEx5rBz/o0u4YbZGsXA6imtslXQxLNxBdWpoSzzHjdUuxuTRSJljyID4QdlepGAR5bdUx4Zw/Qi3fWy84Ws8yvZIZ7niOD5mCH++RMwuRYJlSBmNsLUMLKuA3+N7DEoowebLyjE5gL26oMNznQ04o+QzuP2JXLXL5pZg3RB3Nw81DNk6E14ZQheMKl2tTO+PZalZk4PpYGRc+b2IxFWjdQmFqTs29lqQb27ZBwG5qKaeKRGpHcdaWy+ZbyaOGWzx9dXrbZWfcTQmatTxBltcJuxsLbLuS76KMU32wtDH9ntI6dM5RHFAWCidDqp+qlgEoJ/6a4qLFErgizc9GTdP2FrSv2/Eih/Vy8mW07VvOrA5t6y9IvYAiXalcjhGj91NuJ9eV4cYsBjcuGzwE5rnhYlQdACvge5QXDFeuWwd7xSFxpTWq1Sp4qlZAB6AfPmNJkzcWTBvDSz9Me21rxes97MoVc5GgHWqtJWTMo2X8l5Wd3iFlXXSAHFzonJLnyvJcm5rxcD3EHPydVp+xd6RyQ0drujOwjegXchdCoBOVZGKNuKpFVW7zB9+FuImjfNia0JxV04DMpW7QA02TAy7ktQj3dXQkCNe+BDPWMSfkrWUcVus4wFWrTdEu5/8Lmlw03/6X43EjzZgb/4EE75BOs9vaGU1GVdm4FrQdNvZzLxYQ0p1sPDomuS8rsRvrhPejsu3QeDrlmQwMQVxi1sgx36bq9l9fC3o9vGAdn5rp4lsipT/ic+MHV3MFqNLZ1C05GFG9D888S49T6YHYHMG7GGHTeirepF/O1lLAh7WS5YCwOWRyHkn7zN5OzHA6gD4b6L6Iw8NNe0F8DPYrcevRtrdItmu0pQMil243XKXalmBBd78VI5C+2cekaTPfetwNV/FDPyZ6w7dyywnbnSaID0dZNL7lmtb7KdsKlAjbtxcypvonbKjsSZEx+kvOS2ImICCVHARXH2YIzBQuCoYFXzBaKHPv+GFcwpoGpUe0O9p2fv2pXaqou/SLTl7CSiqzAwDrXy1WOuzuiejGQDOMljelqbaIKtZSv25zELljM/pHhxxjLvv3yTlK85mdPS4DeFZvN1i9TIkkByvR3NX1AUZyw/ahgR+SKnDwA+4JE/Cx2slYuzs3KBMIK1iJeMwUSePGN8RPNJ5s8UNrCa9CEMQQTI/MTATbqfcJWx3/2M0pRRxPCdRQvXaREPdpPy1/3jwIjWHh+R3SnTnR9+5PlxdG8A7Hg4gOwOlzINAVo+JXha/vxRYucsaBtPBCYEtf4/xpLdwMOO36eP4rspVJE6vf6mJLbfdC2zE9qws8LgNpUHemY8IpPnuUU6ue/lIJQBlf5E7E2lZ75w6u2iiG+StXerOXhp/D5h5vLkYEYehtm6Et5qqdwZ266CqH7FFAS/eV9CToqZoMxvvFpdMGSfTgB1dfkTcB7KDq/VK2qsWxLJgHMYTiKkjgVNcmpvwL+0Vi4Bo5kkd0a1aOlPFJ1xjMiHqCMIhHA65Fk3AhaT1VadS/c4bVbj5WMlya7yPTT27KHThq5mhOE/5WtXqjnszMglkQmQbqVrDLVjcwjBCsct9/E/M5DyQ/YsxSKTxj/cBdpUa5RyrNGftWS4v6iPlUlT3PfSPW1xHKPHjikN0kbdd8LkYjf5duKCr8Tp4YDcwOP1tCO1RkDRu8HBiPVZq1gDO63fmZtLefyy0fO9+y1+ag6pWHk/iznxTYgpey5mSRJ76G6U6LCvjOzl2dNP7HAlbGukoPjv/dGa48tdYncUAJGazDBDZpkDDSFlM+50A1M416/n8VmOFLjVAVjcopg2RSX07TqrMu597eGOINi39A8V2B2Klvg9vBAJGbK/SFgx7oWlP1LqsD1Q994kI0D4xKtgb7bNW6E6P4oTeCtIUuRLr3P0cHDlVrzjiCVV3pslAuQf84D5Wc5BI6paBHtc6rh1XMm+Er+A6qjDz9B3bQckpypFg+j+pQolRj62t3lu9d4Wcbdy6PrQME4InFWNPbGaFWEAIykhkfsMxr8bDg3jvl7k2P8owzrO7Vdbd5u9KXsbyJkZOSJ4bQJ9hYhGnq82vGabOwDgXJ9KO+y8J/HhsM576uNFy2TbjNSs+PaRHrlTmXPvBZwHbnP751M1wUeJlKogF/eJLJvv6scXjPuKoQM0JsSmQnRXt2XOs0mc7Q2GC0i+qh1JubcTh4bTHDPxm/OsxlJHPaP31plzbblLWdDxOnCArS9U2OUc5+NAqJ6DltsNIMug2VEq0h+LRdtBAty22Anow2+ylj2hATtLfGfL7952hnf0KuDWJWfznexn3HBWILsL8lgf7fQURSNW7mgyWb47wkB0Bla503chzuItGGoSRNER/Ytm0cuiNZsmoU2MBwhslRQ4AXYk7OZOBAjWjcwz1I2Gy+W/YGwsiL1uPNV0l4CWTef67OVDy8zaPDbYuQYTtxDA6B9M0oEtx6JRdKwGdR10lmmnAkSY0fSo6FuHKgRqXB0YxG/RbeQTc4ldh711AgAcUvnZ0ea9FvJZQnrVeD1h4/bgADdX1ulGTRkJyAJKPDmx+PiCcrBliqXu27S+iDfHvsqbN+RErJT7XESqa0U/TK8UvkoI0Br22S8+/3rieYFk3EfkSeG0yhpBAK5Q4msvrKp5BRrzF1Lc4GOcSRPxGEsRGmyB5U8Ac/NmNCVObv2f62890VhZ/xC+w3ESUeDsxmC87js/L8Gh/kpWBblOMFRrmmms9UPxW1Z2znKqy8fnwgJJoMzdrZLHzbKSqRUQkdBv8E2BQbf/AvMMA8+fZop3TJ2YVppGYucCXvCawNK3l5ssd9lzCw6QM1XsLBXD5GVRxaMWVqggrx03PCx3NxG6MrQ15QjQg3Bl2hQQBzgQwLlSVw0Sx8fNLCAE3odw3tPYHQeooruv9JaEaKN860lm/lLhn7bO26Kbf7cUdkuTtxdvZ8KWm2aXD3J/T+iLoD0881XPlLLNPZP4lmO/n/Am63Y/AVk6AiaXcbCdORa3IfXSAkw0x+Hp/OYnwSI3+BuT9rDKyy6m2ZIeMs4nFwXr4S9KRQTLYWMymBp6U1QWtrM1MLrCA43jLAOCok22ksDZpFsIRI4eWkPrN2Ir7G8JiDeLs3zZHz+R6QENWYf3OvMCVj1EVGWR+TECQ4eL6+vEsU5g53TPTMsOURQ7Jzxfvi9oPKq9QrJzI4FI37NZo+tAPxnu3ZGPhh5u0Ug470DfWOVVrWrA6T3X19lGn2YB7IKrwZAvDmsKYwH/np5NNS9sTMRnJdeQDnqrHDYNL2HihT4Rq5fdyxkKbFe1IJKH7gPdHn+3ikvY+Gz4j5CI0r4wejhEmAyeevxymkMDoOZXrvHjoekHfMgCkBCnL0UWor5DCeWULvOygheX/itFGnTkJKnC3tfP6SYe6ofkafheK9P3vmtVjChaUgm9m2IQu+zsZRKNWAFONZ5DGZxt3PWLf4bJ2GD1kEAzEpWoKN7WVSeoTonYpgyHWB85UfXdIgegLXGpHlZZXW1ODfmssoOsFWVvQqpmIYqBveGbubzlJzPkxtDSn3FLecrh5Id1Z3BQsfDNJaPEz7wGMDGPTH+peXzFudpcAWojVSyvimYChTsnMrT463vwotTQT9BXL9Uya2RIjUvRyIIFUTY2hmCu7PGcRNStz01MX7ZS0rzWtO7FCrPYXX3SNgqOI2h3ubCbylLLiTSweIbxpPRNml0xy/Tx1EArwQ8yPFPFz2UQQAxm8SkaV6alWghdEe23KInfYmV7oR6wrqOr9ns+ISQHZI5G/XXmoQP8r6hLngdDmkFkkAzyMRY2zXdYrtzNOCkSFIYy1Lm2xAQkoIJ3OZj6Q9wc3q17IeGGn0zME12sOjdcyAcm4eL3TFjIlgMHXav/TBIYWLa1+u4LriM/bC5JzQfjuyl2BFkfXFnrfnEyq08mR1QY3lDK+AaG9B1+DfHUVL7VqhpJivl1iwqnjm6sak+Sg89VMVw+LqXjGQVd7b5x79P/Su2pNde3VDTmEI90ge5pydMfLxza9npn0OuVjGeBGf+Fk0ny6z1fSxuGqiUk1AByXgvFJAzy8j5PCzsRcSW+FKeq1e5pIGYNfYdkhW0VR1z1wE+TFi1aLpNVgjhokI1W9KJGUY3pXkJtn0t3BcHiSyh476kp1mM3gCou4LqxuLCqf6E2jp/g8I8NskpvxpffoX9BkIAS2lCipKZQI0Q0oN7znv3ENK8Okho2MSpeHLnAiLJMP9xCXA7tn4oEELqgaixKYBLCiS6DFJXOaktEzBEJRQuaIuDteMuOzQZbFoJ22yW8FrZcgZo+5DyEh662hOtktO1jf1k7Siqo1noP1aXkbAkZIpyPGxe8y7rhfF7q9pJuwNUJYjdI+r50bmTWctTHRH2NqVikLNJwzXopD2WhAxedzGxMfDbasswhsN5nzzAOxVRbNnaJZ1E4rHH0w6r6zW+/1oUR8+/U65yH3bJidHdQO5qYhGE8J+Npu35x6hypTeXbTZD1m8497B7iJHGipRWEVdEjQ5hZrLLikHaBUE0TDixe3DwKJPxU0wDpNo/FOsPTyzXhy1W5+TW3IU0Fy6D2aTMnfJ+wO/pOLLMleS3wqBdp5ZRKIjBO/xGjtTiEoXr97BOM5vC6ekXE3rudgqwehPRq+EwGKdXI7yVI4vCE/GQbwaH3gntnKYDK2vLSkpwttA5Zd0LXPB5+3OrXSetAhwvoHctiTSeBWZnr7+xD3mmUd3WhXMN9WuPH00DnjVUrave2WHKiApVBgsU6c52PtD2ro6OZuP+unD2aqq3Vap9irW4QMthDtXiqxNYJgn0DZilXZUB3mtvcC0kNA/MLZErK0V+fkFJGdxzcM4DZ7gK1+s1BPvSBVnn1m9ZBx8godN8Ixo5d4Cyxan2UVgMSmZWcHnAQL4J2Vxjg4NVcKj7vx8qyPn9AjFZNT8tqr1cm3QoYAYKmG/OBQqQTMTxMYeYPoRGAafoVsEcpmrvvmj1QSV+nY2z+tm6c0LjrvRRwjxM8SQLCQN8SwgU4pQx6XQ51MolnmHDS6otMjvbG/ZzuYTHUY+9KVOE8E8yD/rEKNrjWcj7sdf8UXJNg2NsDy5Kq9Gx5W5iFhPz7SqotmZiEp5vPY1fIYtx2PrmlGYRCf9A3p9fgH3K6Ix96uUf977VmQpYGVVpLAzP0b+0OgONJAwvqTu34EiN03UvMUCtwzcv7WgGmxWJ/7wHyxhM6yyNZnWhclFhsq/aY1Tp6OgK6zL7JjBckIuHRFs7E88bkN8LimtA2AoDvUKiIs5NvaGorlMTqtUpv90Ws7WoTiuupnXeSoTAiFWd8r261rthbZQw+6iUsCwt1dR1zR5M5yax90SsIlFJEiwfGrQUm7gk8p9/3QlGff9EUg/jFLqJkZWWFj1UubywOWJMw51zfBUpL+KyMQ7xxSGU8GW1ghET7rq98rZutfr31qvSY9QU8k7Rwkh77+/85W7qwX+BaRCtn3LOJF/eWLWsEVPYUE0AHa3t1YszuMFguOlO5l8tolU/LrY/5r5znwMQbJNSCF2C9+R+haXbfDKsHuOxjbF7DA6EVm/GIyi2DMqo3Y6LX0nxlOL54dIVsko8a6y5gIfe21zElnEnRkiw9wgWvq+GzSAFkfryffq2T/A4baa0Wfdu4iIZ8q/SR2ktOKivcWWa3kMEm31sT5s2Ss2woeGnsc0rFajc2TO2jfT/ay9v6McpyCTGagBCt22tG5Ir33MQ8Hp5mZtQ59KGTRIEp2KOdsuzKP54tb1e615shVycFKLQnO95bnZuGewgrkUeCLGigzk+AvZOY5GTcpJaujXdJ8mEYzDrPgDz7hlvZxqMk34blPwEFFz2tylAYAJn5w30UxDSxtiwZKm48Z/k7eLkfsi7A+XcTI/4Ccvmxr69Ixfua3igXkhztDFysSuIrQ8Rl1xnqFoHVhTvy5cXeYPiUpQII6itxVRpQ2/9URYwPSgTWn18GtQghBe5v9IELWpwrmkLiM8cfg/Hw/67vhN1aoxg/Yg8Mx4HiOSKZU2Pnkr0adUcrO6UEuP6VqoEVJI/5gFWZ/ERQ8DHYF1e3cCZttuowKw1cLwt23PzmBxSyToDjBs9CbwbZWX7+N0AnTT4pwuo90TXuhzSHLzrxUdGi4xFPPszmZ+r3rQyCnh1Kk5zO70ftaqqYRnvMZVpFZZQkZw5hUgnAmrhxMsyuLu8XHnvTRLbYLoFPsKF1BlqjA+9sFMAiWBvIRDsMp2pSiaxAf+qSAf6JnUFBk+tX1ANgi8KU5YnrcDovVcJ7UJB2BziocX6E10SDLoY6jW4M1k28DmWrHCIC1wz89RbSsNaWuVFezeK6jX54wHxjlZ9JESaKA/daaOIfImfIPgFl8LWDMrMNkV+0Txtk0QoOx0jxs8cSy0F+fS4YzqIvtW2ZoREhBPIK4iCKoFfjfW9JgHWWLVABTUEUZNkw6r+EBRlRfr3KeF9iHWad9Ay/fUQbiss5rET2Ny2C9mUwpJsSFpzCpkfwcOxIqG1sIwZcSCT0r35974JWuP5TgejG7WoNVBFe+YJWdFO3rtE5dsnXmSMBz95HncChR48PeQkaDJLoKrH0u1EfXuLfH8yHtap9gKg3F6N89zuPaVGIJTI5+zjF11/+vaM3TdF80oUXxJjNSDC0cmqc/+TZiZ/wE4Kov8AJa2xCyoYZzgrZYhalR6f/AAq9lJtCz8yvhrgPwBLhTysPtSgEtQdmkiW0T4DEGk9KmcAekVX+s9eFv6edDDW3Pm4GqmVSDw9xaAhxK+G0sjvg/+0Fuj3ZKk9nBHBC2W8YlJmsJ1yQWhXiEp13eFcqdehke38YIXz+NHAt68DS3paB45rrCvA906zBWzTZnw60wPk2fiBelQrrgZeo/JvH+WJSiWXAEp2xVVU9sS00vKWv9o/9MbPKEiUPlf07ZH7sjHywvb0mRIN4cbMWwMff58elF3Ch6Eih4GMYPdpOZnx6qIYCwAPwdlGXFznFKaLYpNi75D0nsi0AjqWKaNnxmtmN1JzOwX7Klm5mzyll4KlHLRPDUekfgPsdo8KB+nSSiShrOf4CpPYiso59anBXXoUrWUwxGUmh1u9y0mx9O2x/8msm2oCAmpa5utdsfgYxNvV5VaXqVFL3bq3zV2hINu9nvUU/QzwtDISVCrFeRsuXZoX1qRBkdp9nulrJ+UUdqOevsUTwMC0mJlK+3hDsOdJMwrJ2D0JgoGuz3rq/kNjKCs7UXRJjoKS/8H6+0gFBUt5swfmAgDAAsifY8fUxuS8UsuJXMvAMl1EaBN1DEJk9yZ45gpBijdwZlS8mHj67qECuXR39wPWF4I4mU3vqg1bliZcpWR3iDIU+wR4w0J9O3ffjGu/HH4QZzF95dIzC7Z9sbKSKIyr7NvEMgAg/9xaKlH7jDSawypdd+nX+iwL5jT0yGnF5CyedaSAAhjrPPXOI+0k4n6Hdkh9+ns7bGXYmPXR371SJe8s6qv11DVG9N+c1ZJqEZNUeGRllGvdFWfxsX79iY2ay+y74llFXlYHl7XImk9o6om0NI6ccfUZjA5PPRr0G1BMB5+f/DTgwHsx7endVImnc/WdMUCe7UriYH7PRe2o9JzT+LfMY96UsBNQ9HzIHMEkTrjIHujywVPWKl4U0YseRysXtnAl8CVjAjlzVLRMa0fclLC2BzPYwRVloGnyYY1TRpO00VGx+dY8dA54PfOBesAXXfe1RaAM8LOpa6w22lkgeUpPtKqmxvh+pP5a5EOzYopdqz89tFDNZb9qnfFxqvmdKrvTd66Zaqz152oTpVopNB7U7O+z/LlQzpdauQICZ00vj9D40lSn3yCPp3lfVE+TqnMRoiJE9N5B43EHwW1rBcYJZidgUSh7kwlfbhsqt76TpcYGGT0lLJW+4GZ4OWTV2YZbh37zPQGhxEq+hojY60UzGqUZ4SPuzS0iRHsHgoexloSladHOGiPYCC4i6JsURCRo5HEwZyeG5PDqzOh9AaBQ2YgDvH6MCB0PZhHbkbNKQWJaOIgByDrK2nmzXsv0Dwvg4dTwPNH6HvbP+ZS8eip3GcJ0cJhYQYU1rVwEIr4TiuZgSStp9G65VVqc0izrWeK0l4yk3sylnL82wNVJk/h9Gec+NDLqUYSYEp0I9VFQIKggJAesPBvUMNNdPgvj94jwZUgjbzHExOayfXaiIm/MHg4KombQTaenQ83tsU7HW24k0BD6uWWsF2Fq6QrPnegLbYTwVjX5VyH6on9NMFtIEZi/+GsI09Hglj4dJrlBHcUALSVDDxyyXsMDc/qHl1MeVlVEe4mYdVmrveM5U59nGRgNA82+sJ2YOCKKUp/g6OwhYeSQKsyEq3kQCb7jh5OWBhOT/3aEoVRHrZcBknV6IxXloAl8cxrbd4E8w7Ber9U3FZYP1oMrCUzdlX+/Fy/1kqmniPPMr6TIAiJjww5HJXYff9KjC9jIQ9BuXyy+0y48QO3HDp9uw2NT2K/vLbkPcvqBQPira7RKS2sgUpU6rXi2zSzJCA1IGjILYypVJV2iuRAJXi+vr7p6osnG3ksRPTyX2xEhm8MoS4w2gExwXbT4Z9l36Oh/X/9Bg3q8ZkzLJOi9K5ns6+m7N41+wlJsEPsmMyJSrrtFauq4TMqet+kUexNFhDT4g54fGi98SnQ2WOatzUo32eSlYEwHHucf5SiXJoWZ0+NPwRocVpgk/85scJctsGFuDRJ54gplJHXG8+LVrBW7LdmfYdaTJ+uyyMvPiXWJlhNxEKIfPmi1ZqbRwliaI0jWVavG1ZvVaJ1iM6BRdwQxQj2a6/R4maUwz3aYRLcdZmnEb4+IHkfnuJniWPxzBF6SnG+LxS8xt+ABiVv8RHGn9h/EHQgsgdMy3+829tuoSChi6UttxZXlc0d1lTyV7KS665Rnsw3iTBTpFY8JoUmk+0L3jzsG/IChjwLwxba4tJhyrJPj+dhX6/zjt+X+Py842hgk2MxNlYDzscvxgMfBiGbfvTaFZcz6ZPuK5W2cQl9urcVE1TRc78hr14SUrnr5i6gXEyU4Wy4l42IEAIRWivLDu6iXtRdbYRGFLlvV3DNl1FiTfOpFOyovm9mJr4fCwaUtcjy9DESaPpyhwX1Bj8vnjirqbqbYCc5a+BltF/3Nh2UAsCZfLTX/UzD2U2f3G64Z8OxHZRt+NcJdlrUI4bg2dL1uoiqDU15YJdHO6nlYLDpvg1GByTuMQphoWh2OqygWA75s40vlGfk36SlOprXCwVIu4dmXT3hutnwB+0WDOzc3tGPmbz8zGmARnQkxHdc2Cud6FkCkzxYzuC348xHZ0Lzf4+6FHPadZOh2nZ4DNYLGsOobFFgosrfAj0oaU1nbNyvZxiYic3sRBq8PzU4pIz3/6gqmohtAKqE5qEUQ+/na+1NjMkBM2NyFzo4dJg4twagk3ZdNWrjg0M/d1sZVjVX3aEUl62W00E6epqlCRNRWovR9m1zhSt1Dl9cBpDW7Jar9Oak5kKsiTTyigi0DQijN2wcWfB8s9GcTioSyJ6/dIaSUtg+FRm8LA3LUbRG/tlRWfkPzG2gSgKBCavF76tINCKff2zVOswTYuHHBbmSHs2RsLkAEyh5LjDY0aw05yFXwzGUq8BkQcm6Y9rEHOY2I06IEG+XQEbZsgmxX3mkGe4F0XivoYSbIq2g2ByeDEL0Tf3BH5+Nm2xzd/vSy7cmcVRMzWl02vGBhTheLtLpL3442s0zfHf680uQxVUzRbYIPOwkwJjydWbQphytebCR8l00v46kDnHRrlghWCuuYW9EZVQArXXuLtL3ii8zjbiFHeHVOblLKTAgJhWWroBUJ+5IOBQufohF7jTdzvHwKIijE14dOBNw8sDfEUFUrBR9YUgTzRgDK8F/RTCkM8aIZg1G8/aCfmrLF++uB1b9P75awvQpgMKvIxoU7X7CF9YPjl45g08TBmOQJfewBGSMpyG6E8u2frbQzw73mLYVL9Gt9bQFZPFO4P9CVPGGJLTRgqSjd51SULcr2WjQiifnQ2r7FsWBMGgBJHimWOBkglwwOEA17DZBTuP8j5H8PnUGo2jKUjz4/B3m8/d+CupFr6GBus7nk3SAboh+BarzHE7NZeELdNobGbgd2R8gNLSJkH02GkKMppEzGaOZt1X+lKaOQEmumxKmikknycsNlWTtbxeUIkKx8nLq7K/Sz6m5Gr2VLujEAw4RT3w+C+FOZNV/kG2PezyZ7eqv1m5pZzni13ekusQ6nwfi0CYRcS/vts/qGeQBeEIelZr/GkmUZJHLIwLHbyumu76ZzZx7T7guL9RY3tsS9S5FGLI7oIXWld4bUixtVmmi3cA9tLqWjxZ7FpXvHfPrYmGFSiGk6daDPvtb1G0yNIqE9s5Rua6qtfIxOR2T2hqUW2TQPotTFBPavp33XJT8LLKBoUtT4Bw9NEiwTcziiMD5ewYKKj9/gV635h/8/ZzzxdtsSUwarCWPYg81OK5pTyPEnL4qX7S3MyBHwbudWEDUXNSdIUVs5Fz37R89GXC1WW2l8uWYmD6QH4HKL8axhsS+Ars8yAlBal3URR1EhsJI7fPENbdr+hN5qaE5LYV98rtr0nvh0xpH2u7y/qTBjZ5ttQ6cZiQ0SiUaWPhbPXUVl5jqmg3rPqhPUI1dIBHEe9cMrLdymhV9Siq/OXIlXvmUt4b4jJpGFi9ZMZVVqBYMmPMls/1CwkcsVmVqDww7G0Kb+FuiqL6FFnYVMOIsQNrHNI3UIfj78lfwTk1kAYRn0XrqlrAs2H9Y2dztHVI2GscUeg648NRRp5T9v+QcR6z5vMA7R+g2OdfAzavZV/lYVCiAgxmWbCbiwQ2FX3Q3QCWpCRtowtNrqNCqDKJtqEMACr/jWvsqrtZ7VjNu2qucRHln9Lr3a36Ve7iJx/XO3tbNp0U8Y7+c78KeYso85EzYPbSW9MOjoV6Lf0iWbNUIlSvs1tytqTZVkvLR/+6VM0AANltzPlVMKOJoNvuiAUBQ76v5aqLpdkh8HLmiQOQYxwLShnTZz7AoDDUWW2znfKfFUokWLVhdQGSLJmM2o0odoROpoMjXrt+BUEordtdI9A8Do0q3eWdXLDqOStbqvg3XFO4grtZRLncXBvBTM/vTXUOoEpLhrGVqob6v3nKU6QwM05MkPczJkVn1UqLWQebwYtOr/Issk6CUr7ctHb4seAuShA0IbfYPOKZjkU6YmAlfSyjtCFzdVZK6zJqZdUvL/5a2EHgKcb3EDU5IXVjEJtD44h57MlbAygmR6JfJ7EtbMxpBM25Haz+ti6kvA3W2w+n7mMLwRvR6oKBcZbbVpo4dBZP1+iblVHrvpxQSxQOiNzmkFaTceLn8QH7cgzHRekpiLvDvurWbfwXCV7B567SMCEG5HCnpVYKzeWaX86y99W0otY8tVRlka/E2CtvSBNx2yyNtKGcCQc3fb//zCwYM1wsBa15o+E5Me1kzLn7NgMrfSUJ2JyefCXgIjiazDWymRjKPvJlYqcjzCX29pNLA/O1ITGVghs71yIfjdHAptAixisPcT7hSrlDbBxhP+G8IrF1d25au+iK1W6GZ/35ugPewi88cqzdlznH8MjuaK7PkNGeDUg0P/sI1NIQFXdvHiaSZw7IutUh1Pzy6N1v/eM9y0teom+vzXuhkwdU4vqaXKvg0PoqrXSgxf30zLtTALXmcwfqks4mzfgJNT6LYcONuLdNuNcA+zVtGiEo4IqVSE2gGP3TFKeqym8ZzOSCECZBzccoCfiWDTma1YqK8uHfcve4oQJxJ3bhukaGs4FL8P6GVhf18Lb1NQFB4GjFN75aVwYFbOKNWNCtP/A28/nf5+ohPxCdOigc2eeiEySEYVJH8Rc6UZI5SaIoxc/atp/FzZkL9/XqvanHEyNTOY7kaZIPCopPo8RCmtBTO7lF27LtNPtjRK2RIfZ2iiQB9JIGce3Dcw3xFlqqw+13HBfMjyN7/59Kt7mIALTHwlgPh+mQx4el6gmywT5mYWpAMJAtTAu9EQlKVji+K681HUk1DvDp466KKxbJo+fvvxbDZrT7shLTPPyXPAx1XWixG7rXop8tqRm2870dHhDBUM5cZwSDrYgCimN/6nYrABZqmsNrmPEP1GBhtJkPuP8G2jd1rm6ryBxRF8PuOdEd7K3Wdr5kbu5OsuDEhWtUam3N3oxHolXmWmyas5+OY5GZ5mgd6Jk7vJmYSyx7ugOLOtl/GJSNH1/rpXGG9WFfWHT+T+bYrFjTikOLvLczNGBciwKWb4BkRZYkDetkghwluS1CXu7K5Ot6IlsczHcoTYOK62sTPELh/q8Oww20TmXGlS16rW97cVt7kGHKD86dOMlZMyvwaelptc0hvx7cGrD4hBbk4MnzHzZzF0nY3K6yAuM71z6JL2nU/0M/dEqIrMl984yn0Mbpx57xtE+iKuZ/EKD/qa1doELNxx4mwH8Kg/6U4xlIuI6T2B771zLYFjRTB7aVS1QUuCNzOFWtYQ1s085t96GHZhpr3Gocl/RdCAecy9TQY0O4OFqFg3IteT0Vw1STyZUlTTZWDQ4rVkkC5fdERSccY0tO7v/HvgfiGwADCIZYA6jH3xm37JvBtHTl5A0XILXFY7QCC8U3PT5xpqBRjDp1tnK1aKClQPm6ibgeobEJbw8URIWf1ZjrNGVqNBOyT3SGwftxFNsEio3QOt79IoNHTow+fNM0C5qfEEkazbVPok3EBLWoE/pzzpDL20T8CNT9sjlTgWfPcU68UeuMxRH0mFCJzondVoAdm3sWG2rlpvTYM8KCNKIyKFIDOg3UIsFz9r95JyoNSCC/+VL6dE8uzRK8HN8mV5WunMSMTR72gBvEN+ToLvahsECmbD+3baq1TNQelRhK0QOzAbM+QSQz3s1oFVIc4Jbc0oSRbdWdusT2RQ7n0+SUlzb5yityXefBj2aJEQ0nPuaC1YDMQxBNuQS3XX4ynlkCqYqnan+6t5P5JJfyKWJ5aaqVR2rl9uBwIhwdm7YHBuIXjxrrFPNwuDAtrJgIClfoG45lDnc25syBaMTtyZmy5bFOuHbDsU4D7pHIVaqBuk/Bytq5330eKyatGlsWA/dyjGGVZXnqtcxbO1K9Yx4059ZyA67ImlLHOz6Q3STzxRLHEJeYrvfMeI/8h1Q64Cqj9Z7O0onXbexvuvAlP+nR5qo1PVq3viUMhbmLEar4me21PMJLBlHfjlOzMSg48+eS5axgBc15VDm2gl2wKm3yxW/2fyAszzZWprXvxtog7w4n4D/tlU1+DfzQv3uV79Z6N0Mie4ScYisOIdLzvssWrGnvYcTEAEMIScBZ+fInm3PqFg8Kh9pdWkQEbhLN5PrbXJ26sC3CZ+Nlrf9Bp4nTRrtvSbTjlDR0yr0YuiMCVK6/XPmyRV+YbZ/sPuqWzNy/KKnj+q1tGUk8RrBtge/KntvrNhlrDGq6Y7JTZ7pK+qCMsTcxgtBLTIyJrT3hjHgXNhifi6pbUk9wDRkLy5xhFhJE8AtLy2FvfCo40gGv+wwI84pOqphK4+LbWJ3J7p+FKT9m6HobB3KtmoN3cd6EwBxkJLNBRVrruSkqYHERJqq4NPtuyP9FnHHvvva8MINr/mjyw0hVidPPHwQlmhe0mMsmoAgXbqiv+yCNHXxi6ortDANw3eikCRL509Clfuax8eLQM0debBSBJE+9DEc56r5GYmxR7AtciiWVLkEqijFk5Hc4/Ikkhpo2T8Hg5PP3toa0utvY1NRbhc1laEUjh2k12erHVxTeDGbUqrQdNm4lePl6JWHePj/Gs6OQROimcmnxR8QlJB/BKWMPQnp+OZWFI6Wu5rsgx9OuUhLgUtkOPQsPjLc1EuO03JuwZZNKedP0yE49goGfyANeziTOnHOCUVp2Oz+hNAL4yye8rIkcUTNDrzoER17ZQGCU8NYkq2GQIfU8y1eIC95+UFUznq74+atEBuOSbLDaL8ZHg86dBHAkclXYwP02fpbG+QToyGGwGkjijBTKgTUAgK3rClnvzdrExEHqtTbPLtuCA7aPncX2UjHwHuYBTB/8fvHRIo8Px+AaM5LXFOmR24/KwkbHSIutCCw1HJTrTttHX6DComXIGmhigZ9J0QDRTfHQW1mzAllCkLEGCjzZUxu+q33WphDsPg0hy0vOtS27IdgL4QmLNwe6EQOEpPcN/5HcTqqzKPkeFLEEbeBepUVdfwXed6UyqcqxBVHtOtMa5uikW15+YuncMDgV6cLFzLXF0Xg1EFF6vKyBtiUsHOp9k9qD/ML7A4HRrGVu0Wx1hPs/A6jbxLhXhMebD/d+T/hFaWnzQwzMdRcj9f1TlZSwUyCB0wDFH4ho9i06q6MpGnyHnGW7G0LYjxiYehO5zaVBpJwk+umUFBB056p8llr5eJl5g99x4sNOB34Fft3Nc5YnJ/Qt11OiyRkh6UeukGBSYVslmEBTKSnPiLs2ELwxDqYNjjCMfBRA/gI/29m75uAJmUG9P6xkLzITIx0BnfXL2RTbz2W6TifXk4ymzIKccREn289BX/CxbUIhZVJx6CmFqo+6lhuc5oILvT2m2uBvizGDskE6Zeak35KhYc/WyfgSPqLsLIEDRb6q7cpcXAhWG98K+3CGZraOpW0rYu23BRBEs5sahpAIZemC/any08kza/lu380+CeMPACmGNuV3H92YfhWR0sEA7K2+fPmdORuTNt3NKtb+/vrunxp+fa60jSrj8hg8gePoYF/Nm3D08pWiKCPn4YV7Ocs58QOk2XaaLRNJZ13ZOTFgbO8OBoZQz1Tir72NXNvzIOALRVjnuBhRKzsWvM2O7UAZG4Q2o3G+LoRHIHqR/3witahsllXT4sCkJNyaV1XuKutP7eNAkEqZ1/iNZcpw/DGrZ+z/Po/jlgiZUi/3usugrvPwmBqS2SKzXUsyaiHCiR6SXBgi2EVKrkpTh3jcjiuY7W8/bxySr2G5BJ8LeF1EoOhbeeyP/uBsmbibVp88wJWp+/5rxj/lfwPfE9yd6GAyYppIz8RasyfB0g+sycsDTe7RhE6sRIGLOTNZbc7stjnMWc9mVSc90yIKt3ZzjrTw46j7t/VXzsvvUlRQ5bzjsK2wol/h+9rLR6Iaue90BMLDpUYBdMjTv38uhOak9qBWEVEaBVE860phTFCpO1Oe0z4mMajOcPqKa/qw0VZCvcgmcALX5XIF+jlZ9WxpmAt8gWADqh6jnNMT27KP4CJHkplaNaEHrK+hrngxvsDBBhxlCVzfHoJjDHXii/cOBjP+Ya5iEkGRllm7Pkhw9kqhvfzR3+Vn2ZVV7fddpjxn2AE4K4OJrRL4A20nHXxb3LCWyfQGN/wKLWGjLpbmO2lqKIScRa1yLLhmE+CYud+5kc8KuF+oKtw76DwaiJ3/uGl13cehYlp84JatLlwBsODCMOTOjpbDnlybw2mTcbZ2nVtpOSFYbLtEaxYin95GPMsoT7IzwIahaGFoPTJ8wMhYICrnC4c2qiBGp93njXxEaabsA+C464rHrhJnpIYsmaXUo+RtULu3dYlfTRlfYfVwQ0oE9H46vvYkeuNmTc5GZeobqG+pJv3NGszCj4+Ex/7Z3z5PpraiPVCh+aunKdEbrPUc936FRxXNhWv2PV/rXVyy6faptWKpR+wZD/WCjkK1oOcs3M1zvSR1g6ogS455H+Fga7d94gpMQX/NvNWCYJp/RLz/AUNsi/t11rP2rVAC/C4eA0m48sSC2+qQjJ6bG8M7Wcv43A6qvi97ibmiLpSmwSGP1H+jzzXl7zpkzf6fsYtdwuYqm1MGos7vCXGjVp52zzx/KOeDxdpSr7d73/Atlh6WDiBKH2pggbVCwr1q+0pdBbbyC125tilfyQkoMVHaxZAjB5lH1JlQXnBuXIgAm5pm9sK6ES4okpDePppuaivY1yFM6gIKj8m6hQjtA+3RHwM8XF+5hXsJBgPTFg38+B+NIEXCPZsO3K+Bg/uJ25KXdeJeFWuhv2eCyUGubeS0dOlMl/u2+jokALlQZWjpt+9KQV1sGq9r7cUMgRO4hVggxXooOQzdrYo41hVyc4JP7giZxOZMLPFEq2NpE90eeBuqBbKSXOEeHmUEItbSJv6M3gtGFlf627KjgwQadXYzsZqi8LrOCzIXfSbGctmWYWJLecYcpy39YIQeBZ3ddcxmEN16NvWkq8vXCi1jczkU/RUacv/IR6u+RJdyyu7gAyYHnP99f1EUFWCqbDfXswrR+pcij84Nnn7yYrup1PAhG20IvLdb8FYGz2r8o2Ncoz2MEcmpCwBoXPLKbsGgHjurz6urZEUlUBDSBpxI3tORLNdWPD+pSE1sxSkNqApZ5FMgs9LTdDxVE/TY65wXe1jCNsjL1kP3yiqxM6v3Rv6rMw6/vaot0B4noJ8wEhNQ0oEL8zxbJezqm57L2bAlzwgbdaqHvPR0aYuE1sV+vDt3NgQHe+dkxVyH/tDsPH2t/Lg2ROhHqPi6vY+zZGVce87s1iFiRloxbzz2dF4PU+6K94s2kRM431291wHQVhrrQ4sK4X2red61FfbM/NVL7kwl0YXhk0N5WknoCvalQV0hW5PhJfzmjHkK6cY8qx7MmwPucDRmLrzspSCa61U3eAcA8jfCFIA2B9taVCf8GWlw+/03fbMSmevKIDuOcGnDnZhQyWlDFMpErHHIL6BWqx2AdtsP0JWL05Y47tkrfdFVhMzypu2mE3PmTkDahsQBcJ6EYhsmg8c2d0Xuh/LQCr/TSLVEIRSfy8Qb/a5wjDOUh8JjkdF8AIVD50it2uKc7apS0U2F4FmdmI8EfO65EFsznts3wV2mE0jHe751Eo7+ar4xs+FmqrLQOZ2V8qGFJuQOd1kFBf2vJUQD0OGVCAEhWvY+zcK2sQN9nrQcyZJPVsfhrgVKn14DWCIukmEefjAX4uKIxx6mFDxL7n56Ddl+cwQdJkp1egPYJbAg/KbMQzkewE3+XVTuwV3Jq4251NvdBce6yIGNqv6KpGvs9yL5mh0UbCV2405X7rOKc+DF2AVYJ98cpYonL2lTs/yON8oy4g7RMRj5Kea7hd8NbIXBy86kzVRXS9LQfVLcFhgFFrVR9r8083zSn8IyKg2am07fRkgoypf/mxUcHs3g75x7IMn/mH53xB4rARNG4nIPgN/rdPwppyCpOanMknqBzhFm/K5lHYFtrfw9r6DjrLUQTQkWCY5d8owuFbyiXbB5w67i3mJLjW/2r2lXXoAR4+iuovi+1ZpwT/SM+gaVx7Kd1hlwDK3yDIVRG7mTvlAseW6CYwCQm9/Mx8dtyXfZOthn2k5WrvOXxmTkv47j+8AG55nZi9WGKu4lxkTE9QwnnsVDdGXVcFMvfLqr1tsNUOtz1kTUryTm3gA7ELGHEeoaz+JgA9bgacU+BwzdV7cofzn+aYcTRQRXR3sC/9kcgzSWxanQLbZRv+T7Pqctuh2+FqsAYRghy/ymcftT+xttGV4zqbePuffgYePGlzKpofecqoSUyjb77ChPuEzB119kWQFgKkUPSBYNXAlYhkcW0ZnfFp+yzhGvVadY76rJV18H7nlXlFr4IJx4dOYagyoUEaruhu2+P6gtrRGiU6VaSIsEzuijvhlI1lpJuZ2baHpIKpsVzoEOWZuk7EhWSzSXUlwU4lwJtw3bRUQ6z+gpiuxjdRRUYNJ7f9Yal76XUJkDHtDkzGW8MRVnoUU9503R1xpTHDCDFLZWNJZ8NZRRaUTGkISMVV+nRogI9OCviXSeC6u7WpBG8/9YvqZRvFRSK9zNAHDWMINCp3cQe4xhz/mecJmipUPOfQY08u7xaOpbU2JNNWahgR3Svwn58Tz7VH1ChZ+ZBUkT2o65LO2zDyYVGV8DsByWHf+d0oZIkivQXS1VMtnfBrxECYaTFiizlvHuyk9es6uAK9Fu0+8/GlDsAO4kfvROc0DPRUfNBnXW8pJv9ZVTBkhU8uut6aB6/6ZsK3Pi+rHN1AkJGzelVKm/MPTpedUDvxvcc9vjzSDFukYnXKR/hVXfjNGnfobW5n4u5MxmWkzDKg9jgszRX0CFPoB3f+fVnFovwcko0Qf5On+EA8Q7YdJdrdXeyYJg/a3/sN18V+QBodefdKzT/qHy19s1jhA9Yij34lCi5p36IFwfA6RXW/HmiEnO98Rz9EJKLzQOkJs+W/o+XKB2CLvcNLYZzpHvFmkVFfaiiDFKTINfNkrlDKgBzZTp5XUPkL4Hq7v62E1bkcxoeukWuKIVnLe0qdlV1rrmoSEoe420JeH01cnX1jNr5eHx4h/B8y6CPo0cZxvc+M60zRf45TFoIG6lg+lsILBTicntk1jlkfuegcjh5aiaHepA/ykcSh8rzEAfPbWkUBF2Tlal7xUWtkFbu+uNcB9jvlHwgMryX27Tx0u2VJZnee7l1Cd048ac5PgnIrNiujkC1De1z7XZpDQXPujebCF4gKMNi96ZaH46YdAW0puss+WLbgcec0Zy6gVIPsP49wFbR3c9rygu8bgcJJxLl7QzHVku3K7DpHGdiLBTWraTSPcmid6xMdOk488iNfSF4zI1voXyk9r5vvWz6svwO90ekdiJw+rkvIdxMzbRWqMjNJpAtt7Eh3w5SWMjsd9bP5Mt0x09twSqLfsM/5Eb+4qWjbPZFTdbnTCAkABsXDlFrqUy6/NwAII85OMMOdsz/dM97Cw6YrW68I5Bm/Y4p59xSBKyHvU+a26cAiBnn1SP3JTMMcxDtNjCm8u6yhKDH6RJiVikisXR7M87vsrMIP5lLEIcwUZWpOKXuq7py6g/Ldz4AFmakcNG0r5paWqSBmDEpBAE3s0ZycCh4bx/tSoeXc82ot0fNTrKVBTbbJr2f/1kQCQmjJ99oPTHpRAX8w8auGph5Gy7BFwstiFfttIKdKMe9+q4hS/lWccsISsh7K/t9bsuDUwOhGl1n8+I9bK9H6VCAZDApyZdfkBOwtSOPBvnqD/RLt2vOYTz31S20VYvoXRIwHm1fmGc4KDBy+hyr78zp1/gYK2ga9SF37tuuyo4a9+Ed8oM5BYzVhE0FVb90sybzDLVLOSHu81iBV+AOeQELIVfe5xITJPNG0y1hNQOLV6zHHMx/PCpGW6m42c/KeX8C3l0bOXLG2Mrq6a7PmFJnDuDUaEnuKxT0cctljjFE7xKusdJy71qgfMP6qARKwBn+mq7R/XIi5az0AAy40G9fTwicJsCUidfGPIQufQtvEd3v1hyWTZ+K4M+QPaxzLSIeCseiHdrec98q3r8NgtcFJCU4zVlgegjYSogVDE0wcTDOPELQSm4uU+7SAb1UA+/v8I2EBu7dSMDQS0TQwj/W0JyjW2nJCTzqXQCTdga0u4OzeDUhEktZ8vRpMkkS6KkYWSdowTQlM2v8noKT659p2BmAqtx9m4a5J4a7ZiyqZRFcrbA8Bw70DgNfyDYfJRR7pwZo+P+TBNUbRHCbNqh5QEL0CiPuBpQVmWAoUNBKt+VLNaftCDi9kp+wgfQFDGcZ0wZdHvBFPDmqyXUZ1IF2JqQuRtThTL94WliVXNMTd4wxz+Xt+ujPnIUB4K0rWzgLbaeXRbiEfO16KlH3bw0PKCHvVCMgRC2EnuBf31pXUwEbcAU3OhATi7VwLVmAv7DuSkA8DKaNjgdY1jO4xC8GPH/WEgUXnDfRIpFd8q/NLKFmGT+rFUDU+VGXZNfkpW4h/zphcHQCkXLjBgUuq8OXS1SEMUDPKVQxC4UeaXUzNm4igp79YpS5KgLq3xE2rxNULAkxXXSgNjfSxHOIIhUHvic1w9GE1DIoorrjyKp6hr+1H7igpokGkevhkgLrSRvWOeCncFXv3xl2B+7jvIEWB29QZYdERsqEVIX9HNVtf2A6ASfVXl7r/KS2ZghOVsGTdYmPF0BGj7Sc0todEArYYqRfFyya6zNGV59HugmaU85Y4NS02YGvTG3SYZ1rcAdMun/9vuJ1W/h12Ub/NVXnABdy8x9+mZmncsRzMWuD8a/gYe961FgTvbcRn09go4mKhtJDcOHk+af7XMErNrMrKiOE7sC5jSbiDM885vYTbh1Y4qd5jJOV1V5d4MIVAdUDtl86hJuJf1ajcmfIxiFgeYwQ5J7XicRYNk7xn8HC1Ni/I6TjmgRZdwXGV/pXtyEjMDwupSMVSryXeHoqCBS3FvLcWwv9i5HRmnZFKmjEWsY58v6NC2FSXnzh50H9E/i9IjtbV9TDXwbyUjGUW8Fw5XIJ/ijJPm2s0f4U0QGQA+U7xQjF4KZY0UGXstdjBpY08Cgx/8jRPX7zj1LTVByYZDGZK72hrnEptfmBTTq60vI0kG2zkUQ0BHNeZ4Jhi0Udxvt/HMxn00iaRk1qQrfWQjMHW7zoITjkevt4EEQQI3kqO3enFQpzQ0F8uDVVJC4YkS44SXqIKO8SutZjgHJqIkYUxILpGbyQ/85pgp2kL3wHSbFk/1YiorHtW49um6MPMDe8fW616LFao/j2DDUhF92TSNDP3/Xvl6RbRu5WRaeepRNj5p4AgYNHMFNYgASDOb6uzJQGHlYN//C+iRMstmTlZo5lU3Dow1WRcDhqRVdymPOQa+Y2GfPCKtsVRsjhPDtU3STBz44ZP8EDX+aREis7/D9PM7K2EX62ol9hDsRP8jRukQMhdD5QaLIa8/vKMbR9CAca/Wgn50iR09HX/UHS6t2+NFiE8G7YVdKjiOVNbC2TQ2/RBtyjNeabU4xiyMIrmyiXcM4kXTzTRxH2modbPeMc4/QuBt9XSy80faoDah3qxjFwno4eltZeVdqWYYLPuaC9UteX1Ob69f67AF8juPn3xfE/kS31DojvfBR/u4Uf1yMtzA1xFY8/e/7ZeqgIwNJnAe/Potl+K6qFd9/ssq60OBn07mykGQJvaCANUAcz187V4NqIcWm9tnHDARies8U8jx89Gzk5Fo/o1q7wpuCbfoN4Gt9PGcsvXmemIjUk8gojM8uq6i7wxAEu2E/e6+ywUmszCsLLbo+DlOAjbWojjGY4NnDZK2GIfGxKGhAs+807D7lkyctAPFu/rXwGwvg5ATSTFdkWxo/BSyb6P+fc9+HlzVHYmfWdLZSc2JbS2FGw4MKQV2UD4oWl3MKUmuuvMdaC5JeSwCZWrTQj67bqK6CEVBr/64tcOFu82a0J1a97b901r+H5C+5WJM93XDMd5PvQdzpwCj36jZIXkdBUqj1K6g65cH+jC1dFJElupvKh8Wh05sFWZCF3EAzZAujH+BLiMjgA7A6kLiAj+EGyorJRJ0LEAdnsqIQnnoZRPfiQti6wPUqnxiIOIv6qfpMvVnbA/+SBGFbmfw8TTitk8Dw7X+uAXzFf3gjc7G6Dm8agYdWSPZ9F9h0Lpt++HIcy+W+SYtonlnPTWavMtwEH/+FUqO02tvOo+wcahAkQvjoBXi95q1gqgIUi4WNR+WwIatLrNE/VvJQ5+rQ+69xehL59732h3VQ0kQl+HuOK2KzuSeAeP8qAdujC5RqzlRscsJuB7dAuNO8yZPKup/YkIyPV+s3rBSasIhKuU+T6hNi+9taGjD4p6O5tCLL9frybJXnN6tt2swrscMlSUI/QdzX4jvemNJkjX2xZyPRFBV+ywodmCzpjsLFQxAshu23erxADwvTcJEuuoek3mjLB6wXz6AakFMwZyGpGqA3lZYexDvEn8gFN3/qwXEyev01BL9EtyamGzTCoGervGSq/WRyy80EiguNC7H1cD2WdpxHIHb0v+4roe6QhHVDbbyDaSRP6rEpst5vivMH8yAQKSEJVFHCAAv//Xmyq2ACr7wjH0aT25iUQARTNAoi0X5aDtyeqd8Uo+yGdLFrIJ3izGy91nN6SPGepUaMDvtRmFhlER3uAzXxpFemkKhFuNfdIhz9Su5sF9hNQA5Kqe8vws+U2OJSHzsT24kVSv3EGzHS9BuK1UNdgz20LdrI6af02YArzNljwL1ODuRKd60GSlli9+oU2774X0ngrzmnzNix2dpMpKnu8polJH28674Dppmqd4w2ZrpOC8giYua8mioxMx5A/1H+8yIxtCT61WRD7Hre94qy9xZLE2hhroNMaFXA7cCucjjyLsg40OKDvLtMDPH2lYu7ypGNGc6WTNXXAiqEu8+DMdQW3TOL4GLhPyOVAubaDg+YdN0u5RNwZA6XJO0d4X7/NAoR8Q9ZYnMXxayANUk4PITs9L6dl6Jf0OKuQyFI6IOkfZjcD2oC22FpTaAwjX7xhUKittpSOwOjYL6qhXJETSxDR1OgsMWXTHATjGUc/+6zDOVG4JzJgQticUKyPHiTCh2LcXlxw47HZXGb8IXuBBPIenhEIEfWcm+xj1ODU4SaZg1kqTSnnFfKMdW0yejxih6q2KjzMGW7AegAjH2U8+uBSlUT1nJY=
`pragma protect end_data_block
`pragma protect digest_block
71fca664e6bc359f08255691ca4fd1b693fb9e1f551f5fc87158a1ea0c8960ab
`pragma protect end_digest_block
`pragma protect end_protected
