`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
ym7xSM+SnOoA+G4SqNoFWQhWAjyqDZkfodFOI0NHI6NsNmNVqTlwTINje+NTFoNFdbX5OPEcNdtfBcYbfxuHaueNLXEGdyDXA+6lUzRKp23hntc6rZhmahvpDagXrI1CCuaq/5rUDwu2a9tZiGouSjlSAvc1BRdpj1+/1TdVGV45CV+pK+A9muNW+wzD55mkfmrpIxrErzDGO+auxtm5/gS50T6EqGJ8MV3PXJWJFfl3dlxNx83aVa+4MSVUKpGYc4P1KcsK5gyLIWQj+Y6vHTULUy3Xno+JCN7ZulBlhGca1WLOb9jfFks0AFnU4MOf6ofOcrxV+x6zMaFRRysUAXQzmgC5SPacbY9QFmDyztOnUZpr+Xy20XQ+R8d+76+A2733H640ez9xCWj15908T5Sy+GkgQChu/v2AFJpaFgVgH0PZzd0QTrmb5GKR+MKr5ELaARCpulasrsZygcbJJczmQ9C9gEHEx9+M5lZl78Co7DcDeClr38EBX22BqPIT8z0k9Emi/bf5CRftDZXu5cV53Vk7q4N1pjHDRFKibptZr//i2rf5tgGBZACtgLuOtYSqJaFW9cl2e+IBDf9oQ9e8uB4jN+twHzu7D6NV/WuXfdr1/zdCwzsmCOIcCREyXDFS07hnslVzF+0G54uKUYEiEkQO2d2OUYr5lYbYL8GuaYm4aHQ1OotRwvPZlThWVeb3SXTKxuljmjDqBkkeWqHtSLkA6pB7ZeCuBA3wbFcBkahHH7xugoB3jR3pVrGJpEQ7uwTCZ2bcXqRaKdjWtxN2oJEvOmxYe26wpk9vfy6cRA//RN5YDtnAQ5hm7tqDijvWvmxVOH6zFWHXEyo6iNVSKjBkRquwdRJAeBvhrfGt+Vi1zm6RAR97GiC/x+jR5cUuc1Vz132ZJ4zvW257TePUm2p2frxhOdI8qtOrL4a9OM7vOC5DByEFAGjHgeGUkFLAmrV5gLKLxewb+uKD0Y5Kn/fZfPaWwpk1lwMUAPjlv//YYI/TIED70wREIfkGI0s03IUIGNePkT6T/t+lZ7tUNwdpRhZ0H+0w8Qqjs/V62FtHYjq7OEmo40A+i6q8a4QaEyRJ0Mul5KWj4TETmJtq/ZmWkh7fo1mR/M30qST/fGN2C53AvVZIy76ZhXBDT++YO2gvahAnG0RMHFZCK3ACKA9XkWNkLnB/F2Pxks0XYUTxDoD2YpBEV4VLrpaUHHVUlRpQtxOo9GDTonbtAPphvrS7iDOtLwG/ZIRw77ut1Pp2EofemDyU3+ESlBMrBOmugQMs4PvM6eXBwfpyVBw8xem5gJwTkd8zHOMUoCeAwmYNRqH0OSXP0/yqNCYhPtM/SM5rE6vwHQgSBoyegpVTvulrSSQiY0ZWNvpyhUzpvWBmYv1qn8tf+EUuZYsTHbHFr+zvDW0XSyIsQxG2stYqd02xSJ20leFzroTFjr89v0koJzrXeCzm7P+r9VCcarVJcDrm9MsbK5kXIbZl5BVWsMl53zMGO8cu8YT0v4SQ3yNzKb4TSQ7mFxUsIogNUHa7iCFnhLXi1nKYCXSj2zq/yxeS6wpkFZK3dNxUnEssfZ4odcFT29lP1tIXUyfkCKQVKlsV2pe+v/ueLaKhr8euwwd8ywQXm+o3oVf+Uq+3i5JjN9pWKyrP8vGUJlk8UYKkfmJAaIBzn86+cGM2ws4+S4tWpAo2JP8YTZHQq720pkSYrsYtaq3oFjXSqtQBimCQ9YAwRPf70beLrJHDOKHMiGI8YOhHFpKcPy7Jyp2hQEebjo8xU+3fnxJuGP3TQTTv9wSAXSWvqrhdO73nAwN/rOwK56LwhxhTv2Va59ER2BehAk6JaNbEIlQ/48ZM/TcUNiAI93qrGqIRWTaEucPpqUdgnn7cgUMJXLc65FRLft3VzZTJ6KAp8j2GpJrNe2YDXPKDMYq1aEr5ng0lh3iDCEPujL+r//biafrssLTsoRW8X09yn2xLJ3/lajB8JIS7tpR1qmfXMc8UBvOPyobKFTLCvyzqkwyt/T5RO3Y3nbrBxBiXHPWjWpOarmp+CGB6sWVv3h3WP5bFpT7899tc1hMzLGALOCDouW6EARH4iMNNXYwPQgnTKsll/B9B1ijeMH1Ff5d2HtqmgntD+X1tXgXLlvhAO8ABWNcWzfuL+3+BRWwIYZUls4embr8WbXZ9mjY3zVjw8L7WJqYk0Hhr2+grCUzpppJqImkgHJuPvWGe4AE6e4+WSGRJJtFvlgOjE6xDGLfKJSAp/7IShic74CLGoUazoMAFBL64PVeTlelOptieHI74Uzu5p6y+enBuGJ0oJWk26Nrqn4QUAZvCLDdKPor59VtTFw0Z8JC8nscuZx2JQkhzlWXgMcsFjfunpd8psrmvXS9KnqGeNy3Z0W6fv77NxqKqGePXD6vt8pTBwVEpCghHMNir+EZMTDcMcET5NzSdYtzFyDc7dX4lnwYnzDAbf2lyApW9iiMOHucJllKPejIVtNY5Py8hXU8cOZtZ29Sxqx4GzKlbsmdSWlNDSSX0/BVBmacKPZkyEXSjYfxQynMdtfzNjT1QlhFY09UvKPaFVygT6PNbgkcFZhD1V8JsvKm6G2sVl41IO7v9//GllQEpwJl0+8+rRWjp5Y2r/fTqS90Kfsdami5hgbNGa42aMdBIAFc87Db2yrK+Vze1fP9LIa4xjjskOCp+wRmBHP7j9yEuTSd36nVVRHS+xZIR9lAe5XGcFUuZe0nSf+EHp7jsttpdIKfrrwrvuJN2qhejLawTDOCUDaDi5PIheLJo2QGRLad6nmsNrXmewQSclxuEuNm8yZzgf9CzPAcfO4zNGiimEcKfKzTtMO5/7VJ+lY0b1NxkQp581KzWHSjdrb9VNM0KbnsiqUKNKqQm6V0A3JDt0gCMzp2iBu9Oga/Q1GsIf0UFjXht8ZJpMDPr5kXIxzVKKfB7RYpYZQH0z3FWZVC++D1GpzV6Gv9LBfUbcEw0FyziGF6tnrtu9ab5ibuCBloYpu0yafpRTkM8mbUaxgJK2DnjDmRleGQrMtnP7Xt7QtrlnO9VyN0urMlvlIIZCRl5eCFXV774r5TOhNSBXlmpyZpiXmJuSncOouzc5SwlF1/haamgxKHV87VRbgDenwRPk7kfb89niAQbR0e/Cf6MAsVrWKrxp+qj8g+U8uDxqDe/A/daNTdYWvVQmrlYtQmYafnPO4afGXifcNWj3Bi41SDavICf+FVA+vl8eUKQQrKuD2+ig4RyXo4YPYn7/SXp09yW4X+ux4VHPReEI9JOsWcRmp/+/iVNysfaR0igLDzOqEF0ESi5y8H57x5jXA759PqyYLxnzMLRC1XmTYvGRPiSDXKV2q4pogIT+8C914rt8UJnjqpy+5ROI5xjpdNVDZsSEW/lmUHG++HPBYZ8rjEZKc3/neGRCC3xp0a8KM7E/E+sUH8jy+ZOXG4kpIEhTGXcgLfLlKNG5IYjNDiF0a10/TKwEDu+FTXjS6noPZXFO/cT6Y+cplt2GuEA7BIoLEwCnTL0ujKtpSXO4wpLRn0Ni/8HedYlkFtVSYHeZLHqtw1YbJ0TNFsMYdTH6rN/r00/Zn+W8uy7IENiRFhFk6QRIu15vzvvPZ8YMEvuVJgvnJLKokHeFOib2Yai8FaOM3WGcxqTrm7G7NVUknvMp3suo8iXceTPMcSnJcW/D06pbKW3ce5q+A9q8U+uGX+ypezrCAAt4Vl+xyDx8IBLLAYk101djcl6q1gypphH35dkQqEuQ8L+nLi0aKMgk1mZNumSZiyT4N8hBNUCddtFy5uwwsnTGsuLtkOHEVEtj26D9ZGOPwKU8YB04pxUGiR1O0YIuvr0hUPywPWAhKb67ixUN0UcJ9FGE+NNP27/miA2EV+xFy8tbxGN94084nHH3JOfhbT16dQ8u5FXrg/0pJBl9DMN77wP5t2KhRW2xIAMxy7Qg6nVgD0w1VF3HVl13zsK2Y/DXYVEKVxIvy+BEmrHr8NxI/RSU3TzwFHf6LxJuXe/q7C42IPL9Icy/4qHaFqL0zgMMIun1BtsIKPXi/tIFKCDvjJvfxtzHSvcTUaAV9Yx0ZRdgAcCDYjPnorNHad3C5AdUBnnsLXKU2eEt0WPyQmfn5otuHPd8KvxjE7Y/qhe1iI2D+t3trll5ow9q7x263gWmqJFVIUo9YO0dl1ZgePO0/SFimtSxPLBFtZNG+hRiiO5Z7XDhcSWsgsmF8iTfm97AamSDIdSyIv2aUhd4F8taO1UkWlVJTO0rx+1WcV8Hf7XfBMayGiry7LMBLrwPDjiuwfWxCArb49HYmemiqr1XsG4B+Fza26cyGjWGEz5bvOlm1qOLYloH1Fus/E8VwmBJ2nDK1a9sTdJW4Fct/XNCLKqjSEUT2ffz5ytFwqCLUPxOFv0UZ9yaPnaGWbflYoEESwzeOfc3gioO6pWPyTnlZxKE5i+ytUDlKXEvHNvJtc4jjmA/WahkfB8eOYj68wqqLpYdHGDJSWHEHVGCeH75Lt2K7xIoxG5wGe+JnvF+g1qv4zxLsrBirsg/jDfyL0w4ROZbxBpR//QuThNyc3WqbQjPTq0wjaHrpdRNTg/LcOrxsqvODFJvm5Im+Rb5C5y6+aD/ui48XvQBkF3lEGqGzXHYxJ6MdnX+JjgH3NYpxElTFLC0ek1h4Hp/7kte9YQ11EnojVlYl4hyNyl0ZGThOF4joolYetmvHUJrh9/RmD6t2VrkbiNcsbJtHQx+OldwfSFzq8g0pNbMuhwXX5LeXrddqn9U1ad3LIMxfYuoOVlQLKwVYP8LUqc6OxxrM2cjFzOq7BG3ZnyQy/4+qczh+D8RtPxJf1osrrxF7aoYtRwaThQ7cg5HMR9rRtRJSIXHnqRe2sXEv67lF6OtAhlQFcXqiuJuWJtGvT1gBHygFEfoBbNGNj0uVVaFeH79e0RwEl9U14Z07vR/GmDJ8MqTTeDBFPyJB15quF/u42P+W+CJN4Y10g7z+lnO6sbAt5s8csHy8pZko7uCl1OcRCLxA+dZaT1gh2Q30o1rEAa1/n4SNJtq5a8Dsw9boxR2fCumqQDZRVFQVOqS0EhEchqu53P6ZjSe/1oEry4qys/pgwv4lCUtGMktXbMAloZOFKC0ndc9Uf7E1NDRuLgHwQXlTe+XRrbPWPWIeMnF3KpUy4WZSe2m4SY0SRRBeKqbhohj+M6ynibELtWAG165pFAzyqbZXUYBROiRbob0hNg6vEHNKbB72DbPqWRhGxWZWwVLgO9djQRzH47D+QUdcWFcFOx3O6teYAiBi/zLlac5kf5p+SgLREZFYLHhAaXt5dRTJMIaJzGhuuIP2B+l5/7QI+RQzMUlubE2W2SjUZRNx8zsttycbjefBhnbwolhv/u/Rv/Bns45H73goja0pxtNMGkDJqIvqhRfks9t8L/ED/tPC5KFqnv7g6Jah6JERJxHIW6YXxULE5k4XuEr9ICadPt2Lo0vo2g41JgB1MmZS/EzUDiRGSxzty3uAbSDf7VUXwqEt6yjAo5MwrU0LvQhRnvfR2pAnT10nHAF+nXXBDCimj58IBOFbn/GN30UXaAzVSy8Rc34AgZffDVyx9ocK5wFA5XCwKpctANJ0PCQk4nm4sW+F2yrp4KSSGbkd+/i/RuK4m4ON1IID2C/2Aifq+IMYitihm2CQPTEArVu5Z4fAPZbHpujzgOUfYNrUiWMXpguXkT8l8l02gPCHSydxerD5jPRBPGoEF7UBdfIAWXTQ/tCgBgucBojsmu9ZLX7HkkKaQi8JPJYBYYitlOu877AGthBtWtuhAGkO77TUdsZiUpCB7P9bI2lJkMc///zBUQK9UOj27Y52RPnggQ4R0Lmyx3gnXMFBl1ZWp8jKQ643oLrLGAKs6VHQc+uplbS/J3J90AjvLmXt0MvjI/NW179JrbmSpWfMa9+7y9iHRp0K3eH4Acv6LeZpaSSvJJctIKgRdsCGDZF/339McwRyVY4nxbyuAxeJ0PN+fIRQK8oNyerRZu/zhQOxaNx/wqR0LTMyb5iPEcEVukwVCwgSNodkNOL2ae9BHDEsf1j8pofcrMxDEQTq3K40gzYSS3vJoMKrlea74LDtwmZBlUiqmYgFD2kMAYqYVGLljkvoHmSE+I7KvZWcfCJKKIi5/02BrnlG7e5O61fTGOwc0hjSeO09cH/kd/EL2l6wCynK+F3X/TtWoBBGg+DdOyPB844/Kw28OC0ULWe8dEEhIYpRGU54PV0xg4JVgLSxTWlBU0kTwgFTkqnztxyDGRp8ZMedLnHPlq2pjLNAQwiIFH55b+FA+vr+dsIyQXeCGd1SEJ/flDAQJcv3HunEOcnI0mZhHvnaba8KU/rc6mFXHOfIDVAHUY7omeVziC/xkh9KZttpHuir0OdXLWGHhu6w88/mH7rbtpU97iilENJg2nFRFa8LfxfLGxlP82Bp0GPivBldRyFdEQEuAUSU5ujI0bjXjguP6YW+EeuND4a3wSziLNooDGCXLnQtXOPWnYNhvDZIXreSlOObm4ozp/idliXSHDvLnhmSbNReWE/O4OnxkW2Eo5A0L5myBJt+D96BgqQeN/dNZQm+04ZJOV10ndkXmhIk9JduEfmqKvCME2JM8bHZoFHLZCID8rqn//bv6xqIG6J0w/xnOu6vVVp9v2X5TYZP/A14qqpTd2V6bXkQ3W1PfanYVRzHMrKHnPyJRufyr+CFEpVG5+LKiZaYp9PbdUv5N3qhH6+PfC5QYo04MH1grRkYTWVyfwohWNYJlOkkxTf+6cYgy3DFSrUq1tD4S7HcHeaFFJ6S3b8evm8bc7gR+tEWY6Sedrk8tPaevX04LD0nuYXKGUpI6k3Sa4j3taAMKJt2GQd6cC5+br/s9FSxTf1Nu2hq93SJZ4hY2lhCDRMTOMHlk8Cloi4caqwVQDIWQ+YXy83wjYs7Wxw5oSJfssrxoqkhnESTUkfz2c4ivu5Lmgz4CiOTnMfoQtCEx+mKU+pelv4Tbo2fXbWLdoCF2OG/7eIjHUsXu0NN/M/1FLA4eFQERkMhhUy/ExJuSo4renDbbm1dDZN/6DT9rwb18AnKS/b1F32xCxZhNpGlusmTvuXmsYdibcPKxKHECE0HtSbN0+MNItyBMT4UGWZBP9sU2/6IIykpwBNpRtedAQefwrV28UZRvFtI3Cup/FkmiaHdOmckv1ZkJFpv2KFeojyAoul2UwskGXrvT5ygcZE1KEHuDPYdZJwCJh3mjMZPD0avRMmySuaIrf7oXmUaWqUgWSoM3iWtWGrUF6oTRtkOzSuCpbGLRXi+gyJ2ovEQ4aH0iwzO+UGXBBNeyOlaZqdDc8ZJzniyrE6nl/VmiFNHbcCGdBioMajdSwWNw/qA57wvS7wL6tcGULaH5/NixNj0NmxQWx2gTmSJZXbCyg8VvD9hJkq2r48k6b7f1N8FF1PR0IKf3AqAUA8deGVOCs/ORYlXhMizqcYPGftna1o+zYvQ5LZXEqH3oJiGt3lO2Czuj4FY1Y3A1bHc5imsDBL7bnqe5YXN4lm+4w049iu6TAb6sPvRoFL5rFOFfk6wnc9FvaP5SsUk9n+YGlD1OaLp86UyaqzVlJ1km+7HPBM5M8UJt/HW+ywvPMRNlW77pe62GEGDqkSVFW+xq4n8uSffwDDjkeerMV/cPGTqxi9lyBYM/mh9bKAQuuBKeTDela2Zn8OEC6HhetaDAvSIYBpoYEu0mFNV8aC4jjT/CJ6q9pCxL5XK4rcyIOq/tL2ZHAsyxfRIPW0xgGbkCuOVjtcCaKzJTdskKdXfS/jy1QLq1NyjGn1vbNaEyVYrqQB80qi9QFGIUUgrA/cO/HDMuYySdrncaazNOsnqzfo4IqlRIjEm3opm+APwckB295GqSpXtg+vzjUpWidFkHqbafnkzuntLbAi6k16tg4P9gQlaH8dsV4SDEnAGK5paxSfQCzYiL05GesQm7bTcn1Q1j8G/KDq9csHfn3/kvHjnDxUhS9OGRtRMkMSatA3wRHgehnnjIrjeSv2DKlXEI2OIyKy4kWMTsp2qfKm/J/ElIREdrEI0F8QUvlznZVONENe638ZCv2uN3w43odlojXZtNuGZSKpjNzJ8+f1Ue+ZgJvy2EYcM0rTBpdSGM4K7C8c9LZ5yIBbiso5io1gu2cvuIT2HB+GuddcYwwRGCY79KU9lP50TfDfX1AwQ18U6foPT9pS006HF/SlJ6Sm8O+93Wo4gnNvnvCISgDQ3Ea75pI2E0sZADlDMx7o6sSVjwxWvV9mG4SZUHraYga3I3P7JDgqoDd8bVcs1LKRwOqA3tR2ni90BSWojDdGOc18g1a6qlIGWwU6aXlEBcUOnCbtOVqNqdHDKs1LBuYeo9H7/ghBL3pfDtBVy6XUv2ZhNHJYDe82BWJJ7TKzdWBGkBq4/6sXkwCf41QBPMvOTYF8DecK74Z8KnZj+8owgk8BVo0TQNc6Km8tXjNTmySzxOR3o5Iu+7NYmWlKwS4+GTO9Ig/NJVZsXVosqM6htaK7fmlOpCdZ/m5LH3PpjmmyyB1lTuVGxKr7MmP6aY5Pb1S9fSeFoaiXr8FHY5Q/+F9jbWx+ag0bRtfMvzgYms4XjcvGgPIPsygCGZ9uZOb1rKzl5r/ipeUr6dm1S2qZjl+wQa/dB9WHhJoQ92Ohilp1V09mv/Y+KvrbxNv3zXzZu5MF6DsP1vcYUIfayDjmY8tQawdgVsoEStcvw6kQAN0rVJlobtOhUQlfgEn7NQ4KpIAEpqYnOP2XZOwq69QXFwJNwZyEEUEiedBKt84b0OELBHZtx3cHUuwPKRZIiHbYUrdWvf3HzKwLZtsaKogOgUf+chz1WXaJqL1Za+5aDEDYwCBFz7ghfXgxl7UA/OpEMEzu80WcLfb4RyyePPt+NTdA9P8jl8xlcAeWd++pcQxIqN4xNgY57laJdmdOja+8U3u+fCLmuAF7JDjttrVXHXFPL8IkTUElyNHUFdqoD5oMO6fP1O5jE5bFNpYzkeUK2kn3oqg5hrLFcf4SsQpl0TsZCORjJVf4+LTLoNrXA4xrLieb6wPm1IE644T/bu3bwkG7jcCckxEdSWQ96kcl49C0AX6ZEaheiQJuSfkZ+HBvm3YF7WjR+APSxsaQQT+jQdXsc9A8JSnHmWA6vGo/0jcD68cZ7kzXdAx60+Zl+oafV22evqaQAtrXkIurqEIXlQXXyzImywUfTizmEGqXD2q8/tuSiWzhtnUKmcv8k60aShQ2faVnIE7atTuKHyQBGM3t2oDu5Y83RX1+KSaYlg+nvXlOIGoW3mv7SfdKfab8E9CZa+om6CXHwfuHrjd/2jdbhvlLJxggM1xctUuJQJ17zQsl+u3IFuwekcRny+GNW6y36kish7w2HkW+Xs2Z0AaDjkIyPE3XvBKvswSohBi9ROrW+pIOhGBAMtvgzSmvYsOsfV4Hk6DTbNEBL2lpLWsflGF6TxZMxYzxYoa6DwDgQacegIr8Ns+eibtRrCd/udIFZlm8lvf+06ipV3OfnsozK2Iw4TDZOCIoHOTphFMQ6+qBWyaAXHltV2p2JFRDSxALBfMCQXX+9cf6kHuoou+Ul1b3kRimeGYdogAZEbqlF7GNUOVKrOzaYRz+ONqE0zM96RKlZItihjEOPp3rzfpRa1DwD8CA75d138gIH9T1m3IFs11LuWJ1WC1bfp4OLLw77DVDUASPj326L1C4wMrJLNlNB6MBfinZwAA8F7JP4Yju4drlUAnKOlB8DtX92hKzLi0Li7kyB3KSy/Mcs4/TuKKJ+zVHFJNkH9qmTRPLZ8xdtDY8YRxihWMMrhhySJ3rnW5mqz+vbFOJqsYUwnoLTrEfEhXAVmajRT3Rr8WPEYrfxM9R6thg44IV7K2L16nPmcnGdlJEiOFGpVrqu43t9i7S/Zae8FJJQ65TQiNoc8nLKAGk6Z59Si/c0LS3ae1VztibEByp50u4MioWhN4fjgZsII6M9VqpH5mvXMCJlKnSb1FPjLHO1hOgKhIGenx/qmw2WVksxLOIFLQUYl8y5sGkNCpCnijHuHSAHMM47yqqmBKpAGSOQjRNaoipAbJVvOvJ9nXAuwEl4h6nqcjdnGEoaMI8qHeZ+gj0XhyFvIzATQ4k4Rz441R5VQbTrQJklGPgXFdcVJBzNQo9l5R61ndMH/a6MqG+cofdA6WygHUoOkVlu4BK504gzb13cyNOjFGH4iy8zY7whUQHrldGc8XpPW9ImWebXwIFUICO4MlJ/XhogkbQ2RWk0D3nrFXLA68fg+DrzbrPVX/2r661EKjhrbNbkUcSBmyfc2lGCZMgnCbXzOLbFLi2lkTsWTKqabfW1q7bsNjc9000oXtN0hJF/1aluyls1kSElCRAhU1Bzfi6i33tfsL67eqO9wDj6IGdtCv+kz0zQrqgBY8DYUXnKnmeYYoViDln2kdw1ZLeMMLk70jdxYl+2grjfvL6q/pbmBANalgLM1xilrSgqb2riKGM3g+KW7UjvPPj5gZWQcaELuFRgMGqK4wehP1EQMCL/Bu5X8OBKDSpmStIlMU3PemKz8rq4htoDYPoXpBPHPptEDZaAbpJBW46ggataXibxf405mFm/QyTKZESDJrUQK0o2NObmvdV+OX4tdoPmq9LxvlZdyLXrOobYqUGr6r5oDgt0i6Sv8VrQvKsYuS4PL23O4TRDm6Qe0wLZkqtfXwf/ckG9HmvD5qC2W8ESh4vGYzSGx1rTk9QbUyZz9YqgrQDPvWmZaAwsInKpKvj1r7nGVmf1QAgd2oKNx307zIVT6+7tZWvhba5E0KXwWbgXfdHKRp0B1XkVcW8G9BDzn0j+sKPMo6f2frDlR7Sj2f6KdfN1yucQMQ0B2L+mGc9YQ5/Or3Snpzeu2d5Get/KUG97Xs8zSevcK6gtFyhnq/Uxwv8pL/DLz5uzWl+krr1gq0R5/25svJYBiJ4CU5OVexR4LOwv/ThE67w5po7T9jva2W/1Ju+Xz8PLVBeHaGB9fnr+NyzLZbFcydFx594bZBNLv+3mJbWtz677VouRmI3jkKZ20xsiBB2WtTookr/QaZs03+eASPlwd/gnyerD/GGyXH7kDUrZY5tMSDykz7Pq6CqVdebIAkcRF/NA4eEkL0FCy/VbLZN/jz6bdUk/VT/EAlgooNCkZ92eFuRb96Lnbc4nql84JSkO5DD7vCMRpLIhCB0uom1NUROW8BvCBDQNI8OrmomJySwkD81yuIB0O0SJHBX9bMJA3Jz0zmEo2GIxKLdLJEulNUBFFEaQmDZTrI18qkCDRIioXLMj2SBAkKPoTzUaVWtbpJtZ41vcLow/BQUL02sKycnHZb9zzPFs0++syf/jNyi5fOGBAhEN3HC2a3lqz4vCg7zDqMlJmUw9vSHMdLsEiWHoWoDWEXOhxgt7y/9oo88eIz/a3j/P1mNWbciW7I3n0Vy61Yi9UsrUWlz3eypN05TUIcdS1Tkx8q2ZphoJI+/8YLFUnES1eE0Duu7mrcO4A4WckqzBopnAUhDvjvYY8WbW1PTLiNSYFNL9bSn36EXPTqaIKR0ENwzgWsyE2Bv+vU2n1CzZlSYk0W/UpJcV/iXfSg8nh/tesfolW2V70kb2x7yvI7cZnhkek2qa1goNPvPAnSR4UVGEFV2nCWUUFOxwOqSQ84UpKvbvm+FAeRSauo9RQ0xWaIZolskNj4cYLv/eIR0KD5HkQwes9Sxir0qSOMVY5KdWqnT6YPQs1vkMKMcodJ/dLdTxL8Zzano2/aMO8XuEjQsGK6CGkxdCcVT3t6m0T7/1Iy9exyJxHhQ1fOYbB81WxrJD6zGWrZ8GseIDD13vmR7whOBf3XDhPT5rErz5eqVAkruzW6/+2NgCF8yRdaM/lq662fvqnjRBmpSHv5hdqi2IiSFD5fTABslpsckUJ8eXq05EhQV2r6OR4GOr2WReuapz/LR3tlUg8UvRRqbnrq9y9PtfG5y4kFg3FMtQQQQw7aqKPyXtzRprE5w0KStGZUTyW7pGT5KR6MjjtNLb2KQ6Es+cfZK8gZnklPgnW+mZLD5AdoLYaz/PRC4AnPvvXZVJkNm1gB0wjlB/JkbqNgNnQpTyjbZ+GpkykZzQtsKXUVpPkehAYtYyDc1lZDsk8OSVh1Rzp4ny7vPCefrDYbYeqNc6az+Ny+/RNXf2s+n2swtfza13HBVYvTILUB1g8DZy0wtJSJ1cYXxNM5wOZSl1iKfrr/5GjDt/vqtdPMmJCnKg+izft7RXw4Y6b+R5mPzASKYeH9ECQ7qYu7wgUxj3OnE1RJIFT+L3YjczkZ64xYHse2iqIrBfYlTz4mW+EB56DGxefQ0vdtZBzH46F18AMwbnI0VcaIFE8c+jSL+yVTNnsRS0H+ef8HGfZcFgPQh7TUQlN7gS99qBV+TAamhsEl+AEkGHPkKWFlydMX4YsGynKDA5hzhbzJDVAFznvSCHiv1FrK9sKSEQqNGguWmJGcdnjuOQr1AeXgdefi7cBY9TmfpS52Hx9KOKYbQqvyMO3AR6omkMnDT2D7NQEWASv5li0Lwm70BNJQH14Vr4EaTHN163VXbUErUbfJPvdIsrjUn2gQPh5wzyFOy1DEVTgHy1Dw8ul0OZhOWXUdAQu/Q/AXfIpM4Ur7NBTUCEWC9uelRSPENMLJG8w8X6wosnlKQRJMzUHS2jyqK7sg8KbCfKD2ebHaPewyeZH7+wCBQ2FnOhd5fHIaAw9XWQ04whsG58U7Rxl3ZSs6k0aDPTg3O4CipbajbRRwRdcjo2+LDgaaFrURrReMTvMHeWt7K7vZIBoApmALKmjdjbhOL7gfgmmCgeWaP6ejisDd8Gatzcd7ggwC7QaJDjGMV3OnJdQj15XPKx/NnEup1DJkLsgCmdvmoYSbJ7pNGDTTLOTMhr0pG+U9pYmBGjxiW3UIPV6Xh4IzEPW+hVwkbhTQdLDYcEA1EaR01jPITyLqfrIZNt+EpJ/wr0pnVSJiaBwhO8OOGvKgdUZe8SprjnF7XTXvXRr8FlP26KOhT7QcmTaSk7R+Sp9lQKJSlQBkxV+U7q6leDhJgJ4IrXBx46Lm4DPp6q6hH/zYCUJAAOpOVpAmMZEO8rc1psqozkDi24/5sywi2SzC0ipdGTYNevm/ttmM9OYruvDzq3cTzG6eukKOqpDOH2QDmIgZjfN24JuPZZcbVfbOUoVSo3RAcSj85TGScvJqTY6+5lYiogIALtYXhoM3YB9j1eW92oFzwQldu3sTvfg5ssfGzddI7cpr9xWO58CU/dfn9XkitsBsU04US0FS6uRn+hNMAj+e7ExGE712Tk+/7i67HzhnkakKyUrC8CTXzrRE1+6rEtCdw+F+3klZS1MLoaZExS561C4O17gNlLXl7au1ZXZmOK6sihXAYrYNCRsrnQwSoQlD12cVxuvIDbvYkeP5y0X+nlY7N1Jqjye7seZTQCth3zt350LZjzc6IUKA3+aXLlpTFqF5Nq0dKd2Ww+LLT/MPCgPqW/pUDvd1CTWNLW3nAzCssK8Nfv4rvavXdheGDe/xoLPy19zMtmkSh8qldfAiINkdjBxMt5TqoTrQqfh0+Dpb0XNBKQ8JOeBXwvBRP0wGHbmGh0yelBQCVTtrnU5IxaCX42a/hWFsHym4rrqV1Wkh7YbtCToqUrjdXLsRsvbNHSp4YQH81WCiefGC+gfkG1WfJpa+9rudgcNrDYiVtDMPBt4/ooYOVGycu4rxvAl7FXRQHcPCjlmFL3BPZUZcypygCCc0mOpy/USHzfKIEcXDN4UEM+suLzyJzgeF5MmkY93cQ3NEDQ0aHfP5oTNhXokE8LLonGAnTLnuOl/olMa8EFdySC9aGz49ChHun1h5MFcMr9N642q43J09r2DTvOSBF/oU4ouCzNvv/xdviu3sivD+G++uI3hM9P/3LdLatWK91408xEFlWouaZB+84kz5ooZCPZQoK7kbMlSOlXbdwhQitkmpZDHPZ1FKxSzYecsiYlnrD8ELj2N4MszR3wQtJr3/ZLHgnLpagHedJGN88Z+L9uaOm+tFHWP9Dh8vwi+sMrZ+TqRM5sddUbHGW1BhTOQiQaT8RIRLYsOhr45Xpk6Q4jkC5jNcPhCJ///E2PRY9NVoQHZbsD7DdhgUmwrJnerRyvmO2cvtZNM4CkRIct+tKGMiCvNhIxrje2XoMPc8ZypIW0bts7KWKTIdLshtZ9EG2z7zTlWuWHwPqFNY5Y339548GXhaFkLj133aQvhoN1NmeUyttznQ4EJaKH9pJVrTG5Q12brlHIjcmioxaRvKeedUegfn1LKmed6DSrauAZRQCVxgpMYZ9+f9/tcj/XeNpZSw5YWcBeCQV/P1qVt2A9Yz3p3WOPRy0wyZ9RvXYYSdQp8HP4GwgNsWTpZOb6qaYKEtVbxNVz4S6RbyrF6ixSSuKTzNr9YDHXpBDOXoUshIxxjfQbbR9RxjY8n7lRJWdDXXbnY+Q4uaWu4dDvOwX0pvIhzLXtbTyjjITHSXMdXxac/HDM/AJVE5+uuqzIjXhjIahhYuVhtM4vutCABdy+XY3AsGz/8p+eI6z/e0CYGEgWuTwB3YHB4wv+XePmkB8wFXzuXMM7FvLEbdrKl0dbxarvrdj3xDFLyvzIb/KhGOH1fyWBOpGJZcncz50n8jvJSvORfhmF8FGByRU+AYT6sVd8UFLIoQ5k5NWAhIqj8vxBtJgmYug7pfAPl8JkgLqaI6V6XRRtZxqJmvhT8tGPBwlgZNepDKDnGPyqbrC+00abR+kouFrw8VxWTit0jxbe+bV0iV4aa1fOCPFON4TpAl+4b281J5FgF6r56dZ1tuphr0IGo4KnmfjK69+96wUiH6ywoA/lrDpOUtnNvX5RNtln77RZ829STyGpvPwFNg8V3njvM7dssCQbrJz5rH3UpV4WeWg0tzTWWYL6lq42TTdW6NI5vMulwZJqn9WTbzy05XcQmzSMpHsC5C8GTiiq6ZOTqoRfXZp+DbfoCq6VAkEMQQs169tyZuvnzH3CF68ShKfxGvZJFPLuEoDuZ98CZoAwp9RvWmdZQDc/ND040SOvFFsnhd1NMZIKzbhgJE4qPOVD9EDW9xCV2U8mRB8NffzVbwxNixHDcY3lzXBJJZhQ==
`pragma protect end_data_block
`pragma protect digest_block
dcf1e0e3cdf33281cbdbdce5ef5d0510d793e470a668971da52b7cafea651183
`pragma protect end_digest_block
`pragma protect end_protected
