`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
CexAhvl+uGlnhUQbCzOXWJzxBZy9dywf2jYyk8E4I0bOyIRkFpuJesc22etSMOI+CSIo5vzEY0FyOZB24/0WhMc5sSCXIYuiQiRXUfJNMGA3iWqDN2rZZcb7RDI0Oypg5hXL3BfJyfF4gjyUjt4eN9QZUj5xXIUdBHxSrflJMxXRLVUr2ca8Z6Y5ZG4QXTpYdJFFllFB2kOj6knMjOHBlGwBJ1M/p05wCU85GteA19DvpBD1NScNFiZ8tz2m/e9bySX/O44sM2SOZthLKgb5RqfHjs1iiTGpGDrsxviZz+Q/PhUkE95G9RFK+FHOstqkMg6swzXFIQ1bbM63/ma2ffPZ9QlHA1cDguFG1esKkqb03GARF/YpcNw1kcC45R/BvUP5U8u07he4e8p0rA8gMldi++5l5NCsEAeHOpxmWv8fJyrD8nBuJKv27vNkkP1+NIG5eL4lFOd5F52wIETSPicLT6Y92o2RK2TSeKM1TnblZfh1JbcxulgMo2giqpeyCpNGV/Ik8HjmvZA+9HXMB+SLxm7dDncRhhJffKV0HhXzoNxt/9Ju1lFRDstnKdJbxRL/QDcxuJMovZ/1glK6DKnqZyH3UgBR+WOgWlEjzcAY3bBFrDIZe2MG5TTtm4aZKyZMemCuQXOa8tNE6Jg2oBu4TqRE6E61jL3aQiRlaGoPShZdDD/OSU1wv7/I2z7pt1xLO9LE9s7xawwHWEtaKq7MAI74tD1E/s6cFkcmdZnrET9G7W1fQi/0Ovumb/HJQ1kIpYwbmyPjniTgSs6a+SGTIgO3eYOnaKlLU+OgeYjYlyaTMp2HeznoXN7wIvHS7Hs6WbS/0B0zyUj02Ryg8n7HH8H56UbtisHv0dzEuWv/Vv8Q+DlC9SOb5Y5AEKJG89LmS9XSVkBk5Y0o30B2Qin5p3AH0yPJIama4BaNbx4hpsQH3OES0NaYMlx9LnHzlNTsYWjpeIhmLiohdAiHO0nD5jOGtcY6fIyYH+oWSu448tp4qiX3n4NlRMm3R+crpJ9/s6Z394/8XBFizjEHgtN3+Y3J60TXD1r3WigNEIyQmZlKExVHbpzCa2ZCwxMwn5VD9ol2RQH4LtVTNh+JOIImzpQKefGKeKf+e9EsvFvO1sepgWjAVk1mSOBAuBzdlCAS3ADCnY7NppL5caIbQNzsO7CLCL4lpvWjVDGT9TgfbK7RzJwXAxvO8Fz92wrWs3jEblICE03o74BbrhVEpzvk9QfSKC5iDz+9t6fAn2Nlq8Mu2BdfhWs6JBZyFOa9qdqV0SRMM2hfRw3Bm4vBW0iOPB08tHS4528r8G4ryPn/PxdS1PqVtvZO1SyZKlAnaHSPFQhBySM/ZmsPZ1SYU4TGcSr0/1C2UPbOep64rPEtNKescnPEEYueCfAc99J9buXxSOybISU+TGmQwj6su2cw2EhoHCEuURxuqirN5IKtQtB1/fv+4cvKWuq6ylYOYbh0OwdWLzrU7wxQ1miwIedrnWRhs/8Fge8Ia5ZZ+PPQFsvtaGJxNRQtkyTPKDBqLQRlkrerK76MM9U6ZKfaYUerPd5T4dxcLo6GGeJMnGClEBKpO9QPZEWjCRZwrjShJHeEw3pL2UgZHVR4AmRkIg++/gdqCm2yX3+7m2YJJg+q0CZDkwgm7gPSSLqdNAaUtC6bJNIR3s55pzBZQXjRheDGrc8CQ6PQHs2eKul8u253JtESVUxO1MrQa96zOIbpfpD7CRBSrRhsRnvxF2Xl3oyHpJ3kSOo+xI5HOMeVrUViMkfrfykEAnpv6mBsOUY5byt0SEzYG7TZHlb2tzS4AeKQDSETdnOR6T2nAo75FjYUeXNgfV7XkMvZvNfEtoBpZxCfTd27+vSpoekNtijlcbVKGCXgERmwMoJyHbpk9YOLpmYQrYIvhsUjUDXyg9cTIsNGAAI6BToSfsTbYQIHumFwTvu5UhxwCbmAwEdwvVw8CeyunaBujBb+09LuNclbh+/VMMfeTNNuGm4TIFmgpU51vOo3FO9v/L/1nGJr8+cHw9SqwB5ECGNxAfEIi6hzdceSFIZ1jQnRP74HzBLW++IoplYJ8E3JnRvt/WnxGnDrZDsbNWYAaX/WLDXeaPS9q6LDyupQDxDW8vH7ibvQsf6pgnZiUC9c2JurUufE3ThJjkZqd/M2yl2ZNJcZsCvflJjTZOa0wTEqGPZeoviA/1GYh70O3f+uKr4aJvFJbu+CAda8uXYBuYLd+hq9yl+U/lneNgdm+TTN7AfoX5NYK4hMcjUkL5vuZGkNx4qncriPdEks3kKnyJULZi+VJ/E9vQ5VqjigNRSPmW9dABvMUXu2gPMi2u/mq1zblYfKEYUD4H3571bpQnA+QE4BgrfnSbs3blBZQOz9ARhJkCh3Mhv3AdGPFmj3mgY/0jpLZWXdYTjhsjywIvRbSvMp8jhxHcxtm4j2HoXUEOxOkksh5QFXEUSj2X/Jm5j6uwJkC4Nltui9JS4EoFdjbxzmm3WrSkTs4Tg1cTrkYvW19tf3xwWW+3XmmimYsyY5JPW9E9SPmEkQgOrveO5oitOhVtHHu/BNI3RnkhNSKonl788JrX/L26l1o5U5oR+dBhRLsF+0SnRJ+sc5TwCkrfMyfnTHnmXNusRsDyh0IQSSLzk1m2E28vlwch34IzkLl5C3iKwOHLSBt21jj9SpNLyQrDjBLD7uw2EBaAABZsZoGs2z9d13CbmDUumvEb/S27bDPuDz6qaH0/nVvyqshJFC3UQ/lNHIxgwthSTkYtTv9KTX8RP6gEd9L5Fyl1Yk2HCZdRmz1CEDX3g+EvR/pqQMxtMUR+L0RaISn1+V42AbyqQQX99LVL/gyyLnmXTQCEToFRX3LCGfAWLShIqrk/2rfYteLNSh40eg2HVwAkkIf5nsrvbvxaMS5GuTmFUDXTHslEbD/IhsVi5Oplc9p8M1DJUo76xHfw1OHojHrpNQsvRgpZTj6o26742jaoQOMQ1PWBIWmSRzR3IJsxGhIMxlthuz12mFSLJxzId7hTewzxkQgZnaaNfFk4Ki1IfBa8FenFUAXtbzYMATmmyat3Dx5u58S2gE2AK8zQtT++feFHMKpTQPySe8e37BDhC+tlmeye2BuIL4PqS6GOAMBuqh/bJHhr4lSiK5QIT72k5Uql10A2TUXu4zz/Ar5Q1Rw/5CRnZL5lNHB5K80jynXY3+TaKgvt7zgHhpOEuZ+cIAasbgFAsArmGQc7lPL13+vVtYiLxbNMU+qaE5IYCy6fyhelm7DP6OKL/Erro71zFhevZq7pa4cgenpV4aEoLljeq850njLbUkr8FL5mPUxmPMRp5+oYQXeIl3bfP2w5ik7ybUR/8QrxLYjANwOL149E1wxfHFG1eARs4M4/D51/5nzyUdZ7RZ+kfQ/+ZnryWckZweGVjwKeyTM+nIyTVRmxJV9hjgmM1BuLuK2JQdX+CWDk+24jWlRPZmLSnPMhqDa9J5MUTHpVyJIK3XATqcGvwgByeuT6mY40bcSacrvD1twDJJbALnGh3Zthnnv6YgaSM9xl12hXONYYWFg6xvFtNqke8swoOtClWWP8eARyWaUIW/tUJ9IhK/vabaX9WLhr+G0k6ClGjNjOfgxl10KD9oePmolQlftS5eHlsFmGZzMnYoQaPi9Zpm4rp1Rhummmw6oqSisKksyO2kui+TNRiZNvoOyrwCH9EeQ+gT+XSgQbmF/TQn+0NUeImImZNyWXxbO6FoxbMbLdaT5b8eUnroUGr+tFxSNN8M18Tfd1TFW0krLcN0bedt5O47cSfxoqmz1SfbkmQE1kXPg1ZHtrLDBG4H5nexMBe4Zm34WCUcNgYF0JW8/ge1BW7D2iizsQnCHKSSh9unj/kOvPCztLa+TxWqPS/F1flTvo9SiCtLIcaH9CRt7mVjVoNyClmtJuKQKAOoK2t/bk1Xo8k0MAzoX2qMxBwuP9HGZvSRHnZXjZa13cj4F70RObeN51oXP/sUhcxiLybu2aTSS6m9E0Ttisj8cchkAOKI+nQ2Yr6Plg8ITa6Gd+fCkub+rsCgdcgn94p4eh/GvWD50UQZNebKAr1x6bY83vBVTJlpa8lfFNgCgn/9qLbRvTkrm6k0hWmkxr8pc8sNGU4XuB2tRg7HU88uuvZrisYaM5cJiBEawxLfP/JdC9frtke84HO9IXovgMUnzYq+zMsIz1WX3RcYO4Pw0F6b1yC9fR40FYGng607mmUGyvXTIWp9ot9GcVPrfj86otmkZ70cNW05QWTi/lQNNbzMjC75bcnCD5RPc+kKr5+7+sN5gv2JLrpsIqMy8kUSvKGeTlla0wApkT7w/koCxiBizzmon8Kx1DqjuIwkthdnqpW0eU77ekcBRA8OPwFVQB338JaE+/Da53Jk8/PLuMN9Mu8eFtLy018/JGgRKhxwIYrF8H5U9deGM8iInCigtgrN9DcQNd7P3EME52ZTyOrTf9A2bsUoXPKd1XbNtgexeFoTAaMfyx2kqJoCXeQgt1yeu5i1s4cq1IGoxLdhyhAaZgQW65s2ax2GJ25ZVtqPZkUZzVgFDBWrHZ9EqeDajXobsK8zRky+qf/yugG1p+yksHa0RZuSjNWexnwQSxGSGTSe4DH6phq+OVG1yHNvYUuIjzKK06snWfoGKt7PsU+cLWfYO3z2yebxhOod1r0jFOagwny1rLD3cUZMxCoT2wPWjYvKCcSwFG9gipMbg+44Cjlh3og85T6/3MxJVEMRCcj0O5BjGN2cMm6VL0s650l/QdtFljXN1Stz/GtTEeNn2lveEtjZhppMwrYLCehnX6OcygMeSSoDbyTE2xwcB3yCAeUO+BVeBTZUHs1tFVS3dv8j9+aKFPNwz0M8qmAQ0deULj6TR2uccmItrp4cHb4BD1n25iELP6tijBH+A+h+qbhd0WtCBcgfO34EBFqpy2cCouO4gJFI5ScmB6BEkrSefh+xNYcPvIwCmpzfLvy/VsWL2OVpWl7HyWuLBKPptfe3Z1PLTlSXor4Aotjk/A/FjH0+NGdSRGRbWcIlsZgdHJxbjWt3gqZl7b3CRFypst1XrwH+wt9mU3x3vZqAyA5JS7IwMDrpLwnkhkiBhKQ7zGQry7EGnekvJkjfSBJuy5fb0Vo9ZKzqfeYFEqjdm/6ks3oS+KBS0WWfNWBpPGgzjRHeTHq5d7IUbvfd3pecQofvil1ZrRjCtW4uqnIYvRjdfBVLsNoPHV5dgAa0AGf+YvZm+ITFWbAfm6DZpea3voa2mCsWCNx2VLV4uuA+pZLIFSfQMZjFLPdvuuvtbT8BA5X6lqPki0vLxrq2qY7gDOxIAY5jWBzbW5IJW3MOLExPJeZhXAIh44XcIKOicH5ZxCzQedlD9MMkVJR/EeE53DnvjetvKZO/Ny74+lX+sB/AfE5USte/VRO2dV4IdRU0UEtLgAWbU8/Np1DaxVolUo1kx9XzfcbE8VSGOgRy4g+KWsw/Fnx6uhPv3aJ3xY4OTMb65BZLsG4HhvBpEee7MapHW1KFGRLjFkWhN8cIFLTjAi25WLG6rK2+xfzyW/irgLTGAHmb4/NeVGPE686lqaE/4wtHTwlsl+7VEhkj0oALriVYFiNuP9CGj2WuZn0ZoPj3tvC3NtrUcJVZCjBzgw46IbOIMtSIBosvTRMijdQl+fcbfHOCuo6yOwlSQtPqSsteZ0rN9l2uVr0DtRhB5kLrUdbwpdtzhLNKkyAxFS/+MQufI+6ZsqrOAjNsLo6/EFUEulAh0cMoei+lLFWY5KcWfBSZPyase5yjpWPdL79E7ocuClHcPt7n3R5N4xw3vhV9DD3Denymc+bk7HNcKpfjunGYyjFbLhut+mesJeU5ksFfDUI26OvASQFKpYS3XIBkaSPSSzDG4EWXk3/mS0ECrxsfOjbs7BszGtwz2wkYlK+El3oqMAyqA7YeP6djwjUFItr2unokLxwGXx0i7EjTxxyTPLCCeeIYs3jhtcbPocB+FCJUgcXdb4uVxOZPHY4+ZXeD3hGibCFzglyyWsa7uj+8OIpUygrbVn61hmu634Q65BGaL2Fn83b7IqKDmbOhTVJxcqtmDomR+5MsuYYu/EQvhbre6qYZIQQvg+1hbH0STGmIlhXN7BRYATtbIaBb1z89zgFlcQGgaA19cmFQnAqAwhYb5OPZsp5Mv00ifSgYxUDedYft722m41H+pp7t4tpcaB1RXAtUoDaZ8y5R1BtWvOyJzE4mDP2+XJXT4Bea259511vhfqFwNJUBQD693p1Xnjp8ixCm0SDeiOFfgTFY5WCCzHPSkgqizN9IeEGHDCD2gCQSrAYUKhz/6U2vLvlX0pvEXBrnnBSLzosuCA9md8LQMu6rcSXjFNggBdzMdXDWv1jO13Vle/lsI38txdEgm2u/86JB/Qg/mJgmaEsXc0rAgnD4tUL0tv3afvLTQdhRc5ypKguQQXzDqxhFchkj3VzLCody9l50BpnT0A6dolaKawEpdtHsC9UmfTLby3Ifm+Bh6c6pcbLqGSDoxCV3r9xxshaVQ8Chaqt7xQXqUpOB2rXln/ipztYNsg16VGJ3ZTIbIZdUeyI9ZLWrse6IWYnyM69c9NEZSEZhOWJVKoA34QdlXzQ70cTH9S/W+lmO5RlaQU8G6VOIV5zlML0nBtOnqTRVFWoXRzkePPQFk6AtSxfA6xivCC9J/2thiEAmCPS7tYPX3oFR00EQ1OCORTf1Q5N4pAFYfrHRwj1A7UU+w0hrtQV2lLBuKtjxWezDqMpEfOHXSuZFRHuJCba+QLCEr3YX18WQfhnLrPK63Ltll24qTREefd+R+DToYMON+9qwJUkocv/Z6p55Z9FdkHxcZoF07btZhObmb3aV0mIV61lNBioROQxB2SuzWx5WJ8yP/LLKRSO5/QvZavRo6tLv/VegV5cZZdzEntf3/ZOST7L7Egevsd0YT++F1n7v1kW1cDqKpAP/13uHV9CV0xXOpzvJRC1oQ2EHV9RR8S6VZ6XmOJ4YrK9nfQXe/eRfKKztYJYlfaZf3SppbVulRscGoJq63183GV5/uC5tt5hgAXCi03w6W8OmbeHwLadkZzliqx6rPIoqIfecleEId5X/O+LbKooPdG7DSt5YGd0p1k/mM5obzR628c6eCRRdFJlXIUTUz83qMmydlQ1VWGVXcCTILQSy7lTcAi5Xezak/T1+3bpjv9y8Kwb1lMhmuCzwkxX0FxYjUsMb6bJEOFfT0aehGNs9+JgQCNoY3TtG+tZ/2wjNbgkN0XtV99LE1R5cOk1w0PvOSkOuP6jibarPVoE9GXg+hdb62k4Fy976B44mYdzvYW+0PKuRhpMAMd66/2G4dFBJbsfPojlMMC4Q6Ha6JkQS8pV42XymO/I2zreaG3zbooMGZWpGTR2Uqmd/+IUAq2WPeKRyur7qabutvWgEtL05/1vdiSuQ9KxWmXYyaC/KSdnub8uQwcUM9f1G5Tk2aMvSKOs1NIhAO/ZhwV4L+tfzg6MFY8XQo8FlaZgnrYvzA9CZhALKBFW654Mi6U4Q/U3h1migXHlcpLJtjgIwjX9z9a3LUphJmCL6nOIBdoTxNI2GuBXQABA9BsUkeyYdF3ssLF5KiTsb+Fq18KGIfiMd20bux9rBllBPd3GzURjCnUnEWpjTEYhVgIv3M5E6yoXgRloMTELsADgLqcS5MeUtHSCOmRGIAojCiG4SVMrQPaGPbSz7M0kf5TPmrNUgA3wsDPBY729T4fbH5jWX66Z90Qpebghg2MM5XcNHzTbestvta69N4BJ4llWwx1kBOmh+ICJgY0ii5aLo82iU00Q6eiC43GrReGwDxL9KeK63NqlnGK3wU1b0PQuJq7Eys+C00IkyL64mENxV4uuwVrkQZjypscu6L+fI8hAX4Wpspsmz384FYVzzgcl5EUnRkBFyeQJeJo3Cy7uL/1y6hTgPYo9gKbZ4zCv6Ni0vph0Wos5uMvNJ2SICunOUHuTuW/X5TDaNFhybOX36/BhQSxKsgtbSVACG5eTgWKt4mw0/6TiiMi86qH4u2zfaHyii9qfbI2Xuq/aPF7df1MdVJ3jT+NS2z3BUWxk5HnnizVuDL7aovcx2StyAtmjcMpeRq9133xAvnpJCl2svnVj/MEdYmzfsbK05Rb7B4TjeMnvenIBuIox6tDeaHMpt/k5fmO03wTgkd2Hz9b8NT32URwKE8E+7duWW14na3tRQ8tZmeB46vMY2NNUpib7p87m+Z9iazEN/E80nHYWwI6bxVOWA7gGguiZO24/hu/iSfuH3tsdBqfOpOyZwwb+49wh7G7jHmlYiuP7Xn+aik7GU7FP+Wbt33qej6gn0QpecjREyuvhM4nO0rGJFK0jqntBJw7HdaicIcuVBZxlUk6rMyW80BBjN/OjCVGw/vTDPSW6rEPh6+6PgQ+/fl54N/hssZzShg6ihPVGcdfNFvOk9JhdKdx2FvjzC9YOSqpeKRawOxZhQdjVn0ab20pWs/ZR8ksJnql92RJi8MBFhMR/9FaRM1hNC2c5Cqwg61z5YShFmfrJXU/MzEps0fgkms7Bhe/fbAHoVKHD029/Si/AK9HYqPegRK215TV5nn3JpYchUXSaS+z1vzB5yP0H15y/rek5MJ+NM0doNLGE/YwvlvPDEBvCSNXN3mb4hqy+TGy0jvvuXlEEzJw5wvouC9mAmTVPGCJFMS+Kf1agSH8OWWiIrP6lGqtFCCxjvIazUOuCVQEM4TFCmFGFGRwMWXsXKyp5GHUAw/HrLpNmjG8rbNK99kMjHVAPIxxweecNyiYe1mSRzc4Np2fnL91qwUVj/zg8vESdjY9Tc7ehFJ7wH0x2jaVd6KSY9NLlyqeBKOFblNM9gX+av5Gfq8nf0+FvZcIpLfQZ/Ez8qbsBsuPElAQLutvlMtg9iGVsjcLfuEAKsZMeUigAS20QXM1upzWsFLC3Lg/t94DB5wFhn6TznQrgbWURIJgwPU3TMjJyEvtF3wrGIAMgEKD/W4CvD39tjyVFia2cRL0ohgO/82u5EiKN8P4OGt6AW9Fw6ABlTJ+YcFsgBYkO95ZMiteIWfFhF9RLZj7QsPaliqIivtrV1USvxDZVBfsKSBvCuNTBH5BqM2MxkC5NQrh7Y4VvLsFVE9OloAr3nhjzmFr4D76G16pF9QPfCO7kKkWANEU5vHAa0fio7dJCcTJ+DNJrkMvfa5Z5YkQqwxWYNwj2ad7eF2q9Wgtqa+2bSokTrpB+oWFV5kLgDaRfKYiFptLPpIHpxByv5K4Qu52d3oYRaW0FxY1UDaBttApb+N8Qgf1Bpoq0iYS1UY7+nKMwTk78DXpjxiWsf8vdii8rLMtf6LAWidyTKnFpuntMwFN4Cs9YioV+9wy1jQnPqu5Mn6c9cMtut73Vo2gvtOFO9RCVp6oHOsVpkxtBHmLEk6nUnfGXOCuhr6cuFP2ZkoW/hvPxa1k1G2pgMKKSEEzyBuglyPts1qC6LO5XAkpNlRoQSzIoxp7z47v5cNQkKnf+DwOmWWUWSXSDCb6rfnbD92UAi/j08JfllL3P6MqnUQ1lnprrlDv0ZjPkuX4Tq2n4kepQjRtqIy+ppfTwAOYnnITwhNYRx0P+QO0XbUmBX5f6iqZG75L/C6jsfeY3i49XQCtYlJXaOzeWDgvzKH/Mb/hSWg3R9x0UbQACIo+vpusisurvNB4MSAzxpV8q4YEKcCjijF9rxz1inSJdJSAAcwChlsBFsuzSyHKl9FBPhjCrFolzibuZan83vA6SoVk3fSKhlKWS/7Y+ttiOW/HAbVCTtrSBOwsIbZax437Qmo4EnAVOxhVVR7xvg6kAYXOWIwPIwpqb9i17rhyJl3AWfe6L0dSKpPIir3ZNHUXrt+Vo7sFZW8hZ3FAqkf9MyNAi+7S03/JObrfv54BIcu/HG37s88t8pwOx63oPQFRQ4RW2JKm38ELQ303EZ64mhMtnYP1MhdD6jSvNLTcFqtW2Goz1dYmQzO2PJeJZKN/WKsBeXkeFkHujgIt3WHBS0zblbUOJxXqvDHL3x+D864ylzuT89/HiQpGJIrRw5Dan93QW1udgdS3JJRO411dq42FQkyqge67NMOyLKTB7wrmFiTJjHfsHxASIpmzD5sj8w36M8CTc3XYz3lTqkB2Ui2LVYZFyXX8QhKu6EwZKfT9zJSx1rtyFrWJvZPOwmFvKgj8OHyUkjWHuTfesjN5azHIrbUR0qfppoH8skQgd/HXVAFA0UUZZCiDEb6ah3JK+0BWnTyp59nvwEUxSzOMc1Q5tgH0a4JdL/vaWS/YPK+QYQ8h2fsavawz11+nrNpLPSY5HhbK0xlWTRqlZaH06nhcrhREYeFwIrLxAff4DwSp34OLTKir8vtu8IqliVzpc5rhNDlkFVkfTzoBEY0yLyBh2cE59oIb4HXuBII1G/fnp8BDd++x5YNCBKcJOgt0hLaagP6s+HHctjm856dwLVeRmXRrw3T6xRoGk3ZpjXzUmMsuJDK4q7sRbMGjJ6zxbhXx6hxyqnkZUkB/X0gIsHiBJ3qLFfEFhqBnFtBwBAGrtH0U5YcePIP7HKW2MCknqtx/jVNM6pdK5HvYWGwvuaFrgVfP+rVZRc23SlEXtV2L2WdIRhof78TqsMf2ggy41f75NXZhcpaFkvkAAKgeFTd9ihTuspMDkj8u3Qg88w/JOtKP5H1AcdFezDk7JP2RRM4X8plAzZ/coxdWPfTuwsltAqrfEqyNYJN7VlQgecE3vWOCULobfpI/lLvOK5x7enD/fhG7qmMp7vcY8aZ0ZW+1NRNQU6d1uBB6bS5qemdKOsiHz2TG5kOKD1j0Rpch8mKnTW4bUWyKww0+yim5RiHue1b10/I9tRinjI/db3H7XBncpkE7M/7OywS+QdPT7LQY23I7r0tSHfG8SyqGyjqg3HX81QOgPylDNtW7vZTjiZ/k2eMEMolJP0qi/2yLxtA7wpfIUAurvsLjScAZ9Fwngk9GehazZE4e+dMCHGeKEhzqehpLd9AO4wSnXhYRjv42bT/eluMa8sPXuAhhskin8QxUr5ImObC6nWcKOypsJroTwWxI+3mZBMr+YEqKb3P+kBVk2YSH/Jtga99llM/z52Tnq9Hw0gHMx+z9/fl9PF9iHjbtuggmgiX8YKdJDswg+FvJMTLASNql6Sa4Xg1D57QxrFl94gR2vew5vXm3nUg3arV+zQpTv9BDyAmM+0AbjgDPJVekTU7K2fKBjz9NRnBKIQKFDGOyOqszmhU1tOe/8iGZDLaTniMbC+O4/hieSlG84g7SHcKf5Z/dB9xT5xlcZ3caq/j17tvXf22dzNCcQaVv0F4z+WbMXccF4EOEGfvB+mRC53S8OC66ujt1/dPbcVoolJcRWpbCf7VmAGbakvLom9KZd8uw95XgbflnC8ZJMSpI7VSoM3TpMdY/GTO/osW8aUI6cnQyTKrwfqLJDoASbma2FZhjXKx1/N2mBw4MJI2Sto5DDd9weBpDRpdoWMNm6Ncat43OH1KdbRj9xKKWc+Sc54q+DSluyCajMaMGQlonFMqMRDxJISJ0j8Qyc6f5dgFRpEQvD/YR2H5L4o+kriUDZybw2NIIDPL26b2G6frdhXApCVnMCs/h7nzxPvoJla7PUERLfi52iQ92DqGgK6ysV/yIbJB0oSNbeG+Kp9dmW2wbCDn5i+V+3A9Xo+fRtnSBompLi0eRZY20/MoOGh/Q34cRJmjuDl+vRF19EuhY7/B8VdjdBQ4dXtHjWE1nk1RcD7b90888kfkp+Z1E7Bs+ofHJKGcy+GD+N4bZQGQUmpIpGiuocOGm3BEasV9tE0sldPXKTPwdRcoRrAfc9LmUPpYwmTgQeee9fEcnw2yFORXHrS+9CP3qF1Y6V0K61eJt2JfxNlTLNdWDbfArZ6RqJwUSruTqU7MAajy+4JDq/7EXtK90UkDguwRbMZS4u1wmbEs8wrskcY52gJ5LShZLdO7Izf7hDUuhehuMyvczAbLJMBFn1hqNw14CTVHJMMpLS+H2sWfDIGjNWyTNwg22MxqSoFg9gaICsKvfAqa4RlsA9ACmlDvShOzDqAI4BMXAgeP/hpGosjwkyDMNp0MR4WUmAvEndzwVuwLNkkijM+jjjnG5mSdNbOtnxPhb27pXLddux0DAgO7eEMzWEvx6nITRsRdqLTSkH4cqSEZpNLpGaSz8v0aG0cN0lCixTrZrigH04jO/YItuQ4ioZ29njooYJPblhmpbxUcDfpZDBOgko7Tg6kdrjzOEFpENxYt2ZOUd/tYPJXZuNaJOY82BIP34xeIu1VswCR29UKUDBBu0Y90AWjshzH+KE3CyRB1vgnCybTjQvQ3bsXyAm30CFDTYzpjHGu/g2w6d9XVnH695rKoX3ro3ecTNJ85lamacE5bNZPIJmLsUSSEzukhb+3DeF0ItMNPEU4a00/OAAz/kH2hTSIJlDFFRd6nFpwZNRnuXth7EuQL4tuS9uoLQ1YxVywTJQHhKA6kqjUzSohumJO1Pr31g6rCcVcO4pXB9C1V0rjRAo8/TdFa8/rX/yF+BF2ucis6Z/4nyNO5CXIbPDEf0g3YkdDO4UNDv/hl5FvD4XQLoymTEba3pBTbtUxC9U0g01UPCojAmcbnRu7On78QgWVFlnnT6BrFEt2hlKOSmSytvkU/G8CNzow/l7G9LG/hR+DqPJJsil1JxplnHOnXHnQEQ9Rx0I0fI4bX2onugKrAEkFlHg/asnwB3dHjaJ6GN6E3sMusebs8aGRxLf7XawgH0VWUFylvup4tNb/SKMpZC9rD8/tdN34nzVK1SztPVLuwXHIGB4NeFYLHVtriXaQfxuVfLssFcwlcujkNYl8QNrOn4Q/nFWQPmQ99NC1oBl8FOUj+gWMpqQ45JbVwD6OA9bsRJrW03O8k5ic9Q/MuItNLIjIzb9j2jdi0wdk+a78s5UwF0AQdTKoveqOrJolDSpy/i0pXvfOVttxIwmU6kG9UWgrHoLGMxKyPDPnwhMU3cVDmMLTRmHPhEE9IL12tOzQTIzyKpdiyjpyo68Apac1tN6+KD7hejA2k9aIg/4f/NiN2chySd4tHCGDd9IW5xddhzbcubct8MDzlpY0V6eowax62II/3S0Ey9dLN1HVbRrTPmEd2GIE4j8lrVNeX62jegCx5id5PspipwKRkGWKBIZOJuvNuHdK25LZPrQx2gKzHVrZKBZuiLu8pzIRboM1Z6tQ4flU8gtzuelaMKic9ZviVISRuhvi76EW/wgEqz/3qWcvh2+0bAg6WMKSphizueAeGXyoDU6NQWM1soXlKNbmLag5ujPvSPODXRpE6MJMUraMWaELB6tMSzuNrm8fc37yO8Jjkb6XisE6ljQwj5kcQYjTiXlkaPq29hRzd4Cjn4tCy5fZfhSVjQao+d8NzQDtfado+QuuH2A7vYg8fSyBNvGFssiev1OBGYTMTmbbOYJsdv2J1v9ml7UmfGM2iX2hpp8ADGRIRAbSdCGxwP3mykhkKBM8mJ6cSItFaLVS78hi8mWuQAZ7C9ZjlJ7afUCghg/A0MCeF+uLeQ5H5pUgymLIyLxH56ughWgUnbrxD9cVqRJitSxvtjtlH5nN4R2YJdZiGLbf/S8rXhI3oPZhB5QAUc2enZwYI6r9p0eJjs8ZyRxXXD+jEPWOjkCXZCJj8ZVb1bn+hfErzHnikKEknX1OVRaN3WEJt4X1FcvBvZq+RmUdRXaMGaR5l9LUDROFw1AOFB8lVOOp9CTVcmyoiiWpu1EbJ34NOPPewQMqSKYZQ0+U6WWX2qFlywWWAKSBCkPI5h3v9qretMpzr7sFOS2Ljcb3YVRRl1/uzuEEksZ2I+uemzPlUVWeVfxmZ32YULS8Y/3R9uRBPkghRDZnt3d4ZZY/sR9B2bf24XDYQeaIvAEmZI4pvhqJtzDBrAZDxfURb4Gk0b6mIonojvF1SW8PAZ0o+JHHCgxC6AupBQ3mtC6/04ZKfTpAbSLCMht5wR+jQXUSkJhybIJF9m4fv0CaTW5vBxaaepGmPdOcfOWYQlvKXBgejCG7xJPGq/bI1HqE6ln2eVlgwpb7j97gKjnASsRFnpnUMt2souNcE5Q/LycnNPUczS6r7Nbz1o99P6R3lGrdbMA7lMDS6rB3Q28NUHPfdSVw4swjlLPSMAiVxbbzSUcA8zc3csXyAxf8PTu3mlrQkkPuHfy9Z9IbmM+5PI/0S2Q9kfABz2xyT7PaU4eW8Z+c20PMd4QOB+SOIFJ9A72z2r8r4fwTJWnbbOKCbYPQfSwJW/AuP9Vtx8Q/HXoq9uTJoSbn+5KPGTbABrnhhtMAvA/A+vftyw3LTh3KWVHzRWlwgiLmvWtS3fDdSTmpjZg8jtNTPHPQzvDexmtTXzMqvoC9e5GECaTHA/O44JxZ9jVYEYacC/r4Ggkh9WfcQCUNMElO2R290iEcNJ1xCP9qTUqZIa34WBftVWgz7KDg24PCwx9jwcECFifNVE0ZfC7GY5ms4hki5EaMT5Sy1rL1Hy4WnDPgpzk1zL9eNnWIgtzAfEOrMKXfxpVKOEAwS9nSYTkB0WPSh1LNlsePICqLDs14HfuMg8nC8J7XPVuN4pgYoa8X8r+sPVbv4bKjmc9ECGKSZMTAHUljYrM31TbxXGfLbAyBTXwFTo1WNpYTlUQ1ZBDABQSL48Psn2Y8F/EMtjstCfVJiMMM7p3/JNjjXR7QcDb2J2zdmCfhxcNxZBHEnDxp4Lq3rEHKIByjHdg4V5/11ZPaZpnsg98FsJhNHqQJ2i6Oz2iuPm6CSFWoWCXk+vWal0CV639oF5O9eGYF7yWuhXV9Jv8WI19KkMs7kNGf6fW1IgsCe7WoCVPkMvqAgb0m/jo1lbCkrikpo8GAZ2VXfu4E/Y3C/54aWbGBe632H0q913Q37LolxdlyJGEO9HgXcQlqdr+/G51JIaYVsDGrmyS8UPQ1FF0BusLytkUhfjdyq9yfEjoRpLF3A5NMyTJk5R9Hq3dvxU/zVJP2GsKjf/MrdVL5AFU2bYX+/+dGPNnt3PjkXTll6teLjJNd1s6TDFcwoNHo7ErkRMisZUxqrtHuIAsoDNQV7pPpfIiqQexrTpmpp2kfjzhrdGcu84T29Atos+AA0AXWYvJTC81JpmvBCfBNgICKuuxJSWh5EETN8j+WaYTS63LmDAEtqEtcZc/1cRfR+LxjQ92mOmlozOOTAomp7Hl4SFzQuosONWKNMyemkliI6eEOx8o/MctTmjlLD8A5fcoOfzH2LYuWnc/EnSZ0z6bpxQf7xBVmisViJsQ7AaKlmfFuzdfA2kmKOKfksCh7QhG3vKTJQCIky1R1uxLmuRiAmfgBXxMWEQgnSBC8/xDzUaJfgtngXjdDoTD0rZuNlsulYIJ2vOOO0jmfrNXAemdK6UE09rgJ503V9sqJP+0MbBuDlquiJhZ32FkjuGVMxJp1LPCPlA4lzLuJfeqSpQKEY16Q8W87lPD0mPOWR9+mOH9Jfy3hkTS3XbELh7J+6PqaZISQIPo2XFXCIJ90JcOg5F5Q7Fm8F7YRzjGYlvXBaBIDU2VB34SqSURlVRovFlpYgaD3qHMTcWgFuKDXfsWk9VKFAZaEyzphYylVbhMPCl7blSumlXHL44EkYhs2ZOLyAaqSrbkWlGmIjavLEc4eB5NE6ObKAp3vVD8DLXZOpJWwhlkzPafD/hFaeEWWXfpfHO7a7mdrQwo6JEYOAbZdbxfmnk8NUYOArWCVGoveyn/tjiFTNzlmFPls1HwZHBP3zBu2OrTDlROZBimlkuxgLdPDDf3wlukhs6UqBCvOicpSDsYovv5HALzxPETA+TOw5Ns0imcckv5jSxi4gTDEKjJmYE6VK3ZPcV1qRmPJ1ux6u/vvC1oEGSHFTJ3gzEXJsSv4q8HzrhhHA56K515ZpeFCrzu/oivxc1Gru+iZ8zP/kD62TXIDHIX7aAzgjLw63fYWuw2yo03FbWUpW23q3v5wSPh3ZgGXG/YxthMxP/Qc1u/JAPvgKGDhBSuz2cbqjvKGmlrbPz5U2tzvHb4kKXE3aIkGGvcObQcTqHSPQKBJ01iGgtxV4aY4WI35iiR/ZxT7y23RL9K43sQEubEJLDq8tZe0aZBB3nIgm1GQKIMwdT1Um57uMnyw+znosdNN+sI15dpmyC7ujPhILf0/dhpnncSQwKvr1XyDkkdugp4Xx8mMI72oprovu0COTaJPYYw8JkGjCN/9im29Gz+uebyEe7z4hmes+MU2k+DW5a2Hfis9R4NNAA2gkM5luUwswgfvHGPRcILsrTyoXioxpenOfmAHIgnDWDp7SHpjN4T7B4R8mNrBWHTYOtqe6HfLG8lgxvcn4J9/++OwNFU+KD1xlp8e/9tZA9KJWhgeCEaiqZVxldiND9Fc0lA2DwyOHcVMzISogRnFH2wJDk+UqrB9JFxaY1nyiv3C6Hj3lbUFQ3TxXE2/A0Ro3YgAalS6ZdjqizUoBPiBDP0cooNKQ/qeADUNLoDWM+XVvu82jHF0iTHr4s7FHh+i7q7ODneQLWk2H1QWiHNpJzFi54znHZKkB5HH52ujaWj06TZFvPfE+hllxzaQNnAwFD6TtaEvCGlDaI28n9UxBf6WjqHMuIQW+WsKhDhxY2AGyco8cqB7hDndSSJ0SCu7d1WyKbnEx2JWcS9HlZdNUCDNgK/q3ci/I5LqmN9+XLaCPjHQ/Bxl4yINZeInvZoVqRDNe044Lfi5kkYeXKiFNhqIi8sh+BtCBnYFvWryI3ZDCVCSKJefryhvv6JQek0nYG5SJi+fRtfTneNWeRQVc1IuOcdcJvUvTyXLxfbWoYs7ogDIbZNu3BCV8tLv4/M+xyiIW5vIT1kezRkjC5dPm4YYhqPlDW5nPNf+22vIi+lkX7xFNrtri//CbOWWIPSIICwLgyMgHpSPQm5Butt9PxPR3HYBbRfOMNRz7DxiddlpQwHgU323bT7AAGkKmebUjNp6OLvjx+78MEw06gibgsXAwPB/VbabNKG+Qes2cGVVy53THXv2kMcQtzZrj23h0MQAmYqz7FIfPCyEqkvG1x33lfr3QE6U0xudMnXevHfeQTUHyj/RtJ84ph7vSOEjU3UyG7/zKLcyYSUsXycMzD/EEqTX1F8N1c392UYwIHLC/hOZnbdnFIrIPMgwdEg0NuAz4aUbNci1asQRps4mj76K0CF+AjYqX8Tmdbx88ZRD0LAxVARq7bL3AqNeyqdjNO1BX3bdLUNoeSbws8zsCmYB9L3BaztNCPuIXeEWwZdAbdZGQvFaN9h8ASpQXmgoNyUWGayabfWulAVtU35BCtsH5R1UqTtex3CULXoBhvGtGrZp/o6eUaPcvgJZe8inJUhiAQlx3l+vxmk2Y0mbw5hUqm6Zulv1WVj53lNIKYh1EMFvDIqW2CUvuu0f42BSyJZdSv5Q4diMbcGQp3BeNiGZCfd5uGBT+QGyBZATO2FRidYEU1EwTc8b3QQe6Ybmq2MJXWwqLRaL7icmJjghBGKOZ9qmnhs277jAVHwGu+Qs8It3xnAidxR6o9lJdzY64qRzSzw2JcayQMy4zvpwMq2BQPllSPfiFewWatkWy56UreUfAAUMmj1E2c6DXxIBXyZ4lQkHhO0XWa0sBkv780KvAhkLO9T5y2XjZ4fPgxXAh1OVoyTmw9OHZUoVg2ZqwOWSmZH8qDoQFvvrwYxZM2MNMmZRHHxnOGWdqTLJrHkBrKrc73rrWhlTnnA4DIiZmGRxF9lS+N2VwGTHcV71ETtfXQRUeN46zv7pVRRcfmjwZ7Z0v9W1ML2jjw2tlsmIGwHSfq1xg6F70dkjM7LBac4i1hHb5a3ddA/as8YkTD/Y/kBNzSpb5ZneP5UrAswpMRrL06g3YttQXNPLtlGZEJ8aDSyjtl6LwlSS0CbQ2OxfHe/mbAyjeLYTRG7OcXCqRQTxMdFynqHXh+R32d+/+2ZeY+VODfZnkW/OnE6Eq737Dhc93ZLKAT/O8DwaE1/ChP1+16H/bCOC3PmcjpKzfTxe7XnR+JZOCR4ENu7GIrVlHumyaWEFYEPH/+8NKzPdm8aLWEhwyxXSbPvWwsT+td8plxlZbGRCKzBf9jeYUgbD12IiYMXEMiOKv78LQQw1IXNvu4e7HS8Ii7T6qZetAR6YagqGbY1DSHDj5vndE33gNSOBPLseYzM+AZIExp7HS/eqL36/I0VmD3kyEj9k4GuRzk+5F39rlD5NA7y9+6afPOyilXgsNOePiw2nD10LD13j2VT127mIH09raxN2OIuRR+9vlvm8zTmSNec810wh8z0il1ZXpulFzMqTMuEBSaYSa9CUd9xk3uGbXSaLhItPwtkaRSNvRttt9AQCU6SBhIN6pxF+WGujTxj+shTEDAkSh3xPohT4CnZ8RlGkHv0mEU8d7B22dGoyUdd0fDlrCrex72864atrF1IYFnKAjVIF7H/t7/doFvuBrj+8ghNQguVdkQHnG3mfESrxvNYz3iK4Orc8aJsMNLxeCTexBjazPoQdzsdUGw9/R5lzLPYMYrn36LKCK4xvfHx9WdFITWh5JylCxOqEQSwwkLxPbxRz9euFMyxvN8JRwnZqlC6Gc9ltmy1Zzk6kwWKdJm4BdgEOXhv9K0f/mg5xnlWTE8J4Ous68r9iRTT7NYncZ/ZPbn2I0TfnArKcZ3diLxfY6bHKcRQl+tcAP75T2CxJmiW3LYzWxaQmiy1QZIKscryFnnU3vLqq0X9B86w+IydWPXfvXxgPeoL07G5vkbxtu0QcVG3SlLgHk0yKSMd0ZSKlwWg6kYOY5g+cZayo4S6fyXUgikhg5WUB6oLEA0fJ3kTQM4jaPo9HQ4VpBxtqKDQZET5KUh4Gv/IahV544e4+/lBbKnsRcgHr4ut/KFRFg2fiKWzqdPeGj/1Z5FAleFTSaSYcQKQd0eQhtW6VTdlaIYHCZlhB5CizkYWxq5ewDzKcyQR9CG66vUoY0VVkrYEMoFM7fEu/u8ElwLx0BA8eHjGeo1jk+U5rolXkTk6Zi6qp3TsAIiD97Pe4W84mYcsYsxt3u7PTanJM+Q3a1c75CLdVGfbC3DOPlJ7MmucN5NfFVxIWESrPPXlypVGz/E5kHCGBiQHD0bEoNkyAmo2rxYXxw+M+6z7AGCcGX0RxOYk2cCh6Pkg/Jf8DKfOHHPALSUXOGZkLnusrQ3ZYv/bLcDdC6ZIvwgXUbG0+IjIJhDGw0A3gTyAU26hxqtKICeRLN/JIEVSjMZRqUaV2KV9bQA9GDvSJTP2uINZdkpBhhG/c/C2qWSuBpkVsQWLOFSrwylYDRre/MpZbIFBwWmVnXNgDpEmKB4syIQnsci19/EkB7VbF6Hi85dfbPJFyZEdSDJyqQnZ8VAy2F3df5RCgjkYFAKEA01g85VKuIGAnf18+kJW6/LY43Zfn9DsFjw52FvjdwxSXzd3G937oX4TQk+wT8KgNwoA0b+WqFquY6gqSdX8pTzGOH1VAOSpEt/1Syz5+NJmMYl+Qf6nMpBn2atlvVPfLzTwlJElEcdaIhNDd7swipvqr4fkZMG5h4no+2m6HCX8HQ4Uc1o0gX9xynJgqXD7bKs2MwncXBG1Ehr3Kd3vUTbq1dhCxY6ofzPM7iH4nCF3XTyHaOXZdw374q8qWYkeGrVHNyPnpBX7Z8/74Jrhjt/rDs0hCC5r4ruMFw34MJvwExxaNP2z2qJ65AeaTC+njeVEu35dy3hG6dmkWICOAjMINFB0PzjLLVmrQ8ePzIFXtXQ12dGK9HMteWi+JREBfwFFQLrT8Xg/OqlBJiNKWKFiK7Bq5aecQpGVrLefUYlYGtfPdp09k4pZbbawjqqE6DMzvfjNGTdeUBmJp6/hRh3i0HAD/a73O4WJ7Sbn1t9hFah2s6Qwe5G2cSqnvmeYiMD01s9h4NYs5Jt8yhhHkNZorzYEshYhvLJTK4+DQwYouvcY/hzT2fWROkqOqhPTMEyG6cg0AyLdxgZAX4BeEMVnHaW/PIKiBpZi6IKcUt4Xj7I62RgEC2VhEUwHhorzixDllvwaXDGCMME6JL1MttER0SOmNKToBtzl3OAriNYcPS1fsVEoptsArBLikyMy5fsZT8nJmH/yVLDeHiDKIwlBHw3ONSwE0v+TdFWuxLkrfeLoVuoMcN/v2yakrX8NyST67J0VrYPZqebszozZPjke/yMcqtl1KK+O42DaF8GHVa//txckQKX8YsJoxW9b2LdKKuyY28p177NILh1sSYd+/cwkXZak04vk08Q2SBvatbuaUs4iEcUCVVjLWeP+UElJ1++dZi08JO8HoVYbSyQXlgy+VsX0TvU9YPT4O6MGDz05CYftxUNKw0lMRgAptnxZ28jvHPG/iXV69OUsZJPj4dSOjt99mQIsLeqhkv9nPBTrGfibhwWbFg84c2fVQ7ylW2VLFmwr6rKNV/soP3fkClN4tZy8L8QIafNwIt8aRNqkGoWKgtl2+ArPvWbZqHiOL8R/L7sJnrO8bL4CLIVQzLFZsrWmn1Exm1c9HbKYNbfgRsH9vCLONOg5H8XT9xisU8Fp9iZM0P/l8uO4lWlAen5P73BhzaM+9V4c=
`pragma protect end_data_block
`pragma protect digest_block
9d7970f115e9dc61743b8a3254285e23b7e253bebdd2336da34687211f21baf4
`pragma protect end_digest_block
`pragma protect end_protected
