`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
rHaoDYPAacWKAw6feolqQP1GJjbX+/IkCs+5YfE9bjxMlUDD2i7LCHp6g6IDKxS7SW2fYamuqNR1PXNBMnCcsmc1hNFQ1p4Go2g6w8Mj7ThC1buTG850uM3PeUIY5w9VcwDUQYx16F/BlOMjqgYaEk5H8GgW09mL0lh8MS+rdUqpvcGDmCdoM012SClzfIV/6ssDarrGYfsNahEhxD5k/BjfKEvMMxtBvtj71weOGWUCvsmWrFuS/BHGkDi8szG0HLY5ODiNghhgzO6rXSfz1wW+7Ypkdvg3ykcTJ4fwo/54DnG8VzyHtuuuHVlQIa/IqV9M3jJnRadD22AADfZ7MISaAzGr4BQAcXcP15csuc7I+nlkwb86ASJrQy9d57r1ePwa3PxYbGmIE3U5YbMMH9mW1gijPnttbak7aueQB93MNZaxbJ6Nqc6nwN0sLcPzUI1sBh1RdWUbWG7shD9g49FAsB/zCnXzCzzz7+SYUSfxXrcGq+6q3fyuok1LQwzFEcTPCjtKg5BuASDgOXFRp7q16c5WuLIrgHf1nUBOUvRyCICxIn+Xr4CYTa6IEOmcILjGmyq6TvO6pHE6junnWhwZUIyeg3/5qGljNIH0+rsEetKNMQdsG6d5WkOtnEZZinNnbQ+9KT09aqumwI7nOEzYQX+zoobf4vxYDqyx7jjL6dx7DJbpQfzflPZMD7c6yMC6TYUFWYkNvwkABVnX5Z2RphIOzBTm7FIba4XefFylIym5W4R4uKl9ZtOLUttbjRKDSw/deKXksRUjf7k3ICxWqPzS4saGyVKlbdmIlQVx3wSxTHZVxWK0aiK22hGxNgP/rJIs/PJ3X9L2cm6y6Act45QbELWYMqss8vTSymXD2kYuqcxse14ac+Q1CRamB03NYBWOgcQi7IflQkkazK6lXPfu2XaUMPhlUU+DXFYod9h4n/CBnSbe+1/TcwUZJuoAmu4U+FlYaA8OYW+rqJAdezmJasIahxVQXdpIf9rTc3NrHhgyRBQBPuSDNpCtEbXgNGmoFtQc8Udpc+B2CXzJT+I7vWYFslEGiVifmyBTpZf/GY6fJkv0GR8A+hICAVKlV3y36vwV0WKQYIVf0M/UTCW2a+Un0d0QY8bomRyjkz1RJ7lV2T5oo+4KSZWPgsmARQMpMGKQ9vZwIUrFp8pZi4/pKG98XsZoIkSThEHv4JM/GyP2KlCu3zAchCnLfbgnmDKarbp/G0c3071sWO+WV9A/uVpn3ocXoyTfeycy01ioR0kBm1usgIk/kn00kkhiTL9trYkDI1/KQM6KbLj7Xbq5LWCjK8aHmZipEEuiU1aC4+jyFU92wC8gLgGVMlPhsgWUncXsNQxOgd4ny65A5WGZdgB1HrkI9VUgZPJfJ9Ts6uqCvyBfwSP3zuAbQDkz8t8wBtg90/JvZ/ZarrkpHxQcly5sabN4Vzv/ruPzXj/5FYEdQ8S74CGXQIbLboGVhqyjJ75xtEWxS+S6H98L6hsayz6HxIxY3cMto4E+UKoDTFrUnoxAQ8e3dFZt0ShN8OWq561eH6XOYdW401idJxHbHKLW7N0Nw6GepoqxfmlghgozGClghP0SdZA6ydTX2MZlAKybjTvAEZn6TXLck4u1gncfRFPSaxKTJSAlREk+VOkKqX7yUFA7+1F3VqDdDpWv9kNP8/J1mhTfRLX/ffNnCgTfFs9Bw7hqrU2kuJ5JTg2WTp9ZNjGtsEZ6OCcgWR7J00ORQab6O0cXgJUGLhspxpzBhG7uC1lcOsuL8a/LN++tyVi+cNF+aLr4rNhpG2v909J09UxSwx/b7GHi2MD8VYayAlq8RgznpCzGrIGEHICWWGyFz2H3OHluSULqasfxtOnvIv4V+7lL2jUB9vqS+kC+PvqHw9CkWL7fGET6YBFWYi8ZFFyBvKZ3MHCLQ34JhiMzwJyeQkuvbSyazozDP70qHDCBTzCDMUdyL1CF4ziZcmh6LgW2GxNG+ec/F+d8JkBEp7XGY0ELH5rpxGZ1/++E+2RwStppE7SkmCaLQzxUrTYzxM/+BhGnMcMmElNYX1la1tTznFMGqXImVghU56k8l5R812JpiWwjwyXJaCnT9LW3G48esSeg8c4CuxFb6vM/m8jUPsFFKJ6A2K8TY0R1Mp1JQfZtHcSt4IsAuCi0doWPhRfXCnaKwZBDqivxVHmCVAKOpv1EVD46sPYvj6H9nYnt09abIPgYLERcjShULE3SbZ04iDe4M5JeztRBW25j0Knxm2UirhXDvZGk6YryoiN+beLJYczoSH5Qa/pDWowe0p0sTRht1bDpkYzRdlqmAkBsmPvFi0v2id+42f5rnJ2JTJbqLWluNZjD2xVcODqBDxHarmKdWdDQ+/FRCKTBbVlTIpHRoAtzhBmNVUIlgx2VEXwDcBGIeRBZ/zz/tx/+7QmUGU/jshni5VfZkR/pm3/+bjv/DfzGwmXE6DQp8FPlSP3LlJRSAF17b2cvqUF8fRMffitc1+q25HYNOij3LuQrwm8nicQsJLy4FeQngFf6okz/YGa4F8lkyRpXhnQ3sfuvxpxHYuO7Aec6v7LGBZnwldz3l/2VXtkHBCic41qPCF94Yu+hR4AjnsNU1LyXrYgBxWR0bJ87y9KW4VjZ6a7AxKga7LJUiBcSPFY8M2Dd8ihlELKk9oYXEe5PkzcHmdckHEjMBtL89xEBOLsaIRbmeEYzI5loh2iLG6V98PSAPOWk6LmPPKxZVP2/dJA19OiClfkkEVVEGygbO3VF1+A/IP9UuA/fqknuy9Yh9xIBHxwr/4nLdv05iUtjasg0L24sIWEG4TzwIQtNFomWcTvoc647l1W52tl+2aGh6ZPWLMDL8zslW5K0+6V6WnQHW45OY9zWdmbEFxXRzrh0mMKFchDKRJbDyi/23UaQ8UDrxFr+MQrWbrKgT/CQylMK8KuqVTEdYXK5lxh/BBgPbsIlkJJ3kgOnspYu0PhrsSRg4T/2My9+1X8d/a5GfDIeKi7XMw5c9/lsrIuiVq60VcLWtbtU9I3IaRBNQ3w+gF94DqQJxl+dem0Vsr+6To28QO9d073Zw+ztM2HoctL2Au1bOQjA3WGzeSu0jBUAAoQPRQnnfR7QgZfgacEAyD4mHVB6mS2iEAfLg8lkNqlHrTjJsFswQevSykg7LBcD6klmwNr46oSohZ5dnrmDB9au9I1I3n6pPITdcxtKE7rWPhWbqhFumJDbzW7yWX4a6UVdhcgQoUE3msdzc8X3J+ewCizlIwBQob5sj0RejWoXr3252EpfUDZANB4OJnT3N/Fr9Wk5WCmSbsa3/jWxpDfCGCX/9snT/0pIIR4q0GXz5dtpklApq8LBcC5MZcZdwsWvNwB570TTKBYA60m/wNV+LiQuuwc93kbOYJWmHo8A3pJsvdCzBqLaH0/ISjyB3MExUi5cALYmgQCZj5wYzKyX+nBphFl8oxS9sRCM5OCvAbbZz6mn8xZwXrZzA//8HBJP+Xe0ac4yzEEB/Elv3L4N6Ro6G27WlTvan3pZiBs0ArveF6RTvq1F3rUQ/ecNpPDqIXyPIZdLwr7RTGjcnh2lc0hbHB73WYwB5Fx6eXwJ7UYGbMOITg6zuMBMJYHrimRR2XywqFabLOt16vCbQPuDEnMjHX9ViNMInvYkeLDEVsv8MRWlj8dqA7rnd0Ij4Q/LSLkTu+kgeQUxY11WyYnEVLs6av+tpTqNaGWiSJdAfvY6vQUytOR+mp4mySH/jhhqMcdJAdt8zI7gllhwilm9Uy0Os50ApqMRxvuVfe7GflEiwfSP++qOZVXA+maHcBTRRz5SiuDVgvwVXkIOgZ6/oDOwGBjoT2R9nG0eQusv0DyLPJUWDi6HIaErt75UKh+C5XSL+AHfuL7CH/kht/BjSEHvJxgWvnXGlgGDHLGAtTB/lRr0j7uz2SV781npJqv29aISGseD7sTb5VS8W6j3UFAYzF2uCDoYc6xlsAcbAxGO3vFL032t2oyyqcaBDhNFrCeGWAH7zFg9bQT6MEah97nzObSHp3IgrlmYHViQni8D936UDHfjxcJG89+qUPgL1mg88ux/mpEvPfi8PRS3QG3wImBuPJ6dwKumPwHgZKKhMFuOR+j8OQnJLUH4JdxPgel27FqlE17lsMKyCM+GDwKbWGEqROWv2pCsHrJL2aXmZXIV0m6ad3rvWsmHiLkfBeyx8Mvxp2OH4qCuU8Y5+gSVuQci0xPiJz0VRf1vC6EKZv4X3ucMSQJWDs2z5JkBRUuUyrAOpItJpX9HPV4aexZztCLI2E4NBavFpLpa1zUA95D6Xj1N7wvalEa1iq4MZRWPdUasVnCpJfIv3nIRf0j+Izl0qowJEJT+xF2WrRuiqFaGiG3O9ZAiglIfx5OuoT8ukfF9ABN7uixreBFdLEhnYzrZLhUaUgfmHFCWgQwjAdEkGg2mt79F0s4b3pCgP5CLjC9HqyVRwIpjhmC4fqipGkm1R7YMz3ToBfaCMoPRag4xWNmCbPjnBqI7Dlp+pxpKkaIVvqnynCy3ii+DQy9RRTaHOjVV608SNsiHbuYL8q1YgdObEi4fugoUCQMdYHaC3deUjWC0eBZn1kFCIdvWkT26KvyrsyH7lHK3Cr+a4Q+Wu5KDNCKEtyFVQRZJGo3cBEDxNLarWcFLdwO/+0vdQV5nfdV7FhzkGgLRJDyqSD1rdEl6K+YmCOOROJwojLGh+IoWIDvd2i+LJHGbjgf1yrx2PMf/64yHDtXYmesZsEU55Yrvy2xxQ9J3UXXQ3JFYYDCpX5Ut3yi1bUK9wn4Gt8PoTfsqDf1q3RzJKDtFgkH6KysHQsq/mFO+Q4cZpEoQo9fZv6uEtK3xlvoxNLZxVdTD5SpLPFGZl9LLsUfhXukiMfRuFzK6gl8lwyDr4KDncL875IXPlP7gJMH//6QVOO3PuAEFxPrTgVGdQ2NL3sSCuSzCibxVJBLR1nuXDA2i08+w2RjkCgA5/+63U93GqUJBSVxGZ+B8nV1nD1bdjrbEACiM976seus0Be4RCJF0h88AjAwOjUookCZjJ2KSoHnlu5vAc8nyzxARgnWe48EG69+LzXlTL9/LvASXA9tMG9dapvns5wlFpFcsPhHW+Ejk8PjJITPOFnp0Bk/kxxj4qcoVyLG8hzh4TJlqy7ASKXPeYxXlKkWkc5pBjPTVNIaY3mvJahLtygjOuBGMtx+6hATxfd1SCCI4xHYXkmx0qz0w97eUO0Ys9fqH/34V7XZoa1OoF3N8fqobvdXyc0P0PuJF6t8kL4bw9zyqDeZfOh2r8tx/kEFNhRbqCWcl7JgndK+TY69e3bNjgjELBoTzDj163nWTjG7Goo1lRF7S16n7jcM2Z9EXyGWVk9uNrh7YRlSZDbZRr/8LaIzxcYwmKxaT/kZ4VsgK3uNSQRtWDBZ/SUnoKIeALsMr2u0Irnd2n5UNAUqgSE2k/jLcL4aYUIV4L3fh2u4bTP3vdzkPRvmvaL78z9XHMvP2yQnLq4wG1URuN5wWtyRejTpVZsZ4Vg3cGHyhwqUWGW+pbqAeW8sMne8DqlRFCKAGGEkSRlzh9zTxk8jbPoR0w7WuIeWkYJbpdvpKDtGYKwVbAfR9mVcpn3D5Ai+7a6JHcyM+lPzXTJIfklyeYi2MqfpBErERTRJ992ZgqSVmeIxiFEZfNDhHWW2xg5/h/NP3UZC6trhdWaNm4reaIqQgbRLFXMTwNu2KTWwJF5nQmpMb8H8bpuo55qTFmCwosCQQC2bu5V2HbzUqWccZ4GdU9xKtgAvGqUQZMy254O8xzPUtbbl9IEdSofgd0wcMfTwfzINq6zAyXH754+KQkiSTDwTyBnezTz7HzOXO3es0Ywm8ylHOsMKbJZQyEhKK4SudnzJEVWt7+RVpslwzqo8tlHrk3aiuZTkGjjLJmKumXQHtNP669ksCwDIv16WSQiU0Z3qOfm9SRrA4JBrPevq/kjj9JB0hfi5AOjqqPB2+wJSU6obNuJnDYkXZaH/hD2BAgQSUOKc+y9YaIbD8DVS6IQ3cC9jNEpeMAz7OEm/no5n1FIbsTqrcwWpSG4gzIVe2KEuL3JaKAWmybKkhXRcCh8y5vk7vDABdhhAO7znO7V+B4+zgUl5zZ+DGEv7NTvIhwally5zgAFC25xx5Nxz8p8JRd7PJbPJMUNDs+AqpPFb/GTE22aUcpD9tQOoUdNgtnvy88MnB6PQnVZIJikrwG4QvW8aXflhBz07BAdzXNJHsYXTKjXn7u0GRlWK3FRkijJ5S89y3zVGiTDqKWd03cL3FGgVreKxMHWTUp3t7lds8ADDFjhzh+U+z9h8ZdWs1Z3J8jE9oakwunbSiSzSYjzCj2WIFrjaBJImDQweIpmTZAref3EaLAR77pe8ec2BrOMV4UASnaJdZ/cmG+BYOSJBFy0GiYuyOdHgEJ00PWgx9gK28cWas/TQdMdU+WXPFidJ161moFXK+nIDzXqbwnsq0Bt6D9TP73z4Dh5HzZ5V96rS3QtqV02ZyCRTUW+LFR2m1GJoSeRcgNmnvebE7iI94jHpGZO7befVnIgtmooGxNnu0MMRhyRnlxAHegI4ElRy6+Rdvsom1uFFdfB0KiMGPMmcR64/V/pAmWW3ljNcdk4AkblR5UIakx88A0fVka+5a0/2z9pHeEkcCFOxnW22QLMyK3VwOxGBaDwUjwJHi1NqljDmEgK4AS9PknW5gVeCwhpk2ryR1jx7KAp09ATnqQlDzOorU68l4ZwOdVQJf7d8noauEXFkdMJx33LBufGoxRFEcDU0zjJImtFrkb1C+rK9Z+4UnaWzwLWL2ldNfI5Lr6KK4YzNxIZfJ+c9UCLRbJNJNJA/g/fUFQ3oWtMhdxxDhd8XoGkiszDtfwkL/YA59SnJhQdCTJJ/tTBE4kve2GFHmo1svS3cFDp6/2mVi+KwCC5emiaE08IENgyeA7dIjy79JXqqS3cv1lij9FEWewEQNPCi5SoHisS9O6fj0Ekss/JdYXy3GCu3pPPoQPPl3YUgkJW3d2vLrAoqNomyxmf3oPNh20rttRljzfEiKT4KclbsWlgkb+Hfj4+YIsZD83Dyrf4skI38TfsQrGwhOFyrZOmOfPRPhhZ/EXnNaTMsU/qIzQ0RNoJvGN8/Hdl+LwhgW6oEHPo7EfzRrxTbsQknte69vqWMe6ki0FZ6kJUzzudDxfrRSr4/tt+/41cUpZ8kJfTjGxUVCDfO8ktRk9h3Te6Tv1y4FFjkp+TC4FwDEkNaAb/M+trlsJcmRB0n9TVGeMCUfW/Cu8D60CWVHFg+WwZzHKEW4TD5KTBtIvgvmsWNPZbVguMbQetM/8D9zndWI/tcMCsCJenGC1fgxX+KI4+5y+FAkaGbVZo9BxGfk7Arnk2hBySVFp6FOE37W0UWmK7YsroQnjpoqjiSJko9lO4SOb5fyPulmJ/543nnBM6sUsUcjD7ramshOjuwwevrSwCIXOGcN5fUL6a8UySea49TjQezAbOXx81V/T9QZ3c2F4Qqedlott18yIu26KAIISpUVBZNL2F7esQcrpadHXAmIkwuwXzZLNZ0gEk2ab1m/BYzJlABTJn62/+GPz/i+IVhQnWkxevAVztGMXZIo5vpO5q0ksrpYO7MovJDRDXQu8+xqho22BwuIO86S3v+c8BTdMhr9zFK3hyV1qD5mplDGv1uUDAWX5mthfIUrAoHGKw02XkTVoZdLSjm53RZfeevmDE6dG+GbYdfn539L/e4uXRYcRNJU72Weu0UjnKElV7VvM9g3MCWPQys9P5JtRLoOzMAjeLNKxE6D2p9YFbg1LWyQ6GNTVa9vIFKFE7sJcyT3O+I8NHMzmDxMce7jmNl5Ab0y3O4fW+r2rjpxXxUp6uy0Kgg4cqVYLQoF0XqLR+HCpzNr9Qxz1o5rfsgbFoyt407b552eYzmKHKcI6XyJdjSmcxUxQQ+Y0KEJhYFUmU4EGjiAUmRA7pUKdllv9n7Z0FsTwEdd9QU2/oGTc0y1LoX1W81njQQdFluR3yiIVLQDUstv8GFojPRVNXzTAlbmzdhYW5Tgr9d1dL7pINQCFFqVBhCbS2/xJxPKhX4TNKgB/YzIS44xxHGAHXD9viVOLc56lZmDhDJ5Bm+5ye3gdEaNuc/3bRmJF79fWpCf/9jiXRJ+zF4R1nVgMJYXDScS61DkJVxrqAlAaUsWh+rNeZLzJabR/jcUo7lrQqqU3DrF023/3tTau7FuxY2ZwN++/k6dhQER0pUIdZ7037AHJnIlwWM8ZGKNMshliahCOUJkoBrvpvKAD4Y0Z0ZN6HG4HLtYpnD/Q2nY4ASIL2Zy3G65HSviIxNPHBGhco69F5gDvg3AwHBG/v1qxKUgYFuTBFSvvE1nkASttMRYV56tQav0s7YfP4WbiT/iyrqEDUi2q197PLMWmfxICFNgtwtSvMk5G0wCJswsaxp4aOKgDoVrSKjk5U32TPdWjmijNzoBQqxrdLctoGkQyxNzs2DWv3od6TQPo/2FRHgYkCK2zJl7JueRCLwo+WVAYlMm4Yf1kjPWlYCH5uWd9txmCV9HcmRxm5KLExQ7x1EwsufoxgQxEbB9o0ri8LVwi5cEvcCrMnuHHCRsefvBmEob7/E486BGK1NPKM3oFugb5Y9rBju8s+TvO9OEF+7hPOB1ILblDducGBhNK9iDmWG+FntzezImERvbcx72idiDdBEfWrH+Zbuq2Bt9NZPbCNx+GpwXA4Rf7s7e+KCwdw0so+2SE7LZKPPNgDbcqvJoID7es8HwBVIt5YvnO8uVyeasPQKeRXvr82QnKfWUBLE+qAm/hNnuAQhTBBD9lwOswoZZH5uXzklS8yXbtyCGxBcHrtybs1eapiPAVvYW3OCNfueHkIMnWfsmvikknsN624NI7ZZ0B8bEtLkPT+Pvf90wy2Acz1P4T0LjLEdfmWPbjo0Kz1ySca217LSWfhI2GG2A4CnDkA9O6hQ4m5XS0XFQLCLUhCEZKG8PLVOMZXFVyV+MTsqO79zvLgkUQhssYKWi5vUf+3O8VJ82UJCnkv9F6GUF5xU64WjULGEgJCcOAHfJNBD08otGL8k3N4F3F0dX5ICS5wyYb+zW1mtnqCL3duZOcjEf9KRiIHNxZYcAEDI/R4vBB5Kg8kti4oxjRBqPgFtlVvpnSE9VsRYeoz23NlGdxm3NNFDN8s+EO4ywBzU09HfAynyM839ah0tAblbRGu4K7mew9C1Fl5rNBUp5ykbCPs8OXgs5fzDDKRvFejxAzcSklNllZko7oW+4sjJhQ8QX3Ks0gOoVHYnIRlvJkGH4I3oOb0s30yPHlhCPMoLIQLcNqBusy8ovNrR3nJxfvUrti6yKijsMnXKYdkiQs0Ob/4+xBIvd0JtrQZjIoyF3XHYMfbRKeUKdJCBVQcMMVk4rpkIkgYwWpo5IeCsNqdF4IthuOIiXmqanj2L/uRDSopMf2YB3AqhwmyJFq+kjlAD+k1Zs0/awWEGlAHFh57PltjleETtJiZu9F8SKXczrX9Xj2ghkfjBTmE9cOPqBUt2zGvN6jGSh8O0T6NbMB3Z8NqgbZJSMv3jrCFxYPxfQ2E2SxNEr2FZd83LxbuZIXbwa7VRwb0d+XAyEAroWMpuXPh5JvKe5C9zfdH3DtLnjBOqhPosESYo2dNigYASDE6oUQlwnbxCk5dSBe9laXHoFr7H/gQMYjp39PRIxjJG1oCQag+ionIejZVIUx+IJROWOoPnAqJxNMAe6zhFbmJhP9k1f3ospbe2nGADRGBPGCvKUMdA3Vh8jtBT5dxeREq9mgZssm0ZHOUWE5Q5mdTl6cTZE45rTmX+X1wDA3vjBZuy1iHhragSzG1ILDZb4qFacP7xlIvhTcSbZDenZrOr1xpv2LEvMCck9M+F8MZAhfRhrMenLEkjYTIZnXLyZy1o9FyUBQG0nQcmbRJgNP4Rg24ePVdcluo9Uf284MDASSMaoYG/e38W7kWhEC4e4T3tDOO3C5uxUQMH1ZfvArHkUFTfkDl2nY2cRKxKQExlw4pT2bAOGM8IvPuYVLNo1kN/IzbosJhqSNme+EDD5BMwivwUXIr92FleoVlD453vwHlOgTwCyo75D9qy3ASSVTyjqVwlNUb+BnqSHW4k4QZR1rmve/BYiPPr5QCs6gOFOcCjshcstS5eRmcBZruvvTFkXBNTPeQvyn/os9XdXW60Eo/0wYPQTSikxqeStlD0bwDE1zpAFemhhU1pgugR/BkCzE5Kqg6Topbjqvb7DhYGiPHLTI4qYKaPkMXBSS1Hi3BV04Ilv2omXX++fvsZj5SmJD88uscf39M/H9BQKLBgjemuy80E4eFq7AjCQ466VdSvv+9gloLmy4FJ78Mvt5JFpFDMULkTHU7avqVDDXGpujELhmbZsO18RfDUEIgunqpHjldVp44eXfiwPzsDyUvQo2eRFM0Db+T7ukKXydjoL0CdNBRUGIU3gxQb8yh3DDssD03Fm2qJuUiZ46AoEM9QTssOyixagf9EcbVOnS+IWlqsKfU05JRkw6b1mTS2/8P9ydCrXyrEyX/oAk6/JV3f1CyeXLU2HTPQ0WPBs/CUoCrZOpKAOPh36qDJf8bBArxHNmHc3OSOl+9oT/XI3ZMEjoKBNVLvYmgzJkTBgetq6HjAQA4atVPze4JGKOGVcmBysH5aUwsNxX4DwA4P+ScKLC2G3g7efGiLPoVee+qhWVFgcHUK0dZIgjWxt7h8wBzmGTJT8sIi2yEP4G+XohpltVADbTswo/cHZuSWQQbm9W3QqTDh2y7w+IAVuhAMf1j0xc1gPlEuJ1QuTk0nOq5C9f67xCTi9nbAEQwMW7Sv+5kf16waefkfKr/VbA7wmJ7ZYK9fGZda3ymaiT4TunZ1+hAY0Kq2vYu0birC0qB1vmV/wEQPZzCMKsY6SG1Q2CzgSPXq2jDeSpAOIw0kZRTDuRQ8z9YjOVpe3OS/u5wT2Ra8OrfCAeSY//T6dqXWVrR9REqTRaFcUJFisk0nWCPXl72o20Rj5NEe+10hi7RDi9Z9djPg3Mi8l1tvg5Y7wxOsIMOiR82WOV+zYvl5zW9ij1NR2IIsBu7Sbc9okN4qFAJ0MmptDBUx2BoUy0VMkDbzLC8eiYZ02bFr8YBPe/EsxiOdT8h0HusTdraVb63k5mGRmr0Bo/OwChDs5R5psLer/wxsUn4jbVMPvtPD3ZADIs0oBTE5G6AY4R8hNIFHg8S23dTR/R/lRDWavXtqQhr6rweimKPhTK1g1bYF5PdqTcTmsHJHz8fHnjYZLz+tRLCy+D4KG+aKUyKFaVtqGbY/SLz06ETrgBFQ21PSaAfiVkZaGeSxdatN7Fdj24Ty6wOA34paBtlt5zDGF69X1POcJsyUcryTQLvfBdWij6oItzyUp7yE/nwNy3QoLiM9YHftO2JkRiCWaGli030EgVylgm7O2TuMbdZYGODE0KzAy+bokKXWJLkA3lN+ZB/YZf9rFA7D83oZ5NxRmwEuQ7rfpzHNYDyVeiLNhLXNpY7fLAX4amArnN57F6+ydWRdyxAC96hOGDUqLgxbwHyzu9pqLrGq9MaVWloe+kyenuavHZeIhDifFGi6wd2TczVZPxN30aRWhALZ6Vcpg+64yWhG/htdb2iEh343J1bOFxSqFCH11wodCi/nkuPYI76mn9/88h9weFA0qJS81S/vF/txbGbxm/yO2kbcD6/TUD/JKn+wAlsvxp/9qW2lYCBCo8Enw9L/Y/ZM1zOPMOHHV0RC4A07QFZlf39BOba9BsPfm0iArw+3vyVb52Iw/I6p9uDA+r4TqIL3fgjpGZOb9m6YrZuPrNdW/djcU78aBt8hSh9+n+49U9Qdw/PfHGVpqZqz9ZF36wO/lUvOzYo6HeBNL3koJFKkxsQsNoW+Yqru614x3rf0uc+jjN8zFCYCzO60D1EgdhY5sxjqi9rxOJx0XIBmBoFTI73wNRQAgmQghu8T51a4TtRY5Cat4EMU/Q/8Xz07UIomL/ZJYpiGXn7udTZctDraGK8iUjUNMHL2+NRgSn1VRmUAi9umBQ3knz8O8fammQcKQ05dNsHeCIbTltDcLyW6JvSfGcP8zY54mV2H/7hv1r5WmDBQ3U4TZ9IHTnHM/NnPFVs+73iwk1shZ6HJh17Br0eBsWMWIYCBnnHCmVn22AiZQRLA48ARw6bQYZ3ejxphS+O6s9QM3ArzbKOI+atTel8pFHhZ46AR//X5KHU33d4mb2D7Ka1qeEg2YZQMql7mRoAzWO+kZ0DazxzGaROoeEFoE476nBupodUZpQgmCEiyucIdACHxf7W0WEGfgdqV8vMJLAd/EbahbRSHM7Qg2CEoTKnbINnLDKrkvLmBwV5ZGmUZpWwGu/7vWwatr4xI1SHdZepDls0FUhEcqNs3P/dZHBEhw8QSY1qhIT8JmJjgBB6cjZarQcQakk3ChPdAY2vkV3wR7Y+x//aKXbhVZZDSspf7oLJNXz6dmZpfOCL7uE39IdLBraoR8+7LVc96nrN/XBqz6flInRWEtUXd3z0jaMO9D5KTyAYui4QkHEjbKpXpYfrbBouzHuR1N48nSSxlnvEcMU5xCP7CGjRH95TMxsengk0YO/9+zGpTSqp8HPyqV8W7QKtsOY2hFcwfsjVDTTiEhVfznj59xhOsyLEwi3PQFFHMQMtB0LM4FUtaeLXtnDNtWrFB080snVeRWXlf8kNzRSHFuYtFDRVL0tFK7ii28CLgcMPTQX6amBpzX+/GvF8CvogTc4yz/rdeyQwQyKWLZAdihNNuIVq3nBKeHsrvtozVxrMCNmxRM1tbhzQPFoLvfAxxOCGpwHhBP2Ps=
`pragma protect end_data_block
`pragma protect digest_block
dba1edc6ac3e5ba8480ed50222823c2bbc1c28f04d21cabac7fd52d48ce4d948
`pragma protect end_digest_block
`pragma protect end_protected
