`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
Rx7ZO5T+cBu77C5pAq4aJAvVkVB+ltUnPc+LawvGaR5nc89aSe3xwTuH/dGM5QeG/5KG4srS6DJWCxbUhuF6GXKKwY5TUkulwQqxod5MGPRXhI1w8DAsBpgS7tQh2GBXa56GAy+lLisvA8I1aAD8S0EE9GWQ4y3ZPoeRV6/TLc0WJnNcsslWhcr/hL8yXOc8gL2qlY9HDuArBcjIhD4RDiPlnhkBpSmbRRH/Q5+BBLhS4TbVRgopDzpHfBBsIHb2SIlI0VQ3nSRHtiDki45bWvbDNYE6iKRk6vVL1VjrtEUW/HdNIGdkcGYgO2pripDO3TZUgU73EJUsGHgERIucSF3NApC8/bFDqd92ElmeaP0nvacNFYuPoiVjLKTq3Kv8SKIRL6eXQcf76ElNYxA5r8PMMbq8NpOOcHsJggjey2FhOy4kpXUAC5oL0xFBugI7Kkka+eWrVGjB3jF34Aoz6Np73SpNfi33ZxzZE//q0bqRhQJddd6aA++sk/ZNjDvhqxir2hqiMZy86J9/uLUQn3JbbXqSwya3Dun2MUTBirrG1+MTFQQwnmc+oLnhXy97RS8/8XcJylzse+mXGI0Fv86I4MFMhUn+BfOWlsllkYEO/hNPX9rX8nOfOz7syCHxCKcxe4FYV6JuB+XLDkidLPxxxIYvXoUu/e9lcUOB85qNbbBNAda1As9Wd/xz6qn7cymlRfucI5t/AxhTDj96PafZbaFakDwijdgqb/E8ZUUIPt+1RClhvU245EiS8NbtsLeuxUu35odoY3+kg/IKrh6tf9ugTnqgE1vxTBUvAYpQbMr9c+yUYECBLlb67EgQKSYJbTJ096FcSaRtDtFs6UEso1Ln+C62SJgSpZtXnfQRi0kJ8VYCWGiwwrouZxWEJuTl6u204VoN6J6U9VlCNhDMnctuJJkIUOxlZD4Gmncn1Gho6YfZK9Epu6S7F54UD8h4Nq6dDZeg8Ty6EjomKEBAautPuF9q6iM1lTQAYvfsWEONyKU6IcGlritT9d7WyqBvfsYMByus9CIXs8EYfnEwfZC3QMfw6IGYsu3YOlsa3ogXGDhVNVB3Wy3RgX7n2Twfj6QsRXpyBvtjFLqqGGudMm9MDzn8zbXekJvG+cEegNVQgd83dclwFlCZ9IaYklH0FtNCXVHrJDZ0S5YRmeaAMnE+RGSG+/36xHPTBbV+Duu3pmgAsAq1tl7n0GJdj7UFxjigUqTOCpxeuMSaOrraS02EfMUEcemmntr5WzLhj3qa2djpbHx05dHxUVG6qshJ9PIc8vTw21s5HYgS5Ng/FMx7QFBNPFqdTlfAZ6ceEDeo3S3A+2IHyvqcgo6cP39zjaLzz0znc1KgPkLcJfNzUmJ4YuBvWQL/+sQk64vg47wfcEcWN3lT8hf7fQWp4jQpC6sR7rOM/K6nZezzUA88y0qVbVV6u+YwTdwnY8/wrLf8RiPX3W0r/wk+0vqeLIfVIOHiYEoaq7P9dk1AxeQDP74+e9lTNHxWwPwLGZy881VBtlfzchL/OIod4s/HKDmDnKlEngVua803kl0GLDJ++dZx0PvO+dQzvMwItaDmoJy4IQmsBRjuF8XmabeNxt05TlbrZVR9FRLJ/jIHOIdU0jLJIG9ncBuWRJvh+7EytkiD9b6gY5M0JCp5aKWySKJQ5yqPGAxYqFFd1w1FxLuG+boLZj6LGuWMZNczVHmmcYkWlz5MThoGTZbiXCF+tqokv+kVYekWqjfxKLMgmfbSjgxDYhbB+rvQVHwvJaBCxA43F7Wj99ZkXhxw+VayZazxq0zfos5dBUNxxGcCNwRbL7FAlRCmRA+rQDZ8F8Ah0gDH/U05nrychBDIIa8UHzGrIyF8bdYpOTYoeCUNTVMYHFmmJy9V8qID7FX/xlQkbJWq4YbqIgiibOn7bAoSKLQJjqt+joDCqpbn17Y7iBwOeWKWvqFIZDeOFzfEquiQ8J3RDwWxomd5x9jD0YYnIrPdjbuZin+uCUXJcMwF6/uakAx2a448QSNr8JeRs2oIYijSnUDETJ59TuqRM2wC1bIGy3xto83IPdMhd1nkImbS/vtxGdUwFIx1Y04uTrNfqHd84uiEcT2EUofC0qGI7VFLIGYCvMEll2ooDTg5cCh96a6Vva26bis3w14jvxi16mkrpk4V+ZY2kVqdo5mrrJzj9XdgrAu5QwQYsc/kEeLBAS8r625kZfNHYOQlPrcB6w0vlpq7mv+cI2GVOFloFkAzgrlnd2886O/sy2eqvIEaB/+UAjS7MHPrZx/ALTcMxsxNX2eOxvETokJBf4yaqKw1sB513OYl2ec7rBs7EpGocaFmZv1VAFg9tR/ikAHHuPSr/LpHhSb3bVmT7rIBbz0UDx0DCkHrcrUmSzKIKUbSqNX3nZHjNKGtATvhHnuUhkbgYWH1aF6TeSy4L7rUYki1Tev8bsn7+6KFKsNJAFS/ukD/iGtEqgapC7eMpgnGO49nM1qo2uNlJCZlt3ddoGQ1tU1OIFfMGP9P9sV9ZVCMLvRdmRtBt3F5ZUzQz3DyUmQqXuU/l0NAeDsnmCS7g9nKDT7E63oontsexY+XYvHQz/r2RZ0q7q3b+u8nSO2WbVvhxUYTSXavqNAOCxTkK2Ku1c0Cj87NJgdzaYg0Syi4mL6eeHSojoIjqWaIgp1C6hYej5T0wZDpes0+lmExRsxACIDjvSuPU/2PJQA7KWJIUcX4EMJArwNTS/W9x0GYIRN9B3ezDKfKpHwzi+5nwX0pnJxuGGfd/27isMTcbp2X0VjQV5i5ktkEJQl3KiJJKEozggOSZz4rnoWQFiVs7iNEoToMeG2vmAsHkE2yp6V7OefDMisRVPUd7+dvOWr0FnNzej/tfQUKYnwdfn0/D3EmjlDhmil7LrozpBFIhisb6/VD0H1Vodt0Hwio5CRHN9XmkWLb2eiD+IdWw1mMtKOZB67CQ1msWdMqoHhumMJKf9VtCulqVLsurfhV5KAaGj+Y+pQfCMrPkGI6c3IEJje5jwbPK42CiRwpEuESODOrna+lzz+Fatbfjtc19i4wWva7PujuJIcUCr6P8PmNS65MwbN44Ap6p3KLcqPK2YssqymGH/AqnnAT3QWnjrwdrU5yBuVHbUphlqOxMPB91D3a+vGRl/OCqL5cELm8tycRLTZ1yLIdclskgcbitbl2zINBdOz52C/NNXAl+K8YW9Cfq0UKZ9yvcMT8T0estBSUug2Zv4IWmJreUfTRdWIt+/8UtK6KzA1si4RiStHmoIUPdWd1+YBApGEHw2/FjmWa3/o9O/TL/6hNh/ChMbf17L8veM88VpRxTOqqPX9m9XGNd0hfbbkP8ZDLNWkzuwIghfzX0/ZwdWo+pUTqxeEloFLs34V04d3A8Tr+y2BmDk9wJzbcjBhnR8mtJWYg9ZcBEZty93XYBfcD8e509bMzKhYn4Vmffzlr8yooqri7wb9x8OBCaEMRHOLCQ7uNwWZfSVZSJQy33U969TPVSLBRr9Jnv68zwduEEGz0xhfLS7ailkQegaGWlzW2uo1SBo49JGVAnJBSMllsCj1K7D//nNFlfuwbaG2ZMOMaao7o78sHqIw5r5EVNL5Ej/85QoW+2Y+axReljyUIKtLHnz9CtVq3xKF/gUrvrfIoprOxryyk1EVQhIBZ/7Y/KvIc9Lhym/CH4iHroYDy9DFU9IPuZiTotPNTF+5c4geeI085C0ktaKr8yHpxnPtNBJSCC+AzwGN7nNn5TSOlo0mjbavxzVlhjDXUn8Hbe6lsU9aEJI/scqlBJ5QIXts+M8zTNBot87GGjUpvKB0FEMw2TXg2jFagXHGWm5VQpIX7i4wI/XMpoWr+6aSfmY9hDNaXJw1X5252q41fl+h1PmQJw3voVGN8a5Vym3mPGrQNos6PRC6a8yT8bNDzbNnVUxGPBZhXo9+QtN/+TrLXxHDz4jlCb210xftDQRlRXjBU8dwDiwtfWvlOABPSzkRBNCiiNlhdabOkaOZnIs8fGsU6ys/AfaXm+Sk00FvDQ4COqvjrSFYkxsj4wU+l0Ild7apdDctX7n54870oEdvqfBfiCA8PXYM2QrnaXH8jRNO1S9CA6YdXsmRUpTnyMrgf5uMlGm0s7U7an5H/uJeslXoRQEMPaoOKURWNvPRi/HmKvCHlKcZf6LjHctdV72k5a0NxRVQqXAughCvOurYfmrrAhGTojgXxLpOMxTI2uTEg+P7eoDJ1BYSuBrS+2kkXlklTwCdZ9ouNI2ZTrSQnkgs68NMEmlGuRwyFiWqzblEZphTaAESNv4IfzGX4O1/t/h6Dpnoinltgzla3DPd/BgY7reZWA6QtcXeop5VmCL9RhA+dgsWlLDXYaGW14c0g7Eyc9deYch7zqsJAjMDc50ooyeP37WRHyXgcrHI3ZBKtCNS44Zlj/gDBSP6h+28+nicisOvHWY9jlwHj5p4bUjPULQBZyuMorMjJOwXHWizrkHyw/VlISBRFmCqe2V7kf65NR7BywytqY+wlc/oSf8SkMWfigDUYQVtZj9vBDHFH0F5yG/u153/6+QkxHi0i4SqxvczUBusvGuzhAzg+YIqECpuvc1QpPvqux1lSTkf8Z0N7vAzBrPIo9yzU4UwGdHBr1LMvXwiUBOHPkTQTqQUlMnTsTo5Qrla2pDUjGVNz2Ve6RUKaJbbt33QvMlJhtFPc/kMwvp2OmE2z8Jp7kU8GAbEy5kA4Nvw/YpmZEr/K023qzE3y+yXmTxOqV/8OM/3OJVInAjavpmHqwhUDCqCogndRMAxczSc4GA141wKtkGFdhzYSnWXkfhIo3LYF6pQ/wOxk0Rb5GxQGR2nL2PTh1qzUBIWksVKzWGAyqmakj7SvqGa0hhT2swuX3o1jqJ6x9ZAiM/n90RrqVo/Xsx7Ewdw1jC+kCOajh77yHdySEhsLkdrrMQzQHZhqAnZBJM+PoxTkEST7zII8LMbXZDaS+bjmdWBXxYLA9omuqraEerKuAun6AQBu6BMpEen5QSDeaRPXYtaDMh1hokMH55WgJ36XYCOIHkkZN0/+WZAjclO6lhUn3VyncS/Qb1EIx5qecxqoXy3nbb/NAr9NbqCmss0uFv/s+XV4BmUQGPc0RahLsziSBcJrWL+/Xsk+dcWJXNlQ6LqrVVvdJDO0gmEotdXFkKy7rSuDMkb0XdUidzwbg1tkJBOReiU5EGpXbY48x4+OSfX4yxO/UKSJuQ0UIz6qqThY5otBEi8sLl5nk1ibU/QMZGSKlvEpC+OO4WBzVKH0+pYXbQ12ClJBW3vKLeSmXQPmuVMFwZNcZJIDrvUCbIfBZAL1d4Eu5cUcOGtRpZDvy0UxH3yQXw6pxiE3Wxe1b1n2oJcweDqL6WVyimHY2S9ynNQlTJ6Pmfbv8VntSybL9ixfJYCv13MCSpsFwYCboCY5nGEL2CMSDAPumrvEifnelcMz19rxcxe3t45SmQ86mqeddmPZvL9h78BwunsNhRwQArVcX98LDp4im0HqeWNf4XQEqfRPwWvlJ3qepUqEm3KfxWvo6O/rLS2dGZzLW0vO79Kwo2KBYGk6nPxumPdfGb5/Jc7nYCT1efYTTX2+yHjl3soD22QdO92+IUN/JkT2per1Z+fEwUkz/PqwUhJ0TRjC3wt1lqtpmfcbP8fW1uLj/XrU/+vy1Uq2S7MLREKSFGt2ejwmR5pPy0Ub92XKweoDOI2CyAe0x3rGqvfObdaUOsGgT8VfndBP9MDH68AN9S9CvLx8xPzyhpPqhLz0wBTes01vCtpLZSJfqUelcSK6amC8Hm3+SEUYTXpxWQqXZCLL5KqHsLgBdPES+e8Efy3b4AN45fjmEnNixE6eNltFZpOpoPiQc7PoPkNWc5bZT8NuKyh2JV+uggstxCaaDbxi9UX5SOQ+8oNzN25NCU+jTwHSv5Ot0rImo1J28xf8ytjicBpoptXutAMuaejN3aQhNvS5LDTC5SyengwjFRBHXuAD8miP/YmQStWvTZ3gtPMrZHM9h8XkgK+QpVoNRD4EeDnw0Ff5IlpWBfRyQzrw77Vl47wR4ruQQ7XkvdeTCJucwHInWPwy8MHgDuODpUpGijabS88hzKTDRlwlYXETAt/pp1PS200p8QVKqZ9c9YGbhp/3cduezt0aBGmSzC22TVWNkICxYCiEDEwd5fT9YQX7qWEZXVQG+O81LVmlQgBWqZoSxnp7jJ5wAKU5xadulj2IQWTHo8aurvOGpofYWx9drE6HPKAOq3/bPcf+y4Um6Skt8ivZ5tJC1940MTiJinP13wDFMr1uOPlMV1tEaenBvaiiOSWNM9n/4fjUA6/6xAcUUKbQmYIEZ2jV4+7br0E7owuPszihoD4k2LO6oNsEGz8+iASQED6wgIGgnocj+Ddkbw7pikqG0ptRpCqhdsOpMrwNRn2wbEyvUwQOVrTZgDNsRr+lF1dI7rgIC5nRggsZy7eQ4e/XOEKmzbkUEcQIuv5it+Li9D7eyUNLz/+DA6krK48zOhWii3pJOJM7IngcAHWFWjc+ZpOsXhMS4+RcCkTNpr5uLqHvFgfoOkfKvFb1rDbH8BzFuHA6UiI9x6LGgh3fcAP6y5/nMdlszR5LoDyg8RENR63O8mngfM/rGU+SBKnfv+BBxxF+J4U45og6rjzZHy9lQjKR/PN1OqMXZmRJq69BrNVMjS0zq+E7CJSS0ctiNbT9HrAPQVxcTTEMcn0gtNIwD93WBGCUwomecTxospAIDu9wR6p7dmlUzkbfA+5rD2IsJeBKYUoGEY7D9CNgufwBQ5Ve5DA/lElHKuTffQbipQ2mPZ8hhc6abP3fH40XBJSso9ZC1H+8RQdr1oFWyOEbKefIaLMIoVoAedld7bBFRFt59F4U7z16qW7JS9D9gTtu0BkiDhE8k7PVTNDcmI3CJSm7R5CihJUkxsMA70Ki4x2kVhKaJpGagKJiApSYLb548u2q0IiMW9is5hsXPN7Bc3uoAMFJIUb6wNvYx4W0Y2eq48ivnBk2iCpgVH2MDJN0SCoUPbvj/8y30AfNqQfTL+LhRgr+2xRTigl6fclEI2r6t276Z6Ght2tJLcQk0+aV6S8l5WPE6vZVwJ37aO64ggniWuINKuveK839fpRyF7VCSufpriKm/rJ1Ntm/cpTjySIEfEvyr3GmqPMdwCN7p6YjTJdCGNd5vi1bQkdTAAcE9MYj6W11xhU8uSQRVN1M6a1NC/t6NgCcxpyKClOwSvVMVMvQdXz3E1GcpPtFuSgiTCJTQLBRwowZRb1SmezIGqx3CzZ0ZaLHFFAsyuKYUkwkM4W7Hgaks4ZtfY2W0DW3YSmzvvMJ0rHBE0nvwlGyiJdkn3YQz3jUvel50v3X/4mrGDrUyWUy0mc3V9Mp+yT3HXGK+Rhk9rBUrnNVBCj/9g8ob0ohZMXwEKOnYmkeryiFb/LcyqN/0mGgxXLmgdnZBRI1FmXIAfUHF1A212FWTumZItaJ2bmOATkto0VpKHXU2Gw23EqfGuq9Ec3k5BQHViaCh7xQp52fsKKO8xADUBpOc0DJqRBwB5jxknjLqNREctjcf/hgYS78O3PEsOXSqqpkw2X1X/d9S7r1y2Lyol6BEgmJ3A2Uu0zfllFq5eKXnh0CvMZVXnDyNFvtuOEquJ4a3Gxp2XPPxcO0D6b1HQkMFoY1hpbrvuzIQKTBSS49977GtXvkcuzdNhPOj8S9EvTHcrW49oUzeRSu2nmWHScjp2sOeQ9X3PX3KwEf8kPSvUyy3QHBXDXSgK1DOZ3O3XdvLXMxilY9bhVE9KqmexhWRnYFoia9iG/wdthI7qQNQ94AIrKZ7+TXgTG/NSI0jQKh/T3aHvNS2uiprYTD5sZmr3M/Tv4FUdx0z8IuVRA4v7W0U2YYEQsR5h04NdS50NBJsVhKAy0FTqWd2hjygpNasKewSDMdDzjM9U6/hwrrQCe/E23zDJRT6uTCPekM+nPHynmeGWNprdLnoOZbv/9m7Nd1cL1WkPwUGdBMK+AYzoqBm+DPQApD3oNNfM45LYEawdVeuoH74sPGZiW9wj/SubsRJhHiTAvpOcGTo/W7brcq35yfSImUVrG3GE7ldNvdrbqmwWMYnKCMxTgnFx+MdXYGTHsMeMxm4hy/FzFe31z3+VJaNtPZ2DhgPdiu+ZxSdqhjlax1l4d2Gvr5OSILPwJJCDGqaZAPCDh3OKhKDSpo5Lh3OsXGZfWHPWZvFUo7XgwNj+KUdLC98hMSr9j7BzSBJIQNIGh3bl6hQ1sMAco5/ZDvAbusVZXY9+cUGl41sBDAIjyigtmzmIAiDQ0/kFebJfsqa+7+ry9yFJy7rKdENGe/Mav0SSHKxyYZatz4myy/JLGhoJuKTTjsQpNyaDGzwazOQsbfAzPsvfkZQRrM205OGGimnXCrpfphe2b/FreFIPYJM2NJPFti9+kJQJ5DieYHZlk36AscbOXgY/mvV+mGRJBIfqLYs0IxoIXqyZS86rmtWxdl5SiWV2B785atz8slXnUcQjpnHbmYQKIL34W15YMbuvcM694/Hruh1ueB9/k8IZ12RLxgUtiWder5qCGZlw56z0zreSg9RHSegJvc5RvIZ+NZIcjEl1k41h1XKvVvdJ5dx2tybnqGDl0l2JF+k98+lfbuUJP4HuXJXOf4Sm29j3N+FAG+he/bwX3aI+RRGpqmevwEGbMUSPOG7mT8nQDKNQWXCynpGv25zmQXgR8Ik6aJGGNPbXxoQy6sNRiSNZUEodqKqSHPrGwKBe05i0+myD1ku+99iAJPtVtDMudekxo1ML0VvzcaCnSb5yAs76JITusB7wcA8Rdk1DMsh9CseVcE8V5w91RrBoyukAO18gmmB4CZGPQ9XZ2vNThrVM9XsyCJiNS+qnCWIiGn4CzCIlYsN1A91w/cBjCN6RyXEJzsdRvzrjePo6OzfOaNaUAhyw0k5cR0/CyOLBTTHN/S7OORrXU3CD6akTad9JZPQ3WY4I66ddX2QDOyJGdBelw+jOrr6Cp8BUNTNHPAi1GaqlS95lUv4gBqqlf1x2SMFqb2kqFUhMcVRMfZJbuPnPZvloLcZ2CHXd0DxGTU80YslbXyoV8pYE87UkQHE3NF7M1o94A8dH6oG3n4mF6zs6628O2hmVw8ZXfAYQPd6fTncrsEDsiuOE1btNwUPNKf5eI1DxdxPqnlJRmyDBn+f9aFHhtD/dKYmSEanqyu4T4WbH9saKdlc8Xuud+l5Fex6RueYSS0+a60s7+a40WcBmEqZbmMQAvFRAuq7AQ+W5cIJ3tzsNUx5B6WR5D70uWp7hcbj2Vx4G43sjVKMOKPmerRnKiurMAV4synASygjoHcgEwuwDDpVu5gkuX8DX2jOsJaNjA5L5AviBhL1zaKDaCcsyIKdmUwWEr2JoaVX1XnD/qYGIVqk21h2lUXAr2hKegmXgyun1nV9e/uRYi6SZFzmkN6gsdZhJGV+AeTSoYvijEyhkFm3VkTTi3YPYvbKAr2lKr6rdl6k2351uSXNCu7mv5Snf0JTHyj+QC84AzuOnaU7IgsIKxQZ9xXh2NYuk/gD3N85B+aHbqRFGn6y8HpV5n5XGt7Dq2S8uM6KcVzWfdL11BcTpqZIwMwujLUARBNjVcIALtTXMR1XzSWcca2V2bpcBt1I97tEv5heoF5pBgK7qApCfCQQVatPqvjAiJQkdhCe5AtEClRxbQz72xKzb/JfxF87301j0FXKv50VG9aPs0AXRONwZk8etCDzd++dbNArM9mKv7sZgIDYo6EbZ1obK3xNC2LVKVYjGIf1mmA4Oyg7GUguNJJmTV/W1UdxfFx5jpBaMuJ5EabbkiaRRBzkqnkU+eG4w1f6e2IXxEkrngaaJNozXQz4K+1blmMBsvxI3he5MFcPUMC5xnG8ckaF4jLYjymK7FidJEZ9mdrLyjDDMR6fH5UQsaKXNjdLCEvUBoB34kyLNC10j1dIUeMEvcCMFCEesY1DgHiHqPwkrGCffLrDzXsWQyrZMCMrN6lcYrw8u0TfLID8cW4BIRjgriAsvaAU8oZZWzTPUfrji3Bk4WmpHITlWm1q+5rLMoNGRPLCGENA2AI+lwnINMaYwqa6HcRjl1w2zONv7p+FFCKckj1SbO7hhfEhz8sbGyPFhP7iSsEqWhQF4eY6hOgy948L9WLSBXDCtlA//Wi3UWmKt0NUaNaU8DUV6XhCF7gJkWBD6zNBLR3R6fQg77YXXN6lzyLLFor+Ic+p/3z8pJpCILXSGr2/JhH354jrS6QkH3zERsrI072mjwGyYlaJX8wkJwNi9hyK6O3vwQmhnffm/WvbfVDqQHgPe0xrM+UgU5Hyrbl4SZLcfirb1NOnx3SZWk15RKppGY98mEdFvj/KcJIGWHWM39l4lSUFetqGSwakkpfsgg9UF7IWaqKJwVte6cs4w9xx9mYcgUja3stZncPWWB+RfsPUkUUiV0r3TrLAXVY5kW/ZBwKadbbbX1G3KXWJtIOf2ZHIKP/9KDM11CctcN9o/VDZngCV9iqBsuxx8mp/f3AYDz5zkkl4aD9KcRYCHaxJbZFX7d15luHd6s0nBrNCPyzmjRLmVrd77t90Jf9ECbBkEtoDpm1Ji7bL7adwwgwDqdxcUtZE0KC7t2LKasVg0wIoji2ljkwFNc6+QV+grWnkMET3bvqg8tE4yU8NyEOLhLhasbNOMwMNVRHyJ2K3ZOc7YCieCb3R7E5ijQqhlkiyJAzVL6R/SeFJ0rXzmL+Cw2Cmzp+eN9kVzhhZF0Y0vNKqapaYoFaytCLRCuQ62Ypv+0BQF0Hbr0MF2HgafJNbtYGcfGtnyUifLJqRB/GaenRxdxX6XyM9jcC/Y9249j0NXky02JAd9MOM/m7rhcWqnRB4D8nhks2Wwl95vchFgsnNUp6U3nF5YCRFbFr9n61DB8nOVRLJ0u7zrRcRpTljKw8QHf2t3F+hFs82r4Gg4nuX0qer5mvcQ8KEfLGw7MSfmqk5Ta9NCpdFUcS5DQDby2dFUxQYl7is9t8W8rZRMoLCcVxgC51c/88l9bTCEBouIxIvukurvjw6RThn1m0PRwZeBN8p803oaVZn24YYLryY7bSURycVCLPuE30DRyO8vfAq8LqQQ+wLQlTb/N7sI1smLtnEdD5neEMEOifJUmXzaaHM2/d1Gqz3/cqz1ch/iBWTP0S7I/Ds9iVr9UpKp1nTSn36hB0AB8smDAcFruwB/ygs/rh+bo7p4JHRXFsDLCXqkBRwYWLr1mdpeIHW3Li9BIzkRZgz4tU4G/IOYUxF8EU7XMqYXVAvhQLB/Q7bW1+hisa0unfsWRHYqvsA9nqMwNOiMijzWacfPjMdm8x773B4Wx/jlqBNHplH80TUYeXpJsj51zlcnWNMpDfZaAyRSOt1DvT8fqd526Sr4HPjH0aXEgtEVezTzGHTtujolGWvtpXtsuDRec0+I04s1JiFoO8vYSr/1kQig/1lIQ3Fluu5xbafO4b6KW5RCUBhvjHEGB1eGLQ/0zsmn9jFMNOJ5i6movor8R+1IofM9Gq/+ml/yJ2JTRSXd9mWFVcA/xHHocSreZn7yaFH8Wx3puS/Am2lRAiTgvEtGThf/7ASOREfdFftpUdki89Dfamg6p393dYeYzagOx1UsPUQQq5vo4Ju5hu1qC/s2lttpt/sXHklxPl1//BlpBI3/tjq6qt/A+l8DAivDT8CfdJJnSWZpqp/lJYSUgapG/7cQfCchNKEMBuMA9+its160Xx7py8yhZ+lp8LOr5aBETytOmiuT8c7jizLPGL/hvnbKPM+YEH9gr8FvUCvci29wlpv0MhauoHTV5updBWihK/WNbXtmPTF0lxpfJJBZwP9YAFleERL/AVSUyAcCi9AlnT+fMqBzG/trQezIGtQaZMyvJHqJTezofnkSZ7Flk26kuXd3KAn4ERSyPTk8JGYaqbMKLXcdO1w2NiGwYmhXAXT5zvHBA0lwcQ44Tu+iXUIPjC41DoG+BWQmB8PKxVI+Klts5KspLan54APsLAgeEmFV2LbD06EyITfsr+/ua2/FqhxaKGkU6GTtyVDDz74VAhGpS/NBv/BkjNhtWWQL1pBP2zLBL8g/MFn+peWRgaAI9EOO7sovR3r+vwqvVIJCBbFzStNYNZASFsyyj7AnB9FRIWQfE9UJPFXdYPtNAYcHiwSTQgvurnGtj2uUkpJuTD20nKJnVuVpV5ZeHPV0ciX14Gt5ukQnNTarjvuxqXxHfDbH4zHpgRK2ZT6Nxjjw78MWtVj9HsEokY50/hWZJrN7z3wyAxC799/gJRuVTMkCc3MMaitI2h/g5MjIeC0loijDVOwS+Eufg6fBThQCEnA15BwPLkW8wxp8KRZHHCTlv4bmXOdg+07J0u4bRJCqDxLpHx3uk6ZbWMwQNXqSe9pDxYpBQwpNJd1dytjbc8jnx+fThHYTfZcHSOTqq/dCV8cJ3x9fjstma88HpPpqMoX9Pw7HGF7OHJ7btBYNyP3xSVRQvIq75CE13ZzA7ikz2IaP0VVxTtuxgjaYKOvguTH4Hw0cuGXo0RraWrgTvEMb9FmamELQVDohnPgH/NdraDCxIv1IrfNE/6slBu8SOX96N8/Ov4ap7VP1xs4IpGtyL2X816fPg6D2Zm6j7gZRSb+tiotoyFuNoMFOluh9jqYcIzcRFhTijR1gxoeM6zbxcZyKtvc81joUL0W9jIBeyrI++MWrGGGDR2/Wt1PskqyrSi4AY/S8oGyggieLY0VX9pqC7rGL88+iHQ1QTZrAb/zCaXl5HXTqRPjSUedSoWvem70skDAWZEk5d1nhAWhVSPTxmUArQZiWQs4ILiBdMA5VZjUYQk9Nv0B4qFe2Xp4bnSlYosvd2Vo7Ipc0q7Li84p2f5xM0FDhuq5sCibcjyXykkmLtBB+VVuXQlhWuYMRMMtqcNRhpsbhNwx1Br+fL58caX48OYZjX0gOnNnYLOFm9dpVGmrH9vCHlbVDCKSpUUl1Iw0WE8xKokrqLOxyP5Po7YTm/l5P4kQxA3z5ji404mVi3dKKMR+fH+L0C6NnBOEt9BsaDGcUpc1ZHFmbFZOqiyNABAVwgWf5jG3HkxIRvTSfUmHqc6qiAqUPpznfATU+KJmI/9IonFa6nNN1+ItaPW3c7301hjHt/D7E71oqWULjWIUrHpe2vMxSQ2wNwJDvtL37cG5GtpRDYDTUQ9wSavFBiYdV/cfJ5ltqRcFdK1RnynJi7FASYfBXbnKCD0GfR16FEPcfVD5Dvx8l4qnhDcvPs20VeR/LwMSPTKxqEftYiSnM/fKjO37Y8ZwmZyKQa2ygRe+Xy3eOwdTw/eGafGakWJjUGx77eda2kjqM/LZKFoKmJS0zK/EDOwdDnngGpJiGiV60/cZTPw7iyLrw8/hpOTr7L3WRRBS+mdkutsreWxMJAlnxFAFcNVOVee/D0J0J2RQcyMWnvFJKY4JIFf2vBC93OPMq1oFbKAqb0VAPH0tXsSozFHCFCjuMvbfRPVDyJf54+JxXWzEbt3R1OkUWqApRsErXm7EkP0R+c2O0bjqMruGbzWdqmmNqMTt4iHyi8xts6vVS3uS+tT7XUl2NlxbW0s4qwQOX3+d6RrC7ckusIl2ZIja5KPivxrLEU4gpDxbQrCv3P9viN5i2aZNkaDW2OExAwDO7D2+ad0Sfugwb3zPVicwTilLou/iKWXEyAUN4sDYfwLvs92VZsBH24FaU689OsBz5eXuKleJDqN3U+k6L5XKVVXBxIgjQtHdoVsOJ1SyBr/+JWd0hAZ60x3cmJJkvD5kZCKxTLbj/DYhcTv5oA4PhEJQ0d9r9EmNqBac3aJsoQFIhP7UCyoJT3n0mjgjJot68k/eNA2FWzCtgcW5CSS6PzAURghLrMj0iurZsn9JtmhoDiUWSGpQesvfakbXf91u3rAuwfUoA+Qnce1mP7FixJI6Edb2aXVficwrelvb5eEGXmTxPYn7pUjFgGmFZ8bXXgl6lEdydOuTCYwxRDSVwg7cQtT2K+Lo500cq7P4t7Ga2zsIDchdGMTSwZHXoXQKkk681V4en+NVgHfG7pv8gAZr4kWYlRbhtHXURNTzEZI6HbVjWl6jR/2UCZUxSyjqYhrmz7BbEHAaOqxp9Atn+VONUnPpXqv/k6iI4sklw/6DRwQ/n1rzruAB65R5qFww3QSoE7GfGCUyvbUaTdt/Wp0/875D04xM8hZbmuic4vGouLmqYA7sgXsNcL9vVxBBBgvwEBWfXB4mXgbl9URE1t4msYva+xBLwZEo8caIzn6xRdKe6t8Ju0q2GpQM5/xOR1vxIn3NExXTJC8Su+4FWGEaCqbvS1+ExE+KQMNvF8xTVZ92aU32+TYR5C2Bey6BLhQETC7/+KqTu1T8fQ+OXtJQHpV++5naIe/enPOhG9WQgy+V6nuZVoxQI+G2rOrhIkqgNGmQfrGJmXf162rkdDxHtHlOVRX0hMBXlZ2Wh3sHddhjjrEIREPApe//IRaRPaXcm2chiFDxvQuh7DEaWGcQHfjq2sDkjX5sleCrJUNh3z84axuLJ/jQnb9GkVLA+HjWTHZ6V0TRrEHJLmrA9AAAkYrOejS3Se3NX4IPMWMwHX3F9FP0FEZsDORN5EnYX1dt2UBaTsuFQ84BtZW2BvycPm3pt5WmwaK/XQTUIwBxRtDk+wcGibFXYkgYkSj/iqMp1SRrpJUWKIuNqxN6DC5wzKogAZbhljGuJSPon7wcK4Z78KS+K1IXyF2RuYWssvOPpdNBMffej22RQ1cSW/ecDIXIx4LLOtJHFWv3/k/vbh6SI4gLzkDgV+KPgxj7e8raB2IvLazxchHA50Ba6LWs7DAImX5kjjpo546hcwYh47cFBan+KYAe0UU8D+WAaveulaHf19jyCv9wo5CikqdTfhehdPPYCbJihQMyN8wiGVk6nVjJg85mIGuYS6V80MHPOcsou4zB83JPlZ934IAuTPAHya+p8dvvTDvTRpg5/M4pamyPwaWQ6yHGEuLlmH9rmwSRZ+Yp4BmRp2wPfwL9YQnGXhdiAs163d8IKZr+Q7rQ5uucqT4uz1rZBTr5LHKUS9eiFFH6BuzAIrNmceYqv/g/MODAfCnL4nrVXcNVVo24VjKyRFi2/x+KA4EizmBodc0ZiHlEto2gQu19CE4C/w/2lhzNOuX+llSROkivlUVlnqeBJfV0Jf3oaIEgYSaqtbZDjlq4ntIuMty7W37DFeCiOiSTxUx/zNvk2/QYoOBRy0a6k7Ur45G+rV6NEMGHVvouwZIbjaawJLJaZpY3LDaoBeUOajUjq2t27LoQ2wlSJcGaK/Kmaz8Kv3HxCyovp74ZpnwI5Nd9IF6o1zYcNiRp++mGtzS7dGmNyZ/pbjsylibJbNY1+m0pxKQqSsznUJiHCyX0ZxMwJcP67pike4G/tLzMkCh5vxvY4GxKDIrm1i2LkKrkE7yTGwKCBcX5AgcGrU8JSMY8ZynKkvHpzpx18dsFXpQpgEtB3K2k27Fw9Il9xPu44wanzV09jyoFVNJGUkAVlPwbQxPKKMKkm8vaCAn8bfqXnQxskIDLi6FR0XoLInYbNekW97ba3wGLvVx/iDbQgi2onuUCpF+sz8oJ81S7QGI5FEwAOFAc14qskMYDb8pU5T1HlMp/6RmBv84d7BeY72ypu6cad+adkFCuerNe8BwHtIYLIErKO3YUZqSlVDj1HUYFjaGTXajo3gbEgi7GR9atLgyC4z8cpRMIS6VnBl2Vn0NnPSubvCP7fioZjDgLhaKhzQaLZd8p/VVWAlFiB865M+hia4i4ZefjIsGMEYHkH8apazJqBaxx0W7bc/lKjSzraStff2Wiwj+0+rsWqg0mv4qbwqJKWaESnKhWobLRjVAPIWKySmGqdFBVWXNPLXuL37kaX6aNhEErZJvhvAOQk5mZ/JKFMXaa0AlMP0uxa3JBjYsfynkuGYkdwh25tcoJAAWUd7+Y2XhbJcfH+mLSvgbIjtVJhNP45Kh+Gl033SLPSjVevQnJ7SzY5BDIBXvzzAWfRmUiv1hNGB6H/BnNq/Us9ms6OxB+SwcbzmWTK9kUsCbXOZCrV2iuqDAolzXhr4KDH8Q7jKhA5fTyjvZQzh9uDKrpmpUfeZ9RPQMMpqlt0Xvd3kOKKEn7I7pHMx3GSq1wckBCshbqhlEKNL/2NBEJt3ucC92c6AkEWfD5gEfA6RID3LcTzg/8d52UXNJZf+lddv/rASJWb1fvxoEqM1WWgR5bUb2qg35k5GLM0dXv3I+aNbeIY9a0gmfjVq0s7w9usQrqW4fVGteLM69NvYku09FeFWEKCRTMOh2GCgfoPXZI9ViReGjLnsomTbu94RNqqsHwCm2Sb14cTqVJqUCnYGIuc/OyVvtFWnsn5ji9J4HZ7H+djdhDOo8AHHyYYTbngpYdrAYuUAopJBjnoghXZj7PU8U8mAk/49APmviVl4ePevsIf1Ei0Mw+ZDwxT5K9oot7TkORUhNGY3zEWGRYquyGMx2uUR+2u4UB/pTXXuo/XJNz/WxbLQOv4kJ2shgfum4zGX4zR7nFxbGpZov1KO4f/LTFnXsFGX4BbO8rtanJyODwwOqB9aY9gRlqFuHDV8DlKEtzzoaD2wAWEwU6iGOMkUKfseGqeQNDLUhnS5+NKx8miRz37byuM4AFMzF4m1hOkNu7dCp4cWUvnX+kG7ON13W2rogs89eiu7OogY593wSMVEzNZKwn2x3tPK9pv9ekw6+biu8CPdH0ytYOPPt9hISS7vdnu1cER9sAzL2KIiAvEUZHmqnV6ubHmK2C5COJg16Pr5ayhUXvxJKFQEo3TMKxbWymhEXJY215HZtH8CXfXmhUele0Y9d63Yqj+g8j7PdZLCxkqG6whyBY5Pqagu1whvHoWAsToYCqSsxgFFNt6OlbMv/KdksVy8p8pAXr4GSCTHhOi8oyiVb3xYcPuogdA22l71JHS2/ox0+tycjJw1JcUVG2trTPgxNpsNv2QSnOzyLIlqvKn0ab5ToYbqYNcrIZdgXvdpD4sG1P6qElX9qPUPu3Fy60v64rqL9HWbiUj/mYIG/k+AsvWsG+aIGj2B83CqJTrlyLJKlowcvwOnheOdtKeIQgCwBc+fRyt3lOnudriHnNEw2tGgIqEJUJHrG62j0S/6JkJLkzaLDbp0chNrnyynT40TVYUEg04FbttoSB1f88Km1LoPKxYSSyWj7ool5OcBSb/M7WTHk3BqKiI/9yW29llHxtuT+GfxXEpaJ0WAmJH0SezP3S7UQLFgmUgK2I+Hdc7/LPUtxzPE5JLPVCsrcpHbP8wijZQlzKM8Q2VliAFHfMb212l4xFJJg1UyOZIYzN4gBv/diOzbr+Qh0k6fEpK1QjvY1ifk2ujeBE/pE40S2acFzCMGBTNFUSMENBqE5VredSqgbIcQ2gHao4QPR2a55+yr85L9kvZXE4WTUkw4osTC8JwaLZpw0e6qhpWOVZjv8Z+G7ygoTJhDszb+TmDL/FPkA9t3sJjP9Klm40ynvGsNSOJOt4JHYJkNTyHKXt8xnGRUiFQvzH/qbt+f9cn5m9dMKAe0hiaC7E2eIjNM0lVNTyPJnfOnYDMVO3G2VngpxKExDQi1vBItujHVNDRAPhSKFJtYijvE0BgEAruY/KEGu33QU0xQV719MRMLFGVPfXnngXQv1Z1AwoTnG304aw+496OVzBXT4WyOuU7QGzWiQZ0viBqT6T7IMOIqV75xOfVq1ULbjYdTt0z1XEqQTmbrt+asSuX6OaYEi+BanvKdfDSIk6JvtXIcnS09OHsLdGllKVYsSTFKG6jpI98oJ1PEIe8Q4pYshrLB3Q1IrI+C7l7DNkJkDwFXkMzLCe5gq0YqOpIwdY68uzZBHpOKwfDkK69XoZnkUGye8tD20+9BHyEcCNkDFkt7Efs0g50eWV8Bv8o5+ju+duHP27V+FuRBIufdAhgVMlAL4PFQ/AuBbzyTEPitkpP6UCzLy7SHNtz6+KZ5oZp5qYIF9m/ACrnxKeBgKWDZOydBQxugJiT/pTknZXJ+YCTHsD7jFKCpYI8tNGIs8Jtdo00NbdzZHueRFDNmsGa0OmIU0V/BLsDPz1809VWKCJC5eemBVdkqjKNBatPa2ppKSAMKzvSGyU+wIvXPfG5RAT6n2E1RdTwPc6FKVZfwxzKTPcohDwlNTdo9PsJND/c5O+BpiAZLsR0DbxnGpbsuA+bxwKOR3BCEFqmIysREtVcwxfC5voCMUcV1qwvbtoe7iV5RRUTRrn8hnYj3d7JyuWSNe/HoprQrdhzYswvlDFng66mpPih/C1siaTu6u2hvoGVjSJSruOi6U9vDTv1CHy5eOLkehLh+i1qEAwrOzQw+9I9BnYYxH1r5kF7Aw5aAR990QDfzaoBb43FnkZU239HgDt7Kr1be4IekLWdBftgaJuuo+gkYsaX9tGJwdPasooeagdElw9OZSQ4Cu7k09YKmgSJiSgbl9qIOrEw7ViM7ZAStxd5ZJKmA5Pdbxzop9n86o6lyN4pjLgpP+k48hwe7IT1SqUWrN6dRfYq6agCIFdBVe8xeg7LGd7uftw6+FIYv+w1J483dvChMZBzF3fpyN0T3eLotQQ2PkcfzOY/9fD6W20MVIKKqFgKmD24WdDTHu6qU9u5YgZggNccvTUXzDmUjwHMIrjzVz/rqK9ZTRKNoAntsuAYylfnKvpMAHeuLTZ0xZLO5EBMXGvf2zLg3gwH/hY6miA03kiYs80rVEwzIHv1wVAZ8kKn0SgNsRoUU7qrAxtkRSdWDLMJmvCjlAVf5N3p/8PyVN/iWmYhtliSDopwSNqfFBQncy4wYqj7ap+Y0FPMbOwwuPLEhaFr9/YYKLOdmU/aDRbd/x0elJ5nY3H6eKQisPnZMEhKgD1jpJW4PQtosOR4R+YNmtJxQx9VVjolvn/77FtLj2HEKS3DOfkIoytiG+zvITEeSxsIKt1dU6JqW4aT2i9bTJBSd1jgjLUbUtvyoGrbh7eyUDUHzTi0+p8/bPJ0smMpHKNy5/gzKWrSC1tCy5uSxkwn4lD8LT4/gyVaZV+9/s7oKjXF0UBpMFNiPqKQCJ7OZ5ePlk1Il2x0+rUdlv9UKue5A/4W6vyfkz9Y1jU66FcZ/DEPw2+UtiLfQHOxQwdJUK2U6/f8SBm+PQxPpCVRjDyuzw99Z/FC4gQ0upa7fUZVShMpYAX1n2KvKEpFnmYIcgwObapOmGpOwhEA56JbTJIFdn7MrG5IfmKCQidafXstgMfhDB+J1BIhLrG0nj75zwuV5w/Qsm7rMAONYmnoKGAE2JMWsGFcPafSDpxwfC0fjy5XoETAeeVCShZHTvH5v02hy0GcUqnAxKtik6dtYfB6cctPkkNitFhdYtmbkqRwvxL8UTG//89KjDCTlt8x7dl2zHa9jyq42/DoUJ/MOMuYdEnj3rl88pYCEMy/BUBMEDCz36/ZHBMsWd+NrgxYs7tclTCeWZSIiS9/ilUeBBC1SgBgXKjvdceLOH+Ja+yrrCRhAw+436kCwQHTtUjfMmYziPS2TFVIcrCgmWSNsI/2Ug00Cwu/IWfgP77MuuGNc3+4VoBVAUTHAKaop0zoG5tnbbglfKCI3SqK9KDjwvf+Jx1zLAKdzJeY+wP3LBrXg4wWxUhClqT+toS7V5zVpPkGXdVU2TAbISdZFUdCXJjgp+0D1TEmuFvJsPsSYRnk5bJ1X8evfXblQS9KS2kZ/foJ9sadZT8GbMWdd+YadDtdKoCXPvqU+4rf+jm44QydjIBaLKPcuAOa5/EWL3Uq2CJrO4UWwne9ymoQ25j+zWXOmLwEy6ZzKqwxCqCcEEVMK3zbpRBTUKrEEYAcl789f3GkCRSxqMGmcO0HvixoanNOh8i+WiI0EtAh3soS8y5y7Iow1G6imJ7OGrCmQ3whAW73VEcnum6nlLunSodaYO6t0XK8Sp4mHed/9ovofl4P5TT0CR4pYJ0q0kG6Erfpzk5PzUZzllqxAvFBecmJS2WkwgLrOqMpkQXjF8S49To23i3gj2IzVam/6VWURbJmQ3vpy5aPPpivR/zWfOtyknJDGKZUG37/GJKNtYoklHO+0DNVxuWDZoECuhxwjZFHmndXPoEYate7IQzkYOz8hFH5tkedTWUcjoTQNQq8JjSbeaIEPG44dCWfPdVIGmcCnrKuK7IXe2e9lIvnGJK/WP0B+FGaAECkeaM3mvC1FdfKN9jCOiLyQUcO/WOL5TqvTBn67tzsGje7AcwtXtW3o7j2BHF4btvaALRmC7lAQ8oqKE622tkTzEZoFxz5a14OwG5mdhIT2x5RmpVJnIP9otjUSDwKVfJcOO7t4cR4HWnqeKUtA/MZ8srWEnk84n5pxtv2Yv+0eewBa9A3FZy1F/M3i+EmQrqMbqRn7zoHCA3Il4f/7Y5J8DcL2sY2S29AfuedLfes8nXnY5kMNlheTt3M7BBcCSquCYSjbV9hIRPYDFG4SXmbmQ3Q4F1R/DI9btUd0CI0EI27CxN2+hR+eBP7TXvGvG2+ORpdmHC3kw4IvyKckBEFZdCBEqR0zLkCSSW571PEH6fYCpXQOSXmo=
`pragma protect end_data_block
`pragma protect digest_block
48afc70cec801479169e09c479e0894e4f21822ea9b240f5f2a5ca0349a69a36
`pragma protect end_digest_block
`pragma protect end_protected
