`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
UBx2aFDcGuLl5f5Ik8r74g52kB2kd9EQ7NHH+Tv+aSam67UDQN6veNXH+FK0puNt7DQ+7e7PIjmnANxHPuW6ih6BJOZ0TRvUtdFg06pBB3qHPaFqujZiWMz+smaWeU1WPNlJctUgKuPiwVKzfaGp5UsZWSYXmdhX0DIE35fvJ3AQTS+UUVcyFQSqGT2IG5YhrpwbS63aDOV1kmXcHijUZ7SIIjajRz91+ZrD1YFDO3rTvKmoTnSd6KHWqnBEbNfw2WZ7THtsy2ZvUirxv+Yu9Ljjn9xTVGae0LfrrRWJJ4/AmMH74E+cWcsNq1Un4UpPnFEreJd4fZnctsvdNmB4X1XYTySjsHxPKtB0+YL6+0a2TAfGjoCK5Gc/ZO/ijcILymoh5JnTf2jcRlAkprqw5tasn1J0T1Dtme3GBxoRm7HksHF4ue5M5IfQpCE+oEJfRSjkygIY7fjyaDAUwwo8fKt1x6nN9DPJmoxR2wAzx/ylbasxNVcvA/kXgM1zA0CoevV5+Hx/iC5xpx0DYEJovYfpMlFHuBDDHmHCZZqzQEhPZsFAHKPu3k+9vBuVMZWojWROsu3Sa+ejppT33ERmFB2OJr1mjHaiYhe2NgzlnAanxnsvZNJ42gKLNtW4mD3zJkAQt8Dxsw5aXPbeSq6bMAUTrp+4F6wA+WS7lVzyBA5JCMAE+EedEuS4luytdGbu+xF0I3m28jjJnqZ2I4M3m91W4dz4ZDbGoMl7hknO7m5XIKQy2tPWwhesR7c8CR3XLhB2fCVyvgPAxZXGv6ts3gj0SZdZ6vRrJAGFKq9efom5NlDTAlI0o6+cQvTME0ZAqTugMgfcEZChsVAegu5RD6aibjCNChDjvG1ejD8KU+uZGnzziaoMeYsmioA+DtzFnPnWd7wX3HaExiCgc358afvcJbjDJMv0hT3RnoOiElaYQC8Sb2FnOKMJSub/ipjVvHNxvFxm6qyrNgaxLXQtV2jJqOe1db4G3OiICuWSmPN4nfrydp2zJp8r68qID31d2Hme0b4OwCbge9D/gYiuIhpyjWBYwmc6F8bUyp2no8dcDTU99WPEhbkucC4SMwYN+BvDtrViQakMswrBcIBCLhRm7q5ozvWjKV76PJDquis6y5Eq40obmu8rdxb/2JW+wPyQDxMt+KQjqzDm+zbzM1EFyE0ioKxz98d7iXx7w9LZd5zOy63Z4vigq3naNM7atdBsgiwhC7n30IL9jGK7WlHBROlqK2qbChA6GEp4133RCnxgWfSerKLbXJM6DtZ8/bNuTZyD8dgCxDrwk0jzHHHxwsAq3BNFHX0oE+7xc6Bd0qsW2YGOT3e0i5jOE/58QNktpKBHZqp6BjTPkF70x+N/Q/KSfNdHIG8i9/QDYwROhVGD6gLxa5r0g4ubKIrNb7frXZYLiDFUazFhWfdEgS+Sybdv8KXQ3TxNKk+gkKY=
`pragma protect end_data_block
`pragma protect digest_block
501cd789e2dfd7e50856d2522dc54221e3819478f73f9ace1d89f28dfca00f61
`pragma protect end_digest_block
`pragma protect end_protected
