`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
eUg09GUEcSgpLShfcQDTFl52H3QUOr/Eaysq8LMp9goJjx//N+OsK+vUPZ5zRkyoCDnclN7wnyFugfTG08cnSQBXDaiarVaelS3YEaHjocHl/GynD5gYk3wFqSbyoFONyJg1qWyOGoHzJrKP/Hf0+eWnO9bwlypMX9xKpSWLnSjrr2LYex3S3lbXzvxtPdDnfBSDNb36x1LA21kZS81QBJT3z3vr/srX4sa8d5npF35H4WuPO8Z40miP0mMqO6j6atE8kC1qpLYIh0ULU3oPu4g1ebEOSwkzxd/n+yXn9hx5SYJneKFSpXu+p8O1BsaZDKqhF4ErTAugQQOvDaxbc+GmyhDaGRoaoXb7gm4xOBexlrngbmOjEMdtKIwMLUSpVug4yXV9oirwme+s+e5IOxwcM6sNA3TBAx+6s6CZtfUcR7P6GhSV0xJq04rZx/rb9ArB6Dl2SAYHk8ck0Xm+SpmUZRlgvFmsGGlZNGN7suyYL19oW33TW+K+dwCarPRNUDVrozSkMCRC1szXjFGx8FK0ALlMugyoFBrD6nGp5gLCnq9mLPllXxFWKJdIurnHfv79dIcBKWPDIGdVt9o68pyI01YWl7qTdun3aJWgmqEDc/P+laDTCXdilNTdJPphm3wlpCVWVMbfWsP/xVydx7NHlkJNP0NepnbZU1ab+afvRBqSzbitb3SE29dSfClOhuCxxV9AT5LqwFd5QDnhtH9RLm/HWa+grY5cIRjgT2aSHM9cGtki+bdXEs+NL+5Ha5piXs3v8goUjxeyQAG0s6u8JmhpShBU94TquVgLXGBpnR+Xgk9tRI51vws2HeU7c/B2KKeIib+VH339xHWpVHluXSq4POgOgPKL/IDbTXZEX0eUfZH9f7K6JXOor6q0Ozj7VkCM14Bi163FF8GCTyb6ZY5/aXSIX2jgtkfOnUuCWHFJdA9d9eH9Yh9JE/+FEn803TzYxbjeSBhkz/Q6ar4nhK7gmefwcZ3R4meZ9BGZN9I6Pcd0VACnRhid9CFZ9YzAGNhl8ly5pz/ml1IxyXWI9iG1KPiBaOYQz1Q03GIVY0oIBw7EQQGsI2agRVmcwD6zxN+TDdGGQUosGoPKrUoTIILDeKwQbPMBdPB3KUw+qCwwOhRScmXlb6oD+y2WWjAx80gY3S9P7r1yjZVLnEvNw294gNHtIoNWdrzJMpTobB1JqXC6ZinoFJvdxkrx3yfF3RTeWss89tMmt/Qw2hPOqrkImkS6SPQyw8UsbMSx2XuMZe4Ex7b069Weq8xs3Fkp7cj8L8ne7GfrQQhc7qLHRdQwlmCL46gyH+p0NrNzAu4Zgq83rKRKRv2eVDpsRnX/P82yiHMg51y1/0y27MzvXqqNmYIQIqnSyXGBTnGyAs03Fx30SBrBHEeNLj8vkyJ+D8iQayPDB/pqbpNEU8ByK364RR8wCVH0bnCS02fzdxUok3H57JZYAVy7+2mwnnACHlvSadcG6pHd7sxrzlPflGsgWL0OJJ8O+64mFnjCSdjUHQd2sG39RDWC+jbpbOSwO5fNTfeWOCsf8HyQFLiZFtjVg5enL9ymu/RKg1SnqrPBTioPM8R2PCXFkl2IPtjyjK9/Ht/PBD1OM0OfEjtFwIuZWC/DW7c2NiXD3jJnNAKHxPGVLIstCahk7atgei3jMCVjPkkP8hFBF9VFHQ+/IKCAAqBx4+9WZDs8Bj0vykiKyypqrPsaTcLcN4K9rPpkaOgBmkCXeG1rq3RlUij6G0w6MO2VjZxV9WW7QuUO+Ez9GXMOSmUkWjlJelhV4ptGYROmzQzHP4Q1slIKga7vyFJfY/J7/L/xprsRdT0LRnoeaHc4n0kHTmVsJfJhy+7pElCKinQXiKoqxydmPpwRNoYNlbsX4EiTyvCUoXWLm9E1kyRLeSLT4+0CjAmrpr+22kSsp3xB9hbPBJ9+9jwI3N2dBd9JWZeBS5FhbaOSrMioUkM81vsqHoS67fCiwfklZm1G2m0XYgDZhflNAyucbEgb570z9k7CgHTDxuMgw5jUUfw+Kp0KE09zmgIhEju+Hcnza59fjs10AdmKo4lrH5TZymJ1JO4Kk/EyQHFgtxzhasfFzdeWvQhcbpblp+PTDJm0F7cR9MN10+KTp1rwekUzWkyGheAKdfwGdkeU81PJKeP8RngmMxqR4eQqagVtM0V5Uw2Wssgv7LVvsLqlaqjEFK7UibBuojOJSjp+Oq4jLMcADVFooiH2+7OY4vyvBcc/qVi4FZxOqpVuaI4zgM3aulb6XRk7Y6GyyP2u1OJgGSMM9n5HE05Ge8j6UT2AOjweEOof4mz0RGA7JTNKynNsU16yShif35MRj27RFlpTGMBB40xJk4wgxpFnK5r8M9zT77VyZ9Ag2VapSDDu/s+QRG1BhIP2RTeJYUa04+moy311Yz32+hxbcHljsYzwJgVD/OL5TneVYRbkO5AG6kKpnlmi+0XzI+1u6GdPwhd70mcQVAeF2sQGXADiYTkIeElDaoP+eR0sPjbmsC7oxE4TbmIwuEoiLAoAJrtbYaCiOPZKt9vzXCwxdgZnDB89OqLPJyN6pAJnFfzeiTIaTIrvY4Ix2GB/zaLiBE2zoSLhD4UkDFQ1YJ/eUhGvKBrAbJFFOOhPCEUS8rZSBNgYMANPt5I9LK79REE4Jxy3KyGy6Ma4hNPb+b+kjKgHJtyCfi8/2bFeHBfAnc1bpFP8v8qcoVBTo2kdUVuphWMBB5iLv9CoVyrxKbv6q1pgedIkPS7rfXIEMlwNo47oLSvNUGRYFp1NItJaDZma9YCRPqIdRzcfnIvkZv5zL507ANtJKW4acvZTJn5tTTr2BSwpaLq3CHwHEku6BK+mt5YlaSentY+2oI4PH/ITP/KlsNr3AOlFun25wEHnrS52yD3OL3Xc2Liaa16O8BG51MROD/4YsI1cXFEkw4Vh6wnf6PYo/954ZFfbvEMa5/b6s6B/uTx9LC5Wy6N66oBRIx6gzuHaZEkfgiMXWOVKtz9g8PJ2byseLOWzoMXADlmDLxziVqGP4ggq653zgS6XDzY/tQSx99sYydI4pljIDfphF303/Ju+7dj0AwhPSvZn2YekAkk/bVyU7+eSHZVy1OqebsNFDhlePwamWGsHygllJf5XxTDGcoyEarqL4eh3ZTy8SH5CLlaGQzdySxoApeEGtpoAG/kBBvivSTLYbhN+acvCR7sj56s0FbzpdaGTMoSFt556Chyk5QDYalOFy23QgW/bVD6lr1jkC5RT0sFKpIpsHFv2ubb5W0k+Xgq0rX80c1z45oUJtqAQ6QdcBUPbpMzRv8dxpFsJlaTi3nHYVR+Nl2fOYoxrqV1qUZKUtdu4gJi+vNQ82PnmkstWyPB4O+4fMer2Gnaq/bqWkt2Jj0Pldc+drypb4F+sZKj0EUiZ5G+z5Zbx58xYWBGSCGipYF39czTGl4AAasrh5EzmfF9y7sc7ftVYzBgX2VG/5V/4MLCwL5kOGc4maBUZpwNOhE5j0ZNRbN0MGNQCq/hpTxEY0stgLSOh9gEgHtBoG90OQ87mXWswzPeDoa4nR68OsVv9Ccosy7uqfO3Ps4Ngg9MLtUVA7LT1Bs0B+4CvP2FF+k9xLsC1p5W3McsQ7Olx8aFfdb3rYG2MlEMOLaPXlYm82YMzqeMUoS5/WNnAh11JOLKYbbNgIGc7hJX9KPmM1qVG2yl1ceaMqOyr9xWOSO9ikJU2VeBGBlkPwR6oF7kOeTaFmmyTKiou8SeTApTNtAAkyqGdlqRjemsuK3JN0oIm3Xlr0NXo0oAPknAEhU6rqkEDDtzgmjwNiVjIQlXEz2yv+HLy9idOBMSkfOwAeKvV6KW+pOKJTjwy5/tELV66G/NvITaabhzo7XcJ7QoWe3OWx/ZdSihXMJzOhWIMlJkauPPL3jZ+v15QlzcTr9E+eyANFiagXEKnSpNbANW1Dn4Mgoq4DBkH5SemhCofe0b73NKgFvAnetgMfeGo0+IB4KRe98ZF6dvpesjAymXIy5SWz8FcaSAhTwl4oyr2UucEdA5LSukyjtjU/vcUysvyCgZtdADxmx3Kvba4kvNgKY1rdZRlww8dUVGZdG+mWC48kIRnWiHM/sFMIdLo9BiUwPMLOWwb8J0oOFoqXZ3zCEo0vBwBXn3M77+L+bRFZt7L4rJ84j+l5iPkCL8ETu9qPuVVeJgppWovf5HNQanMKzxrseYU6hlwYJEglS/IIC8CYEsR4i+IG2SGZkVgMWWcMKa36QjG6M1T4A+WQ06Of/GFyoHCCRWX2WXiXcNETgQvUlmnyYUBvw892Ogq0LdQPPzPUksXsZlXtQET/6sjyvCwhUSN5a/9oVMcNsno2fpLeov0p3ZzyLV1zc3PoDInGPk1B2LdeXZKOiSsAIh4IYNOPn5U558XFSuV/0C3NqUYQbdwZNa2zCFBVB6N+9+CdTALghuh8yh4kpYfDHA2xhfHzuVyAcYyucWB/h00gXGOLId2hsDLji8N26oN76XsojJXM9XbC/3XQN7SXRklqg19CnI3ekTPgKipTtsP0ZMYIAhinqs5kxjijH+Jgof9CSRHaYN2Shkxlw09wvw7CvS9Eb56+VndCc4VD2i4RInSuzrYi9nUGQvPl0yiIq+lGvj/CB3UkkYAHYJFSmCLB2CFTGBX4xQVWsAuOU2w5W1PSXl2qaJCa3RtjPF8ozv5U9/AQGLifXR17+ibjRqP9iSGpd8hSzGVl7CX22ViifuBwZCt/D1iu7C4y1qmEldKjX9P4UP7QM773zcXbRhBV9jgbV5L6wzTjZDoVk/ITels2o2jtr8xYXNST1kWUI1OOM8mraxPNVL56s9/kcLegAr1aUXm4USW59PMo7I+bSBRvIQ1NTl2NgxpkADFtzAi894mpSVKceajFhetY0i+cuFzMU5w3Ua7odAcvHtIvaDPe8aWJoXhAdrkEkR+07Etuai3CJWRd0D/YGoEOV+4F8ASHpl6z/wPdXElkC+VXB8ua2Xw9u1EVJWbeS6x98oJBDDGWOkTp/lckBlGncolFmR3HywggOAurCZI50pApNp/0NxE8rwArLdx5/jQTyNzjUxlVEop6ipbBQZ2/nqFzTlzA2/fbBdts8Djx5qLKU6y5vJYN22dw8zGsyxNtehxMrJSFphm4u1Koq4JifpPsHQ4hR5iqYV3oOjExcul6eD92pxJHbspmFnnNsNDwBEa+2GUlCG/I360y3diKBn9li5LCRVaBsscD1nA/VcY9TYhpSSHQbI/Vz4G3uJoG9orcltoYCcWQ2WjOk58BE32Ww22ox5A1zMV9jtMMue7h+LhhyNHL/F2bBHwgKNp+ISJOeuzS0ZBv5ecb4mMlLv6iSQcQQkzPjIPY+v+EAWmY8Ke1XqiApjNbrG7A42AgDjcIL7D91dA8LPa1etPCXJ71qk7kXXlKZAX2d2oatJwgeOlzXG0kMCr+sLfXEEkaW4a+A80cWjwHrKl2Nvvmu7alg3yuGuXYPEqGyUCnn2z4dlntpgZcCf0I1KeSlCuv8sbyqvIMwrl9dvdRDsHPeh/KhO4qUVP6ZKiEqiQXwcOnEmpYog//AxbKMG1BPOhl7RdQI1JxoV72FEhhb5sYD0nM9bmmbD8Wavn7RcP3mi9+KMxpD+kuM8mz9+H+T6eTxRr8UND/GRA1NDgZaHjIpIWtiV+ipz1exrYps2so1jZuqArSn/sfCTxEPyRZ+JK6hTzdl64bG48xo5J+henaBzWiVrKfLSNJ+sXCzyHKJwqrpMIMIZRO1O8z9txXjNZ1po+StKMKhxRzGpBqyzEZqqjhSj1oMzihR1ua96VhloFAu5jt9ycS5AetFD7bEdR9rQL92Skuv3p7ajePeWYnj1MkggxeKQ4rR/ZbDCYv0RzMax6yvWqLMlqJPRTzaJKT0AeAR5gY7PucXAXlb0yCIyZGXwSaTMWtWRnWJsFqXlrUQXp+ItLMhEbRbuWGWKqgk3ld+O5HTo/CYB+pdQWY2lOf7z5j4oQA39FqcWRL7xrOhkdjG3yEBkHZ2FD8HthkgUus/0Lkj5KypN8BloDg1B1Kof4f2+ffad2nW4O83ft+GkWg0af1IrvBOP0Eec9cXGz2wvCvo+zekcmVWIr2pyf42hD4qmJed6Jxnl4caxAUQddPeXGtH7sXARskGOOT+rxPecyAdivF8k0XruPb119L5eS24uCaRQ3OG7vM0G2s6rIHkPO8GXeXpYfs7s9g5xLWGX/+WY9nXweXtWz1cYK+oEdU0/QC/qRFfN6Mj4daJONbWJsbY/YkWjL3DQx/7odDqs75hTiYQa00ApJme6pnZTqr2WzjW1uLBe5bHUA/OBqvYv+YdTzZHcb9aWK2MTGiLMx7vyGhN0MSx/TB2XazIi0nfIyzuMtgaKULFGOW9bZGfjiKu91jxQtj39I5Hyab4yLUo1OQdK5i9vYvDtKnrAe5jP3660jpRvD6Dt4/35ymcHPTfUhUVW93SpgbdHUaP++/TR/PtrKbtkTf1oeGMRatLVLaZxdag4YDGb9Oi6en6Wbs4FE6AMVptP6n17fRwtNfxUVSkDyYn1D5gXagYiqKt5VH61i1SF2zcAAl/ptLl61qmvoeAVgd7z+aWGx3RQwqYhA8kn/p6z/yXbQQOWLf2ru5eqo4eY18+PVT7hr2rfje4QCFCAmEux4OgwNhPhfNMZSyRZ1EEVTEyLF6d8mOXOQQZKdMYRaQ0vfreQIw+wH0T54u+3YOxgv9Xy9B9VRpF6qJx4Po7tKYbJOa5bNTSHYZBarBZHq+G7PbTAYmXntJaj0STVMsbWi5rXqin7FTb+iUvhQY0i4y/I21DaVv9QWht6qGLBuXkAVYCfIda1DT8FXynJ10YsCjL6/YeYlYRa3yFkBYa2vyw1mP0v75MkMuETUqwUNe+CmnHfCYXNhepoUSDHmjC/DPKUsaQrTyOOFDSFhHWEQoby4cZXOJyeNpC2eL4Wa0jG3uJkfAOjTEmw04+qS+KP61WdWhV/lXGcqkzwGpcNQp0yjlnmItkhcBrmFWRPS85eEDBhqcf/iicmo05j/ObL0OYUzojOFll0Cze/huY5kOeKYKLTM887PxBzWJTE6HNvNAaSqCO78qmpVcJOcLzZFRij3z4kAXMSAmYMQUs5V2InGNkyIT1IDalw92N2ZoCtXfsOxPZ+rEns0KgNZbucHMkMfQn3GqkzHBLIeAEmxJrsJ3HSofxDyybDH6NPxbZDKMsKRexOnG0qUS/eyilb4FmPKdFFwGuet014RJXS4LN5l+nT4b+KdUNF5XciCnsq/UPqXVnDrCUedBcOtXR3XUjfwMQPpXKV3x0mp/X6h/G15bFTickfYNmIP23Vrso7cxRD8HaT9WEJTVU4GHLKvMXuSPNzprTMG8b8zUab9ifZ0XsN/kQEzAJIW9aJxTML1MYz6G1Kx53dNEMoTPkM0AgEp63AxPhcdGqr3Q6GQacroNWbTEwR8FiakA5jPHyjYmAJJQFpOAlU/6eLG23GKFNXfI6h4DQdzTiEPWduuuGhDKao+aTJ3Am6A2hdCfzZboRyeDxKDngZtK38wSDlShNQ2D7QehxrNnrpRy82lc8fTZO2ccw/U7ztlfkgqfGTg9iC4pf5ZlaXuORLobUVCET4022jHhGA1anefZDzJHaM60+I7JY6Wk9WOtEZ2yq4relOgjQZF2fmjQ+w1QHVsIOW/K2c85U2yw2A5Y6PqeBvlZ5lmAmHD/j0DEAIrd9rTfPN+HlZw0CVDxqCBzJRfKCHilk6pk2gJ0RcxwTret8Q7LohegvPlZDzoqXqQ+rEcM21oRBSQm5hHp06DENWtWA0VJDMG8aV68nvdGnHjmT7Whf3zgib1J5fb5arIQb56mRbN6IYyT84snfkGvY9HNNeS5hzMbRttrqjOzj9s8A2M3bk6MeYpLGZwGudgLagPe8PA7LQtWJFQ8v90gQmlU29pwzW4Jn6g9rBIYzrXkDy+G47fbPF9+umQyTWaaGqfR00yMnAgrCm4UHX9LJllI2nk7hKWNGMSYaDYBHkF1DDOAiy6Gm/QewBrkHCX7dEYJ+gBaSXw6mswxb/RyNWfVz+B/wY4+tRynZytG/zzYjRO4fMbfn87zpaO7muamAuhmVkzsK50L31gr+EfSl+HMoYjpxnZ2ED7GUVEcUqy5jn7d9slhYOzNeoYQJYgAVKlIGzJ/Y7aoVQQj/NUDYsmqY/nXAYQUArq3luAMkxZU9WOEz1IqrOA29LLZVFa9T6/leFSwhQni6jkOFyNWEHiraUoW2D6YBk25xF7tEsTzdWhBRxST4i3da9pPfITCy1+HbrC959wY/h2KNbVR8mCDeBXDFFzGKyYEAkHQY2+4DgssPmgJ02Za2kBuhEIROljlnFVQz0OnIxwn1eWd0FHlKZdMoFDl35LraQZGA04sznzTzI0hMxxj2NoUo8/0+vLBm3y1A1FgTojyrvouBXvyr7ZHQjLiN+t835pfjqfCyaqQ9A4I18eo7FRXfML/X96AiGArBEUk/4Hf+IYYWyjM/NDQQ9aqmE1tJaecISJ8D5TjPjI1StJW+5w2697+9+tafgokvIadarp+j+s30nsZoJqjDRo9GhcN0jM0Ovd1AXAqS0RsQvKohCRvcS01k4rnhD/O9TfKm3wFlCGooZcNsBoMZpD4IfC7atfLiJd6FJalMVShWyltYyPUYX6nhdu/hKVm31W+zpQ9vvM19wK9VNCPlABm3x6r/gespNlWwMfNTqdhKWL64CC2yVimgdmaXZSfgJarfnstunB2mkDRYiVe/Wmu26GVThd7kPa1q7Sx0pJryMnFg6Uj3fCnxxYfFzTLd/cozjAAD0AK1QYozqkQqG3mYRJR1WHptl7m5k+gGX/5pRqA7JFGrjN9e68a/c9+3/jQfOa4xh3mQrv8c2PrLaT01rYoPzE6TA2/ec+wThYx2EucHmvG66LfPpav87wQPddVbATrhN/BI1Ga0HTx73ddppBfxP+H3Ki0TF2MxD5iDiDogktkjcrCwUoI/InA8sgx/tcLWyXdbIeQCwlmKqFOZokpSKmqS9zMRO+CYb+FwSKevX2dezRKQ0GYq128MbXubookyEHEru5D8fLVHIauF9F2vsPa/xsTQkhzjf7tgIgbD6AGWR3I34Ln1fYoR6AHQt6UzfuYqkmKUg+Z2Tt/xzJHukOLiQxAoto5deGB/nUqYqEo22KN6HJLC1uwqHC5f+9RyukDLWTT0L2gU7SkhWUunYz5rUxoAWYSOx85KCmKvyz15ijGNoYNScqlGQdRmk78fH9aDLj0kY4iIpB5DmulpNt03vNDSsqNQc44LeOm/XAODvIWm1BM4DfcC+el0u33IS3crs5+HXyGP9sxg2YYi59SXojAyFARbUJ8BCrSu+1QzbApUo5XjMpnr/xv7mt4NGftw79F51SSiFfvSw4p0qLw+PMEPk7oM0tmoVNvS4AQhFHTSrEA3NdlPm1ytkrCVQhcKM57F6iLhCtCq6yK5VykvXSLLAmmtTaRa5PtXlExAXuHpn6SD4nYJdMyyP8kNG3IsVU5fiCbwOWGDs/om0iQm+aJrYN81BtpoLXshpsYahUtzFxwc42AzUclATZmOavaD97TQ67vKMH3+/Qj/qBZ8w7So+RX5r9TKEW3x7RfGkPwVXmW9WOk0GabVe6dUZQwnbTfxlaH16Kp+Odxn8zIlN+D6uQTg1G+Cx0y1Mm8VYez5klJK+iQk/hi/zaytL0wvVuY26ZUcIjpMf2CZKZUm7raQlVIsH6kmIHz92Q+VnKs5C27qCRpJX2x0eQlKR04nMlZqRHdJHO7k+Asfc64lt4b3LzolUWyhjTi4Fj+QiCYMd7LozNzytpXBEDco52rzhAkmgEUVgotI8WsG7XJBIy9bpvNDKo43X5RfCxG9mCu1Yu5MBVs6YLghrTTStYO+A9R9sTA6h4JLIOepnxrTiC6wCyZSf4VuT7GGUI1RttcdweiralYguQzNB0ll0Wr6AhG2rVPk969OaxmX9YUtGC8S9AR/7zmyndSyxyjrosibd46t9Wihj4bRGuzDRqpWV/F3DiLkRwYR++iA9Z8Hx0wpKWJEYuEVz2swS8CetW1VVaRMOmJLdVii+NRQv836I/Yu7ocxO4GUIRTkERzXc2gbWBjEkZv4HcdXNyTgEMMsEWZqTyVc2u24ca04SPsD/H1lrhjO1pf02605i0Un3tpbYa6M6VCCxnZFs59hDHZzszSNtWbCIuxa3agQuaMEBU3Yr0BqQevp1sgvUHRPJaHvvKcKXZ9CjT6/BQ4m2NcaVo4WyS7Z6NGQleJ/EHA30zyOL9PrTB9BEEHvspzT5xm46gCy6I6n5UJsrbrKn2bkcJ++H3bu229R1meCpkaW9O4nqmUBDxFxuH5jNQckj8GkjyqzzO1zXqtURfBHyLZaOLKT5HSVJIMIQ0nDSqZ3bMfjXduqXzFibFHMfAYqKxCpxsCCgd301J5QUYfIkAA2ANfgBPxgppRFClH9JpRkMN+S1iZCRrtpXnPsKphWrU8wMA7ZlHCdDQHh282c4Nh3gjKPSKyUX94QanfIFiFWie87EXOIC0GaXVFSdqbDvpsGJC6sfKryeMZ3Q93rN+5+Kw+qNzHFhrGhmfmJDFN/pAiDi98dzUFI9zz2Bwv0kgB02K2W6zIK9M8ws8WbizuEsZpBtuJ/fs3hmhN98GOnpdqPI8R2a5VT7GoR9+b9bkWTuuR8P9OjxmzYuNc/ayMqBFLOJE0FV+dGDuevqbMhpTE/ljCkzlihB9oGHFJ6kXojrU6F+gcnsLLWk9k2bdEjenEAVyO9Jo7obyTeEXXrc75hzzkSin53iFZBNMTNrypXSwNlCECSEiRTegHnJ1HuDq/aPtEcH06L6No9Bt5zBGjH0JPzkSifP8GVetQBwQoDFRRzftnLWxC9N8cg/Gs4WNcA8Z2peb2/TSVhKjNGkhNsAqApJC+vNHk/7qnyspxtxHGgk70Zl+CpYfHrLf7jKPAWIsUQ4kkUzCWyrQpW10gyWZTT7K3j1z+0OfSS+W9Pksy/KSnlrAZlfmb+TIub/BG2r/UWk0z6UBU3soCcycJVNzxBOEhCKnQRBQmupAA/z0ku+04Lw/dCpMM519GS/j9DHXKofh/J2vCmClA2jNNjxj/tBoZGHl9vy9JZMjg0JnWc8CIPiPFS6mRhYGGjOsND+Ob387CWJjKXwZiwnIuXpiR+MZJCSOAdcSqjE6EBEXF8FBHggAgs4xbqNAAeL1dOAx0rI9CMYoWp66fYmvhqORKs+J7hiRIDzN5JDy1Vj46Dx/56jwOAdJ44vxfEq4eI/+nny9euK1WfAc6dXXNEzAHoX1lCAQZUdREn1TcT00P6tv0isd646UtsRWMhgl1vihdMYwPa3LHHE3JNHps7R/q7/f3nLaR+hw92z4Ghi5tCMPhN/FIoOd56qretpsvG2ARd6sWct5ik1I474PFIrwI/gWWT9zda14+6+zTLDRZkKSWhwzIy05i1qm5EQZFHNM9oABaBTjN+QReQAUecrZQz3GHTcjh7VbrjaVY2VJk5K2LU7bitpjh8NsUm5IGTjPDRKSQ4gfylF1vBOeG9NCrKBfx5W2gnmGHgwAeOgA4o3KTH+8WnIpW6rn1Le64jTgqNG9qsoCSesBeagLYRH6KjPI2OMmZxnmE3COg5ZwQURTiBGEgGImcorTgIKWVNJL89/g/yREjjWT1L+r4uTzUrcjfxZDMmCJ+/ZbqQa+JzoReYyR7eRUrg2zBl6da0wa8ke6KU9AELL9fe91tB0nGg2CKWstBYksHm+HQDZXtpYYtV1kLPmBPSiQYy/zkL9gJ0k6GtLkOlXmkw9+v9SRHZvrlxu5aK+Q5yWo1RhBmlAeEuwhAyGadzXzObrbum2EMkXVCYlMZ6xanHyMNXueIfod+KKFw8dmE53hLMMmBN0kSQVrxFST4ctXK/Yg/JX0OCjiOxSXWteApDx8sXFf3zTSINJePDD0JE2VGQY487qiWoDefaTVEzZv6brSVqxtmTs7r8TkB1uFbEfyuGbFpWdq80lEOKY4itKIs0HQ3CTYzZ8rEbIbDI9e1Pv8WhG+5jJpIfAZggKEX2MeLq1gbZxVUJhNDABbfs42FpfaUBYwthcAjcLs+cV1UKmLCWmn+GgIyadbmvwUyr46toBHfAiRrVSaSnWIdtG8pZMbQcEalTwhfVL+IZBdYQ5PzDdVnP2K3xHONNH8G525afe4nY9Io1LTnGahJ5e5c0owzd4pvOdK9yxksa7mN6vKRhxsfT9ZYVp1n1LVjWyvyT9S5LN4AZN2Z49ovp2rPmMKtTscasuBsu1KlLC0SJG9JIssfkEgpqYFgkLgtNviXMA3C7VFK6kII3HDTiWBnaRohYsDdIilQvBhZLfiGLzWr2fojMCtb2v50M2gKdpRSZvTWLUKhic5xQHsrQmVUtNQ3TYPL5DGy9A48VFMvLGZ462v3HJEyEIG9Z6sgTjBk58SbGyWfNuaAGQN880LQ64YVF3lKRlt9+LQQLirdbydwYfSA1PzGWUbo/vcNJPQdz19AMd61D5A7jVay/LZ3kAELdOU51TPa7/ogKRYsb5BNJtuTQEeWA2ladaTZjAozrJljnXjuJ21ZCKZaQHM0rNXkK5niYyGGfhJbGZv/cSqPpuqKa054HUr9HvlTDvTgWZzt5ZQJSlgz1oCqIL/mTTNYT65Bs9u+F4YAUdWPfXQGDpA46Q3s3q3JqODQS9SDj2uFydfjrxFI26h/Ptq+aHQgYagBfKOaMQmlu7WURobNZuh9K9AaSe5ZMoiPEne9U1L8HVivYsmFDGH8LT9nx6todKdpRsQgydmfDQhVS5ULEsfjUQgfyUBDx7I/dgf3vCY07pysmtJqiuCInBq3Nm2BuMLvBEn2hoRSbOT9Nq8K7M58uJjOqmkzWbGG7lm+Ld+YFyUo8XB4S4Fx1u/yRQTQHx2XgX0Hl25YMV0wnkJx26xGJvOMCSFX7ydiRHYzDLVlqe0IelMQ3GgruWZouET/3htViLhMw9F+qilEKXzvL31JDXTNjVFCjKwq3KSdTjqZgZnA4flXYyd2M8rciDw9rM8eW+TLEX82TLvI5OmMoZl6vyig/rdfirdB5HlJj074DCSROaqAQSV3N62/O2UBE/dkM45qrMKLV49WgQteUQoerqtEEn6zjIFSkjxNz29JoFf4gHwcakCjOmItoJnaHsBxJ5YQEDZ0yceIS5TlIXNVVw2zICckkxNMBGT4pcMAtr58ioGisS6sUQOc7EnYHp/gOQyapJbD7TwPzD0r8oqtl6mx4vQabVxU4u48ttt3C91UBfrxVBzksHwKBeEsECRLjKLA+ppI0Fni3mrD7MYO0D0sS0wbxXxDvEjPrqtoUXOb2Kqb+7i5mm1W4r1j8JpP35RwU2eHZXLpIPRLMUp+CQu59TlvqNGLmFWIcupuKrqUt5GS3MClZS8NBQVqRRbuShHcFxQKE/bO6Dd+kKcJQ1X09otFyn67Lzcf9mGFG7C4UpmyrmUN/SbSnaM0UxRhk0faP7Kpqcct1edn72cO9/rWOCTl5UO2VTNyvT+Qq+j7baT2kYB7/hSn22irndQwLLiCviQM/ciAKOHT8SgplufD1QFgaclC3hZ8Byb9w+ypgHm9try+I/nbytleZ6Sd33vZLcnPRk+gnDdJhjqmtcCTvLC3+zEuVeqg5sw5ZG4vJ1Jo8/GZH4EuaNAaSR2ircwUGsW6ta/j2xbNURYfLcTwG9Vc/LyFl9CVVhcpDlfQA3UgB9In6clqGGqtJcLXG3zKViZEQ0RUvRWiUwodLdEfbJy4F0IAZ9X4Hpjo42uFIjJYzrjpwszCTZAekH7BNi7D2T+Pf0ezQTK9oUkVRvwphicD22zqiegV+Or4jnXjqpya454zliZ70uOdc440h2AAGAp353ICP6leds0bWBe2zCUfdJ+X0QHzUk3fZWlix4TW5trUuTIK/aSp2f1xincaP8xPLabiqA+ahy74GF4TwaRrFT55XXlgBXrJA7WzY9AHmb3FLFRwFwXHvWB41gJrD2WlksJ5SU3veIgP7YRPvwIuC4XMB+1IKbc1K7tKkaTa2GlL1n4NjPJagBUz3HIJaxvPWzwLrhOnNBYXZQREe+TtNr2iD83NPPMs2D+EmoEFiin4+nQVsUnIU70aIcsRZ+D7PMjjyXf9sGLvWEt3QPIN9VKqZc4sO0qZXVWhJPvxjp7e5zpGlyLev9Z6E8bX9hOv7N/dDqp6fZzQIpq+G6gW61iJo0v4lkYLe/UuR3x1ybisiDGAIbxiJraR1EK6e4lCKDv807+xfHwGJfv2EB7DH3H0mQgVaVpGJwlegBcS+RC08zfLPrhq718Nt0zZTPXW78FXgkJsXJ3pbw9fBum4AokacF0f5v515ijQCI+6TzyMGJk6j5g1NwsZzfXNG6pPXEJOJnPt+hnLLlA48sNPjtOdt/yLW8yxOjKbq65V3d4JnERKi4N9TspLlStR9l+AhyZbTnKHG9rPCqBF7BqDDQTGteR31cb+GXvhoEXhNXRRq883+sZg+aLxpI+D5eTNh6OdH9BxqjgT0eWTdF6Q2dJ2CZ5n/QtN2hnu1ijER4onCARQtbwYNDRrIJIk1ynekP4oBjobOv0M6feEfBhKD2LZt4g+K+zwx7HKikfmQ1BqATxMoBNPcmYbuGmg9Sk3b//gwudfoYAR6UwiEAawnZbwdLqNmRh6MHiYZF6DHlWK1yMi+9gYBkK6/NL6585Dg0ZUqLfhMexMwQ1hRPUFnvNyf7pNi1e6azTT6Qplv3P5ZLeMDroTmzoX3gs1UZoaqHMolFxxSSGOrfny+JkoKAjsyco6jGOX1w2ISmrJmnut67Hnb0ygbixMwkHDlTmBZ/zU0NcFKaoQ8w0COGPzJPMppGaTWrVRa9qaN7UhUlim89kkk3mKf/HS8MP9tjRvSc1RwOdREFQgC0iuoFPTV8Wp9Jx47La7mP2sSRnCC/P7tboLeKcFxi6Dtx/rEsqkWVkAPJlUytkr5zrzjXa8rTlgDLYEOQYVjvrMzaPQuX0vMqzEEMKRUYFwsychgtvZaSilHjQvMr/kHOi0qodEONpunYp9Ct0probI8lTJem8j0Ld+xYXLh0o0AN9+18T0lsV/c5vWqJLHv5wv4e3ycyL3aNjOp/Akqb9OXOIWJ7Uziwn7k8BJ30VVZyywWP8mAQUW4Rr3lKmCkxzC7bAWdXc4djvfQzPtt3gK9WwEtg2WsKEiNOB2xIEUpCFCTvAS4/B6d73NV/r7LldK2c21wFXwZXlQHmE0h6CLmvDJDc0tozcXdMghVLO6PwBrmHCdfekRDvtuZl3ag57U6sljhJ8gUOYCxcHNUNm5qKUV2+pR4GXvHppZ26qEnFJoK/HzkMrtoCCZ4q64QxRfgVpZ6uDRijT44B5n85+i9O71Qc79HXz4J1ezj53Y3tzsrmGBdIci4mWakH4C6QbFWzMKngWc3on1oU8dObtCoIa1tpmzZ15E6oKkX+cuj9cC9Hf92+y1I/XyYCpm+BDggXr5PwfoCq7VDyBetk3p0OTxD5hmK5Bht97qCDkRdMQE7r8ZWPZFncLgAAKfQBLINshsH7d8/I1i0N3YYwVr19DVdXq54y29U3Lu+K+CelqGqsqz64tcRlZ8z+SaaAqvGDfkTe/XeZPYz/Ec0oZ13AJleFCJwnrcrKjxpdO/fi1EfyxcHjNZmdA4mx1AAmznazAjCRiNPd90h6K4WR1qlWNWAbp61TfN4igJbYlTBLPfWMgPS/R7RlNO0yuGYiGZ96EYEzdUa3HXoy1dbuFrM+Fzkc8lzxsdifpx8+yXMqm7qL2A38vCGznxT1GZJD3tIroAz75YiJnl4sF1h7snRRccBYP4cuyURa1XPKk6Fw85UdkU23VOAljYde9QvKgntCi+Ws4j0/6GG0RlVTA+RcvPy5tmVQbNLgbhPaeJztGizCqlLzCfoHvbv4e1jUgAN8j7Ejh/vJOsiy6Gd4ubCQ0inIrJdKXYMvoRtDQ+rWz4WY2e+YP6RjbeKXt9mZRMqcu5VabK9Zo0xJwH4QkX8w51Be/so/C5GmL6LbmhQ4Wdz0dQzclqosbUhIBzoaFDNkobqjyh86s2mLMianxc656T/xBCzToVhnpydz3IzZbc/xj4SBWAf6Ep7FGfwyL7Yc3XkXOThoHhREqAM4D+WnnNCBRw7kKDJnalMWovpk3ioubTait5LQ0mZVWH9qXGNFUh4LFtRUUe+IaOXVocuTM2fOYLfXsSSoF0cdxo79KhkkM2bAkLz94NnIL0WsTzmXj2SVX8InbDjD2npxdtKsr9dcvJeSMtdgzRMrWXl0jJ7wVU+l4m2lMyKs1nfxxybTmVd63ApSA3mGkZ7XQCfd0KuZAAoyzDqjoQADBzGeXgPwosSJhDpEQMSffQTvn78hAPDFxO3n5S2zNc5iyMSWv9tjdY1gP/lj1oNRvD9DYtJwGwwe0ber9Wff4PIkAM7+frJYFT9xwa2XE8+1FS9xH3Eyu/OvoNPtmB0ZAVFdA/a50+blqRZL2nSfAX7Uioqsl41SfkR0jfZXrPgcFWUwbv3L2Fm4Ibove4Fii2xRB1FcYCN3oDV8lLtP+sqCdk2koP81CK3qeWxhGZkZ3bw+oH/pOGDJO812G/P5RD1BvMonT4LCmvgwx8hJCvTtlBlH2X4fteUtS4ZN7AgzjoMMd5FpFxV93hVwk1gYoE0pbxt+FzBvEjMYKtotwyIAycsGiy7dWaxiqov0BAs2Uz1XbkjSUv+w5aoZYqVXDuWQxcTMhILmffgR/j7ecnTbA96NJmIsPCvFCD9HGDsbCJIxUONvJn97ZJv5yF/BgvWQs0nSw/SYIg+l1HjxgOEvDJI/ddTgjOm4Ijx5xtzQrTka/UK4hMcaXTJ2S6QF5ri+UHJALNVYnXwXx/6Uh+QTKSDqma28FEZAFIgNZcRN8b+G/YTeA8j85kt9pS3cIv4D68r9m5rxMI/ffW3ICiv0a4crqOFyoV+g/y7OEGJekteO0GutF1H3z/9j2ZJ+VmjPBZk9nUdXANnloLc/6FbZnoTSi8RCUTFBzrErr1I02p/GGxrB82crXDc0prVFt2RMG4cgarBpUcIOmEFuaSh8F9aCD4v/VikPZiia2V0N+PIomUymcLet0hOxroeSoRxbJtkhKv8m53WiIJ87SmuaI/BTGWm5H6P9VvAjaUMJiqAoEV2Nd8AtxuH/0p89G22QZb5VgxLqKzZxg0huLPRFc6VjjbuFWjTHo4ReaSFhRs4XvPXdIYw4i09xnlgNnT+63Xx+zy+i+twlOnCvvWRFuecP+HoqNH0D/GwA/iFA1yINsTiyZN1TLVSp5Ze50hJOlH7nIfEfYb7wJ175a3q/FLvStmJ30X0RBJ82qpR9igBG31qlsBTflxUXz8Gwfbrv/rMfJBNI/brPHWc2uTmWnPzV29QE6yhz38xH/TEekoPRKfgrT6Dqa280mjLneHGgiIQ2Vcy69mGkQjYyg4irqqa0HQsPxGcakQE7aa7rI3gKZ2XZx8Dcpf+Scb8SmdvUEfvzouj57JsPQETte61LoVKzvYKz8nxv4gJWOly2YzfiInF7NCQRYf4n2U6StiqtJxDuVbnju4T6cQ5aQM7tGwEJckxMnxHfnMxJEJ4tGJgJSfj/mWOLMkE0rc/fvmDs4nnbl7htUFtWtKqcOZWh+eKHuwv+QB2WYF6G5uXa7EsTYQch/wEnB/xt08HKwRQRDPEodAiRd+VwOh4GbCgamDdqLXaFNeEwCGqedEdskoR4GEY2b5WNNiAs4b7OxI8QcObXOfuEEf/NRjL2VkL9DOi6usP3q6d8N37SI0SzD4diP7S5GbXT15zzPc3mBhqCuMqHcgokSc/VhH2+7eXKdFazpwbN3DJT4tlF8Hzv/Z9kdIIxcX0hGdR4YbaDAd3ILk/G3ljnkU9hu47azghaBaerpZm0PPl/rTXWVaU8siGH6grmdW2Th7VTs8yVWn5UJF9Xb6q7gmdd7EaFYdsdL1KIol/L5hw7uhE+QBFDsh+BuVizYz8JLW4QUTI6sJHB9nr6XeW+QoX8J68CD1PMm359RrXukiDaQ2L9659LOOQguWjXIFRawulwvyMx2/3RmpDp74qTh1hHtmZO9wvdl4dQBf344Cl5mBMhnGnInJ1otNht7P/nB/wGTBb8hcgJxudFQhAJSbbl8IMULYxTrjYu41ooBAyWfssGvgwlfeOmGGWLsG6+YxgouiE4aeh7KntHxsx2rWaPmJUPKLg36zd4F++1UOsTJjJwjGOTkWnvSwaf2++9KUshkW4tFGst9N6YgOlFZo4B78teleL6wd8uNbr7ffAgQrhC3RoQ/WGZgqzOfAI4aBAZorz9jV7JzNjoUNhAhNRFzlYVwwD0ykZxSHiZT7qcBXfQZylCUQ6cQER/dKbaVfFXbABGJIy+aUJm8fdvbdhDl5gwLyhRv/6eQk4gK6hixx7QKto4B1ITnKXqltBVIvOhqFhLEb3qe5z2tQ60ehtMVWZMuQYQMl5Ti3MwIWoQWtFrAcn0bOa1CBf+TfKO2G/WgbHsUgcj0uMUO1Q90MxjferjHybHfTGq3vURfD773S2vRw6k+iEvvFH0uFwbswukDf4IbFkSIIgTJ1E+5M8jhZ6MlZZuM9bCEBQEPJEvYRDi7rO9aB0pEk8pVhtzVr1y9FBfaXmJBcHJSp4vjCH0JPglbcsyk2dgGhk2WOTuEI7EOAdH5KNTVn9FLT9KPcuHMVYhfm5VSBqdikwQ3IHb4o4rOHS9qNcMEE2Js371syejuQcZTt8lLaud8EhtFpDneZMYTyMb3puJ1c3HgQG0p8kS4Fa/7luqvCngp+JpKwWiMnBUGUIWIZTqO45+uDm7cMFVdZkw5Lc0DhL8t0eKl2USigp4XP6N6PMqssc/bd53BCLAOSISTGLkYzWMsUJhRbanSmy92hRg7piLByrJl1/qC8Z4lcfg7B+Dg6uOuJkEy87G+bzqSiD+qyqGfT6slZ80I4HFnFw6qPm2QIJMK8onJ+Iz8q/wwChTdpdpG0E5I9dkNhZ6jQuP62tc3354GHJmBhpSv08lfDU7wyD16P90583jvILhseNWXPSf3SvPDCWNOscSeg88ZRTEvQ5q7riYss58Avrc28kAarYSh2883Q8nns5KcwnS0wMphO19TCREcBytl2AaymtI6VK4gR+RKVjP5JBjltGQXpTrRXKO1mxrMxaOy0uovMWI0wTNZ/P53/fdvN72OSjUQgTtb5IYfl9rt28zudjvevpgH7wiLJolR2V01u9ZA0f0XXDlv8aelpNzioI3Q8frXcO27A7rX8DGQf41MQrDL2WiFr+wLBejL+DFKlWzO0P7+S/FRHjQS2j/DRhwqdJ8lubugJcTOFAw1eQgMsn63fKvW31NVAa3M9u6lwfH+p0nNJHpu/NxbIMtjbwIMJ3920ARgoK8d+j5g8pgFEUjRFCckHXF8jcFxuLMLhMoKXyQUj5SxgyXirNnOQZzPVvLW6aRKagkKo3nzd3reNBztvDrsDzgAx9HD9KmmYxm3YgXN6W1dPd7XzSr0JeJmG+hsk2EsZpZUCEij40Voif0kLDGwu+Ok+vr5sZynVXUghoPEN6Z0p5614r3M4uT9lshyJn/EySGC/YmDxm3s/TjYqHT6BoUGIUzxzAp2RE7ekNU6inIDrDB0S6mfdqz5oizGYonGcJDrMR8g3WmTpVNxiXmKIaIq1O7yihu1EqU/Xwp5ootSsPDziNjalhDJmBMnvP87GeTz3jnxtX7uuzjzuoehmjhWq/py5f7u5cFtjhWcfXCNezn4p2AAjKW1vT5wNvinjENOTY0ozzWwEaE2cJ712qUWau1RjrwpuTpU5014C+VWiGF9nSrPK+bV9+yIQH0KA2RlcPamZlq0CTdmvLqocXhOWEncQsaIpVEHNo0K5/gpgiQJdbP6BEo7QVZRhkY=
`pragma protect end_data_block
`pragma protect digest_block
54b456057b2619a537e34e1825859b63e1e4bb54889a5031fbabb1443f4667fb
`pragma protect end_digest_block
`pragma protect end_protected
