`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
hFw3YgF7lx1hQpltoN2jbmDDE5jfEVFUhNPATssehHysOu6gncJdIR3dw1qBPrd3pA05cMVOwgWHMI63GoE2rRLTlZWoF4k+InuesW8zJJeBkOgeCgQn/a8p9gPTTVEqVVjIHPZj9/y6A3mfOc6ebQ7suXA2jj4a2z7DiYNtp5MG6RJYRZyiAKfmSnY4FiiG1xWTTXua/GCn/Mtqs87A8trpGdlSnM3oiJfxbgjIyyjNcP7ndaCYllqHBEM1slYTfMRlkr3vVgPU8A9Rg0itoPbtjWHpCzYf82GHtMSyldsuDQyx6i8Hl2kpoGVkvnB59xkJOWjH20LMzgjOS0WSZ8a3AqtU9CAP8r2kHZx+TC/7VQdUAEBy538Zm5blX2ntyw5HdZRtW71/CE30LO2KSHU0z0q5KQfd97dsy0hmwLp6TC1ep00Gu1uiaGojTepVemiyXEmiPI2FS7CAVVYPjWj7uQpIMhX/6HLBRL2NEeH94j0A1uwvzE30d0O/jAkg+PMfT/W3N76xjDlplJVGzK3MqMgIkrg/gQN//9QnKAqkPFz4+S6c7vA4Dl2l0ynON/7Gtpsfh2OrOGAZyDX/F1W8tLlTG4SruqrXhac2e74mdf/KTnzqVv8YW1EGKsib03zuDD00SidZZ7gkLKTiQdywJulK+ZUt18i/6V3XCcDJfprmxyYCfVyQnee0FOAT2fv7REZsZDYx/J9++s/ba6VLwLRXXLtwCfgqAjlU+5HpNALqk25IEOYtwIjPgnBM5WhIZ8YNSiaTlr0c8kmYLQO4XpQjWHIvbIHTw6YTY5dR2DBXhWEdDmBZAP8x6BEIT/FOwmiYzjGzasA2JhJrohdAzsH5AyBG5SDWjrchwDVPffC/hvaN6V2pvjAFK4dzTrTz18pzO0txmwfbKPmCqS60EywgDU6jX6LU1nX+u126EHoxLcfrUrxSsTy1uwe+A3uUQsurDJTH/biDya77am3bnd3Bjk1wTEFWzZZ4owmZkpCbvTIIzH3/ZzLuAD9T//G+OmD3X9Q6Vtb8xhf+7AKtki5MYFr8qMMZ+w12AiQwaFMvSJbbgfMacb2iP2IXqqngrCevswZ5NQSlJo/rvMt/0buIpwDiUyekSu2lJ+lWJSCn53eOKCdSAlTuFOpWgY567cDlG4tqDHWRiAimenqsdcNbo8BXkyFXRrgfhdpQLJMD+4wBLfvNBC8rcK3dpQytGazoyTMnI7zTsAfC9yRDfBJN7b8T/RZArtWjzyV62w959oKTrtph8Eh3+yftBjWfAnOoOENMKxmTUCxM7KSzz2cHh23iGdNWcForOsQuOKKIn3Rjkb4s6P6/FxbB2HTvQpu1209AC2xh71rewIzsUo9JGa3JbRFw2zh2OothbKX1W8GDMAh+twhSyZp4L837cGlzYw9pZc/VTYbel9XgVrhRGhoTR7/RVyj7o2SJRhwgD7k3Obd8/9djh8R/MZrF1Gm8gVsQ/REaJA8pFgTGW61L29+VkfDwqHLENFNctDg1FZ9f8fi+t2sKFdTius4T7HAw2mgjCLIvr5gd+CzkumYqaPcNlfbtK9IAhe87w6b3JbXmc8/cQkLrTAEOdbX3GcsgTUqR+Tv+tX7vUy0D92pgcZZKGGGD699D8qdVgdLzid+iQylCEEiDWbd8sy6ds40s83HETmISc0SA82a35F8QQSOmKraXSk/beuAng7lq+0Honkr4Sjtu5h4vuLoGU5iMLm5hBD/U35AKMXzzNnZ+q0I8RlYHylGDtFhL6KZR0mgYRDk7ekhOGgZAFTAjD5ZroOP1Ux0BZzd8qZxCl456laqg2IDZeYYNV9AI3JIqtlR5fANOJYMW1pF9S4bi2gPFdXtnNAQU215iYCJyYsLSIACHgaY5kkC+vEOZ7fBfb8D7fX+HRkuekk5r9XOzZ4plS3hlKgLp8uszawQ0emzu9caujhfoZeXwo0GX5Vq31xhnZ94MjENg0YphjnahyAFHSnZ7eanvFLRx7d+2k+HXv/BdI3Ook/SCsFEmguGauBHo6Q+D7uSWWIyp2YIQUCizxwe6UKn5u7SZXzEUq6f3F0f68xZYPqFlAXx48UWeNxGjvPDE84CbvpXWPCmWD8HighUIja+hnUNiqBVDo/SLPQa3yE41ElNViVCUOtdm0RaMviNfDZDgYQ7ZJQjsGPE/CmuM7ine2tq84P/5iO/XChGRZRUd2/6JpZcFYJZ1dK972TILTtF5e2ZOmnsOu3AZL0o/uRriUnBct7y69hQGpkLO9AIR4pW1ZnYKhI4IRyTie4gFuTBJ6Xhgt27C6gdtarKG8elGKYp5tnlSrlFqRVGnXtgv0edVFeRAq15MvHikDwwGVNa2OQgRIXAEuIu8ZVvw9JYAuuefQ9Y0wh3P7Lq44aw8a0ntRRnHHfSz9KCfCSJJV8NhvaR2z4KX5QmJkA++UGmB20tYHuAg79D95QCkAFOUN1Yr2HxfPmR3wSeJfeqXc4CYzimVjRwDznNzZqe8Xqh/Z49RFbG20VyjsH1K4wJ8vpGPlzjqgsTrFRks56nfnnRqxqd434lI7mRxhfkZARWnxbu2t1XqBitihfIKarWHx/yJgByIPVD7OVTakaYt6HuJcIOJ6UqlQTqeMoUaj9lUxpT1pGlVJZ+o8FPpgpo1sn2Hx3KfzWgupEDuBS0ke7sBkg6tGXKY848tDpu4YElBejl4dAlQJGF86JStjw6FKDgXQSi7cy/cMfXWA39k2UeHL/oAxa5MHmlbkxEJJj+CqPkUaw9TS08SH7mOPDn1XUoxMlLkegjAJJWD0lydW4fkXbF6f1tdSSiAZIdczNaw/SCxCOo3megTUcDP54lc4pQ9mJ5CuT+Vjz2tkPqadf8vNh1scnFOipoY9ngP32EH/qSKQ9xOJt054KMKA8hy5fGZpex+m6mI7HvEaQA4nn4BrvlxsSKWH4OhPI6SuFlNivwTuFwvJ+YLJMKbMt3dwQK3rV+xp0mLE+ttcJ3EGwmdrPyMma7+y3OKQps+gkN9FGynSJqDRL9EXBULsQtASAqQPoQssrwtmd/ZFQv4wYYObnDvLaKozfC2JlnhlnmZa7Z7I9McWwIjFHpbRVdvWgd3kEVwwbzm8vl/NikCPFiyj21Yio+rAZmBDbdc8+mpa8U1GBzi9GN+YsnAdRq2xV7ObI27tENhV7cFcZWN4/OvL1oAYsVsgW4Xn+6NIm7hm/piLKVKYtO/dtzJ0BXPibffMlRifNIZ2yUEVvonsLWRExnGZiRz1ptDbFABxvan8IxiYC3Las2U5axgXba5v/gKbjn8W8n+P6Y/rLBT0IVFGV40sgdX49w+z+d5V3B62zldmNf8/5vJ71WsCIbeyYJgZSPpcTF5+dXOwUc0+8vgFQL0VN0RKd2gBT2YPFFq4/HvrpUPf1N21FxbNlDJ0fkg0Ip5mTTklV4AvbhnMb4XHrqV6XWun3vsLvQ0rKIFckOmNY8azKmr/WFIjebQ3iM3iqW9mkFUhGe2IMO7Yi7puFb2A8co7P5R6BXfFz9PoYiS8ah+fGNtD22bX0eBFfTKNAMWP1kGDUDyQAO1QV439kaeJDJJ2ARC7to8oAXYGuu017h+2zSswFZTz94lQ4ZD9mzsx+Us8HZfE3hRSbDVYv0FL9Zw1fZcDT4SF5rp1219hOjWmqUtBeizLYq8euWu2S8pI75VBu8Veyqjp2OTnrUw4SDP6zpjY1RTKa/2f1rjWyNE7fgrwhPzPixvYSprO5JeNTI5HEURdKiTSf9a3ZQOkCnVblTm7puevjPScDV3XJ2LE78w2ChremrQpos8WfiHBa2pFkKGyjYl4YgtEXqF8nckDgGQHoXPLh3/uACrdCWaRdkDTdOGmkXc3Sp7f/9ZGmnYmI6jcOoxnFIvxycDPrWkctM7Fn/rSR+G+gmCBGGyqiH/5dftQ0NN8flbLbfS9l+dKeCKCZYuhLFk8y5j+9vpgxMxxgs5apcyAEBe07/a9S1v/xuMBZaJMnaEcrQvnt6kk48Fs326B5UZWriNnJmMtYk+4QjbSFPLtD7lhK5feIxtUW4sdX8QutmU8eyKQds9MOeb/UxfbpMqf0VgciRHStU6Ad2w2STP02qtPTsDyUZ7A3bekqJ0ezR0L2em5oYXnqSHNtgJRk/KQlYjVZVtU8Z/5DrbJ2xq6LJhPzmqAf/WwhGwcRVelqkeQsf+AiV7PbkolOqJmflqOdwB1XeLEjgH3ia/0cn3+I9OuOKOR/MNTGJ/jQ7W4CMrFliGyFhRSx7Wq0hCapceH4B9+ch6GtCGaX842dib8NUWIbNo3ooKmlIZwc9vHulVCVy+W9kGEoeERY97lqRx86jAl0ggCLsPPQt4WoaNM8zBFe9uv1E2/5y2ZedDD8o8Hd9tx9ncpCpBBLv29mwNhHchbZw5gBR1oai8EALqWV29qqmEMK2XxFacuyfBFhLmQ5ziM1cHt74Kq7gGfTAgh7SG+2MN9lT72/QC8Fdq+sdNsQk/vM7/RKyds6wT5QRd9/wwNH51Y3h3Ovq6UbjQi7sP9eupm6K3AISR+fioJSz047dccwkgDmU0DvE0y0BRuI0sGL1FjTNaIZOWQGj2RzdJcKoX1nMkJA88v+O1CFgSgjAuxIP94Grzwid0V7K+rGfKjg3dn7K5WlNJ2uGPPscaR7yJgAmU7hg8zJpNLHTcMWIhqaLai7771VVyUceO/ykr3MqUyzPsy9nQBS9MWkR2QqMAkAW3vUWdbTEcORJGLd+m8cTovCJ31pi67Hba5d2/rEsuRUC83osbT44GJvyRo/g1rw6wN3pD/ZMO1BVOoSl41ModeGSgiAnIaW4g/JaBZOR+mKaxeIEIcOPvpN3L5JF8jjhsiEIm5pjXZ4zgVNcxh6NdzqDmMbQHCApvxfy9ZIIwsTfwEdDjeigIqO99pnOJpwXJ3Og1RiZ2zZJ5fmzPEQ9SlxKF+pLIEKvf9qKprd3Z+hNkHPcrM1rlMvT6VRr+xFUY6RVdGB0m3+MN0YdWASHUoKJ5+43zdxP7JNX35U31Y4DrbI6std8UbFln/0ghQczabyX+TBw3ToY4GyGKS6tdUN6P1EQ9J1dmuUkFORybwgqdGmLfNgwgj2rpSm3tIpVvK6UD8wQE2b7VdAs97lORYvPzLAFujiex4WeAe8MfZHnnhLTcicAcipovAv9I2n9LtwAPcYkvUsZYI2ivbxSfqDdgp7AWO5/aw3mVNO9MSZSfGooFHBLW9tOeIq9je79c37vd63joqjnJZn4HCPT3dYD75R/dXQwtoq0kOr+BJ5hBpWMTKpVeHUxfiNrCBnHBQoOx8nWciLo/vUQNdy6yX+leSJ+SsyZZVUc6athJ3OUrq7ydwXpdvW7joybNnPDCapmT17Ua+2NYn5+MESneRc6PTaE19jlTXFgfHKrZzjd5RWjHVtu+Tz6tSj9V8hCjQJDadcxYEVo25u1mIjfIKLbz9HUZmr2T/U2YrAhoZd4k59l2CXi3EpMgQx+rUQgkloWXsEqzObCtMvDmoBSD8grVO3pO17kLW+WW+0h39d3gIslr0t9M2ZUqQ22pHZ7M0NbfE4hzYgQL1wvSEjF18Sqkr/eSDbiHrSSSjahCGgNg86IDHpfD1k8/++jRrvrC0XZvnkpBp4QgoE5rmCgRZZkv6Veqli0qD8cQkMpya29z3iQFoA/GvxbC/9FfgQOXw7Ao5g979+Urg/v/zwLW3neMa11pi1d4ZLey9grXQpXfSjBC9DHi6kcl1vfh2bK7UuqDrxF207KconjD9nvlete67R/TDjmgFCjFXauq6htngY5KRedIg32yJbz8fT0Vk+OohHqdtIv4hHSOkcsedDiJGW6LNfZRNqiKuLBaDyPHwrmsxJ52FVQzL5gWgAvWM4kT7T9T8OQCvXjOvTlE1vlGyAYQX1cHV5zLFlqnS+TaQR/ojCNPfcMEd7U1JR4IWR3qF8O7BYshHv0VJv3BASm9cxS2OLdkfijFykCcbMVFyjCcHFxwQffWj0rh4yKc0qJBwT5HrRbuAimMLxmMYJDeNNRK08K77DWMVjOYFc/0/kS0ik3Pedj7qStGijSlHedVTuTvEOvriiUaKUpA7y6NRKJkiTtcEbMtmCqMkuV1sq89cm2ZXhlz9Ap5fsWP+j1Sg1N5ojR28yzf3VVlnYDK+DdaHNFVTByO7mLhcuaOSBfNdiIBNw9K/lQvtqo4+FgTjTNJzwMvdLWyTDrpmD9mt3u2Ks8BtPnzZCqL+oX50XP1WkzMF4O/ZGlw/SdIq+9Fo/qKK7kUXs5CTigRB2qo/bSuJ/hOO+TGf1tWRdd+aK8ueIvZtoh+z0F2xw/p6g2GyNDAfIZ+DySfj3CknVl5bP5Zg6rAw8lZruo9KX5qAZaAEC5+uj6AvmjYy6j5YFRcUr+kpcZa7TTFUw1Mi9KvGLe1iVJF4CFtTFiFB2OgJwK/dDVXnFVWP2WDkMXFyEpTwICO6LK6Fky/Jnidmycm3ymWS2msSNweMTwNY8dQISH0xVkSQYeB7Y/swwVFl0Fjc2oEyBQBIuLVkQxHesbQgp4vV7JO3iA8qUWUGLt++Dn0W/9ImOHRv7FypI8LKo0Mw+lJDUTTI/2lG8+q/tniArJknfEaMEJbk/BhbBw53nL5PXec7tV41W9ZWW1yi1udY0NM6M6G4YeFSkCFn6VLKNaHsOT8QZpkuSyQzFxpy1SS4xlobVceSKaT2txho4nOZFXY8yJEH5ao1bjix99QMPendgBir7pku0LB2wPuXe2KqYkhhGUPvF3IKLlQoibn5aGRMRVLmrXsOs61rDpcBvipL+3cP5KQ3V7P6PbQwDVC3LRj8/KYInn/PvGXc+Kn4mBvJfCwaPcX0nuBJBDbFzZVvI8Db9Idp18bofbZDpTAEZxXryQJHaqBts1FynmGTyenSKnIuWu2Xo8ULp14rcnmWw2kFpwxW1uOxDetuEBGc4KeiSzcN9+NbV3reCyyxc8fTFhNc1JAkwx6XY7qkHHaYtIYgchUB7WBE2Bo1tPJhuOz7bdjdPr5puFz5oOYjW1FxPBvCnZ1x/t0D8WP+4biMW2kMeUyxKEZulYk7FlvlTYIvb/mQ6nPtgogQX5kg/2rooveFjnaX639Reud9JlL+RIikNOaHbl891ktNi+bH9tPYYGeMcs+Akyy4k9GorCCU+NOpfDz8THpPlVbq3PNigm9rPE5Nkh9lpEJz8Vo5lXGi4G47C1888qdj4xc6pb0cmMC7v6moqqSq6mUs8APTb71GEZAH3gxJeMKZstSXIXm2O2mBy8dgKI7vp1SkuBkhaMSh6gRBB5tQ1qq0WWW8gOASK+y1ag9PNYRjri1IsICbfPIWiM62ErI+R8YA5vfVk5vVIdqH+nWvQR9M6OfkRUDytbBumXy2pO/CBTYYViwLVCHUxiqPNT+HM3WssFKv3NS1Ul1OaK5G85CK8jOPWgqN+0Bs6LaflAlijjU/BHwfm1i8U2j1ykqjeZynNS/IW3Mw4FuRd9RVvh0QBh+ZRR4OD1guZ37OMyX1U9vn+cWrU5jD0Fk9sSlIEh7K/zgKnfxEaNuFa5axCT4zoBqWwqngo9YWXd4rqBZHRZ4wwyihhGn7knmlH1t3D6oC8L+WSmZ+Orlq4kIpjPcgUqfafoHTQjVjC+3fiiiJ6YFFIQROJCyYxT94Rx8xzdc0BdUJRYOTrq/6lheTDxbb5M6Ck8Ko5QHfK2lz+gz+4O8Gs25vGlYGicZxbnICR8ZzdItb/8IL0cu+uMmuBib1KUUxpF6umswoAkCYcSOQkspqTcfb/dqoWFlV/81o/De9+T/du1p4yXXSjOUTzBPKCNMNr5MAPT97rGuUn2IKh9Maeeq37nlMbbwk/ahp2SKJqaiN7GgMcohybb4qlAKTTf9aVDv+pEfM8UDRTNpBVL2rSVtVSuVWfsSH7/fW2Asc8MxaSAID52eLUOWn+DHJf46LaT7TRYsWF3spizIQ2vZmF7IMlqvXWLytvDOs5BftjaduEgFiqaDHyyIU8OwZss7DOisN00iqSYcY5WKYjANPlT2xSGKL7fBiEEQZ9zYFriEdDnVGu0cxZsAO4aDN/YW8S86z6OfenDU8I+a5nrB4/O66BrpCuYlWv8nqrSl3KNfZDe0uOm0tsAEw4On/PVXdnrBrGrpXh0R0n6+eikTPD0SDiqgnCsqfADYkbe8I8vgyL5Y88Fuo5yANIqyeuDWY9Ek+jJbjPWOkwEWW+UgSg1HpYvarsxPoDdo9Y9Oj5+CdpM46kq3NAfF7kHsSa91cQT1txOFw8iNF7BwIiI1YzlKKtXY0aUk36M/tFtEZcUWUWfHUG/u79V6B70dQ9b4ccCNVotuzU71p0iiX/ovAP8TbmaBaVqdvMjSEPotPy5FLPYnEsQ0UpIh+kZO9pD/UiYXAQGIlTf+YTGRj9GMx7d1soydV17UR3dyXUYifj6zh092TX72t7xEUF8IpWleEiLHGigw0BDn6w0eH4F0cx8hW8/krl47yQKuw2eROZ2/rYXHqy1EpzBygGCC5GrLUUDj/ojiaJxmFGl8qyIZClgFDedgyGA7LabLsTFkZDqJqxqvbImgmoBr9MDAcR9gBovbpQsO68Q+0uhIRZUhycduglcFm8CEFzbDFP2sbVP2H5tjQI3zoxCoQdD/aCzt+hexrC09QU/3NWqKOB1/qH6pOWy+tqBja8sBo3jDjh8EueeXi+Lsywnmg0urRggeFpJCJU9eLqL23N9ndxjtQBRK+5QtKiOmedY87Sbc99tpSWmNXjOpqMYuL1t8AIt8tV3yfemJO8u1Z3r2MW+tgIUjTUsea6+z7aAFIFwIqmsfCvbQGAlT3j2EJvt1tWFqrsWhBYDjigbiNv3/USl5mVrSkiNSKFzqhKHQFD6qzzxcvPKMnyVOD1nD2yDJg7+3PlXZOFLltNrei9yQ+LVMumdsoIOOXYV+rHxLFHoX0COVjTtu7uIcBESqLmL1IBK48eMVQX6EQaAgVpzrh8zl8vN1xa9KnMMd0kkY8WghmXcpM5hYUBtWlQD7qBXj5Y3ZAGfArVlMhGvw/qxIqEmJDmienJYe4agfSDu/gRkudQWaSFVX8+9CDE+gvVD/XQ9qFSMnDGI/GeM6/eILXb5KYIY+DeP/h0wQQ3PscfjZ5DIXUzJTALEkxYDtUNE1AftcuXcljcJLOegxotQ9erOAXCWaBBG5UaAT26dXCn4C4zY3/ATIO3Kq56JzirC6/aForEgV5nLmqF5kRDTob+H/0gsnoGBes7IEyu+vQcXCkP5EAC1w+B9vB16AbVj3Hfo9ErEUY8c/itxUwyOBdrRIAzsQhW35Y71e9AjBzKldbW+tCcrKijCxmH5tP/EzX+jbh2PcZ23+KJcJ3qwQIsZxcoW0/fy1vgSFNi+xk2xDYnLheIy4cRexvKAmsga+RbNATdMTtr3MkC5mWhd3DdvErkqujZksYogoStRQS6f/E/TJwHmtfI7XpbejA41C6AqwvdppaGIcrsCVByODIDcKepguzCVwagjwaJFFN3XKLQxNv4PIlK2fQq5aD8xGzCa5vo0A6bgKj6zEAvtr1VihUgzrJxHqfEanfmIVx9bZkei4kPKgcB79NkxH5DmmMBOHA/1eu7dMH4XTgENMoRUk41aF20zOka7A1FpaYaYFwp5kDW6RjMKb6qwwdaHTjgwe7Mvj1Zkg2pOvxVwVR6qstnlNdd8Bs6lu38qI5BGnuUPRntONWQ1pblDfwpPAIeMWozBRDtj/gUFYQpx3q4SYmgsVQcOT+JiILjzuvPzK6KpFFH05oStAYd/T8/znP80I8QJmGWW44UNZ021VBQEMZs3vKvcMg7rBuXkac3v3BCbNGpwm6nzsRPl4mCYkgf3x9++EZPSY1elO4ehvNfF5FI8TMXVuCkIV5U32vPigLVr6KQ2nvvAKor0jTvnPLGiVfmK0MxAR537E2Qks3mDeNbYHKpAmKiZg5vaGcDcKH+vR7fe0ja7Oant2MmzTcr9pwMr09EddoWMeBddovgjiRSmOHfIMu/dQSLz8vuR/n4G51DMbwbqgO2gkTJHSedAMy1HOrcr970yktgXAvDel1VRtCdoVexwaEWJNIBkLQOvtqzuLOKtC/8ih4qrAMl6g22UwIFYJB8xdm1htzXT2UmZv/rRGOwiIM7GUPaPyR2aSuV9eYM0d9R48kqdkzItEGo9Vyf86dqTN4LKYgm+xUJArEmM8FRoxDdlowooP+N0UiTkoGXk6o7fGOMAB+ZT0Mk+Sc2SmL0iUHqT3/Qsv8Kj81texJMDp3sYAaJBSIZPljZ3CmmM4S0CiMvadQs3dtYfv0AZD+XLM3zGZuD3QPH4Wzed3uc6RW7oqQJHygKdoTlAd7Uj5a9zgerxN5PDnZVIRjqKbKyFp/EVtUg2LuNGOHyX2FJ0gj8R2mwfFoa7ahJz05R+JhDxrmN0lq3M7LjHbIiTOM7JLA3/WTciOgseeHHwHfRuSNqOXoLhHk2qzhQtL7ESfvRUtEBRTxl9MVDnbEtop1NhBpFnYvAaTJkssZ/aB0PPyrsyXLNtNnnPtjMLSXjtTzEwPMZkHXF8htE25Ly0PgcbE6UiZGQok6bTB6bHFm+XveHB6pdZqLhvup8TdfMNFYJTFgOkombFGB+b8Wu04jDHFSn6vrSOXNlzsyPtLHujzbKAc6u5B8J1AOiUnRdD7TVOoLqcETLEtBoWyGS9VAWhKH1iDx6RHgz29FY9sqcnUwtFCf9gdCm/KHwff3wsP2Z0PqlWrIxWpi/LlMFHwKZ/qoeQ3/vUfuO5Lfmf3ENEMvkTb93dTrgBUryjIVDQzZivT6SSzcNy91NRgJjkyWzgbeH5pgT2nFEkOqrOJxprtKPFy0SYsXbDvL2OybXQ2b42709aOslT6D+eW56zcGSIrNdO5m5Qg2Du1ZGbQTVxGddBWaj58GkIhGwYj0ZqXN3KqpQHl/al0WjywTnRDZ+4kIB0TQfbK/h8/P8v179XkwXriD/WdrYe70B/01eacmeJmHcvK1FFRJzJRVA0mxhe+kyZyGs3Ja6698hdR0ABB3uw2qxJVNx+XGnSy5Iyog1wgp/VhGiz4zMQvbx2Y9pZTzAAkVvZ9+9htl1/VCtLMFojpVwdf/NiJqSqqa4Nt7icaHQ/44FZcwfzr41eo1IWVWQgS2DAdDwcbJSHoEMa/kelLxmzxDWmI8pHq8+CMRdTG/jUHNbRHb2j/qyozZ0wZM44P7LSeFAIwtqPRkgEfSm765UsfI2eUIdu9KComQAwWAg5SC/rPV3WXVvWRg6gGfLsBIprjBy+Ra3Mp/CcI28N2zWRSJ5YFaaZGGigzY4xoryx0yov2dAn7cp7fn0NpPSqmUB0ufzp2q8rOOhuPB11IeQJ6TSXEk199bmhF3MmlO1rw+j/SQkbC+qE/kqJ4jphBpjYQwVCvp1Xp1sWWxGR6go9FYrm12sjRgcBxHiI7JOEjmYyAEqm6ieun29v0TjJlpKrykcpPaqY3QJi8fiXQRJw6mCeJGG4SwV73iRL06it3W2+uoc4Q9bd/ICswVKnGi8Jv03S4uO4oo+FN7ipKru2Q6cK0RcIDr30JqMjS9TeaMUgPPZe8/RX9tbx4lKIVnHXAG38nkEhop9qf47zcVZM3RYIAUTsV4nTr7KXQ7OH4Hgd0m4Tl/7GpQmEqAbzsugldxU6vM3Snf9tUWSWz4o2uJgBzStom5Eukp3MbwVVjEkS/AljuEPyAJmtm8i9MyKdlxZSjHYB9Nbq80pWB5mdG7ezPYJyjT6tCV+QRCzLMyfxYUj+ty2BSrd/Hhz6319gl+sR8yXZPFa7T2GEcQWHbxS4KVAoitOithCkvNMKQ0Vg+SHlmoPEeaKqPqbFFoYLtYm0sRwj+TiUSvkkKY6rbuS2FaxRsAKM06Z05JQ81C0ZBIrB4OTXUEl5+u7m1Q4PQYH0NPYGZocN3aCzEcxSnMDGufgvsbG6zKvF0VfWl+xrU+vIBMiVLyJiFaJijpLi+OqWTrugcuWQyUEcD7l5ZPT2KyXDci+dWM0wffs6cVjp/ngPkhpB2WjS9VVvnH6Xa5KcWrRUoujP037crk55I7UbuTU1s96+0n0+Xip2Ulf+h4Zt1YFCXrW12kKzef5Dy/JbIDHjBNnTCAXT5LttiQo2bLOLpacPQLmEF1ArzHeKPIwOIl4HWPzV0drAbqmFIH64GxATTq+28M5eUqh8NxoJjF5OOnU7n693ezhcsu4uWb4fUiB6RPtlAIusWojYh0qNDfthMe3pK+PQirTSCtaPwGutsx9BWR3OIJbggQCcFwJm4GPImcONsD8lRxojs5tiRnhIFX7GCM4LLOR/uwZLFZu9cnVe/XLB/lnZXDItsB5UtS4v8AMg1mgejpgR2eEgQyyGL4Nf63au/IvSiop9AKO8KsAFEKcCkYJmG/5XfzbOaTe92ajAFZDtO0WnbTjTO4f/9IDVnGRveIa/wVU/kKagqmGQoQ9cH87lBfQ4fGnJ7Zhni6Q7pvMSfy4iHgA4rq/DWszrXN1QukFX4FMEotVDsoEEMijqLpmapF0D9iatS6slnrj/Eb2dYR4SGCcaDghWn+tVqbQbx6GbEMeFzpR+xM/0pwjT/rUUlo3SSgNKIKoe3/CenXAIde4aHzCKRFyPXZEvvfMvD0bHR/3MTqDgJU28O0t9sQAHf/sSJhhqjXO7g+f3hJ9OdJS5/g7CGTR8Qcr9jP79ma5rA3/eKiT8CRNJ+hpHqRuGunz0FeToI58fRrepK/Z0SMQICmYujH74tqlY90C0KZ6+Fy5v8b7cRaHtoNAeMCup7+1OyrZG2eus=
`pragma protect end_data_block
`pragma protect digest_block
589edc2d590dedce1c03932abbe2d9a0e2e84656656c2938059017fbefc80c4b
`pragma protect end_digest_block
`pragma protect end_protected
