`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
8naVFCLfZ8F9SQArN8VIj2iG/cM284PRSi5MtfKhv7finIr+5EMFOv9Mf2LP2SNxUGf0/uUkRa+PyAetjIQH2R9lWNw8Pvc4i1szyb+u1a5H7zeho1jcN2Rh0sl6iMc5+yKSFuiABHA72VO73e/M6B+T6kqEFxor6zW2Xok+VLU/miXaALhtiXeOHx6qxuP5rBCtxLnpTkKb1Ld1IFqK+qs7zmCjORUl8Sk+tt/9aFY+yfZvgy4eTwqmcU5wC3/Efa7nr0YhUfGgrExsC615tHw648txLTNxxyq4uIAIX5iu7zubJAxFn2HiY6SssaczNvBw8b7/7z8tm6nB6ipb3mRjJ2MhMzc1o+U7gL8F+73vwNXaMSK7mdvBMHInIRdWYyvnbOxxuYpRVl4paYcEDiIPSLJnMUCVET+mpnGa9lbTVp3VhCKH9CL7jx2W8mAQlYZMv//vCv+6qvjNxcWLtLfTIJyUVU4JgzWqXCUPU1cf6GGHULBXXQPbeW1knFJk6ne2gK3m+FarQU+4rfGmXl+SnN02kR70+ibl19NwvJ2lERaL/AD5qWjXIj+2kXTSCsSvYIMsiHpQdL5lb8vrmIazMIqA+liKYk2fTmE7gqGGWAsTeP7CNRFbNgxbJRsH4gJk1FU+Hf1+vjQT7ygkXvGDPlqr4cCtPRtuZFf+8SLKy7w8q/ZPEoTr1ge5qJJ02D51f0bnkvJXbCr+r+aXSGp6Ma56c0FhcZXLc5e4x2Y9PElPfvljzYs9gzzVy2+h4b1UbYSir5pmylZ3t/yrVWax+Hizf+TgRFqSnwPL7Dzx7s+26VoQrwH36PY2JNqN2Dx9gEA0ZlUrrvYndE/FvB5nyma2sfGLw7AN1WvZrblqpuOjCVBgp7CSy3wephw7qp+uZkJybwoR0k95MeaTtzlYa5NaBtZzSnE4THPG1ESQQRyM5tWE4N0aLEWu3q8yOrqyamI/FJaOaTiwnlpDendjhAvgPTJw9VS7GsBR5/6erF18tLE5ow1kcxJwinv99zxCBfl1VeCyNLT0/5gWU4D3Tjx4VTb/1GLfhkGfouSLIKHiioYBNmAmvOC+jmMcoHEOrEeDp6ILMZqru3L8mAquFZlbxjZKUzJWCOnsGVGKFtP6SgfaWNseNiyJZz5ZFSEjr/0lbRlC0AQEoHFfLpNSiTiMt4UQissSi5k/EJXKra9qRGKl2FxlBLtZQrAdcNUnI6pyXkfv+KDofOpjya9hybG6D74NgMXmF3Y/Vu6EwcjEhnPui3qou8pxhJWxlbTxu3ddF2G0wBQ+ux3uBJxEqDSfIeKMLM8T5AON/dq8cdwHy7UqmbrwO+EHgtb9UFZddMIkof49ynM/aXCshzgFDfLT365SqN5DRU+4QXscJhOEh2KlY+MiBzqEd9eqMK64tC2BWpFDT7oHAaoDdOrDrbPcszyV4c8AKCZJeg+tDVRKzTEWbl0IReRU2ZO0/LAq8e+3LppwP71b3OafhbWzfkbo5YawLxKeYxvzksHGL2NkUJ+QCFh/HSZpyHYlutAeuLdJRfc0SmyDo+Vhb64V/GmBZaFZADRh8uivlLkNpRtC2xd1VO2VskEXkoBJ90h7cFg1TQLm1xmuYiHVlOH+zzQ/jcbLPxViDrg3FmL2lMSIVgDx4uK4mxuX6vVIjWPLm0xoyZQEx9la3m7vXzzvR8zQSTniMMwyB5PhK+NGcrVAJsm5JukPUfk+zE49r1bvjyCbE96eEufF/8eizeAjMZRVJV3NVK3BtZThzbUq8I684UQCgzG+gUdovfnuAGn2fUYbyP2OImpuuU5s2P1ynKh0C2PUvdVh43o2TVVneE+EM1TU24YRyHMkPRaG/mXOyMNU3U0e/ktffyAE1lf95VNHNseNSYP07iACnyiwEbET6CYxL8wg9jimgRCo3DkqoW9M5Mg1/Q5GNqpkfLlL+d1+A4/nObqxEgXcMewIvHG09rZilpHOlIogLin5oI9tsQqqZmoHxkuZQdHNy63shv+n5EjsMA+8lgGvmCqMm0liRptxlVOOnn7I3IQIBCBSP/DSU9C6raNWYcFagp89MYfCMQZiTfjUFTDzZbtn6ikw6YkgpoxSac2CxqgnrABuPJHMX47cztdL72i7/PhEeioy8uLlXGVdXlc4UUTe0jCofvFlnN4Wg5kDYw8E25tbunZbrEIHGFDieHhEhjZ1DOwgba6gM2FZc9fu7D49gSZeV8/Nbex9K+2SB4VOYpYXurDY/WQoDzgTYVq2nkAtmrzJgXR65eIseyz58eG9hx+EMV6+taCl4maqhlr2SvQBUhh0EoIxPonojrIgfBIerGWo4o4kNa5h/DyBhN9KeVBhkclJrnx4g5DM0okN4+yo0tlmN7CUuKzynEFc+DcoDCTalBiFJp8/PwSJcbSrOkG/JRkvVSo6KnOciUuqHK+N5JY3laWJJWM+MRw4RNPgYMnW/iUzh1aRl8yYI76siVlwTP5LPgsqASbBg5956c/MJQh33RRcaPCLFtZPMzHhx040hrVyl87f+UU40Xglyx8H2RSZNH1E0NtXNRHtrQVsLNkIaIxmFo6TqTnBjtEBOAeuRr4SZFo1z+5YEDmj0y25fk0xcf6jma0q+mN4OZfU3+K/QvaPq9UvqllChOZ92IzPk3reAmG/9vz79zZnp4/STBf+L5BaZuxU66LU+XWCfsHYX5pMa49REqhxm/Usz3AkfP1ccylWKD0HsT5DXLT09E7t71T5kqOHeaui+iQ7VhKY2/ayYA0TJMFcWzWqC442edfdlhRW7lFaVfys0d/WRgwLO4fAiXdzGjtDRd6uAa1tzrV0G7WC+BX/36rlb3D6JaaDuEMHK9Ajdm9PKhrddeflrhz+YvBkyvRw6cQ5M0S1rKd+UzOwr6gHhbarQA+RYLHCyLNQR0tAQ8swCTMwo5pCBZ0Od9yMF9Hzu48R9Tc8+7EEGlNvX0050/plgOsaL7LPQJIjlshMyKtn1fwYjLDafd5kDjHEfEIK4T/Rg0ZwMrUtZms4RCRQew/cImISzitjEW7QmzrY7O6m33oqLeSu9GLnVnhqTxcgMLtFPb9HN9+nDGuiMp7FKtdokjsGQW33f7g4e6kOKQn2V/p2mGpbwwp7oaTjSNVkOaTFVzVozQ5vkESkD0jCsZ0THlzb94U3+TwukKSsYHS57jQjm7BFy2JdV9L6Uky7aHtVRKuu1Cq0jTXL1L0IieuOfyNZGblGrqlLUkjVB4MTf6PKtNgRf7lhZprvnPYTlVjOjqIOuGrtM8FuN4GMg7lmOY5z/Fh8/hlb4f64U1EH6gdcP/pCzELI0e7Gs78PkFmWerOqZpZFv9zRmupZLbLAy35P2JGbYuVHQJa1Y/13jeS8/PXAH6VUdeTScqJ1tyWY33U3OZlV/VMuhM+0HTWTLmorC2ajLzUU5uXhSuh4v2O99aD0r1FAT441qFG++7PueZrjsSHn9iiHLGO4sWmZwJZwZza4H4sEIVzFqb9ugoKqkMruTbFGdL8X9+R8DIrdZ+xhK/QnicEvdYhGnDS3Qkrc0rMRGSlJT+8vaGHqBotqnweE/I1v0goHSKWt2nPQSgWwK2O/XHX9sedu9W+63ekc46nm8nuGrfJIKSryTQ1JxxTw714IYcILD23ZEC2J3BkAsfsiGt55rwAo7vWbcH1Zz35owu+wvQx4+NGaUOjXydS/02NjZLNQcCCjDfJLFzco6nW+TdzEiqZ4LKzY3Gzhsx2s7i0TB0x7Wt43O55bj+LAsUXZapUTTWpGgJspc9geceAMcI3kmsMQdIcQ1dD6DBxFAndmXTRpIMXbJJYlIGOHmjwfN7vVcrT53Lt4nONU0qmAaxee/uTit8bSGiCh+5ysJKMQ6uqYveq+CYE1GkZrK8RCbuz940k/J9bUiOwta4z57ueu86l16wUYyWvAoQYku94/4d+I6M1FiE3QkudgNWh9tHCtuAimwP8/AWZCnwakWBNKx8PbA9Rtd7cFh36+UuKuGyVrDN58KJYmEWJW6TI73G86mmqdiff71hQON1ZBzSe7lYM8gw4gFG6BUCDy+JhpsqI9SO79/Ez6qFkqJNlg2M3910RIJcmoAB+DwiXg0P++dj43XHZPNOwuTNPCF51AVyWwvAbwkv0kg/dh2/JpLrZyG0psULiCZaMCIMB5QcpUnvF18xVrAuN393WfsgZKIgf7xIUTr1J4egG9l/p7x5HVcLif3YyeGduUhRLdgyc1qZU9tcEWanrjAMD1KVXvIblu6zYe7jWuRdC4Z/hq/mnJOlAO7lDLPDVQwh6r6DlXpR5YtH91I1P5mbGZRr3unPcr3wJtg3RYoRgIodyhGl0OqFw13hmtCw37eZJs5wm6rrDjZgz7GjCzxmZYH6FS+j1EHg6a1HvAfgIO7cV3495WxjsJNUZevnwf7yaYY5zjMtGtVvUp6094PPCGXGlsl0JZUf3LR/l9t88G5ys/F2vt1Vx7I6rnza8P4A9Zy39XU3AxX5B/kGA8oMiDmGH2QiNjhBCz2bW29C+V7wDa6vYpelk2Lm+4B9boFAqleFZvBzkQiJUu5xzhoOo98ZllykgW2tgPUVGgNq4flwf4OLzpGSn2vEGZSoqeXUVWkEexgl+12irqG5zdaYyinMrbmkmwr2INn8ydUR481oHoVeRWJUFrQm7CJlZjudAHFoCae/fmv1hWg/5rG+VTFzgs5amyb2uTI9sIIZeH3VSO/MUTNi5brvK+WPem2OVdudXtGv63mZVkfCYyRZLfBmmzHGdwjEhGNWMCFZkUaLtGyEWgKqkWLx1jleS+bizUVhN6CD7olkvhq23XWEj4TbcU5k9wzetFgzxf/rBGJL+X6L6LM+KK3h+YMEDNJhj7QPZ9SDHO5wcBnZKJC1qXkN7pqIrsg2mqf3rfWLlHo0QwoT0emyRR91zEGpl/ndapRmaUz0Ygk/AQwDlOBwaZE6XlQ714V/Jk0fA3bB2oBmlL2HSQQ331NoYNK/X1mZEbk0htpYk7mhvftSWA+q8+dR2B0hRNrP8tNwq4//Ge7pwqIg34IP4IPuVwr0NkKE6vQfzS3oHkGI/5o0i9ep2tZ8IFBrRPuCFxu61ruV0jRMgnIgnvS0A2J0sQqocGDglue2M1kVbGo6UX9SUuzL1GOrAnON5X7kMTwvBtC6s1k4YWeyPReLwsTdurHfxkYY1VDGEkpisFLZFcP2e0wpEewZUwNu+hY555n3uv9X2Li3aLh7EJsyZpERcGnxKZso03yWjp7eYlvy19MvR+Aa6un+ZWSiMAVjp2EZ+wNcpmDdjPrWYVmipnyFi7IHecVcE+mV+RJo198WfihnTApCQZ1AsiVXYZBQaZH7HQKZ01NBTdkLL5FxpEknCR8kMOB26gXm2qp+e0vzrCdKWIdVDLe31ExQWBP5BfZSxM6RWllhxUsrtI7++f/BDW+lo83xSevXtLvAQmXp3UurOSFxdVAPC3noSEFLoSMdDsUikULtvNUYJhKifOWy+Kpyue/aZzKPlhZPd+84slR3yLz9hS1p9D4SqhDhrB03Xc48g8xC5JZ9jBQe0AhaKLqnuiTzJvKcMv9shN/oxSYHGJ/F9c/EqD5UQ1hMs95IEMNRkMJ9BSl0XRWPRBG3xFTpu8jEvsCcgmoroNei95dA0DD6T3uxRX6sA78Z+7zRFk4UJ15XSBoIRQaZuhvwiDq03SoH4HpjD4YreUm+w+cPovoqr4IHIFcSeeG8nWVImMHczDa13+8aYTNVaTjwt43M+6ubcOlIHoX3EopCQgcMyh2n3Act9bdbLhttKheMPoSBlDaolaBWZx8TrJeOXoywsP/JgxZtv5C6owaY39y7y6ANqpTLvZs8FPYvBGkaX/9osJvN4NaKUoSwZ00GPUujlpOX08KHY2+qbAdmXeOAKjsH2M40hQG3DXl2qpVgleY2ntECwZO8lk6+xOG/Ypwa5TEKjjEWgF+iPZcyZ/XVNyuD7isSHiBm0bdyL7h5jyqf2T68qdn2p+zjqQJlHX7syKmyyQSMTCVYNDQmcy5o/Fo/gHZYZMg8uh0da5NXZKKjAoy5CC4NTh9+qkuHYET+wNbWfYXQ9niVbB2NagkgPByx+4ewfuo19gGgNrRUY8tet5YRA0G58WapN+NX4jhESmkEE7/u5ccSbz87+ptdo+TWXLN4GK6dyszYKtDL53xj9sLTdBkaHQb+N7v3XXUO/Rw+k0D2SDhBRYHYQwY8cIRehkfDPhQEVUkNyudNJQ0zCyYYXvO03GiCt4orb7gZ9Axh+RcgV2Zd6AmVUj2ZbfsclY0Fb7ZRWCBeTaoVY3WhB/CrKCcV/7biOSWtOoodPUN39uobCHDpS3Dd++YRXuPkmcY19ajZf+U1fLs81F09lymIVAgsFT5jt+gaqn6pTo8+sh6GXDVnyJGa+hlEUiXGqmtK/VGrKA1MQz/vWc9yXYj6C/1WdnPlVbDHpzbJbmQvMIp/luwEsp2uCnSyDshwVTlTaOE9tDgQttof7lmiMVN4TEt29N++2BxycYe2TCvuU2jib9JJCWb2M4BCMZK7uLjdawrBEkUBUU2M61lMXs4p/2o0HuZwj9txyZrW4yRJU8FZ09/dqDIHC7tVOG71NA+x+eVlGz08FCyA3ttGdTJFc7ZSoZcApn2tsGwQiQqfWu9B/M+mUZRVBauwp8w9cIujnOGvqJ0/vm0HPUqGb3dbKbzy+qDn753O2+w/W4lQdKFJlg6YqUJMk6qrQupOTcMGFhaTho0dBPBXF4G2X1G7KfVwwIFBfpBeMbP3WCsP2EKhe5PdiarTFjZlqrvqy1V5OGhxOez3mfdb9v/HrCj6rfQI5NO0fCIvlW+5Uf0lm5C8pfLK3LLxyxomN2q2DIF1fPaI6vhpdzrxkw7ZQfirx6T4YXfjAGILc3mclunFRFel8v4sNGvHK8fLVU7HacwEc/ATGorLNTN8Metx3cbQLhtfdZG54VywfodJYyI5hmcZkbN0/lSw/Xrs77nGQJx6LdGqsC/wf3d0YZpYdgrav6n5o6LCsUTSDGo+S+Nk8C/B7jdMiw8tjWuSB2+uLFc+TCZp3asoo9g7m0I2T6503keUgbuOCfB/jXjHdblajZ+mFIi6TiU0TATomIkP2qyYw5xAWa2Bx5AXB6fYB1nZo/bZtJIGeLp8yOC1+zB3RyCEdaTzsoGM0WNkJLn1/9yRxo/u+8o0mAXsJYNaSAhriRmal8MlaKWzFAfiBvbFHTypP7MOxS9BDDCU7z8ILNFCQ/bSTIC/Wax5NtdhTiSo6PlFsvWThQNsY87ry8kA2E63VNMgxBtpFvNpWvdNWADnpTy+83sQL9O9k3YqJxOeSPJkwanJ4JMGd3GzSKGiF8jcysqbECO7u2LBkmPS0qDgrFkSn8bWt3rioBZeZVlkqXxl1d/5nGdTSFnKlGKi916kjLOw6A6Uda6JINZcE0sy6d5Zc3AxHHpmBBCgvLXNNR6T3IEJhXoURKgX3+ZaAjpT4DDfduxbfXmO5ibW8WfVgEk6uZWMWCNPMe+uFmxkhqjD8+DOEio2VJ1WBs9HZMdvrtoM9SzXqjpkOJzSgDVvQ+7LBaZ9ItOE/PKGoDSXPRvpUX7wzQ9YM0gYmdfzCUUqW9tTKqRA7x/gJHKSSTLZZF22KBeLQcugjhMGX6r80CSTYnYiPB6MR3unCQVK+L9XLBKf+TKXG9+jknPvQ0DjmjCGbiRIYZR4KKDZ2Ax7w+J6vepunOcEki/N/uRdbSaAtsq0PJU0teieyaaOR5kjtXtQfPzGcTN1leYjxwtOT0t8JC/4CRCmpuek6JzmnkGR664lBUessC+7tVnbdLkKLLC6g16TUjXmNWYeA4eZZQb3maW+nsSyEWJLesD/RJHgH7VTISkB2Web7yi040LjiU8MhdSuwpScMBY7HOtdMhQLEAqlYCNFBe8SqjJrckdKkS2xsbnmUFs02S72+vt8eHSTWhy9jHwRYn/bh2B7UBYax4bfbK9bAopuFEk7C0Kb3IwpckN86UZTffecmSyk09o9IfWru+cWnCm2OBsnWAx0UmWCH5Wv1PsGMenlE08v8sOciceOQauFWsRrl//IHP85hkwqywm9Ig692SBGMOYddVBNBKU2/iStrdPbK8DCN0VL6fG+jpHS95OWLvCYOyseL6iKjkrpKC/U7Vmp354GEUMRRWBc34a+S2C07XfsOO6bicz8uv/wN2UfzphRZwSN6eUj3w1UZszL4IMpaq+xEC1RKNkjxXZE17tLZ+rvdjPJE9XDtHHUfqEsqwxp8N27aHYFuZP8qD5m+/u/kGZ94Ms1AGjwnps6/IfHrSqFqS/ayCM0SrWk90rVwsoQcf5ZRvjJ1lbgrvqY+GJqQNk+KTRJL5bM5hZg9iFQ/gEMVd63ET0UCatDFi6pxF7IjdLBg/HH+Xk88ICK6RR7PJ/uiNQj4FIpJT/h1y0NkUQIWJeFVWV4N1EaLHHqgrV3OXEcmmWOH4o3hOy8dEbTRnEuGMXyUkSIL/nehTP6USw83bZ1pD3Yw+OWDRATKjY6ptclFu5UfwewtFxGDfP8HKWU0U16KftgbGFMM0KeNBK/1tjTdZMWjGD7NtM8D1cA2lAAHCiz4w/NdngmMD1X1AruB2GW93tUMKfR2AX74lZRBsT5dDSDj+EbtsQWIUqYEvKTa2hpTp5dK6WA/bXCu+6ktYDgSquZgPOWMZyPNOjm8JXFoIJi5e/kNfZVuapAEl82HtZcpucUMsdPqqbewj6oLBJ90N4yh+umKQw7VXioxVojgcDRCmF5q6tWtXXfdfuZv26n7i/hukT+OGPOTB9S4Vssw1Vi7PH3/U4vrXavnvz0/G1MjgbN9Y8XDV4vhGUTK9tYLXGgJc9tRGrPGVnbt+5iJR7+ehzwr1AHX0bTfgzSWrMu/RkyEofAntJiV1GNsMDObT441waXxmYdmIi5j5wmCPMAIiPmPIlBtLSyra3qlX5M9p+pGBr0w8uGwMAvyv7CS9UNHZPjf+/QsYBf60YlfoTWzKoCzBoH33GsqCQPwxC9enViziMnPzl3by92AVk5t9mv1tBLIq2WKWNmOgtbHTAob4kKVzZu2lGnMyKQrh54QnGeq6Poh31WoNu5Yjo+cvjbUY+aG7QqmAVa3jeqRTsOwRXGRaXPYKyAKBvvDZzCD9JJRLHn7Knx/+aPAfATZRblyT5VjCebIjRWZvBA67DhUqStiQhS3oVoqnYZQ/109riraERnwarGHe31IcHlhaHzBYu1by+w/sRYIHaUi4l71GQnUNBhExhCPy8D7BD+IqnN4Vgl/Z1VVANYsS2TKMWVR16SMfEUjCz9O1hJ9NoqSYgvpdzcqwpyPLA9e8L0imGBtKOb1/rdYaDyA3w7sBvNyjwN5x+mEUJIQ5W5zFbJXs6++nQmyZviwcbq/PazHL1D3HBE0suYjxVZB+PH4he8WLRj2ceWvqVcQha15PRfD29moEkQ1wsyjshKKot2t40W6oKVZkkXlgNETuX1VuSY0Sbw0RUu5j7sT6u2EtBM+Zy2XclGmuhW3umpfSsJ4GwmGw4FYXxgwCclU5lIjNcRBHkhUd6WJ4YW9BlQcJD7CIMR+NOeJ8rqIrxFC+4GYFd6tLfZ86nkI7OzPEkYeTzg59Z/9QvWU/hkrT7PMKft72vp+OSItrgUa+hokT5SRLiSvBfJvy4eaNlpI6asBgbLfsSBwHJ2P0/5Ye6uc7Fl1ElR85FDZBNSs+08lQV5QGj0JR0pXjOnRYG6x/a5Ogv3utmFaQqAHjSx392NwWvRAoB8xZJEAkydY7yOBRziFF1tOSrfAU0OsLol1L3Z4uDlREWjP357DBMybFKY19/oXh8Fp4Vy+1Ysz40Xy2Q7QxGziBroXwBTCyV5/CtBQdVuKqu+kRexMEfSZgtVHDnZiZcZCytZJurrP3620mt3s1wSO/Sor+RZqN7Brgt9p0a9Mv/7ohNgpIubQ05zDC5G3GmIfTJ+O3Y7T6vgfHpPxNXY82E+eGdVmpw+Es30Mq9YbAfdFwVvqABRxijtHf6iU03EIRVqkrjwy7javH8dg1KQjO+yoxBd95UNe1T2zO+0uWMRsPsQVrf7cHykV6PQq/ivKkSrjfMSY12csAezw8IQxwn+dgyzFOvtcl05E6f3Q2n4iiyqDRWr55ct+90bR51nP6HRBDnfEXES2wCvVaaakCtG7651Bb+0/JhEe8ZDr+4vx3hEc5b6FqzoLizLUM6w2F7lm5EBv+eSh4vkaJlqPH78ZrkjRd5m+jIO9YH8EiF4JMB2HWL1WQSTtDtOp+PozCjCTw/SjmQw5xQTSC6YZkWcPYVevZ1owSl2B+hZNE+plyb2iDI+AUL0bbfop8bmh4sRbPuy+y7T8aHTE4H7ymlIt+A+LMy26RiwzVooslHCQ9TuBc2c351NsdwN04tIGvZ2z2kiOs6cyyWL7En1/7+qW51g8f9iIpjuLVKCOuV+P96NduZ+LRtDEK1tTLBaFbDb5XaXrNBInTgujLP+juzPR+aKxDzYJ+EnUpCEPnErHCW9fjPt76fmY1EZz/WOksK35ydW1pGU0MUddZBE5mE6VAXprsreaEyyebJ55W9iuBdlkDp28wC3cyNpIGbcgIRxWPMVbxq/AUq8PfMMcPA6Icl6/p40XyGHDLKtyzzs5l1cKj433lsb7sFKWqTcs3B07vOjHazvKxtMRdZ0bzX+pCdiXgTVKyw9dc5shvSR1p+He2RwQaY8cdXC6ryMp0ynpk5vRIqpALIKU8zp6zGjwuEQtdogaEKTVPfMs3L/NWEcoapPL1JvVwuIvAcYh1pSt9lnRhydjW7ktAdQW2uVIEKsuHquUtOeFqVU53ZyT0s0IvppbxWAfxzifLWD0wrVRcOE80/gvRs1Rh15vea9vAapSTalryVGSj2+9AvAC7ftojMrgrRTjX6IrjBiHfcbw77fr2qPJ30DOlGXSaWsGlvj/V2H0EsGXhX6NKTxVoTExTzVPqVU9MwkYE2uZkSyzpnSXm2ag+UWH5ILeBV52eKOke2eyBmh4SyOu07UqXbDthnzWCbtMnG7G4ucy6wNEDATWEaKkVSOiFISNc8E52S3GC/fz5bJ2snhMSCCBbiOToayXqkL8DEBWercHW6c+LCi4AIV4iId35p+HMv5/xyKx5OyGWaEgKXCWUUzRTd5Oskr09juXz+qZ30AXjh1nVJJHFNEACkUAxsCuqfI5ts9X4taBZmSDxVIIdtlJwncQ4w90UgCMIpalWtCp6wvXWsOr/IlsqTCv5UH6kjd7olso5b9KiQMvlgM8fqOLK32eToX2m0aEtNo79VXozuQ2j+FLCitiByRtKdrXMk+t5q+wWxzegvCwaJ2HqO52chYPHCsKS06U56cyzEn8ijL/DTjZzKM8UoBO7nnXkod0XfGFprRJb95H8Ul7uM1FX6fUTlU22n1lWbZ9ZBfG1V2Ax0Jv4hQEVFROAcT2/0aKvXEpyH4EdjJiGc8m1BHmCkIottRS+FaJt+k2rgwZS43UWWmbZ2bKEkdVJyReGaPZpI248as5xn5daWbFDtNxSp3d6HNE2AnFijGj6XcHSXLXErL2o0X8OzpKwkL/XDjW2w5exEyt+h9wsp8mgP+iNmgmg5SaykWXqdq9Aw2Gi+oq8URxjK7Uw2LyhurK+1iDrEU3PlkP+nTLPR7upOoOe2NFPWbxLFiHu6ln7iFxuvxUXBEf/peQISe5MnG910gcCNbZht1u0qol6NPjY7BHO7MGAQiHYUYgH9nu2XelfSdqLLL5xUPXVOCBV/gsDDP3PLsgdZnmom8hNqoDsQWcGhSqnqoSnku0lmWlYuZy/pivbcic/qeoeT7LD8qbj4JAB9jQlW/Ns5dXyiAzY+0uR0TtgezptZLpFcOzps5K6z04Vcwq+ozj+sYEf3KJXHV3HWcHnUpETvn0BbevOa9xNNGjmgIwEMyjWtitGndt4qyzf9eN1k0K2VACMnn+PNyvZMKdDFpWiPL0U1citQZCvr36/oNRRo6L9BPoPaSgKPzcujavdOqPjBJxbvVEEbEzWDy5jhhQbEMlD456ZdtMrqopd9tejQfPWYme2UxVAlo82UcRX5Hlxish3eHXiT2Vv/PCIj0SEf5zNxXymZ+oyQlEPcmXHWfZ66yGDAewCpxy8mtfcw7taFnokgMtVD2pI+eW7N/veeaXeKNc7dYiVjZw6nb0r20xLD5MczCKtBGqfp2ZPFH9Hnx3AH/gez2MyEnCn8sMBAf9QOWjLkJSu+o/yG1vlTIUqR33cEKs2TkbzxkTLyuTrsVPSsceCrgWbXJuDkxbof7B6eJHg+JDD6Y4gLDa7bVhYrM4ENGGKX6ZY+bkguvvHS55mU7PVA0PYQYKv42c563kv0jYETow2OEuRPWGHfoASBela33bCksgdwMsjc+Q7IDTQwLPqhW9K4HmHTfZdfBVv1YTidyL2t1dhrMp4w2Z7JuBrqf7idLu2K4g2jPt7NdaPOQVDEsU6tTI0Npg+5uMUlzojthkY6UrMlW6D2tAk5KACCmM/Pn06e02gIgRItxQCDm+e9R6KMGIWoOI92kuGj8qCvPf5Q/ZWXqjHZZ8D2ame77S7A5YYdYA3jN5jUSDIEIt3TcXc7rXDHey3GHR9EMovXI4FsS/KuRXDz/amTH5hTVkEGRHhvG5GR07j4B99WmYM2+ob+yIOhNNiWhH3nW/rk0U/Z67SMESJicaDsrY7fgrQyJ4g1hug1fi3+CBchYypmnrnauwnpF4d/FAT2NnfZsV6E6znrNB4AFv7nzQUaget7+8dOqg/Yi5aysYfKKFrZd2Z2rkO4AkMidQ9sejdK40Y4tgx0mC6Q4/DAGCsPTIBOmGRnn+3Mi4yH9+Pe4oFqDPnFPpJHGoUugpwI/WAaimxmMB7dQ+RF28g4XTKgZLno49AC+mBrdT1/mx1/kibR/b6WbTkNq2WkiFGTdrLsxXOXNctaZFQQ3oZTm1VgMQHV07IEvoAjxo+tMfC66qFRfmZ1dqF2Zui8SopGrtyY87RsDeBNBWoYlJKzavWyU8pWp+Ogi48hq4n3eZ8j4DZZHpssiv5Z+B7sYrQZkqgFZYqeZL3eNJUz3PF5j/JpQxmi+1E8VGn9LV1aBUNKFV78PaUMoZulcBswj9WSADnmzOwvv8GOgQ+6aV20SZTSDQk2Ch2DcKxp7yIas7i8TfUaawfXWcgEaQuBdxDhuLrQpNt/vTz9TfEUy3eU5PdVafNWA0VfBByhlechhWNQgjqk7wUnglHHSdx2m6CPONyLl8AVEvwBTWaicjxlfInZDqRh5hYe46JLND97UZivhY+Tgvn7UiZ7ySVw0lyD5cJ8iCcwJ/XPvVb+ofZJZIxblMcT8JHUJC/vEv05M0Y8InhPDXkYWNF5V2mKTV6F4UeS3rNMIMzplxRQCBJO09YwKx0ydwoaQho6FJCdJJ32XfYGTurgz61I8mHn6+Bs7AC1AS8+JI4NSuWakr0X9EJq0QvHPMlOoqmWG4Yd+HFSoOpbU4NZTSAzO8CCX76h3GH1X8kqfyLCQqK34Bkkm9vt6g78hlr1U2F4MXSDiPssWIKTT5s42CLV9RClRoZ5WV3uvGxG3OhnIxlXcTm4qBd6eWo9N1XQo4lV32xtrkIPvgTTqIZeFbTOiw7a4r0i1fBj37ZU5MeSYi9KUYdjeSQ+0TXC9ievIfEOWBM4PxlnYbJyhkFDuzkU4s2ZB2kA8/fARkNIWBnoPdlRJEM/BsTaqbPCqugz0ffhlQV5+OgTWdUX/1pqIGqcX196h1QsBFMkSivg3NPbuILdwz0TbqvU+YbNPFZYaeBd4elPaw0h5aB4AZrOpm5LDIPkPNteQuiygUuLxhU9vLcRCpLQQLh+W7TZjPxOz6Epe80NfPNOkhuzvW+6uEdIufimuxwZt+u7Z69GoOWEh1Nk6WS+HHEwEshYAs4fIU1zeT6WlxHwCxt29QrNRUeW+4y+eqcScB7k2j0LAmFaUV3YHPiIDsHajuwqsxtlnlwICQVtr+2DQc+7P1HU7eTyWZ77BtYEF3f7vhhLzaKqpeTXQrCFFH6TkQrJ5hw8atIW0ciq0jduGaS6hyGoxAl6kiXLGDXGbSaxKKjLik2IdFR/EoyjMwDwzbElu5fCbCqmt8ybX+sGgJ+xxpcTJaMg0YadXSI/UHUK9pp1ntrCMYGwARPST3n7kTMmnPcoHrPyC6bsf0vqEG7SmaZBljX8X61gqXSJxSHY9Uln6Oq7G4e+IfBlvPbE3FAEEE/rsktialoSa9pTbKsDMd5509ze0Jh4epQfik3ogvGXCxqGMBcELBIaeR1zPCDcnDj6xpBo37/ts2002/MlxoIohXP4CaAY8PqYOj5LAdqGlSR1Na2I5N7UA2raMc3aJF/pBNIG+06891JX94tYV8iy2NCIt+D7ikj2eEq5HXypPdA1fnLLWa9ebJL8dQysRnVzTV/qzbaAQSYFx/P96jMjStAYxTDyG/5l3GWurRRN+W4mvkcLGds10tDymWs8VbEOgBp5yUfqpe+L+YF+9iozSz4tli1gCnGULB9fU+TaRV8BTMiFEd0IDSTdTgGTLLpZOAmsO0HPJxi4HqGC808Odyhw5jpVIqybMj0aJZ4g2fXI81i+saoy4KdYeGDwf/JKdWjTQ9T08s4OYD4LInoTGrwzuD5oa7orUyTr3pEmtATsuPf3VEOSXlYl27ZRbke5o/7wOPk1BCVfPD/u/1c5H5sKqQQWeiPqXsYOYw8VmAb4lxmz3EErXFxYKYjDJ6AN+3ri3jKGUfxXwLhaSyCQAIao+D2phmIT/Ji4lk1znpYQECrKGjHB7zs6npb2U/nB0oieQ44yNsWxRU65ohb5YPzQNI4zR2XpfyN+64diGMlb409eCGrfb3Xd7OdkQ9AlTdQtoNkx0u5eauF1e8YKKKegAB4iii+98U8oRO+ldr13t9usLhkWvzNUwekVc1qxTiYLJI4oyiWXvR1V/BnWel4easbX/C02VS1navBkMnBYSy5MGdb8Lo5+jP/sPIzmkoqxYYje3axdDg7fr3IUHuQX0FrxOmtnOLM2AyTc73CTXOMvyZexRNEmJhve3RZ2CJes1mIXX+Rke12y8uMEmHRVxiANgJqrKiRvFT0yqczakdSHM/1/h93niViAUVAMK7aayzUi2/ht9HQ0l+7AxP02CVm0jRd3YJ/r2DZmsWN/INcAUp3mTgMXz+rpiRBRS8awD8NIHeYuTM7gqqW4MMi0q0pEEfvDc35gvpE1DMXhxyMbwHpg9H/z2u3tEtut1qDrJvematmA0IVCxZC7gFfZc3ck45Y5QzvqhjKhVSqPwjnwlTknvEnscU8IPF6W6CPLxnO2EPdKGnXizmNcIsL+yYvkxScrWJJaKpgkUgbK3DalU3w4Ff8QYc3jFl2qPpruqZacRtW4A/2CQU9x2GoLabdwuD8/3m1RCXxQ7hd+8egrj854ZwvXzprx+ogVqcZtL20uroqIGoaIhCxvabOVDKt74uWFohK66PrFLUEnUebqq6iZKUBC553ZRZJ70SWeh+y24wJUjUW/4IJJ/Qm7v8w3WTYuiK+5xGVcSSm+pe3KkWxoRb3hmZiFhKM41oguFbTRRp/+tavELfq0pFj9CsHm8WQDa8GvbL2drkbOfjmyaZYORHXosq6XBW05BxbZbX9KFi4XLHPW4Zc5JtZZ4ugUQLsF+rrp+fvf3RFivtV3U6+oDrAQJIgVz725h4DBiE574PAWaTq/aHPWWTx6llr5fxCgHM+kewwdvgINTqaVUTD+4R+eIk/fqim0texk7xkKxHXfngx8kp9wDk5zeZVwptwwtJTFL5sI69xIU42LYJ62nrT8e/ztCd32Opel1zkyTkruNthrakpqzwE9YHAxq6DOGrgGOAMxO6s9AKVTdW12UgRqx7PVXymW77NXk/T72zNIEZcvlo5S6dRwdPAY/zcnvlh3KGt4KpR0lACbEvo9I6y1ONNqZiHIJ4lGWOfu64jzduHNvblr7S06eM30hbshcrmLAFi5S4BIb+RoTh7HZDp/C9e7EQiXTIlStTNuk4PiJ3WSMpMKZu406EKAVuJzLM3nB8i5SFmrwFnNRgedgRFeSZ1MuTt3DVF7dQOoWFi1OnQqZ+s4GuUnfc1TUxGGcf4y40NCDbVGb+i5bBz+AjG7VV2ymuFwpFbWaQmkqRMe4IHGF8i6L50417fmNRV+cewDV44mrGzETLS9+/dNUnR6WVfQ10x3vbfNSDs+M+Mu/87VuBqrYoVlvWrJqyRWk3vUBKXaRMi0wIx6iwFQal+/TiGpiV8ijbScvEY/jbQB5apvH88wKe6N7oG3cMAZTaMr7q2H3zgZkp3nMfl7tzCSQ2il5RVNAYO2TG6v3aUAfuDIXB5zlUO7ARWRuTVtKZc0F5sFqnL/aAfbSmfjBnpVaNO5BKMfRhLATejlCWNwSHJwx0gvZH9248Rb3/nRoszv/01apsoZh0/SQgCvJoSiYadp84PZff0Gqv1RqiLtKUnBLvZy0oZTjO9i6mvYmvWU0Mo+iUkoE+39c48dPDvOEU/8YT54ZabHR/nPAXc+ZjuSivY457CIQcarMFEtayOokUhgh8RzcC9U9UF/wMHHW74xJNJzb5+3hLLyH+QhnURf+B4ejJdIpMCYv2fYCMPq5CYBozC+mUDTHEuN/3kbQ1Hd/OItrLYPhMJSmDRiu5MHHAnwLdnQh5SyNkYAXWf50WXWSSMAfm9NwVRbXWAtR9LcfQYjW2AIOb1HFGvDJHig4fCofQp4irpy8xX0ms8ZwI3T/LS3Vygrl8FWtp3Cfn+6kvclCGX4xnGFO2UkbznCswXOZPONXwOB0l0H6Gq2XO2KpESvPCgpK5XvZGdrItWR7K4Obvy19NG8V//4O7iZW/qpgS2lCOjOaq4UYXsPBRHWp6kZ8wat6u5RYedbnmjYahNPpaGimzkUtL3iIZsiGEoPsFmzUtNHnYy89DtvTiV3hmvw06wQ2KKk4qvO3D2t//OqVKfOO76ZbUrgZakfK3GPM8Y74VAGN19TgYUseTAsx0t6fQzC14bNyspsBcHAcHmbwYnkf/GGkeekIcm9ZzbXYeZYJZeuvWAQEDd8M2WQ2Jj27xE33dRky/kVDjYuJWF08qTWiE7E5dCoTZAhkq8nZwztqzJEkKGHioskt9GzSSUD5GZKiHX3q1W0uZuvPQKVVG5h1EXnTIp0VgWCxN8MNeO2DXkt+++e/jxATCxCNoXPA/VA/R2jAJdxTMNnp+4Z+3xL6ozJ+q3LlmgQMTMbTZ4/cm70tKZqxZOiiur5lI5o5lU3b/7HHIq6cMhv8TZKdX7U6+PdAYW+y/YAqKk/krZIN9zCrmbD0OlSax1+FxpY0xauk7eRvQ87SYlTYQ1uWXp2ejh7MsmuVhqaiTty8w0NGF5mZrBHcqsHS1Up/2k2EY+ZSv1DEO0KRrn5XefBtfzAx8izJJtCriv813MZD6TEwIlN3KWd7dggHN6gB/bPNGU1E52t6uUPLplu6/PQYvMoeqSabLjsAhwbEXY0ykshMQMkkdLX3H4xVlwCknIF6fUTfdQ28BlewMgPbetm9fXGyywCXov3CRpMe4FNN9O3+ccLXOrs1p46ipSKJK3IGT/6i+HgUao89KWVJp5/K91ZtVRgvtfnF409dBE9/yVmG+VPQp0whpCWb0BTbYoVEBNci/zj2bZ+9GsqNY152ZGSv+PYQDOj9hDHilbJTGSFSSWiTBp+OgQViuZspCpbyDl1lcJE7PAW6Y2FW+VDnAajDA9UDH8tfU6zk2fVVigePZdz4yKUqV08lJ8xq5Rtu+dqufO/jb9tDni7QbEsGjbc9c75PFq2G0DW4BKAj4+i8dSoiB6DNpBUlz/J1p1TYUPsNgueToOLYYO5A07b9XXxbiXl1T6Jn1mPwQuQoigOnljb6LZbtqingpbvBgY5VDLN4BqedVAnHgEM6jd3KUheFikIGhFzuCwuPA0GlGVLtYrdCtRbQ6Lekg+lqP8/paLiBTkPMfFgibGrGj09Y7En5CVB2V8OEwY7Z6eUYf1Hd4UXkFWPfrPt8bwK8WHvkFC7O4s3jlu2pmn98UMBYGCULulANh4qob9GAg3Y9P/NpuYci0qRmG0KDtETYKNWpxWnQLMVkZr6MMSLFNEaWn7mXPA40ywsgCc8NdEZHU/97wW1HscI2d/ouFEHrOKP8k0cPNKZoI2cslK/CqrFgpu/wrIgFT0y0ZyTCtyE/a5q4fEm/rhcA7QjQAkC5YDm94kjWpji8yuF/3Ttu41ffo/MsdjpqalWJ9px8Iw1ZuRGNbbh8E+OmRQdCEH935vCOrFTfYEEIbqerR8PpXqYFPIP2bUSY/RRfM54CmzrmKCaME8k2QhFOd0WaIA7g5RnCu/eyNcR2olfdwO5EXe4IF2ebv8IPKA7mJYcACv85bTNo9sEBZc2B9dU5DiqN8GFTskgdYwFhEGnf9RpjxfWFfGhY0PjFbsS+hJpgvYDK6FYDkXcdAReNDSz/PLIli/vcmf5YENX0hGhvAVCYOMh6ZNNpblCkQDKt3aW9xxPnozKO3QBCd3yaY50z1YnIdvlGHUp8V42ZMhoUCErkwagAgLnIBofVjSrx2SaZy1TcPJniEI05xG/Ev/UuPuF8eCT059vpP9qpLBaF/hF4poh3Pehuj54kOezM1iw5DDvs8Ky3KBvOkgXhyhxiZayHvalWgQWpmEoglBALJzkecdDOEJ6bpGkklp+/VoMynBSjv5hOv/liiGgfVsVaDt530go99KIMZ6LlefjncT24qjS6+seGRNaEkoaEgD1oxze2CWkuFALXF2rFGz+H2plg+BMoufv4LUeTi//dmZjQUNOfOF/y6MDuNWKo65B8+7mGXhx9eByW7/1b+VCu00UWL2uphV/ejZBQSLhIJCyqy3aWwnvx3/j7MGVPAkDIyQ+8KR9YU6/NlmlB6GwCHNC9MFpH9GVkCOECdy0QCFVVVHfbzmFgnmychO5tuCUQ6lE8jsfJepIaVvD8b/EsiFKQCeQlkPXl7NS/y2Wul1KNaWEfS4XFpYeesnlkLKw/bGgMyrk7O1utMH/vI4E8iKJdhnDpTsTLGFQa2VIjDGtHdppZZxkWMh0Vi9KXPpu1rLrdzr4LdXfgbsMMZ2dck5JatdCULamMeK6fpXwuWZvZUO8cjZ0iphe9YlF/AlnW/I/zEDruQjQeJr3l9/95VC7G6cxKXdUvxHZh0qOVdidZiB+w0mhibdv69zbycN6MxM16V0XVuIksRqIwyrvc9Bz8t0+sHMny1n5O84EjE9snoPlIOjLBrtehg4VRIZySoG3QgNjhyoRTnStqghSVAv9DQ4RvsEerTJLelb9l5b73Iez2Au+nZxhJ40jHH3xwARquNESr00blWhiN4rAOLVDMZUXrP7+ALjDXT9vNqKzhyXFlsk7JoSewzsNonBYWHzRH2lQqTQY62alXMuK2LifwQ2u8mniOs6ZT8JJyme7en7MrHNKyHXfwCp6fi3V+WcNsUslFy+QyKc6kqVGdABsoPRpIcSjdb5r8OWLI3Ch3PoJK1vpIqUjAz0fkZEODGzCoKaTmRtrirJinFuytStl7iIe69ap3vqJHWXIzuN4cSWZ9zQordC3VaOVGRDX+dlclttGVJMNGTeV4oLeyXD2hYzJ6R3BsvrrCyORSMabDcjF6RxG84eaC5yav4ZAShpLf3Zkom9aNRs6oQ3NrEgXVXahLN7q71uQcJLZsaFHTGTw1khiVlPWj4lCWdTS2HDuBEi2IA1gWZ0h2xikabJ2CKUa0OI1Aio8NIGSopfMT2lNxbe+PUOSLp5uFEq6wsiMiJxx0WdHWvPEdTZz8hlvWHB6TeQqasqKpN2ttKr42ujGJG+r3Tc97+P4SFeJWgxukjmosVHfdH4afuYTjHhfE6v89iUX488vaYAXvrSwq3OAoOAbQk0eHodf8tpfyZGoBUL/lL91N7h/nK78AsjjEzJamcwnx/P31ch/5/wqfPQL03O19XgqaAA+i4ZMhm4NKyJ8/zLqUoiOcB/kCzQK8XrPDlQVzllJEpDnDQscMxHhP58w9DuwAeADD7geCPTGJ8J8nKr9vhDw2CDwV7Bfmw2R2KHOn5oI5SQXIO95rys+frGgjP2x50ym8Lnatayfi8qo8GTHvxk1dHTnYhGFa8l5IR+ddV60GmmOOVg8e/kYc5cL0U82bXv7gl9hToExYjNekyLI+t+GhiqaeKpXbysx3Iys03r8QoAPlaOfY+dRXvKegDfUhwWkXeN3HtVjbjoC0lS8Ndf46+g0gLml1x1nmYQa6GY81T5vKRNTLNKRblgl3p96SQfYhlenqflWuAmEZXwGCk5OTnSIX876HFescqP0OSsDPeWWFWkmCnG/cCkyPklxW3H2QmGXldMBG9CXAvJxlG5XuHbL1jQzyubb4OMT7tnVtjKkACNm9XrYYxJZDBUMc1B9ZaxIltcbYl/QyE957VOCYftwlHzzerFFoJ9GkpxjhdeaH7nelqapWhG/OIuHUldNwzP3qJkIPgaZfQnVIel4C+TP7AjRfX1OnsiBx2VtdJPaDI+y22CoIfylQuVRbzh4OmL5CJ3hwj9g2Sp3NqAmwEoTV3hSR2NfQiXNRWTxes7tTyxlVha7Ekpj9cv8dr4gyd4k8ApF09z47OVkMEACJsb9AlZ3soB0+299usBCEK1M4rcby1/oHzl2C/uUO5jLR2RPco1iGiY0DCHSbY0qT/XNwDaRep25LdiqhsMfULZZEzapvfB2cXblCYHvGXWuF9mQOA4cMlmNBSRcinYFUR2V20OaMXbzh+Kzrzaj8gJoczZKq0mdkX933OIeulx06NV6HifAwiCtzBc7O/hwsqKeQ6H/I8xP6lXKNRYyjdx1WMyVZ+z6zOBufNnftuwwaT4atViaJOPMlOM+AOgCyy/xIHVvCj7HGELXIzvwMkfnjmjTmjTLa/6nP0pH4dpH9sZtnISHYUqDRzbeFIzmDX6flNjqfbHZ2d6XVhdlzlYLw48KHWJnp5D7A+cH6aexsmoy5BIt/NvM5XRKRCYGNO1xgxj6PwJJK15tUSLXeuO5WVPBSDm+jUnmg7qtqbQ2kEugXqeJ5qh/WyWs5RyzB1t4x4rYUoCeOJfE1oqfIkBnoEz9Caz8JVsz7IEDREYveemAGL1QkMuPrByaCpUasGdOPYTZSyaQh9eq4hlajDbq19JJfW7m3NcE5vcOWbJFhq2j2vxNaLoFK6/fOOStwMSqDCiSffiYIZ4Upd9d598lC4cr+fSBt4Vw1+El97ekUyox54FGZT/wfPb3WAckhLW0jOnT6re6rl1MNBg4cpJcuKUHkcAjRB6a3gFXh2TicDYoDR5/wjy7fYjIOxTzvNiE5aZzfFll5F45xrii57RuukxNBSutkahPbXjOlON6CMng5NKokSQk36uD6aa4/ocfBZE3K6nwlgf9rG8chBvwMJqymZxpCgF46ph+9ceaza3ddf3wSfD4TZ9YxLb09ZpmihXTZrFXTmBe8R5mpipr6j+h1wW+fwV1LuuAZsJKNQ2iit+FIEe+PL9XdshkA7n1bNybIEiWHPTbFhkbHriDEOgOYUacAmZ6ynkykCZJ7nr4mRCyMeP1ZTiXL+Q9EganbD6LCeQaIRou7XJV8Miq5ozQ1cKUhahApyC2DmifjR41VnJ7dA9j4gyMDOzMhMhCZ273uovt6ovjp+qPA73FP9cYYbtnD91aBvZrFlur4YspAw68AUc5hr5QE2lzoozVFW0xtrSqKBiClwUuTzN8yxbHr1fXSCp0xzXdhl28MByfHvyEbMV/C+NLoyGP5QE+O6buckoh1xGQr7IqyT4fXJ76YqxwWbkIp1CFt4VClHMMGQRW7l9kMDnlfwQ8dhbeh8wSWGVFt2OfcwIHC8eP6vn15qxOEujnNYtDQvZgAw2XK/NlJJwbeC4Cq3GnRke2Z9INkQR5Tlyg582tm2OijHg/biNM9rz/MQZjTudZokH3sxUjOmSvgcOAVfHFgHSuBi58Af4wztarLFjuom2TBoJ3C+bOMuUxMVkyuQvWzM1Dm2MGjbEW4RAmNguWnZEMgA9LhpIi9r90hInIA9+gS9esbJCQI3SaiKMguSz38M2R5VXvfNw2iMHdOzhndZu6+FDIYx04JqYwlqPXkI8ePvaxzBASnLqO17PwAlLUDB2TtjK3k/O1qgRzCuE1yaUQJ2QjAYiVFMVy8p//Qeba6WKKQI9om6AINR3snjBhQMWYurxC4i5BpuRWqRs1qB1kugVOVboxMG+EbqiOD2cRrDxzkZ5d0eV91rhcvWnk6i6D1yNaLTyBJfwdN6A8OPfI5flzu8f+7pfzEuOwlZBj2Dat2ZoxV9Z+UN3Ao7pBVN2r/8m6O3WLZDmn5NudkiF6Hv2A7Dx+dQhfboOZCnJZIInaf8yPW9ti7sKBwBKYwmFmWhO+BuI4k5bynwO2hqJkYlPYbAZPEwmXYReiUcCQmQO+lCyeBnNt9lb+xZMCZaq45sdzPnoNYt4aSB+BsOghf9mhQ3jc+MBycUIN2AyrCICyhMT3db/0LCrVSqh/gKse2BN+kBqHsXyXLwpMUhDt/myFcvSq+pGdH1/u1efNArCMZ9TgkBu1STH71gxr7BvQ/zCd7PAuLEmLz86qzCQXHDltLftltsSq1yEdzbDk95uZ0K3ksUg1Tm9zbVHD8TRqyW2UWDEwd+z9gWCZgKxTFa67XX0T3GPG5G0KRTl7O0WDKMQbnqp4R5UUrcZKhEp4tE91HwS8u5UFonYYVspDUCr6CYEaXbXo7MRqy+gfMN9D1714RzrBivoHl5GjEIwKj4EdsbrtqnKK88vCYf0PsrodBLh7zuS2Fv++g74HJjl/r4rRd+5d25gepa+b0bL9N/Fmxox8hQ19ORtIBLR80mh8/Dcr8cNQ4/xGrogk5QQoPVWRz+SH7lKE5fvwbizvP6y6T46me8Q6opekd/KVb0pUgfVCkK8vp3MCyNY064Z4+J2FAvMW7TXUhLSez8WiixIO/Iwu4OR3QIik4QVW6Zu7WlqYpvaTW7CT/cfLmlnIeBxPJWP0rIpqsK+Qv81fakVNo0Uxdo3G455z7F9HIbjC0oxGW+pgd17MinIpsonF5tCV2dD4PNywqPMBIejH0F7er6ctvgPJKMAJqG8UNJ5j7+rx3wBRaIMhzGxUFtV1bBJ0ieg1m3bHEh962S55zU5arjMaiRlwtbTujzwG8PatWlX2JzgnnCqU58g4aQ8po6+DnpZMmrWb+UNspiCRH1XfgF2QShR1xAd5sWy6fcDgO8hnu2pHihoqU/GxXYFDSjLMhMgvArpMdRY+t4OOKWGTyH5jT7inEDfMpDO91hUKlJShRyZsgFSaLMk48EErD8BS4RzTSaWueo0E4nKSW7EkyJJ5ooPmh3CqwlZVxuzBz4Yn69s42q7nNm2lqYbuZSUiU2cB6ZsS2V0+CpgeOajyjQNi/efLlg1Q9IHjLqg3OfF3TXYDT9SvR7SShkht6gtWnvJHOA9urnRWr7fiUOELAQeFIPomg7DmRwOAm+YjwHUDCv+0q0OaZbGUinbeXCGnizLv+r2xtcodPQnQJXdLWx6V/JueTrN2AZCss8f8GnPEA62sBDKz/EEWSDR4hqmgoUa5Lhp6aUWtoXnpov3XaWKzZG5yfQ=
`pragma protect end_data_block
`pragma protect digest_block
e7131c8c6aef50642c4e552596d545deca8e65e56267ed6c2f6064fd3b095cd6
`pragma protect end_digest_block
`pragma protect end_protected
