`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
NF/8jHLpDC3amTDSH2FqQF5UT9OO2Dr1A1DinNWpHz/Z7Lm1/ohsx64S4JPOC+CLf3Tp2JJDRkXsNVwl0yhQF2uak7W9WyCDBA7WDL2R9TTtvGYYrXJHCWktYuZQcYtekL2KR6Y+DPb24TPoesBAnVp02tfdppU05Ayv6OPZ/e09Df2TxDppC9wgBEzJ7WRY9IBD5hp3NpAzF6t1dxKtggexSOhB+jwKi5187mWBupsym29ZrWQ3Bzp0N2DVX3LT0lN0R+M8/JiI3pWRhu4s4pCSvpp9EcNjsw0wVFDNFnF/RhjdeBxaGe5WhyeMeY/je1WdeFXt5yhj34iuaJJEu6CjW67OcYuRjLRxfoDLoBDpfSlpfgoQFxyuj0tAGvDlmKCUuS3BysaIrwBp8nVH9JZYdILLrTuL+MaLDdQWE+cdXAh2veVIs20mw2eOFNPk/+XdNoP0fBzwDDGLrY3GYgOQfcMt4OOcEgo8H9W65mTmCiaezYTjnCaaonnmFas8Kcl2Rtknw3V8ZVUiLd46nlRhIBux3nw7aFwWbY7SQXqkzhiunHq4Yiw4FKGhumnZ+XwuwkpzsxJbBx387c242g6gXr8H5kscdj+1G9HrTAp8xq+9hKx9OHa+6WYOUzl4ncAShzThfvmVdcuEKI0/BlRN8uzCvOtog+NX2eJRT9EkfrZsPZpj6KNgg6JZMSpp9eXjOrfu1HF5SyOWo0Z4/iPHcikmwoyjOKt/H/p8Dbcohn6X2/HBRfIkDnwY11clO5fyyHl+V3SWc/5i00CSwsCHoNcdxn66o0hW37O5tE2uadTYjqpaC011w+PDR4i07DNyVM4actRf7bxMyawwPxvYKna+GVLa4V/sR1+0weDMXhKRQ82iF+CCJ2Kd18pD4Tkteh1ednd4xJ1Y0U4EUURyPMi9kMrw7z0kv7PyMQqYZ7BgCM9v6DyNezc3gJ2pIEcCOam3AB572SCsRH5iW5iDDORBrKx+LMvx+sMFse2G6fyu7roU3PR2dk+Mac3JqSu9xfnAwYg2StsHWKTDMqaCgUDUA11ehlmYoc0yXQACWl2oi7T6FAwu3MpeIxHuybXqgkipygkB6siAXRZg5ZjUZvp2NOCEymEUwYkKUGSb9IvJq8Q7Zm4i4NtJKmzPYoPltYusxA/QVtYta7AT6/y2aIfJ7H0A2pZRIEJqQ4RcPE2Y+F1aIVhWeILwYm0AN+dLM6ic9QfvZbXmRslGpCyg7hDaPTonFMmz/aqQsXh9XU48/lW5RTFiTIqD7Z+bZKrSb9e7o4WGIlcftUo5wSdj1sPQ4vWd0sUNwKxtoFqu//A1elW00zdNPoswSkXdGRailbfa7s6HfCPU4wTu290jMpqhsvL7GJEL4T1W/CKMlHSEj0XG5Rz+lvhdWvnJCgXmf+RgA3sBSFNUZ4E8oSppw9aN4uvuGQwOB+XxO7E=
`pragma protect end_data_block
`pragma protect digest_block
dacc2752a3ecaf8e5e37a652848546b7d091b4409b4f9a23fcd9e1b58126cd79
`pragma protect end_digest_block
`pragma protect end_protected
