`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
jmBrba9VpzoMWYJkyZLovfn88D80VXjXzWkuMApTqZ9LTxLwLvwYnDgvZIcHUKvpcUWUgDnbdu3Dm3qbrK3emXSjPP+ctwIh8L0A+yOYl0U03+/MvCz4w/kG9t4HtAAvN+WSTyMsdV9MqTDcvPBI9TTR6ejXu+zYvkurgI2iQ/VNh8WtM89z/P/58Oh5/cOoc0/gre3rLpdAb97afcm6cQxnTrxNgCX+qKcb8TXYhIvkKjvJ/j28uUDZbh4u1zOBTIML+SslfED5E+8MFeW9pEiLXGhUtNkDgcE8sfGG0pubqPr9bwiSvwhFzsEnFVHX0ulO6dbE/+ea8ecF7soQW5gdixltaljRzZkpvORjKU4XWsY7wyKa5oZTvFzZl4mczSPuCkUHko7dxVzw0h6qub243oYkkSyKzCqVLpaHF7uZ1uyXvlgTCSX5WTMEFUNEpRY26yxRszytIzMtt6kAGDkZkVPV5IOCjva8BwDbGC4vpzmmNDRxBx0YLPRJyut6kpCCUiLWHQAaWzlyCOIpn03bQ9bhIMfxb3KGLr0/nIiw5fzVa0YM9t0E/zri/+DfO2PL7+8ZllGqGgY4PWD5N430yC2+HLaqYGt2iI4oKi+uX16Rt+3v6jwlq29446EOdys16rkCUK2NJ0qnRMLrRONxtFoQgyVxNTt4AGqqP0OJDeFqehAYUdMqzkq8ZUSHuq6McbE698cwi2DKJmc51Jrok7amEg03fbArzcdDAfFv2HSWdGBRhc/7yHU8UqmoWCdmyJ/wnU4p1OrctgbIQf+t1oL8OBLFmDaxU3/rsW6nhwstBmBFUL1o/KDIwHg0U4UOqOq8+f0E7wbqruUzA63jfQ0OMiH8qFkOPt513IDFE1zd8jzIRbE6dTZeJ5JErLo3e4mGNEG6zrqLkBLE9ZydXzS6QKN6IgOocZVqdzSN+dP6TuKsxyZwZ1hs5AcViZuYTtzSNRAVJPWKgjszkABmHPBrj5JyOQc/jDWV20K65HwPCqHL5OlDANpAH4voGLurbd31hOJY1tszg3JbXNuAi9QcMvC2CfFyVypsK4k4+KGqsWEwcOf/1hb9V3/GOZQ8eLyObHef6U1sIy7wc3wZ0U7r3PlNArn18XnBy1hgef+wBn3dFYjBr2wkwJOvCoyuleDhYFhFL776LyjX7NjbdCBf6O6vwXRRjHsTfy7ZPL2Y0/EaUxbQFIBjAruIzkoASq19eST2nODG9C0mhnjHDq5fHKZKbKtliWdtvMRHRIUmVjgQSrpmXzQEA2Kqs71BE1VyDe/xoZovBQ+mRBSCaGDxplNbuHd/Oujhpme3fMF0HLpxn+V0UUwBWSULShj4ehmD+cg8iP8r3tq4FYbVUU6UJiEN9Lqrb4F9w2XqaMUALnyOaKAGEi5pA/aucs8c+ScsVYDFt/23FUy/nvmhVk6lRVqPtgmyOUxhQy5dPn+w8A9WrR8w/DKe6N8JDtUgDbWI/5s0XxshxPKa0VYCF7LLIMs7DwgJNQa2jCi3SNmRS4jlO363m1HipYUL+bLfEOTJQFw//d9sV4woxGKq1LWSpQPesc+Q9JrT/YlqqfUpw1fM0iCWm8u4bRuL0wVXj8KwzwAtAAxZSlpvbCGqOrxAVQyGPNOIOrfT8/Nj9zfjMnsy9IWn5ocYAB7AoxV0Wpm7YbVlS5o+TbaxalBssgbWd3STb2vBM4HHJF87iuyuqj/d38IrsTFTI6v64STiuhzq8OHP2ycvw11xF0hb0MMbBGZaJo7Xp6EZBlgDjCrCvFwmSdl012iS7jfFCdwK+rXjdlWZZqa/hVWKDb5Qur3OMyPC8zd9klsyIoNaJYExS26fFpjQByCde0mWvbGW3hQ9SnLPDzMTofH+UnWti7mt782kthYCH5FWaMDqn4YrB3SonJoMBjehYj4GODn/RMsNuHBdBfKTY8jYjgxoiWNs9dARx+68KvxJXJAjNEcnZS8089h1AMvnNSr6UxptdFCbGLQvlSgkzvXNmnsm4+5GciAuZTY6n43h6x7WY3mU2eaOsVWj7+L5X3VTy+4sc/Pfke6/Lchqgh0qDco2Z2fqssyfk3fArkkDGoQxO5FAnPwSSRdkWjbBGITV236mymGoXxnQcRzlaXZAd3a/J0q9cSGRmfnMRbAGNZ++iKMaKR9+FigC4xUEAbD9zjmPGFjGVIGZd70vZ8F2gN++99gPTiTEgcYNl4yfFYK55Wow8GGpBCmtKfsSLMnuM86biGpB5oo67W41bE5XvnptCrpZ9YrT7qTbEMSS1E/PDQBLVnUvP0ECe0MKlLprI1k2BJNvUn6ebz6PwXbf3lpLnc7rHq05/ceg17hetunDBh6uxtvN8epWN41QXxyLoJezFFJoZxeUNJvYWNbJVNIV6BlQeUw2QloMhGjK1JaeKrDbS2yC1hmkmG5Pte/auKGb+KdYtRQz63AZiAVfqRwU5O452BYMF39LKO1WcluAdBa8aERQP7fOGaynPn3GQJjAp4NNEVYojRFLqIJGj8tLmMEjWHQicYI6KZuCfRKjG95R1Mh0n2cK9WwkedS4nAQU7uVa3v1WNvK1Bi6h06QyL5As2iuo0/KIOKbOSHDy/2VInuipU/KVwAXoHesmglBkp4r2Xt/rXeXW8CL6U+qsUifSVza1j91MKDxjYFf8Iyi0JCMoDgH8F+HhfP5yYEEnzEvEoZPbA+hK7UzIQTbt2VvXGKtLPGumqW+EKcWQ7LpmA8rqb365u4VPEbQ85XIwmAF5qG+lUtxUCld27qfW59T2TUgpvfZSfdJUeU37wBxaWyzgKSqyPWdOBkuBrjrPZ8HuUTadyjsUzO5TYC4ASzFjXfcML1w6AtBHd+tdHoyFmU/CNM6KIQPg3gtmG2xy+VF8d5hPvJkTauETSIEQu0M+VbG+CY8XweFz0GHlXmT38dg4POhW3dfDFvQHp26XUaACGIb+poBsRO6o3gAZ4QI7Ve0qKZHgfJg0benzznwkzW2Tx3PEcEc8zxXOieP8kuiin5k4JTkqY+DoE+zAUEObtSar8g3FYyyoy3+2qOIRVQo2TBtds4tc0HtIjc/Vd2W1F2hN8r/6/XR0jVioCC/OvNLVEgXcZ/MXyDcaUHMmIUkLbVgH4HkrPwl1rKjwuzgpc+wtCMNLy9mmnsZx4hNQs/EY85IOzsD4DsP2SYiXdUe+VLQqASi3r+VxRAyg68QYYhJ3+TxnvPdZHWMLtjc4vwGoWrqSo+tUDai0DUe6JjGBAQh6PGS6j4sF4gUTvup6C3JcTOGOmTGU+SQjOx2dQAaSUDpcqFV3ZlY2nr7nU0/6iykTqGHF+1jmLmNwlXO7sCi86u9UehhEJFN1e36jRSyc5nzI2qqVcAY8wFDDnirpoZOhdTLzNhus0wNYi87Am6qK+wDvzFf78OEXSIgB6RxM9UXp9SsJbffrMwa2Cf/KbSoKXxna5CtohqLr8uQGLRL99b4ETal2OP8L9PAx7YmCdPWZYW+ktFxIyJ2phkLXrd+D1oDqw7cP4Hloij5OxhMXi8Qlua9o9Si3szyXQW0JvGEfFYBucvpb6nPcrqtd658Nfc/U+uEbCb+L8y8YOsFatiZWT1OCy1wXCqgbkMk9NbwxQ5pUUkKkuBgUcwxQ73uq0NCfuAWnxrTpVmDq1ax/3++pjwAevW3iDivxgKa0vCByuwcJQGXqnvZMs7EYVDzdquSlT8nYBJhcwttgBrvIFSgHC4nkxmfZmP8jioV3DVDJfjErKxZHHapB/fwQwOKMhFVIohROPSOGAGFqEThq40vl7J9Ho9ke9AaZ71MOHxEUHqvvL45iu7bq1dc1pniqSrlfATGKfL87z6TawjX+wZ9aXduiO9J56dlsPrN6UhyPGJbCnwNsaArSWLpqeSQs+5vbnQTlkPyVskXQCrWhOmt2FT1lTVtxHjdvq701ZlxdhDzXLOjHl4cqoZ+BeNQSajgQTE1rPE+0NdFHtarLk0dgCNgQgLWBvFRGIpKOtmpp3KY7uQVS++BnqrYcF3lpxiXbH3rBE2+ib6Xoppz7x7pCgYVcG6Lczu0F+Mdvckv4lVT0dvZF+9jWzVvyzqqL0te/YjzEG4n0OFSYG6ZCbIU+xkVnDeDRBbvxN/XPAhw7S5AYaZAuQ2FrZs+uGuImo7qZhP1xXlVtVFVwidQ0PhkOCSPk1yIy0gGzxfwOzlpoxERhAtjuscxg38YqIC5pZDFzkWoDctMvDbZtKhFGjlizbcQGgEqlPGPj+jAv3r/2UUXpTpW4NZ7GT7Uljpxwu242BoiCEnltKMuiBeLjQXHh88MQq42yx0bkNEIKXr2vwhv55s9K3wHnaRaM+n0ojnoz75Cry2Q3LoM0zEq2MZs26EbAUGSHPAPBWVfTSx5n26fQBueuwfrRBA8POdzrLnQv0sFhHjiMDywrD9NuscjgcnMyrrrvYvfqBtpQdEK8dAvyUJuj35K42FncqpPcgsqqR9uv7zwk/o/GzcF4ZYc3LfSZ/LgSvsL7ihWLF3Rgt7bHL9w9tVqyP73ur5bZFJPzlXFsYqESi89cNLmzFU/62wJ7Fh1IQxzNcJ2cHh35AxCLdUzhSeaA97HmJ1mMPGbuCgR2ukLhj93dDQmcnJ2dJDAl/+hf9OiBhwqGT19aV4SsIsxK7wCbRcD7f1VdAVnTrDTrGqFCY1vgNelKo2tn7M4FnCkdtaG9sO5LjV1bempGgZxltb4s569b0HkY0rQ8IN3J1x51mcAfgqeHguuugeFTAwZ8ZZi0rh2wd94rXkAQj4ADmztifR+fRA09AOXsY3hH8jnHALo1A9hEZATTyHpbrj0QPMaRAXi/Z/lQWaqvYKIwTGWl+wv0m85yQ3Hcl3CxYcZ4hJ2RS7cMUSuSCSutcQrRA+HjG0eTWGtTuyqde9ONbQUV4CdgvyCu5M1bl/wlb0CsENSkltWawMcCFkA6cZ+ETEUShU9qHykhBCxAq5Mr4H9KXt0yWmiFnG2HNtvgp3bvkFDENeN5mqZzjJob4BPHElrQcAwYgb+NucXb93qbnf9Ftkc2tdeJcHf5kWPQtTt/PZBtiPH2AXJb/T1A9qQcoWwfIuhFF6iPcriuz/igFv8FX2SgoVKLkVnqNru0Q7YmJHZNNuJAxhgomDt/rY/WFSNpPpv801AEA7naOqKW2yC59mb/aU2Brz9i6RZxPLI009/zFQdrgXu7fLXi4PHb0O/x620jM4dTDD2LPSrTqVQKXiX/PhtV5W4E2a9b0qpD94qRu+h+GUJOFGaG83wUwd9RV5ns6YV+Ho+Ixi8PZOzMMr0gs9dTFTaw8zE2yAbvnU+5Nj6nxStrPRBZwKUGex1rabLhsWLLURAF6vXsi7GYmWEam/sNMT/X4lh6rCrpoJatUM88Tg7Ivi+NzjNX1UG7SpZqaYs7/3JJgKX3hOaN1O3c+vaieUiITgXL1yvRe/oyvpjBymO2lkVrROOpXqpSsr0Yr+gSTheC5MURuCWv6UEFflelHlKXUQGNwlKuTLk5Qn6bZ1vKslYX1aXYSJHxJAuGXUHF81CNO7/BOGHPbhj9wecITDz31Bk+gyo0Krz3y8N3W0nD35mnomN2iGWvL/3jlys7tWjAYfKgELJW+kO7AfQ+u4R1rxH2jwLKJswaK8NIvRsb9GC2DeBgYJm1IB/NO8DhuFjLxMqMsnj9BtzFdt1Y1m13n1wCDu+Gk8ObaznabAcWgTNxqhgW6Rces30O9lA4qLMHpeWddBnheyUDPpS5nt99P+e6d3JF9vuFSkMp4lQn6u34CPttlPMwrAS4/xwygHVtmx9THx2CmO0QCPsKYpImO2M64OB8y7N2Px5VWkGTn2SsMTgMZeKOPTfOBe2LvKXL1bTAoBPBGBL6pmKlLGndXLCqTK92+xFGTnP7Obtxm59JXkJemBeqdMxNN8WotmLeEGiXAhld9pbPqs/5548gHrmvV5ItEbagkzvU3ZwVVGrac6MWaWnPE8MuEmy0yTx0JZm89wAwKFXK//0vN7T7aKmEvSWXaj6u+ebWbt4WwI661ANFOOg/RXKvBwrqJOcarTMY7bjZGVNCBkorGodemQegyLd41E52JQkBmRlwAjV9eAHprjmihal9bto9hegSjzLyQeSArR2o+Tb7tV1kY0jygYxvO5o+Ix4WgfQhiQfkLAJdlpaeLG0tlQlXlAToYWFhgfZEVJHPkqWGiKlzTukZ6mBkaJ3jKzUtr6mrjn5J+c+qBpaXPTWHr/6ySsIlzYH1VTaWycgGLDOF9wanzwSlSG05JEJmgHpYTRHFvkjBIBExLdA5pw/fz3DnESi+Dv9WvOU/rIjVC3dVegZ9AMs2HV9zp8750EHzBt7mtutVrHdlejN7oRxp+luSqWeVmj/fPcpOtbv7V/umUzL/avoJ1DQwIRPvdn6/EgHGirvyBELO2vBrY8rQRFNC8pxO60HRBoO68SZv07O1XZSzfxETGVe1yxXcBwtPfkAR7UPt5OLYFMX55UHDGjOsdEZ4V1Q1J8TNQhBBvcOin13YyrzDrbYliRGJLbe8wFa9Ryj2ElIw7xdRxY9puj5y26NFqXITk6b0VYeReuXP4VBzrOhW8yEvdN/wTu4l+rlZs2aRQbtYHAB3hLjVLXgFg364vkBS7CgC7e5mSf7Sl2XSVxq5B39vH0dqNu6c42B68cVeWCSO4w4qNC8XRqmFHtuGbW0ujUKALpEhAgnS8wVTJoWdTXt7HqnXBFS5ekQNnvH4OIBwZW6ivA/2TP4HsEPGOM/gGg0b2ymbeuPRKIJW2PSIKf68MzH3F2D35tmYgHJiFXxxEcfyGVeE02S6FOwozW3grYRROPsUFwcnWaGatyeF9FdMWMpNoec8HXPMeyqAI3NLTvmt+DlTD6D7X5HJohVoZMJ6SCN6UJKuF2ffJVelzvFBymZK1oKDyVvjNGIHYAAmD4+E9ByPwI5rM+zG0cX+QZdjTZ3Pv8qzdha7m2CoCE11rJ3lB0bYEFV7D9Dgu0jkeeCtjvjdcDNrNOEeEpgi0VSlzzKBA3oMSyNu0IgrifvUW2GbnNILndUD8O3pA/wZ3CmiEXWbUteH9iZ3R3nbXLMMK/W8L/jq+k4OklozICOkHBpdrE6XUKsyB/TvrpBOeW8oFBuDJSPBXg+ayPxqd+/xrcRyfAo4kg6F/Pb7wwFrZYoSmTa+43qJ5pUOogLDP5OLf+PWZM52Fyb1YPJCVjjnI3O3C2Q1qnk3pZze5/CyYUqOaHmTwl8JQ4tvqseLFEJWpIJGBjdSJrHG00YR4yf1Q4RWrR/4IRDY0Zj36O/Re9OS8zKB0q1WwEHWstA3TUQn5ulpMwx5RKmIhVw4Oh+kQumuiQNqX09VYLu/0C5KPFIsWxihHgjVBUy4oWK+tyFiv+IsMj8J0g0ehjl4+xpmMY1ESi+eseibCyxiSrlPPwVbON0hkjHmpa9xr4QaLA5JxPGgLExIA+/QvWcCJ+9R85Kh+ZfVeGXO59edh+sOEnvC/CigOvE+CsXPGeKqOuTAPGfqGTioK7EGiFqb3k8XixgzI9Gt6L3P0c/AQlQZCrqQTxSNCyR4VDst7CEPskRITplr92D3sB8OMRYmE7I5RrE+N/SSfq0sx23ha8v5rQMe2DZmUd1pbYkgmdMm4GGMwsH8+8viRE/vWS9tZFwD5zQPz/9fQXOau66vEsqcyby8Kt3NNrFrbkEYYr+ZJAlJxCZtMCWzUBWysiYAp34f9HL0FdxpFwhFgW6DJ58CUC6k5UTEXMsruYqTHydHr+qAWjLYsW4vISWeZsWymjKcgd2A5QS493xoVRVtqZWVTk709SEAlVLT+ZBrxe+VrUNeXXZgNuZvRl7a4FSY5hB+arpVzaeMuq0+VuFPHmJi+k9afaGwz9FHeRKltK+lQjRQhbr0VMptzIWnTyDJaWT8GQwqpz/tViam2ZXERF+5OUytc8zssf7wyxQPZLMI9qPHZPPBBkY7q17QmvgV+l+8sMEq/8ezvNK6qy/8ODi9g7wmzsAAyFCYxOxzdB7QyrSALxuLUs6ZTJ6ZuF8AAE9f8R7DBeO/wfo+T2szkrLGvpw1Xa+S9POkEgb4PdzmylOnEDtkKzrkCWrX8L502SR5OEbPV/aQrDHtjWzjhQI6j4SzWMTkh8dAOvY7EoY8Mwmxk22slfCu6b2sKhZZ0QFywLHR1mGnnhmvLPIoFhE95fL74iAy/AmdOxVUCNuCHWQkGLzvAtu582HOAcJEL8BUsrZzavju4OTgvGRIXZU2EtahQuRMRgjHrnHqeOZAHEfvC+ZV9INsiMK1jGKllzmklbvNUhLic6qPGXVDaymWtu622SfOt2hyEuHbEugx/7LAfmlTi2bzdX7ijocc92AflTQhSIZcOyzl6utVsUWZRZDZwqvqvf0lGwOCSXu0npZbL4yBeB4Yhvk2e9UvjLyXoVv9cp5gBHvWXEn+2puJBhG92zAsCfW5hkLg+hH8mXEMDrJDFkHQcuhD8ZLBhasWTsO0+g0X5DzkPxVzlpzloz56YXtTJ2akhbWHzV7DifSXvsolMP/SxN17m3oZCTh5NTfUcVkBnHDCIGuL6lIVL75ElH9nXEco76H7U+VO7Lv5nwlRxhldz4r4PBk5EP1bXjWU2oBSmJq13oG9wUZ1lGO73qZmleu//qno0/8/snefwyrbKiTOUK8KKVfU9uTu7wxju8pDUW1Rn1lF72MVZ8A2VAVBHGVuXSkHUyLZi/s68bzb4IBdy/04IqRLyCabRGRRget+QA/Yrzq1rFmi+w2s/jDjYbLdi4uhIx5W2SO4ssx4gnIsOoibqE9ICseBkw9xzXpCWPg1VWOkyh5ivJSs3HrBuhtPxDUXqxEi3LS6EgqwSs1C7uTqSCyNaBzssNKO9OjCYXNR4eI7JSLJiXPrjPKDsSJa2lrW4hWsmwhADzkVWwoGTWsxPBPoDTimF9tbqiYGCyCnRwpNFi0HzoL0ZEFAlynOssDjJIoHtajatm9lxSIFTyOedee1kgbpoLwZYjMua8QKpQSrWYmV9Z4DDX1QGvRO6uBJovQZxAdZsBBV8QDXqfnKwWsNwS+QTqJTPk6qJRh7RpGcZZRsuQPECgjMdTd1XfBvMSrKj24dXXj8key3sy6E9H+eVVCiMSNJkxJlCI/z5L5dqR4SD205/SAXupp1dJb67+zyHa/AaWjGzFg52FPOlIIs6PISWiihdJm7Bcwk6yJB25WvYJ9UFTzlBIYHgMn4NR6FXZpvwzkQAvXeQp/rE5QyrzaR0v6IqcKXb6DJ+hwcrOsujYRWcNHNfb6Y0YzJtyzD6fPjFPME6pGSnMBwhz0n4QUjsLp2MPJiWEvQpznQyx4cNEnBAR6diWI/HUPV4rWHVsttyfyM9aqs/la/nGPFKjsliXlX11OLq19y9Cu0fA5ri0ghDVUrPzSHbNK9RFGcLy2nvSjeBB8hYxdQsVPRz4U/T1EX9GBbNtaub0rNT+aMLRWuPmOQPUj1YO0llpQDPkwBxfUcuGLT7MiLGvzEW4/wmWu9R7LxmDxf3hmzUc5GBXInWpn5vZAYszEUXZWyBbY4VJt2hRm56CPZLDi1dmdZ3YflnaT3Cyo9LlsY2dZwkrviBAn3iYHqg1EMyKcsOZnTxGjgHUPvmpXm10vSBkMFxtca0KhxS030CtNlveBDBRECuGIRvv+xIeWKhQqj3SWzpL7ANOsXdihGrVPoRj6SAOuOQTFwdEVoPZV9/VcEYYKbdNZoOMYLpDQNm4WLkv5akDoKWbaO9fXBK9gwY4XmEFDuSOHrPOs49sd1bWVZP8Qcb8shuONbX56uwlsec8LACAu7c8S4VHbFI4z4EDWR3iERDeENxLe9Yb+wYLJpT/KYjHrmCU2Z2PbNXbkl/P4y3sUQvnQmt4lScrqcwqMCk9hl/eofSRRIzdY/46JEl9HhzoKKpnRM/oIsATQRewD7Sd6pXE2NTAt0XyrINftyJzQ6F6+Fwd8oBU3WTIFSmU+UFGjlxNAYp8Mt1UiILZHwCwog2c7DWTfi6m3AHIGCto1r0gKr3AH+yAE5Bi+pYesnA2PQdJX2nyy3j0oQ7sk9rXqL02U548jgKIbcgkWgd9qR0rGOgVPsbYUp1cOqfVZGNgxfucqfPAHpK2NDFyikSPTKnmBuUqyy8op00dZ6TRzXN1lE+/BB+EXzM3dRo+E6m7B0aYIiYcnRpI3TazBxQATTekje42k47NVaF4FW5go0KsugjT+ncUii3wfIJLg7FNkBOs4qvGqWyckUvZkOZc3K3YEnOBs12OhFBR+9vMuw+ztc+taTINbOaiGKUBxWTEse6iFKQkX+ufi36e1qDQ2/VwYn3i2DoRsYsU1uQqhR7GakaO/iGMmXfoHpZQ6mZZ4tZvk81sri33FQwz2j0aEPKl4XwkeFKCT/q/31LvxED4BwXHg8gz6F1TgA5T+2asYtNGjAi+XluazrS5L1Q6vgRfNCS5lEIpBrDiDWZIXqgYk3mt/zQMBqHFwLmT5UN974u/ZjAmqOIDPkvtHIiF5omBnHGsp/O1q7VSX6JrMXKv+2BUpVCz+X0ezVbNqVb2CEItMiXXeXFRQ7jT2IOGYQoB63dqQomezrLnz4JefD+mGRUpWjxVAXukEVOPNdpI9Ur1oxqfGIB6q7XPXxnJm0malStXeB20j0F/oLAgNj6DuyuqycIedvMrhI12C1bshkVMsC3to3qJi5OavcjxgZBNnJ9pfiZjBlULCQSnexjG9cUKn/4I8WZrw2wlgGy7tPhG2Zk0G99N42Eaj2y6ndZf02nw0ZkUWM+eYD5EZWClSu2MgjmTDlLhZQCVqGbs/vEDKrshy0Liv7SYbMl/UgOOOOCkn9/dDWgtevlBhDY/jkLgQyN7CuHgTr0Q56P74oHcjDLRp2DtvLFHmwoA7t2RVNL7LUPNK3CVyfluPIemHhx3aCzxD5Cg70iSFdq7gllPHTL8pg6iQ770BL0NRxV0BJKfkvjEAehjJM3jj2Q4AGILqkPC7GSIx/Ri61abYOAvlYqQ87uYT+q0BHqCvWxlTbMQQWuuKyRTHjKJ2RlJuHNh8QQHqV+8D9GR/Q7GgpP5XuOIFn7Ui8tWcWsF/9eUMuCUPLe9dSa+ny1GL/cqN9nNngzB48qzOHnwAK78h34JAWLdyymtKdR8H3ayQFLs2UNGoi/ZNCczdk6+0Jh7YVi78KX/gAB5V5o5yfKhK0b+aGMB9PH863OY9cyummyxGObzVDYA2Oo0hPFhai+1aD47JPpSOcf3NSkWG7Q+X/iL3DnKFgI8qBM39MDhGu/kt83JaVs+bISgM5J9OwvpV5Xm/sNFHI/EPLyN592sd8TcmWvOawyCrRlhqIqp2bhbvxQ7wPk7aRFSbcUTzoqH0a6L5S1Lc6MDskSHml3rS1sw4RcPxN+yNUncwJ97JRE2Ph1hC0M91eIoZ7lf1bJarFoeKKGdtAbsAmE3UViz1I+GNpjFH/UmkNMZH5rDQsIDWmMbSUceMiIzcPbX8pyCMHLotxT6gVFy9orwVWxO7AQhx6GGb/SsSF/wje9+64zfmxyvTTp9PdMHbfzdFpsJRRy2N3bQb6wX6A1Ne1AwVaE+KRixCnP2/PFv0D90sxHvPip6+ALTNFwesePC4UPkT/t0JyLGtzT3H7dSntMhPPDij+xRtAB6a5KxW89LxFxt+zR8TDwaB1xDuTbk3uHbIpWExwTqovwXmuQ521pUZ7VWlzQHU9Hlsbh/enzQckxiLkFiTucQyL0rp33WEQFL/yCqNfbKZbJdwYZae82puwlLfFzQdZIaPDHyjMatXZIf/3/5qWS/rvvxiYFBOLvOyLHxD5sc/y9xDATILNysivYdBe9SsONfMnD08h3GFTrvT742U1fQpu8RVzCFmc1txR+75gtSD13t19B/H1W5OPNEpWW22Az/9fxsMLCLWY5cR6zzzQSF/b7U6ztpr409U4eP5VYoIPCx/Xe5bmmnsApDKZWmPRoNvddAWJPMkyxnz/SAyRWoJT6cSp2Pr7OS4zUeZLHTbOIZ9VWW0t7FdmNwtWN+jBE5mR+f2I7x8EKi56xzI1bH/n1UgUgge4ZQPNrHK0Xnw2fWx+XtQSQKKfNBn0k80EgVIwv0NfPs5ZUl7GBxDq/eOt+8G7k6KUqQPIp+/p6DEcg256PZrQWLR9EC3XXxpGRYUZuCzFn8MiJl35XvPgc1VMFo/hHmJNFUh3lzqKwwVeQY+XY4G1gxSs09iMtDf3Ygv/YFXk9r6alpmy6VIqrGeONlQrvd4jy6UifkMNoNVoyDr6/SNCcqP5kD5ngAzB9GD826tIMzbW/NI7MgE/0O+5FDH1jDuxF8rjahkVXSi3ZKnv8Mg2iTTyMPhKCCIMt+kCvtJBwmzFlw9EhAexSbrgTrTpOVqUylAcWRy5sQHJGprcscpHI1SqfQJhloLtJ2rV7a8/rH0pPeBfcY1KZNpNXqHVFALmiWCWZCdyvPRk/FUzFFxGdHJzZnEt9/mFJzVCp+LrBjLfdeNrgMsyXhB42+2/6uIpJGzyUM4o4fK0JCw6x1uPVdj7/jq75amLceGqsuVghNmH4HHyZzKwHJhNXQKPOaYTCk9lhqjB2KYTZuY1lOsdlUggniyCnIlcAqGuQ82qVEnY09LvQP5plsh0JJHi7GdaoNQbn9RWz48UdWClQJhk8Z3CEVRwLz/2SfYXevY8a7UlgfnElclwdavXK6aKpWXyPec+nL8EQAI3AHURpfDvZcy5vMSEP7GxIPvLNSseZlX96LMA6GWzyOv9UKKYez1/JqNG3f3AvIccoCYUcuJAdHa2gI0Cqa7013ge7z0dgy3c4bgSTVt4NaA=
`pragma protect end_data_block
`pragma protect digest_block
783c50feafb301d8f0fc68ec190abd1909f54ebbc1db1639ed7b1bfb98e3562b
`pragma protect end_digest_block
`pragma protect end_protected
