`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
FeyVm47Xy9Lk3std/ffC4trBiBkOscIET8bZq07VeYjmFEt/IQx+nhRTkYIEX0JAi3nsm4X2uuyIjpcDFeu7IBzSgT1kANfrZztqlcrYtGdiQebkAZFf0WeG4rT/mBgdEB+OEfddlPqdTdpQl4X0AbWpEkUOnESm5HL9YM0+w++148HqzDCj8jWBbOjisluBLD3kmiejM+9alfsGbY9fgpbCM8daQlaKd77fl7yZW01QqOiPX58TknMLkMqK2wKtE4NAn8HgXLutXxbEf8HMwv59QlfefQnbjQYa3s/f9DSyNQvC/HJAMr8x7KsHHnnm+9pR/Hvlab1g92n3ixnM43AAYlOOVzR7z2suxIjEZNkFRBLbXhjky0mCpl2LIHGGmeL/P8BLjax7tRkgYLhjEjS2ViuPVG/uZ2a5zcztWVaWj8/nAyJlTlbaIIIniyKspUwszQwRcW1vmZzFJtEJBNJH6WfoDGb/d0DjrfekKkwmRFgqYBHU7kvB+1YKXKtI1xRZWxEVcQM38CdnmqBztB8om4G4gUkViRwWwCaIrGFx4CVx9X8fnAxqR47OINrCmpMQs5cwj22Q8vCzP1Z2ITwPYXWPBaw5TV0utRFD4RRzqJBGb8Iue/flXfwrfu/jNmSNHF+/pNtEiXqYcRzN+DeAXIqzBNpmaC5wOdiGwwtMn6GYU6/MDAuOUSJNiqDMS9GtUbYXr/gIwf2bDgOwl50Ik2OdM1uyg+MzSyaZ23u07WbzO8ZHRoEVcIPE/vLpeoGF+OI2Q+e78jthsx8fyDmVvW5DaCJIBPlNc9C017fBzw+oOeaNq6WVKipf23YGAY7ecoL4kq0Dqyq3C0UceW0/h8C/zFoIdDwib6QJ+rZWTYTA7V239FhHvmCdIrps2DfVwFQkyOey309sXYjA5b6WvqhalKJBW/ldSDryawCEHV6NZCMqWY3mWZfATfB4a5W2/mJvM4SdpHq58JxtLQqjAv7L5Cgy5Ydm+x9LTJcIPKRGUvrJ/BdehHQHmohhmcTaIP780ZCMKGhXRzyHYg43bIXjpXANkIBnSVbC6xe98bAqa5ieu9GiAr+7U9FhSjoc6HpDpkoQYdCsf8P5tpqxqub8EmIlaTHqDmVEnSM7M/6GEPAfNFd5nfjtKSd6QPHDnvqhs86qzXtc3lJQVILOep1+IupPY9s0ReKI3W9RKKGrI3yEEb9iu6cmkUnEtzQRdBtxYrl06f/pmaXQI+p33hGwfsuEqFWmRjDOes4TeMZxPVE8ss6Z/Nsm53AT6/8XE8JDTKaUsDirgYKanoGyX+uAWNYX0nb2uNdaTv5qrhJddU4sieCKd/DlEvjhQ9WqVCQeZVhEPba6HufLOPBAdYhxiKhnntSrx5uugRFnUknW56DfXN94+jOAJ2M6flmyIPgk2wLZZ/kcv1vvHG4u516HrtYGPqV/ydNDN28=
`pragma protect end_data_block
`pragma protect digest_block
3863b83de54c23ba8777c2d882aaca7862336850153ba07065f31bab811f7b6c
`pragma protect end_digest_block
`pragma protect end_protected
