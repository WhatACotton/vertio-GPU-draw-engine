`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
vd5wlN6LGJS7tHVrYVgH4rrfHPAhPYOsgwC4HzRGoY9fv6ZlhyxWjilhUUABL4llx7TdIOPIwlI2pLnzUhI+fJ6+sfePw18eTxKSuCWtMfuVGns18/6a4DjnJucjRBlFOEbZh9Vyp5KLlsQtNHVNarmM62qh7HQz9ZCzwD+5/l2W95stnok4V+5zok6DUJ+2d4AoJbOW/fwj5UNluV/de6s0y55vfwxruTE1R8VVESiTDFgQY4tkHYYzt10+ngIqrxKwqJmr7toMeM4jEZH+embr5kSfWv/7sTvQttDHgZXXF4Hq64mafi719M9qL9WnGs8BYWAzPD8GKUz1mpI2HbK/2Oqs1+Ez2cnMzqVpJQnRvPzSoQ7sbUemGb7JrYCRrepLsHH4InuejlENVc6MUfdnJlyCYHgFmRJkd3V2sUlGDO/2PAu5nEK0bjrVbe8D0HP8r22FqAELSN++FXYzZ2xZ9Hcacgfm/ft3z65K3hti5izPzjIzlJwF7Db8cstv3iSY7wMNuhB/MY0hcuVEp9N6wqUzMvAIibwQTa0iY1QVLU9eWH1WunOMxh6DI+bZ2Ij6cAxEcXaFTzAmp4tg1mvslZ4l8hW79id1k8hYl2R0kJC0Xp9/y7tCCrqW1IWQPsVFJd69P8RYbdOkh3EB5fda1BwZVaMb8083fiaxKFwDxJnwwuZtIsaisObwgu6tVBLG6S3Cj9Viua0NzrhQ/DGRiOwi2VSYLOEis2KmGuprue9dYXmtQiym7r10XdNZ+flze9htjujzl5QN0pNqcr4xhuyLgeEUMMc6C8iYXn0uqtT2ypUQXyY5Psk1+4TOch1A+wtViOhnNSourejR+yAYkMAsKphdAqveqEfBUTGAOAsut6wT26/p3MF1MNE7RUkiI20Jg2/hkhqFmbmRuEaBWTzhaNnZc9NXHDcI+HHl06YuIMJPUHoLxB2sSRVgHx+Q6gUsf0Mjg3BaPpbxy4tBpTaEZaodHYpHbJy+WqLgNlTgZpGJ3urxjR+z6xzi/Vfs5EnHAsH5pRbZpGcYLY3VlJKNXBoKTLD66Kn0R9chv1hT/x7aHlnD5QbIJldP9G+PUqwIgpk+2ETde6++RFsbBFnSu6WSaUm0p8uHOuXsBroe2s/mV7HCybJFBzLZTQ+83FuIKo6QYhPdWMwazdEMDemygXtTMDOIW8T+bYK2FCXZVljUT5PcCjMUevcvwzbEdkvFqpmYx/SXHEgsZdqbnZceDEFJkGMTkR2OxImWuzOjmN7QZ2MXOZaX7SFFUp/tMRdWRYNgko8hD8Ut0LMGQTJRiW+tFbstdpJuAUdOMJpXtsDR9AKG8QmPQuKJ0Vn2gEuvvfXENwFZ9qNj72S92ty8gOoZpt94Dwa4vp3E+gn8wC/KTfdQUG/ilAUNmpv9Y+IoUKhKAei/4asJYL60qgpNKwSHg4JXk5fiApq9wLau+ePEmYg4F5yE4OOemXuSI4gqVx4rOwDzZOMTUXmcbYgAQlaWZw2JMxChxtHtYEoKDFssdYojTqr7cYjZxO96cIJ2S0bbLkyjNJKOIlg2Kgdp3HAhqB37T+uh59JFjzqVO0oe2RTQcQ9Ybj8270NKhoDcOa6hrpL8JVAgaEFMiYJV4Q6fy2E+tAbz29kleJc4sO3XBnaYOjIo5A7UmmvyZiHvQz86GBWQ6jSysgzpfyGIqKFfuFS3eF2s+afiNIu86sLUOFp51dCdwZv2Xz1+SHSsXLlaA9SwTQbw1RaynzcxGm3Bga5BK3HeMDtBY+Jho669fzg82iifOhUMn3RVhARDA33nKk4HNVxz68iFUIF8GaHCfN+haqerUPLEeFzFD11Hav7Q/S75PO47ZHu0Zb35GCWZdAafuBii+yfxlQEteQhyqpA/1a7BhSfy4pbn1qUwd5MW3sDFzshZ7ojq/UMmNf3hn3JQOvfFyl3hbgnMaUQW/j3+XEL+YbSpncvoFIerNNyZiGLuDaKconxIgNzfLr5ds+nIkNUyceR0Ic3pHskPmqt1HdBA5Zu+/fVNJyQNHZv/KTWc1+/r28MH/mAHLYrRxAbDmHZuiAzVcvjjWntDuRGwS/Nf/6wV8xEg+q2GrK3Wt3pZGvPDLuf2PSrCo1hcq+ZrYzoL27NknIpyWFuogbLgQAaqUOL8tbi2D2jlPvv9dMYknMyD9rxgUAcHNDCi229jUae56W/krtky7ZqEBN8yg0xZfjdzzQqcZkRtbIKNXo7UYDNadc0D4mSIxtdAzLCGZvNEHXnKCQKhStFMJXIfn89qTb+q7DgkN+XNjl/hQmocB2rpuZ3ECpwK8xOLt7D+7gK0NqX4yn1qZiizwdDeE4S2Ayi6+xz30dt0L4mA8rbYacLST3HbTbZkHCcDr4kzTus0Uihi8RagEVIORmNdduWHSuzcxJX5tqm07P0rEhrVj/Gm8o0UgMY2OFcOOw09BUa+gcWk9i//6HrEvtd733z0pdrWkZ9THnDas2WCiFYSQhpjWBSkKAYrAOPhHIsMC1mn2UQOEVslD3mJ4+tXs0q4W9toMZteOs+rVLl3w4XN7vCYRqAU8C7+UN5z04WHnMp9yMC6LvOh8sZ2vt8YtMI3xvy2LpQvgxGNw61ZMJ6erwcoonjUELpA8KA8kPPgMO+YmxddhmvlECgXaKpexiYjCiGyVb7JEK57bOBMo0jcsFyMzzYT5rZd/mOtq4f2rMgHDoSicNHGaoVRUNLaZvuvVKWBjf+OXHnEPfW6kABk266DisN8ms3+OzUzyeT7E+GW3aK1QPHPY4VfjfGYRVjKPdwSYiKVLrlJlOB5QG35GcNkUqjW4XN7RoPCPHCCIWENgWTFAfPhKtMzNA1H2dDhDlHW4YpR84HKtMbYKURkgyP6MMV/TZu+acrsYExxOwAzR1lwB8FYaAvosax2uLSrxz2y/KHUZzrwQLFpOVNsSKKRj7+JmS+9SMJ4cX7WtRSqpbh3UQI8wwg7n54BawbbPy+3NPO2W664Oh1rAMUPeLJL51fqqRqHQqvMbgwIF6w5L/O57QkMBVqvHbuLngs2WKNvO+KxXRqFHqPH8KOirn/IJx/ECw/gw4lWI/m8IkwfyxCWwzb2Urk8bqcHNzWfUEhzNnmUk7ii4yZRkNSEuJwfhevaHc25R1LGrw0zGhtauVhvbkmNw+QLcxVaTUg0/S2LaXkwGUNA2U1pvmzM70MRMUSxgnU2UdCfQZoBvxMcsWuBsyJLiq3ObI9RB7hSnMd+++YkN19JsOFFNsqxgJ2WeczyuPJqRyYKJXyn8sFGKppfBlterigjRcNgFA38rLhX9MB8MQ2LyguY1QzKW1fIU8bIxodIFs0226NKI/V9XPDurSWAZ78jWgzxNQECL18TazdgZpsBrEeJ79XhKfRIUrOsgM+qMzlFn4MGoX3FMu908XVSV7s5cBTFXHOdoqUfW/MwQ8pvxE9L7jvJ6CvSk1OaKGw0MKObk4MsvlCP3XYbFjifJybxRusxmzbuj3G4wW4e0UMgfWHq+hHpo4+v3SSH/WVm/kldhu67cVnQpuo8qsYJr6evYuNqfW0u6Zzj+KrW6ww4ECbOthpXlTONDRiLnb5buvKol5loTLynQouudgBTw4rHJve3hqyjUfT5fne9vetTFaVCOxkLUARmMqQOzW/jTg0dHLUI+FqPkbaaoM2b0KcvR3XztOY1vPy38QK+FFxyj3lDtZlvmAHvb12iPplc4jcw4oU6j7HOLKQw53shBllfZWrYbJ5UumfBhCcwRcixlYONtGnIq7u8OEwUVhGV3v6cgATYZM7jZoBf4mvjRJnMC/5sKOTEUgZQK3AlOHQ/S9fdZlB/U/tkIrec20hmhHr9ieOGzEzT4aZ6AU+DrshcXwfvvy11UyTihyEf9ner1OpykuQcRjyH2HO7EEtI+An+kRk6Jx4TFn02mCaxIkfT6mtpMKEgUknM8e27K2mUQpc9MnmsoqacmrKDvVVjIrnKTHrAfhBZDkXdtEZ1iLfkVnCXJhabW+8gl3mujiiMTz0x2/+zeo+vKOnBRJH+QiJJPpabhIV93g4I/NPiUdJTUVU9JE/n8kF48XqXXxzPSLUcOmj3aCmrwhEQmsYSkdjVPrsUYtCa87YTQ80Jyws9VuTCEl+p9soOSi19HdA9qpprucBo+VubIvuw+HUYaRNGJgcIDK1m8rmUDYioWjlB348kgNmu9lwuqVJpIjL08bwlU62KQqCrHLakYjkZjfREXEtBV5Gi1yXCNUmluMbADg+QSdAVvm9/Ti9ZOWIZ0ur193ZYa6k3c0uWdDCofFUVbqsn5xualNTRO4QhDHvqPM2noZbKNcSWg/z60JGUOzQmfx2yMV27BR+s2bdu/HaNaYFOXwHVxElgbLEbWE484dkdUgTVUNUU7vzo+BgMx00+B2JSH/u34vzo/ACWM8Q7fgHKgdVEF2gZBX2aG1uPpFaImNWGCfpo3P8TvXNnmlUW9gI8DNn6QZI04iiVAj3jNazSBRckavYbtanFf8SlZTEnfhOwytYp2xKUT90yp9B8HRkg2jkmwuDo5K+zlYqKsoG7vD6Ampf+PMmPo1ZT3Gsi0jZt0OfC4APoEJXrrdI6KzNsjp+/B+EQAgurLM+47HzGh6KIfIXsZcRjy7RTT547xM+kAc+UPHwaB9lq8TaG4vE3qoipSuRRFpetTiijW5kTndaEgH28wckyc/D51/7ks27COdl18sNx0x9H1rH4zH9yFaDO0ka8LTF2VE3bauNaeCiHG/oLbe7+AL1kqzUQGgWjy8khfT5xo08/HJhjFKtALpLFUjxw9Wn3WGoelmsIQbWEcY6A36m5IjcPr3i++MkacC4nbn0URr0h6jtUdXQTeue4KIIBHZqru1y2e5X963lbpoVGQdz+qMedq1di1xcjAnyiBrQIjEkDPy1rCk0Uz6pat+Tto3jXDg2EvZXnxMZhOIAlM1WVT8aSP/4XEPXIOqyS36s8aS5XVDWvKKzCz2lf1jWhdHTxXn6AqpnBWPlhgj7RFXjAR3Ig4rj/YKdG4EXw8zG0LcMlZprNpoO7llYta4nbYOHvVmvhTym3w9cAS7auWmrZIogHB3B11iR/FmP2c/r9IjDE+b6OLaxXfjS0MZZX+IsOejNjc6c4KRGObocFdaZ3xYInQ55c2KrAkxFoXhWYvYyEnFr3nT2YnP4naDM41kwEaGEHH2wDwTXu9Ie1MwgG98HMWe8sXXWZTLwopI/G2wdI0kCcqejxQwKXhxF/ysilrtjngY4Xj6F/J88HUV8q86I1MJECzawb6Sv0a0TlmxWLQmh21vWiaaujtEF6GcUDoEk+X8ZOFfbsDORSMnrF3R8oIojGz0TdARdE2AZZ6hcMUL3G7xKtm50QCMP5sdEeU1qxrFpDTCui9hFRR5LFH9z5GrRgN6N5sGfUsY3bUbENWoX4fXdAnPYbzGS+TNswoQFgxQLQ6TPskxRpl/gqk2L9NDObHFKSyg7eBgN8Rjdo4gJgwWJ6Ec77aYJjOC7a3vWYLqvzNKNvhFOiGbK3UHQORNj/43h5aYhbO1ryejwS3m06Rh3u9w78NKAYUV1G2KGwx0LAqugIaVBmfdxPqR1PTr+aoGzjv7dHYxyEfbdjRqIkFmoh2RKpArQzAZT/2RJlUsmgNzpIa74Y+vg9nCEVVWMvxmrmpkSOAFNE+QzToFvQzBk7cStahi81v1n4PE4pLL334Vhd0gbLme8zkIf2Uyhan/UkCSPrihtz7/IhShT62y25MODv53GsRMFmF2zHV6SmzhlQm9GnwPc5k49umXw3sfwyEx4+iVRYdpDHZvgnpQ0nseq/wHA7urhJGlkzsZ6MtrLjYMugetL9X4O4I5VHxMB/B8w4NVM3qsWshpqH58MjHLm4neS8SpPKEz3M1jb48+UYGrTjjQV49qEleo1IOvdOkwwBM4piPkthAxtS1QnxXyVO17GwUWh5/vF85fxj2mgttKbf1LTga7sg5yIACztKXe0T3yYMVH91Y9bTvguZKpPZGB0ENlRwktBHGkwBm0XV6C1HUnrN5L6uTuGVcvN+kCVh51VQ25id4XFhqCnWtZVU2enC/IMGRXxweH/s2+QAN2FhQs29J1VQng0++ej7lGrlfSX51cqiW5YZvIL1lvuMk9DNyEpLwxYKNF7H4w1pl7qnOvvOxDaqBdWZ2hDhK4zoCGsmBbNqT/Qay+leA16Ao947eXTu3k2Pd0clznGqLrnr6pnyPTmO3+3NzSTiJhsqRCQutr48XNBkPYiVN/U3xybH+T24XJOmYpGe4D1dsT0eASw5oO+4LVMu5/KT9aDx0cnAp6rLFCw8MT02UBl5biqHOcw6nTj4+YYXlrAfKqKhae/ByszWG+dOLaDs5JP6Rp8NMbMSvNMaRvZcutXlpdqAJer27vwlOBhVmk7O6bC0LHAstdyiUpUvXQvBIaaXWlS97Z87RATjj5bHb5JK87S77/wFPysnMRTBCkQkzqynr85q3cgpjRpDZvbsPuV7BC7cEml60cl/VZ1x53Sq8iLosfKefutPSHDDmIvqInJoOTfetCxpO9iwezZm9A6qjsA4uAGdauq8KHcg6l1txxTd4mShbRfFkexu9mmpDRwj59z39dUasUuNpetBl/rr4klqKP8zVCHUJbFnSEJZSZxSPXaTb8lXoVpt2sAgFY8mvZM516ohxNd7KcWHWzPGTzfAPUCEJ3XnnYOPp0EDx+UN4TM6NLW548XAFbI8mUbrLN++vPSo/XlwCSJudVUU1Ev89LHaPx6mpwmjW2yQzz96hWXqzk/kExBNXPxrkYB0WdJ8EgnoF2bEjVLROzOZ7WXH+M6s/ixBN/ylOeXirqwP9sxbyWDcFW1uHxUdjIia4adaunfNzDe29FkO4cynBAGLPkRoUfYPDzJkJBwPBtPHmmPXhHXRzIXMJY2qxArAtypqNabcdw03SHlWCcluiq9Ce8TbgTbbVIULqoCg/XS+w+WpQqhSnqZi9+T5+NoqQYVnlLU6Ok7Sm4PcO8cb60gDjEwRvAbqoI4Q0EDO65deZUHX8HpnrSqupzLLxD7DyVmkQA2Ur+L3CVWGcSz79mgd3I2nSIuiBeDvNkzYGx58num/lUw7uI25YImvpLT+D+9rT4kDgqy8ADwoNelMu4aoheVIp6T4iSVsWJyuFoLKTmk+dv1NNBw8MaiLshELXadJSUorxGUVHfTPcJeZxQXBN+dKQvPKnjuIzCa1UwRPG9lo9Z2qU6PV+y2R0Ho1OWHuByXD1wPhoevF7QRUJj32BhGihKEQwyt9A6ZsKoa8qpbbN7p9LiMtW/O7YbGhfGNNV6mZ/7EBTVmU1b6703PWyNazcMCI9kcbpqP3mlFh4aHpu0Klv+JF80aQwGkrkacu3jqPqByFlKylzqGYux7Y8QTum5pDiojf6r19JnljJWk0h734N0Fc4AEozYzmTQgRGrdVykLECfBrLQEah5ECKn/GV6NpnAZRB0IkPiqdUfFuXYcRAtc9vpCasrHnHJ/KN9RpR1KPr4VV0+zPEe1zhKE6ke7utK7oQoqVVfR05fwCzHU7HU/a3Mva42LHm+e6o47mHiR7udUSSYVTXM+p55tyVGuG8swk3ooMrjQnQEA1elzi4vDCou3dxfxi+SSB/K23wgnGHz2+n51Z3S2nLgB7uZXeft8Sfm/Uk3rKGXr+q0NyCFuJgB4VP9FHl0CuJjCzznMZrhsAXMaWbswcA1M64oP1wp5lReigWRTnfPvLy6NmHOPfx6UExOyaHCGzw7dld99mo0OHBEwRqXkcSoxF/yUU2/ud/A99qazZRLeaO7qJ2xjZET4x7dPNpesO6yzihMO/1xUN49sHhJc3IkKKt2VSZNUa6rv3H5KE/Ls6nStfhxcykJVs3GY5DJDfy073e+7TrDyni8jkJFTpvTpZGMJWMcUkdQBfRSwvLo01TrK9CTTER83iCo168X6XqfLMKBmggP6xgiFQWqMvxKjb+nkoL/jQH/U5yve+JpVgEW23Fs2Q6I9meawOiB4/lGuXGRO8JnjTeaM/lnj4cABKlioN246xgEsh9wElnog5akhPzG+pMXUGypcrb6doZxWYIrud2KhJSotG5aNAJmCzwkTX30f+r2G4mmKf3diZtiTUA/c/PdxoNBxaZcNrsAMnQ+7BaSKiip3743+e3KNRiG9uagBmRrsQj1zOyx1cTRck7qhGtOUIOOG5/K5GNV7On9O3YigktAA/qaZWoM2TMxsL15Fil5YygegIXik1sa046j2Wm9g0YriwrA8FQPuHqTxGEHgvuRmcjr3p5mX4V4irBZSrAyyUmSs//xQTuff5YrRmnFanXkQmY+GuJU2SsuYXMC1bgPtn4thErEBw8HFht3iE11jgMsGssw+ve/GVmg0o4p4lTOu1CW4mOHz7IvtR41fWJAl5Ur7fdeb6DwHxYlnbxKttkYBvoO3wuzG8/oB060C2ZGK445iWcuXoURL3PcylUwwIZoag1KfgFUM8Weg0tjx7Bs9qBbifpLdnCkUaUIvl7ZnVv0dCJNzSGb5PjjcMRXIeYA13B2lzkJZGXkoFSHZbxuVoYw8a0LQlb6R37FmgeiBCViqm+VrzKP9q9TateD2A0FG4UVwyk0bsoGot/t+u0XJsjrMGOiZt0rZ5VDOzO1scO1atOKUhtEALiP/cDSz4jiBFjtYBzOl0e7G753jev1nbI1UAIFJEzm0wOjiNFYG/aMxTKUcoU0jKs7Xvk52jPiwd7e0eRFK1ypdFAieIyjbVrWY0tfjgQFDIiQ8hqVCZcJdTF4563FP16hajjvVhY4HAVKbrnu3GwHKfyqcc6pS6Vw2iT3R8/ErFEGH7cS04g9OXqPzyGKAci5P5Y64jKV6e2lVj9u097ohrVS7MQ+P12LIj4S7UXTQQjZ4m5Lj1AKMetblSPX1ZvI1DrJFXG87hQlsSQcbFYnODMrErhBvWP/7mOkLOLQ1L/VIIDfRvmEYQip1TorUvAAkgWnjqb6b4Z7jwg/dICpRvTfoQefKgVTiV0eqdFqO+V64ImBX4IjuWIwXyUpG5JMXLXWBMkgFj8eWy1N6uo4e2WbjWsnm6kJ9S0Tyb7iGqJXAbJjnjtwuznGu5B6hnMsr9J5oMSvCcu15MvYmdeUwH35dUURjaCP/nUaQAo3/mL0DHn6gxO31ewxBT4xGrwMoUL06BfpSHbkBtxKRuAwe43yEUvIVjzJv6JhkESH36NZs5RyZmG2iAtjnj6Q8vgcRGghH94o6PDfNEzsVC/NUoMbhHtbmlOOSrhSSKFJVyx6aFjoRMVwHEviAQwoE3vuUiexYYXcj1pExPTdrjsPswKgTYk0+Wl6xubkY/PPisXDC8pYDnJWY1OSwVsOEpyjsp1SszZljif+wN0PpJvEBBn9OALYXpaOFSGTQ9F+4NhsWUubGxdk3xv7iFhj1ps3rjEymEUAMkWb3DhLSAAagTF2DSfP5Sdtn/r78js1L1WpHL1ocO2QuIRVVF39rm2D2GfXWY1BK8d0l0eqgFVmdb9nmA2WGMGG5IJz7aAe4YJVjaxXPXzSU16jn8Dy8sFiZBVRCTkQP1Qi9fZL1DoqYWZ1AVnw9EdsusHCLVsv74E1CmZmbkw6CpzDTC6JQIN5tCm8/iH5Y4ZhXTuxF6fA+3h4dUvZqur0hNWa0e83GSuay6RuJVoXtmvLHjUqonRbM1erOlqv9Ix+E7pZrjPtKtiYzu7mLrXjAqC6keelv6GrOdOQGDs8yRkJmaqmhJL267gdamBehu7m4gEWZ6437bm5ftUPpBdo2zcLFAuzI5+UnnC1IVDuwQWlAR+GO6XNzh1rVjNE3Qp28ocuztXx2EFUb/VFw6PA2EAx2eQiyeYRH0BlsOEfbKj7iN6X5dOU1utT9bTgDblZFl/7VAPQyP8P8MNF7KMOMRuizWdg7mvrEJoc4xZ44FVUmkMGYB93Iz/mM58dORmxFpb3p5vnHg1r7wWPRBWmLYOSe8HK+dJHxmSWDb21BQx2ltSNNs7xFN8v5yT3RtP2Nwr/bXr+Z6UCH1gL4kq5vBRPb4QZXiKV3zKsuwaNRW6NSShSX1YiVCDSwrmGPhL+nodPRkWB/e7ik4orr/QDtYm3iqtWFnF80fUeAsYWGiEIcHs4fW1vFyazqxvxQSX8BbuYi30JjQgqLLvrWr8akSdX/Xhc1bVBtWXJC2CVLg1/l2Fu1jLHx4lolSyh8Vzi1W3nM0lR6EoLuBY4fh48KtxB7n8KJFUQp0k71YoS3yE1XQuHQpwe9qAPHX9zz6EvU5nxqm0Ml/nCrgt6Vdu/f/GuZKxgqrYBLQEfuX7KfgFz1RXPkocXDurMBcFlhZH9XarbELTUU4YkW9hf0sNCS732rOmaIPRUes6W9aJ1VYHwM3y6zM+8Hn4lsen5lmTjf9bgdTr90vES+IAYya1whAxuu7iHGhgWaIQ9iJ5SDVVXjxTW135l7sZnNEFYpXIfprAycxgyfnollDjV1ufolqnMTP3Qr5NtGPJqLFVPRj2Qi+7e9tdW5pyx1N07/F++7efpv8R86mOZbQrkJxhne+2iaBmuAJhe4MC/JbQ6cKbz4STqw0PbeO1dQnuLL/Wu1b96AUKp6p9fJQMLWU4ouEEz7PuBhkX9M9foPIIp+usWiquAUDw70N625zESJw9N6uYeGRazIeQxa2Pmlwb7/cTmEOrtGQnNGLD7wH4NCVC+Gha59p0MWbtwyPSMhhET8q15MfU0z6l+LN3u7xV1bRJ8AiGg47PrPIst+W6WLMV8jHn8fgSbyUFfwQBIgwz8cYlpdJ5VZi9QCazssDniCRoLJR8H1Wk6aJnEWnG3HfyxiZUAawnqlU3I19clDN5wzFFIKyjttfmKk7xVdGKRUTj85I2+mTCCwNR4aM6ckjZRVt3/AA9LCBpOyz/du8FO3oLhBXcewTas330fguZgThQjzQIx1wX3jCcR0effmnoYX4yf0K7B0r0pI7LzF/buqICOWIA5KUBVHbupBQM8GicgbJZZfr9JNqlDmCRjFjw2IZzAxzBklSL/RlOEpNWlS5o/RxJY/76HFTNjn00VdJhIDZOUyCGp7NaaF7+Uau3DPiyylRQabcNi23Cl9eoJx5IbVZ0eaFwK4MrVIxX5W9CuWnWHDmbwhY4lcnQayfdFpyiub0wxCZczH49NWM9HQ0FT4aVWz9mBOLqs2pWGeEgLcrFnecQqfClb3L+dAZ/MDhJha9/FO+khiFWdE1hMn8kJziFhvB9hQD50UmJcB/g+PE8d6o9s4r6gngcDw/ZUaRnSC2mDssBmJrzQQ4gxQHq17I78GfAe3jDUZCiZfSm4BqXN76hLynDy3WH0QSOgPTtANTxEIE0hcqiSAVGreKwBk1y2n1r+0XJSkVC7Fo7oUMpnCSTKvURYsmdNlIXfDbzcyXxhA6axUNlVGLGc1KF4P56tqrXzq/GBpda4YsJu9c95L5YadS8Jcz5hWeDVNXIiIvT6Zji6QeLjbLLwRq+1rHfY/8DyF3jFivsrdgLjcytuSTTuJp31SJY6AFB+9vVhM36+qlZSD9inl4tEz1Q0XjVPjLUp4ztwnJVP/Oeopb3a6dPDFQ4LxECXHd4/PKfDkFOOQfXyoJQ9OUrg/+SpoKa4PFwicmJZonadDlokKImokrih57Ucv8cg2kqJ/Z0HHhcJ+02cjYIYOsmg7bO7ph6Oy+JzL0Ujr0GBBCUq69YZSM+msEHEhIYYNUrzahunI82jHsWHer5ura8QaPTASz15bc31uYJqbO7bzY58bC2bR6DMaZDbWGtdALfXogNMDjEkA7rBaQ7C70gtGC+6ZMlNeuRx4Z0y+yZJXGU3QpkF3Tt8cfeHHeXyrKlE3qacFPeQBRqt2JmvqL/iVPBkEVGfa/55dSiw2rhKoEDIxivGNSkfNerR5lSyNqbadDj+M9s/+cIdo5CLoOedEtpFX8kljQouNpRDI/s8YugREAunOR5tWFxeUXUD15Z/TAQwpmNMvPoB1lLrpHzr8EHHmxi7+mu75+OFc0+Nv8edssO+Hnyu9wXY3ZJocJGGK9ivafnw/c0APhsAi7uYpkwgjuGTs+IAqUta7S5rjgxb0gukfmdEYSDd4vj0fD/aOtFzuuLJVk79hensctCBz2LnqTOONEG+IIc3zTGZxMdeMPkKVGDx/nEnYU6Xt/jdPwguHzwHwg9FD6sCA4f99Mre3NOMgtCdjMLwvl+DyCoMBi84HkcvLc2dOzqO+cBNnLNlSgj/dbllFpFgJpwh8p26axyEVwPE7Nuiivaqwlv6p6M7TQx5Ln8ZpmzkdQ4hBorzYmIotOW5Sugin2sxpV159hmUW90AIBlo0jekLZElqTUxWpvTfbGDahCzNY2JaSqSzuyklKIeYJL6RQY1iN+n5H1XzJ76JI7nJ+yJfqw7JDMWmtuygjIiPahq+VthPBbQfd6dSvBDzIFEX3ErBLcgAjssXZqn63z36g5oj2DsIYnP3ZfS/9wl743MRJhL2bTCUDfrn/b0jbfCJCh5LMHoS04AIHvVAYEDJFwfjnOxvG3w7m9z676C12tK+KTzu//DeJ4Tgs1PQ7+5ZgIfvfN+Sv2GaZVcVGWvlEQKISUnifeblnmKfxjd+YXPDcsBD7XbjaptWeV/7HzCjRAW8uPTIF4fm5h1fS1Y/jkeUMAmWMUEG4sl4Hi1Z1CaNC6FFo/A0XuWPxfFwyRyxPn/lEAdE64SFg52UpiIyMD3QALnzw2ObGmU9ywPCq8LllHMjYXQN1Ft3M/y9a+Dad+f+3tAdfZAvlQWYWCmN/9V4wUGnXJ33H+UCR+5FD/2OJhqp3u6EoqyaVBFwuXDQcbsgTGEne2odFNENpXFEbLOtNO7TkYnDOEiXqgo9hTQvnj9a9bVVTjpEsdzhmcUHnx2oDGRYwywtZ0UCqhNqR4f6QjzwIHHNyvoyZxhMLJqGoHfkxoiO02Eg4BfuUnFZSfum4p/SGu57wtRjOIQsOcK8nBgCYv7NHKtWTO/XjWn744G18u6u5FR2EBMWCRPoZ/PG4/dxHOxM3Mr04xx8Cw9gs1joNB0DLzJ/1phRGqTZm6dtUzs2LmsFe8HttFUEo0wixcPBEU1oxwk3X8AnPiRcmFObJ814TL91A7s/MEa2MLma7etIJRempkCFwSXJUob9g6UEl6vAfKRtU4iWU3WOg2l619NrK2UPdlGXo8INRBMrrzCAttoY903StG+u6zewNSN9kNj3s3xDYehyWBEENAyO/HYZMQmsRIYpwG7jNLrZQH483wOouRzdnJRW1mC4oAc0JuDocxUkMvT7NA7UUntrtNIUPryGU/cGZywvD1LFHpuQwluslmcv7MiP8cTwnZpasuHFpgoptJFucgg8pXOrUrRhl2yjiaEf1xYgzkoRw987vgrkuSSx9XMZ5HdBBbuhucKZ14jQ6yjVEERhxwQFdpEMyDdqEqV+v4mze78s1IYaP+oITUCMovkwweJ3HVoFEl5uf5ZtaYKS5xtK2CFgQBVXBu8RAt0fexGxVwefev0veeJSqMKws5JjGbdXnBviROL0iSWGCmTxG0Qk4mscVBc4hjEgyUi/Fv9rcqXxvjoGNrj4ZKQKY/ySFaj2MbhkFPvBD/oY+Ji4ZLN6NW8rEdPMhBlJ5Jaqnjq9c1cGvvhaNIZyWpxx//6SIVBBrMQKQBUugS1ncHNbF9djUMmpFWiTlWAt1LLaJe4G0uLGZD3+ZQ3aW/2rjMm9wWOXJnu4xfDd35jzV9Datsp77FHUd8bKeUqd6w3JBcIOQ5bGpu3fiagPV6D+Z/kc7ppq64BM/WTS/oMTgDfC8upeGCvVz6H1XWPJXjGAiiXam7JvuddcDaPNJE+7z1Tm7CfOt4328hotNgDaWd51TaXHYDvqqE5oEBvJu/keyCDQBUABCex89evf/8TBoPmi/Cp6sDXs9VU8mGaBFt1MYkfo5yx+C4St0bzMroqsEzFUvfOKQi8/kAE7FWYrTIu0ArgxHGAS8xvZ7YprmSwagcdSMU2kNpUnei3WXJs/UR0O5TzFz+EPQHcAf9Ftp0MQLR1r8/NMNz2uRNBrJXrfnLLK+lqIc6Wl9eYPsmrFdVG3izrv3mPixhld1BNbVpSs0i02+R5epUr1/sN8nRPJv8u3ZGL1hE/CW5DHYmPVy1UxLPXewoP+upZjQBu9Ntlu8jv3m67qVv3/y1njVNuzTnI3WdNElOE6cwgA4SfoNFnR90r4r7b9RFysek8e4iXUz4qMtY0QTXUzzmLky6uhYzdjGPMQSXwVDvzEq5TZItz0xDNos2lalqxl53O4Vp/YyFOy0KdDAKGYbIkoK2gLjnTwmSrw6wm9mTyIOOrnx1CAdLwJqFwJq7XLafvGbhbnaRsEsGLnaZVjkOg2+ymSY1xBFsm6pVdumLq0Dd42mUaVJjgf3QQeobOMsecxuSI+XYN4EpiRXj9A+DcWmGGIKKDnchb4He0MyHjIbDvamePDvtz6OSqaXh19l2zM91GUYfJqWWxENa89ZNkwSkIyBxxqqVLHYnyIuOr78M0C3F7MeNXCFM2oIRg6GMj2lowpgbt+QJ52KMgR5w7dSt1DsIuim3C8tqqw+k8TeLQNT/F1r7G0cI4LKS8hsM04c6NRxB/8tG/BpQVBAqzzDhDz5aWc8+i3A2vr63UmqfRds9KZKH4L+27d25ZKBwLT1wbcBGjPOCTGdEJkEGHkB9UwlRcS4avzZMDSgkRQxYH7pHJ6AV45A0ZQO4NrsNvHWVUpuqI6CAfwb11LLmag9TpsaTNNM3bFU6HX7rx4IJy2rQDCDclVbeORCqrmSibUnP8LePEjVRSEAdWH/F4ZpQAHuXGjPa0bHSJYptZyuDPzSJPYknnLlByDNpwWmyN1IfiuiXNo5KVzcd7B6mMGX7aXGiV8U+/Rsr37yXaazwFc+zQIoxP+QpmgwgkclSOm/lluFIQ/3VgUQ8wX/r2Kn3y67UZpj77CcxBfflj8Fm0zoe4wne59IJventHHXTPerX8iFx8p9RBI4lsnLmbf2MHstL12nmTmVyogJKATrEHGGeA143/EN/sM3iE0cZckAFrdiAuFsDGBxVjfCgpx4/4HxLzh7HHUpvqs3KmJnT5Yr0EYPC8kE+6g5pBqiVxsL6P0pgvMKgaCj6PZ63RiJILUeQD6Klhuy8RZ6VUvLUGHj6j1uyuuVf5vaNTF7bF3Q98dhIVsmPnusbuxrm48J4Kqfvp/UPgmvlYMiT0u3ld4yFgVM2sQUuMyfNe1GeWIkIaRVonmmlSlyoMm1cbhA/8WmDzPmmBynA0QsAzfVSEKW2r1j3dBg2VJknpET2NH0Ac1eN88DOHZArA17wP8zO1ZwvCgavbvJutnEYpAcdWO3Zb7jWF1T/cJWTlinuCHcmqE9/0JtY0THpaXkrWB9Qe69CV33Js1LijVpCtqBm3T1ZHePdNxPRgW0Hyr0Hb94fdmaf7Cq6IuXLtMpzg7E25UXy55Dz6OjaWufi1q8/RC2dhQjy2zAKM5AL1+eAkp80agbbvugtYxoRUqtieR5j4X613WcPAo6ac/AJGY6UowClbpPosmgsCNzJU/1I/WQ76QgtSrsdt4ZmcQHmP0mHTytXiUotQ0TRsRVMH3GsiytbeeyTUZVyQln4+i9WUqZbipJIVXtPsQa36VZlSsYRAVh7J0wxGD88KNPMZ0Nd8QKPmOdAHTTO4cD8wXl3x7ijG0DhyhhabndTNOK2NdpDfuxuk88GfdjeLRaZRUtjiK9pWzwUIbhDyqi1rXRYkSbZCE6hoAcDTykpV121ZF8tmczNj2x5RpeG2a0Zj/2sBHj8+c/UPvesMpLIwRdFMdXBr80k6UaQf7iZxwl8JJEfPOIFFBejbipXYT0+jDdTMqahzGizwQ7cYRwKk9UcRM/chxV3YsJVmlT98p/VfnEIRLE8e3ggZSNWWm8rWyqHxl5pmAR1OWVh2pI49my5DfDn/J+hh0Q9TErzNDJJNAPqwKLKHG3X3qfQA/H8vABB1Ykl8O83TTxWA9QDai7IWrLcOOmwEIUeTbjymxWayk7+Yh+6sdRedCFiWWvEnSGIhNsX163m0peXMNyT3YuLkAzegU2DEnot9lJoxp1fkACkKAlnHrkPHAHWFKXNC42+5xDElNeHlW51VypE19R8B4GXjhT46NXJvpYLpE8QDwhuQUfhh3saGHWdkpP3Rils4VU7/8f9EOpMRNPEEwXfz2JFEnAStUgNmaPum2LkJ5Mde24urHXSF3RPBhsS0yO9sXRtJeS3SKsybmvBIoXed4g+l40iR5oJXXAed5plGP853C/xYv61hi//M854mMiQGkAG2CvEKMOe14W6e6rSBsr7SGfpmEZAgJi0FIDf9fVJQZxYjsJIV5y7riiuB5z4D8bDzTBhxFFOh26LtpCdW6f4EQZxKy7HV0jta8nk8c/iDuim+rLp7c6RZDpzCxgmzHzh6pI+Ao/Dh5WPxN3X09fLKZAgxZeDWoLbXSi53ceFJmNedRSSqXPBil9UYswyVyfDwYvOWClo3ORj60JH93VBu3Zb+BlHqMI2ytPkfe6u5wC6AfFta408Ky6Wyu/CA4FDmH8RDPiGU3DraBJozyWuIKNuH1ieSy6yMVuxFb3JhBOMu/YQ03cpCGU8298Q4jndcw4OyKFsINW8Rm4xFLUpyB/6hHQ5Ow5F6DS/Pe9fAUzzeNUhQ/kfmwb0yAbWi0ZoQ8BNqEq0EI3PirTsyvzG226sVke3ULJURkggvW7aphZjr+Kj4X2y/XuZQHY7Pg7Rf7IqNODvFSMDZCcDnR8OMe6/2WjdBOjSm87igsO9Nfu/iR8sqpkTEDaSbl5EJajoiYo5hwbrUpYWfpNE7dZRPKr80LTT1DmQ9LTcadRgMFIuiGmIqNjdNWA7Guoi3NRZrqcbByL1mQk/Yu205H3eNsZv1eJAVXGaoyUpJjvuPb0KeBXNZd8QdR1q2zPUzqAN/dbBsKrjCtguQT+I9KK2ccGyzvkJx99TQHOfqgZISZOPhp2A2INmCpyX7XROsVDkstfLh3NacYQgmQbpf3nBVeGad+slXsZ4RkbYSePZHKHvfl50VKTaFnstRpyx5wi8zjioqbKM/PrmTbfoxczBdWewU7jZrhRBk/amWfxEgXFoQMzn5LnmpQdAJqI1byFgTID8n9/JWlwn5VDvvIpN7KkI1hn66viy3fb4Pt68/eYuxrvdgMbmdiYDMwRqWAkAXCdxg0ZDdsxU7SBMJjDq7Op7gI5QpvPKnIAYJiIk7QWKEyVdyggtQpiKzU5D2Ffd93A2J5IJFAVOATE5TUR0BuzcEBOAMGhWZK1VkxxpMmtVWIKcKztEx0CHdQc/54TB2qz01I9aCGG/va3mmZz5wvvLUNAyqSWWUuE6kWbAU2/cWnXqBF1x7eOw9RYLNbmn1PDjS7ScRAt1BC5yj2hrPq1Gp/8AuhaxzIFKuk83wdqhDrS50ube7IacsqZWLK4/mjNQUPFcDzXv2l6BlE0MQknTf7IGx54QvbtZCVDLJ0YAoT2YLNHjsMa+e4lbIq9driMUzevIP7qjkuxD2MBZRcYv7PvvGJMJ98kfqrZr/U4NhGDCOfedg12YxXRnCLGiFzpFGLrs8rUrD9MhNHoSoKkg/vo8Amen8wM1SHVB/tTl0fVrbiLC31ONyPGbGu2fMf/HVy7mEDCUlVqO1tFs4QK87euAgMF2Ojnp5SFdk/sZj5g0zoYR8nL36YWA1haWeQIbN54sYS2WokYZyrINH8kI0k8Le7N6AfY0HdqrF/gZOvHk4Xr5Wv8mLPy40/+5DX+VBAKIXWrFq5QBl69vBuhIfzQ3TKXz9MPs+4lZNT8KIK8tpzTq1NZStd5nPBEqQduh3AnJHDw0xpWj4nI6qmhC1KFTVrZwHhaGbj641LUXUEuiFGw+QWrIIESGnZ3tLb+3P5BkGJScCW0yxxgGuiHnhPOYMPu8mNNczwcy/NjfKDDp8tGGEFwmYwEKc3cs1pjuXxgAxRpjfaeSRYvUOUlRgOllxGhTmSul6l3luxjkk3B06eIHpU4jHUzfAICWp9zyyQw8iBu4hbCP22h7PPmEs91NOspXdy2xa8j9n7U7lodGMqMhIYX3aRrSR/Qa/DGL5DWIo4iYf1iTP2SKv1PjWDXsNml1L2xiQxU9daRtLCcYzzU4/4sQlbVfMJc2KubyfK1Va+otbTZH+pUC/jskMe9kzqraexIJANfQOEUsXXFgSKyIpGBvYucuP9O1uv2S89ekK7rjjIQcTo4fFWkC0SHf6Diho2qHetJTlly1qFq5O4XSKJe18LfhXLG5dy30QFTYmQgC6vBTOP5azokGPWAb2ex/JIQjUyO+hs8PVtwYOwYWdgvO3BxmrJDewqa9IkbhC7CHO5rXDYiQYqgaAW5Oi2IGSQ+5JCalwD8d7vkoLRTp8e4fYnab+V56OM+C5kxMo5OLYOr8zUaOzEwBqEQrpdS4I+yeDYq6KLoBH+lg4AC1tOtDTx7PhWy20CS21lBiWH9g3bFh/MPen3jQYNLeHvt0Bon5gAfFsfwO8Bg8fR5JjMWg6+1+BrLPLLDZpykGwpzxbaH3E7/JUlXbjung0tv4GICgevqZo3dMZQHJAD8lKX4Xc1G3C6nJoWQT7e0MXVO73A4LZkH8d/33xH9g1fK0U4YudhhT0Pw0KdvRKrkiri7xCWNhKLWGymAUbsivI9mIYrbao08vPOPzXRF7aMC9mzjNtcOx5pvjoVxKqo3i3jAqDmJIYyMeJxdePfM0t+/syNZFWMWP7hMRQEy9HALEmFecrP/qQ1LLJa7g374FWUZ7nb2EQm+fZIlWY1uQorqY3hCw0/UAkEui5vpq3eXak1XXHS4Rut/BpbRWNCF2d3afvSbk8mmvCUgpxi1eJoslkSMjJiv4Fklxph7Or6EpYfO5YzadNp2OfCARdzW61XXawrYBYwwqhmKJ/QxmZcjtqhiymNUICciq0dMUzqSDJH2Fy+HA02OUSjppD4BkqqF1uHGm4rJyd6mMroRMxHOIuRKq3O4LCXt34N3h5TSWU4Iq5JBImH774LKf8o1bGogsNJ/fanEHvuxoR1pIjVyFeBxGYQmGDUFQ+e06KT6eDIVB9BdXa71CEpKlGPpqXl0eNBPIcJin+JGPyk+G4tmAAMjfzkC66Wj238iujNGW3UaO7c61UG7VobZ74UbyV9x4Sq+8NkewUAWAT1uvR2hCqjZbumh6/LBjcXeuV+VZp8MCOkksfSOxXzmIb0knFaK/wLLF3lv/IsGcYD2GJfPcFyqcBq7oJhpJrgMj8zqtteG2NN14UFiMsKkbJzOnGpgl7CLDFbTyt85oHDQ/bfmTRLP7uEGtMVcl/ZruDuGLyF99mUn9WoDqK29Oqn8EWFm48r/0L5Bn9WEmcoeEV3rxerwnvc7cFcZiGzdJnpMZr+n6bMmwm0rHqV8MmWyD7Xim2Vo0JyxMg6g1TPsuHljY00/Q7WxhThjtQWCEgmvc7RqBl4wBioIy+EJUhKs+FouYaVRVIvwmGXiIOeuwWSvqBOH3SPO451VJpKkjXLbBJpXHhbIEvCdjPMt774DSVUN6k21ltYNyCJoArsWOnTaOUbTkjyQsNjNdgg0rXsF8KKKE+asCHYqwN6AV72cawoqYOQ9qsWnWQHHDj7+IJbZC2lD0U/+Uv0ARxmjIHFsC1vICtfUtYVC9drfMcdLIQKhjkGeZpHNgCU1dqijoMr2zbiSVwcTVFkV8kLHKtg/QFXCY04/6DCwyw4OKn33YEZe16DdkajNjCzqxJau7zzLCKHwyRwSXt4iNIBFBYnjzjG6ZgJNmy72Zr/v31tXY5QBuuAWG54NKmn4Qyl1EwRf6ygEWb/hQiFdsDC8hgqKl8oXOqlIIjOfFFkrsQpWkPrYN+TbdKDqdQW3ZzPiHPDpoWLOI+jnPXgqRNeMR9QfOzjxhIutOzBMMTh/RbyqYGZltZ/tq4VXIN7n5ho7+WYK1N17Rykw05jBAit1Bh6SHjucWIN1rUpNTvo4UgUQZzvV/l9Jn1cS8XKGkrdZ1/N+A6FVUdpBJk6fWrhBa9EDpxV4T41c5br/sARGx1YWh6le2zDNhdkkoXMdarnRfP8WQvtPldWBmNIt34ANSsXQXgXzx4gmRl3cUyKPUF4BnkzWPBhiHt3fylRbFkN7sJOMdYgGqDLR3T6xUWR+ee64yTg1XmirHnQ1Heb85qM08MCKsJW5RYA6dsPpUl/JEjwJTiYev09ulJYvZ7eT0AiqLws80eQ4OplXagpM8KoQ6HZezsy+OTuCjeRuJjp5BLxinAkVOghOC1Lpq8pPbddTNamlGS8NWiY2RL7ERLmsSv5wnfuVceBexftCn5DFO0mbPdLGb4Qr38Hhd70m6u3ixf7hK/R0HsB72Q6YeUjBIG5p9l8+tKw7adOvLqFR3ZlIt5zoSgEDHLviKQa3zHt5pE0lzQRnK5gq0V1IJRAu2swSbNjc7IHljzo60fw0YB9mQEHMICtJhABRkfKmfrv1ZfuPQYe3ukf+V7+2XTq1FGCK+TSsIZATTiJeDb/sWnVNJJduS7UZmCm4vsUBdMT5V63VrIAbyjgqF92EsstSSHCwxKXwYiZ0LSsm70jhVCb8kutIzdhQ7ZYA6qwGdxalIQx9A4UduhJOaZnZxpQgNeL2Gm8I7J8nofICZqRFKy21gQJnWOwug2Kaw6XXWaQbB4O3jhnZcJ2TmpcMa07xNjp37XMnMSNn6bYa54nMLyokoQzWm3kVm79s0+ObstuwZO4yk3Qmk6BlyjCKDvAvtVQmc0+V16dukXjuUYv6pqmCLqbZ9+XGETAXP5kaT+qBq6Ne0RxMlaP6dECKd38cIzqJvr8K1XpzoIV33zX5UuNTb2FFoCnEQ4LK6LbWF2HWzj+uRsywvLvlJ9rLzbr7FZyWRJHEvI2Hu+KovH6gKNn3XNMH1mQry5P4uYfr6fK9i6BwkWd//rpIULMhS3kbqc/M2bCKaLZYlgTZbkTiFVgncrYI2Y8exA55GxiaI40iUuhjzgiAYfWyq4F78clHklPDayUER0MvXGHFJ68mEDu62LT8OA7mlfxZVlg4ZYZ4gHN1eqYpXohw78jY7StdiuAyfp8+/GOfmUaqnxyw4zAeg4J0woIQnz2EHuXxwfdqdBNdUGwzhpoSXjEreXuG3hYSkTjGrAEWoch5uEvNz0P+NSRHYFKeIEwgOR4H9d+hvqo0zUPXWSommr9fj14XSHroWVz38TFj0onUOqmzR6+IXeSe/HfGfGeM3WEe6KR3QOTJc3anPs65CYHf7R5zuRt61k7lNdeXBO4GRKLCW5YtO7w9grw3EXFI6xRHZ6nDUh67c3fyGEeIrqPIF4PmxjqgAQfSUH9G0Sn0IEGrPam5Zeoq30lN+uRzNA1ogeFdJpqSuRlniwGDHGy0DWXEI1WGWlHjk7vRvvpAUG8uEAKuxKca+xEByFATFq5DPWPnrqm6MRGEigfa0tEZDuIiyc7ViUtC8A4rz06uK3YBEtCaiQ2hBFqaytz5ea8kUeM7f4pgyNlSaqCFmTzmQcyFncZJONFGoULVx5lla/Ga7bd2iReLuUvzdVMiT4rq9Nxz15m5YIIStxX0eNHb6f7nMuHl8A02q6NQl1+gTMDdENxjUgbgyyc9e5n7jBJZDPHUFfxhHPql1DVuep9AhLZ29/F9YiNc3LuUieqsyOt/bnnIsRWz9+zxvk0Ib9+ADeIb2FSz/31+jVDF6Eg5GCT5ZEhl21QKATuwW03tbohlPPvc5BsQaL2mCfTrCIUti0HFniEja4RQo5TYuW+9Iolv7G78r+Vtf0zN6PwpTJWrQdZAHX0ntplFo0HLmhsDtFqkrBu2OWKnELS8QZgBDI4ZEZPNXZuQPi2UYOm7OWuF0aLm5VbUp0n7adQQAoNAHJPvGX1UC1HsfmMXig/+4fwtCOxh4qCo9s0b8qwlQ/ZrjhXBbBxWOP8OgSnAttMlWBd/rGJBTCB4J/FpYI1MWdybpQNPtESMio28yI2DBQlGNy1j7rHVEgSVu/NwoSr+QhiFK426xUtn6MDflQ8jc/EZUbw8aVqiErHrpFJAHHhXmxLypKd+mWbijBUUAUkXZN4zLsxCkgYVVbqASApvrdZOhtSrsKPTymVPET+lQKncn6w+BKQ0mTjRhkJ+AHfnOC/lvD8AKSmryMsvrJX6b3HY69rVhVDI7rGTxI46Ec7R68KDvZTrxqpkUDHR56uxG1E9RIaG5vM0c1a+D9giXupmwnbXf6Ojkxbia2DI3WGfORrSF5bRar0Sna9KfJwYmuzqXO6U2LStijmHVRIghpCQok1iPWwlN6+iXx4mzTC3sBC+xp4XYee2FAZcMHgWyCQn4GLipWOlYZvypJRcae8m4fmQNr5VIBIn2YeBOWsfvCfYBfMIW/wpqJm4Mi5CYgDcoIMIRnAT70KJ0AldqjC9fRmQRsHNTOUBfFM7V40RbkaLqPE4stWvnQw9WgTW6EMIMRqD9iraLABdKN1GFlN7UqQTw4vXLAMlW108v9V4bjgIlUODJJt1NpKwCPPn6SuuSLMvdVY04S+JKxnl8dk+tbXyU6Mx2soM9GTc0lWoLbI1+6rfDG4eSgolElbpeXzLi/b8Fv8LW5+l3wOnclc5PrS+5J6m28v8smbRoOm8Olyp2nxTJuz3aXosoyOPynTlht+jnPL6qdjZOlBvsUETYymwqrOeYZxg+QpgL0vQ3TkNEFW4oFikSjR+8KOhYZQtLTd52iRXNyGKGfqp2Etm0a2OiY81VDtfsbdKrUjv5wPL43/lp4GF3cbsbJcLmcgI6/JQn5Ox8j6ZLx4SHtTaNwxlGQIcsrCNC7SoLCsbAhv2Y0f58TFu8WZF9ysCAK3auDAimn2gC4zs4Z372tJLKNHFhIy5JN5BY0X81OqWdJaneiYEYzJhx7OsrVAiykLXhOXODMYo04w+HK3cb7t3FLr8mWSqD0myGMax2NPeVRaGD8cHxg2Gn211oPusHDRLePw9Hy2MrPM+Nt4Yq/65XXfAZNSNDs0xBsuSafaZ2fFG3WFw1RiR7+aDm3wUspUH0cbWd6NBTZng0C/7SIetYIIvKNvhW849ews/u2HPqZKh35MGAoUOKXvjl0ZcJO92L0W3Qr2fWGy/eGrwe9m4xrp6h7RRvlOK7bLj7HIc04rQFReq3b1zr7FXxCLCZLHTHS8AKIsppURdi/x+0NKDs47JVc02mwM9+cDrL/jCPbhYfxLmDkpgxg0gTy20Qj5ddfEhOl9uAuaVZnxv6KiSXHMY83jyXEU4L02KfDNQ2t4BsNmcVrr2qV385wkRw7SsYcowLYChyyiVdwcDZCIfW/kmVfEVdGOunqK7X7ujEWtWA8gLaYQzidGe5X+sqNsa2DTv/3oc+i6n6JgNIYS1LsQWecdXtvjmqKfZgbzgbhiBfNX3C9wK8rQX+aCT+iFd7AkZ8aWN1rR6jSZTte2oALuk7yiOLSBxEW7mulmxvNSFY0mPObNaCfNnxJ9Fw2j8jSGETm3BsXQ0QGsZskQ/vI9gfU/ZrZIo/ueY5V91Z4ybXxkRuyDl6uAdpUFUKK0UHE7fpmftWQcWZ0LBCP8IGznnWk4vbgcas0JYCGmyxB2ph8OkvN92P3gcbVnoiwrf3qVskaKsV/G+gctxVg2QuMCfyuJi99ds4FSZpuN71Qwvqnt94pwdUlaO46/0RL8CWyNpJllPgm20gx8oZfWQbZ1+UxaqoatH0VZRynIXmh+NT99rJ7akL9PfXvtVH1vEwgVN0H0Sv/Ni1uLL4ixXchiBqMw2ZikcyERAx0Nt9WH1UTFeDblWLy8i8XRhw57nVyaWr6tTg5gSx1REL8I1lhEGEcGXmTYy7Wyd9LuQg9awjpR4d1D34EomWG2C5E0lc1yvkS42e2nLHNdr8XkMGKSzsWjWSVr+MLjmq7x2VH4ZuRPO9LsYrsoG8jDJX0qjeM/jBiCuejxNgxOoKsjLmGRMIK3WF/qhkYM6chyfxC1rBHKXsFB+ZPablUCy/HjIkB2g+5AQQm7Xq1NO9nOOwevS8f4hzUWKiNU8weBJSCn9Kj8R00lNqRrQag/gLQC4rMfmUNjG9KM/E/cFlFdyghbwbVISXJv5Rwowq8cWWwWRwpfhcPPg2qaD/Fx0AFOBawQC+e+Ax84+b37ZCpQXdoFHFhR0HgBb3cEuAaE7Ozi3bI0qGDtW1L7JvEYM51X8T8yaeXqjmyM1GxCtAOkDhQHlcsm+DOo22SLFjTCCb3WJ02d8lLTmWIPPp9jkVju5oDIB5ckUcR2nuy2IXsn4JkalID3fXmrw5TACOp3A8Oft1u399OyJ4x/pGSbcLUwitKqUaSbGJPTq71v2LIq8ceVeqY4LVkrEk/gl9gXCqKK/0PCrzFzuu2rO4TbJp5XOg+xVUGM2fUPC0CscaJanVkTeKnlE+uCASLGixD/ebOJdondXknvwrqWYLZnVq8tsyLRD+drVV+6INZsKiCh6NWYCCToMD/4jPIsbP/GIcq/nP/heb/XNMbUsabD1FNJxenfxVPczz+mXE8eh+6vodc9I2HeggaZDztEH7KhAKbg+q+TCePIqEo8ekS6ye7FojoCrz9GHROynD6cjHUDth92wXtLk/mc/vUrfRM+bRB3IcKUCJmERoOnz+CbY1qkADgDlyyLqIZ9rTmV0yiHynEOBQfZjPNFTakMYhkKxWBLiyK8Z7tHIfh12G9SmUu/LvQnP59ww1n0MZ1ATFlw25LGOvN7ZxYTiiz3bjVIoL9LWmISTI0ARnmQ8dUf1640RaFKBCTcHOs4ny3NvvuD83hTJDj29VH/E5sF8IrqDCmdRgeerpxbA7Yj+mqGRVk4XxWAQIAd38ywNsnniUDuyfL7mbdmL9PZfLyeaeno1UrcRn1ZqoFHX/kQM1w1BTmYVNG1WfOPWvFMXJPDd4CWgMkJXSmjifBhwVpcKFEoAu0gB4PTv5NpD9iImTRZ1LS6W9vUrv+Vursfcw4lmam/f/Y0oRbsSvGQrGDORzNotGm9MIUYK2p4CvckU5unYmIzr1rp14c1vWWYl2BoBp1iOMX7qzE/Iy/EcuvYBFTTJomxWwe3kgjxE+SLqbwdDnZv6Fx3t/55v43+QOZAceU+mFTFjyuNVxPr1TbV5naxg7eWCrrZMPmpIpZ9E3EfiJObKIMGFGP8JLGw3PhD0D+ApdNHjD6n75aHKDkekqAfeh/qBdYh+xjOofmX3jMkk4sECAPG3IZH7I9fHAcn9BP2rQqBf2sCsla6mKbIzW0GBZ3Kz/5LwWKR2DmNP0NNQdjmFxZO6UHn5VCVhXC/X9vWs/4PacJklrzFohr3EV5zxNbRfjZfviSecB14DAGjjY/VRnU1R14nRLdTx47YnyLsu8XQxX8PMLPlbMxyKxqpiZq7GAUPfEI3SpMjmoM2pEbGT+YoENyE/h2r1bgPWVqpLUYb7jmifSTXzjvRfWVoSmJkZ/PIanDY67Ofs4swVwk6CZQGah+6r/WCCOMECLvNPPGOCmBiYn+AndHGhAWSwCYpDzfStv3pI8oLrCVxi+C8FRWPU+uSls4lzwKPeAUxM0sikTsKzHiNoLdoshK7ProFOVO0ISzfU3F2gqWz9QzKPqSFQcV+/gBYlqLwsXL2vcPm1KFrUdFbMaqWeMf+hSfpk/XncTIKQZAIk5sow3mHEctjvHeD+8Z3vsoZGx2abW5VYICU6rFZebjIsNu5PFRnc6xP+KKggTWl3be50ki5nR1Xz+Cl9eyzH2h7E5EgJI7KRiMl7SIj/e36G3/5oRBewJp6HwzHNPx2MmnbFTvO3IqAvlN7t1ps4o+qHEWBZfpS3Sc5YCfxT7tx9mtwYXFnqJQZUvXXqsOza9uWs6t2EPRVNPxtePQeBv65O+BmjQ6amWC8ovXt/Ok77FqVQ+GCwXnJgjs8Xbk/bwvQsF+r+FmgGCbKFrfO83WxRGKiYfbWS9C94+eMiERTOOp3a8tqzFL84Z85bHQ+KHWW7IfsALKzcifJauO5x2CLPrIm095zVx17g7lD/dsonuXLalyfK6YM43TopkXoOCckTvwoVp1fMGCv1xRzJzyKjXPk6Y1wRJ4a3mY/dUlfdVz2XquXFnr6frdOPR3SdC/JcZO98HESYSHGV8xcH4pnmrV6h1XoTVMyUa2U5tsg1HNSa23gx4NK55kwzBg5Z3xPkxzkkZiPILyjeJ2oFxwnjJa3FgDjgAq1GhN2i0+ir5MyD85xJk5B4KEs6qdlmh6zKC/d73dBR+rlko0P0l04KmEycrSGg/XbvuSa7aC6DkiwlLH+yL+pyauj/di+bu7sZLFmX80u2KTl7zG+314enbPqXSRYCgQiztV8Tel+2yZ741mY5GhhEEwjAwPiU0MyFKiNOsRIhZ2vRwgieVFCPkbNhQ2yGY+pCZ+X1qjftcsxDPxl9k7PC4lEaAQjnbnzu1rpgO+DJUHe38842o3uAroYn7zT6NDuyV06Ye4xIiDbIGbr5JPeAKh+LbfuEFn1etW6oddTni2EdNdj44d2MvWk7hRWMZcIAzU1N8z1JCvWfwv/p2G0iU431ebQuwbsI9A7AxpLnWoswYJTUiWeeopUO/IlvtXV0WAPHcvqzIHdHca6m6Cmaa5l90t32pGVbacU6dvg27ibk+Tl8kPZJBnDVDL3GNoOTlSavVnFPqZa+QEzcdKAr7x9FbVReobnGyyjN5yiFHOn4BZMNy/Ldg8tPU7CullFa2uTfOB+R/lSDOo5uH1BoA3goKDtHwyPHVcAPoWSZmBklnxY/8kdP4q23ilCWPo0UOCVH67nUPi7U31gH3zvwTHrdEYsXL0itll41rh+Uqh02FV6/3UQyBtjc0Ygl9+CFNM9Ts2VUTCAbRuQZkWekhso10sPcj1s1LHOqYoz/6FaATdOubCN8RNWB6ieo7yFEsF1eXx4imDDwy3GFFIadulUmFmevMbLzKrdBEOaFihQBtdZpQFaNxWQng/9aDSa8fZJoA28l3AWzxxo1qtH0zFHcSnWApxZg2GkoBOexIQ2cIMsBXN0qaIxkutqGAmsj2cvEsuWDJS7HAC3HSYaLDmqX7VSem44WGcAXGpZsw1XxuhlbOvfy6+ZLG8tD0xILWTKuGBIP3jjpnqgsQB99dcpBcqksqX0qhowaI1UFvcsxrPakqNjgpIKByQ2TQp+L9p1rhU0KduPWlmN3EhrjD6Ik6RFIIoEAXBitlT3OA4oqJYOMMBL/ff/YKCyOr4gPs8sbymRtn9hi1mmLLlKHChGqXBJqRVNvpZfOFaWuG/HdMActt4T8KDrMaQI2BiPRJ9kGEK7A0dS87hKXGLqOcNQUrnloDwcQFWDjUdLKIIJbfseAeXnkMyc7yNr3Q6ZemhxQT5ErcfZSEqnkiIU9ymV8cAPomxyw5ItELkSHVimXAkr7wowVvyfLJhS5xTQz1kSiygiMpVlGRxjGKZ2Bg0r4NFR/BRf9sTalEMwi2UOnYfEMYAC1y0g+rfCvMqT2g8sts5ixKjULHHuScY74KYCr3KwhOkdpP522PUr68hKRmLeqQq98LtOM8O0JICGp10uPe1Ws1Fb/UN1YEh45As3iy5BBgSRZm1y8s/7BjcZOfSqeWtytXo+7gawL/W/hPk5CHhwJifC0vIBdLFALOlxBEfVrVmtRH3Rm91njPpSZz5JzkM2SQkI8mqfVTR4O0ZriTCt99oDGJfpyWBevMuRY3S57svVTtB6vtfXl26B6A4aH8EFaKbCIVO7PN5Xxz7imsBxkhuDkW/9hX56Zd4lmmADs1KVvUUBZQeWX6Lm9arGoL5dvtuV3rOVM4CNF2qnDFJe4LrAhRkEDFPSJRuMu3iH36Ls4NLFVnO+jBmApZKjafg1+X1SMXZaHfUO3CbfYd64LMjHbXNn28T9LKGKEGukJJqAR0Gb1d8dBU/uvkEwsXb5+zQfPGyCaPKVej58gdiPWU+fO4DcSxPL97kIqzQVNe3GZyTVwOROEn5lfuOB2eNvmss60K7ZVY08U1bgIpadrUX7tnr8ZDKMCFaKDkTO+0rCX0/mLWVrjDST0pKUxgTrDJiYGlhu5k0aJhFLRThjwYG92Bub5DYTKjVZxj1KJ8EFXUIvbfjZoY9S+zNEJBlgCLRC5ImgBZrQyn6QzQdzvdnHx4sEkN8TAQ7vLu2KDnyPdQ2noehCIqPrv9z/37gvB+0cLVeIYCKhSKmR9/py/pCJ2E5zNgHM+1C5iJf9zl8R8uP85WuzS1CKV/BNNbGeYcav/pY10BkUwcHYVXghtfv2wanQBLzP7uUmungP1eHn4q68E+RjO8JI33G2LmomtqjgQXhXzb2rzmOIduW80gg30WrNrp2wvnDSUaIH7lGQPLRhDylWUVMEMkcsrojuDuQLOHN4TVHImd8QDUIPUugP2YJK7OTnG92TgtA51KWf70MNf2D3A8M0Bx3Yr1cNhWzxMo2nQv9WLTsiS5KV3HNjZJBlAqTuxGEZC0YVE1hQoFd+ArK7v3sStcWfHtjOCfYcXUl+nK3Fo/XFMzQkM3CiJL4Zi/+Jg5iFa3mT7IOdbW7oy5IK6CtiL4l58YowQwAXu3Q1Y44TlS5spEXKHRkpdB4abx7XkTNfzaThsqvPeVguw98hd5DbVVsC5t5Dq8oQu2Er+doVkf0aYVZFcL851NWnjlmIJK47EEK0wTsWpg5tVOoHD6tcwZa5WujolrSUe6SKdL7JK1/db0KJOvWssBaAPiy7R/517ydz8F90MgP4L5v9P3sPeLCSFAOVg1WzoZGnHPP0X0l0DmP+j6Hk7aRJeH75VL2+XK1u1IAKT3VqHXqiAngfT4MrV6MJcJhAbdNKzXUB/jJUV1Gx+r6TjQ1x8VOBaedkNWGRn+rJN7Y91sQKKUi4O6br1HZoLKPhIPsY+pbxeKoFRJy3YoLTi6ehyBpwDYgY97fOLxBcA5hhVLBhVHX9mqjgg7HlvUezEnoXGgYx5K9zWZbk8Uedk+wowiwNEwcOC4izJRJCgkkA813EabKxwsQ4+1ne/WZpBae4Pg+jN8XRKXPde9JdBsw8djwCz4W8XrPoS6injyR5psANpue4XiKTmm0mRzCKdMhvZtLby/jv7KNW/Pc5DfXLp6HC9he5V3dYImTbumYsgaJtH3Bk9ij3hHp50KUCQQ3x6ARr/Ubo+wsMTHkJ+YOEqWL0/rYRIcSoU3fYVhwgTC7gwqYshGck2gEWHvGKiE7WcIh2EgFi/VDYLLyr/kscOfBb84v5eA5Wkcul0JehAFili16GWjb+5LR7sUv5TNYGWSfjswqlEjrvnU+fmsuNX3jqlPHkWyISolXcXrLFLorJUaMGBF7CX0dXbiCqvgbNR8hwYkzg4YJgvUYdIcjif/E6xOnjFqjyQ6ZYcymtmSC+vZCVL5GmZ+a1ejMyTDnjYVa25nGZyg2AGxJrLvy4xYpmAAIFOASS4AsLG7DW/yH89M5ebFk5GywqmpwT63mLOeEUKgCalzApVSCnb2vwAhabedEKQ5h6BUOMkhr7tc3oyyggtk7xlGFk6a26i9KFr4uUOw8KpziHCUpllthG5FxqZPkRI/SXN0vRaiNqiX3u+PxPtLGhy9LJRKbt5oZH4ZyaDbFsL4b+gQBSPEPN4ZslC9S2aFuZG8SEfYHdfhCLC/F/Z6cXJ7vm7sfhPietcEneD5xfHVcZaQ7oAW20eWM0V3wWWWO8KYZ7yvLvu/7KduKyxymjP2HuUd6mE+VMHT5nb94O2Lc5o0L5c0zCV3LycmPlqkeyAD6wHAKDs45YIoE3A9GQvmpk1AYxARQn8gN3Rid0WohcC/yybhOmM4TEJjcHWM+tgl6HrT1zjP9crA6yfv8HhdyI52kSuS6PhUGokwj8AM0NZoiLprpLkOL+ba+uSzGaKejMH3dTxk1cunwYfAxsI5t12c1X2I3DgWlTIMNtxeGg2r7wWsubKp82q1BHr/80j9RMzG6QxlOh6/d0IjiyGn+5GAkB8+5x12a27x8W1kO2VZh9aH2bOqsUtQTqrnt2C3zqWijBLOOhcLx7uG600gFAzab+q+8UNkmZAHmpH+RFYSUfiuXU90ulIG0PzQf2C5QGCj8+kyGenOFIzxSSl8PinocI/z719idOuouExH5AtGoqxJsP+fROt3cbZo4XnjFQvLfO4yruVS/YVA2rg+5wavSzoJl0cS2r2ZaC+3j1erYcBrXzStxA3S9DE6v+xYuJSwSe+EtN5GfRk7vMqsyb+NyXg84j3AJuv2BIhXHg1CeoItsgh1LlB2OsOyakoc9QQJcb8HRV4SKB3mtTpMpBa2wIdmJmptnBTb/XcyE8+kmawdADbEHYz8Dj9Uj/OqqChFPw1+4SKelNSjhTeePZyczB420UL73lsOkgph79ZEyag7z0swqVllMY04OFLfUXW/soi3qVtxt+4PNUD9D+Z/tf36erjEOEGHq5gYszoR6eDuEdHY1XhWepEc5yDqtl5fNOl0CfL6CeGmtd5lVpaAhnhtIKiZriEfWI9WkYQINpU/D0+IyJqC17kDrNMwnpUMe7ntV81qxaRyua+QG/vZh601aAVErvsPOjobLGlZBvf8LfsS4AD5qwLLu9KYXrevHvxdmO5pTNdo3zSE6oEghfhSvHYsI/vAyXSlaz+QHmK5i12gdV83BoZqonpwr5FAc6ZOLuWWI81XUxBxg7UOhBGmC1GAm507WAzviGipfVvfPtqf1oR1Ucgp7Njjzkv//lkYgXF1NrT3NvSdR5TkLC70orPiTOXyKY/k3yQl9eqvWdVj3xFYy/S7Gkh1+Ardlnal7RNDxVn/LjOs0RofkrptrVdSD9ons8MqdplL+XmVlVyx9ViT9OvPsO9ubD5C2jY3nJ8prIzDA857gEFGQtP6Q3aj2YOzGLEUPQWuFBSoFz640b4T7NKrrY7BGEOAEj7mxFt8hJRyx2P2NUrLcb2dhvyN3Gfuc7y+Xkm8RTtTNzuNmL2bNFumO5AVUlIGrbQtEsSg1jmZUbo69EimkdzLTaUA0xQsPEVI1Fusy7sHa7aFS6NMPGVKaSSl/c+6J0n+GmFWyb04+Z6WJ1otJVhEHC73KxqApEJcIxl1UhJ9Plh8sETpLYtNo3ARTY6Q8bH50FDpMWFVhBWN/AJHNIFM5oWBpPHJR00eT9DFSCNvJmAysWjGsIRdPomKcYhF7EWLIvlS7VICGjRcfQNDz6Mh1sjP9HLC+Ju4XVul+FeZ5hOsAy5voM0Ec9oaOm3NaoO4h4JVpGpmuAWK4KFjOtIjoNI/vZJVTqYlhnHqsqYhNf60FAaJmF8PmZkyHEGlcdGUzWo5LPfFqZYo7O6bkERu+8qS0WL4yZUweMHuKHmmwPHFqdlxY/XuV+VaXOQSYrk1n9aGzGRG9/DpY1pniYQVQ+oCb8adyNjxcLXh0Qxi/JeuCs/AWFpBD7qdwhtmNTWmbS077outBQ8kKLAsp++45yUQ6lHG8aXivCR137BFj/5fZpIzRv21hCJyBMhba5mkxFgk/NCtbILvtcYVjlKLa6JLf2Ib8nODEyTH1pOJOyzzL9HvzC5xUWXNhnVXt+kmZcwucC2/LerKi7OQSekBG+HosnhTaOeHnJVveHkB8rMvg4jTd1BLjal+mzyXx+6TRrUByz6rTeEqMMtOIfT1ZRIhIADcc2wU/5DJzLp3+uHTpBd1/xC8c6m14V7W7C5EZI15Yjf1NTLjztnyBFZTDy1f9t3arD9E8RzbiQCp7cyzqjU0g8HcCdkyTCDL5QbIhsvdfURDR7R3MiIlUSMFJ4ma3eYz/KHXceFvhNyvmactz6qbQvrLBCBWLJZJftCu8iYGLuGKeRvoBDzZk9nczb2AoSbDfyOm4zYLidUX/lLynPhdTqvoaPkrlhcWur6MhdxCuSBbP8uyaKYiX6a5V8ZdmNmVV737ARgm3Oe2kdiLhbzLZ9G9N+BWzQ+XASZI5CHiQLK6YNyiONSuytlEa8egfMqnOSkf03b6/Jtw3WQWw77DajahtyxaPj2Kahe4KUt6flJtSaTbTna1waG+yPLi6YmWdCZQPq+Yh/aVlOnUwXp84/0loOS/stAWYa02U8pFwihY1h0eaXQDZIF59Z+60SwcJa04cH4g72DrbXgTDExrJfRcmQWYFjFz+T3Lw7nT1gwCJ+lN1q9GjgN8Pa/5qZ+0SI4AuXTHZMgOgTSHoUmya37HZztPPiIG/jz1v2J4BRdLafFiwNYL16wxxZqBaP+6bGt4WKASknE9T+KkZNd3PqLgo9zNrwDRk0ni7CO+rayq7mM0UbTBvXP/sTzk8ikQwSqVu62nf15s2D5WinejevbZWB2khsbEMKDPt689hzHscgVk5KmcC2SXZCXnIB0y2SHFO3jlU+Irf2Bpms+/1fCtFJOoLLvbbSNqVYKG3nKUtFgQaablaLPzmFk5syMf62qybZ50P5SBx0ebUHXYoC2PnmDrKOzHee35gmzqW8Us7Wi/RtyBeffEkgNEp6zgF/fybPYT5b9jfq4+CcN7YqYPfKLF/iaa6lchLGUDXEF9qetu+G0SvRZjAwQ0NL7Luh7ftuMC+Y5bGmJddJPz00raqgb4QABdq/f/FT99A4WoJn8vve6n/qEUtEs4VQl2mookOuVLx7fjoEmNyS2eUZt8oWY8WnL19WIBb9FatAMTsnNBuT3eT0TEciKJAvmEJdwpPpw6HJMkYLWYMZfPhdNqA8Gzlx12ROCuAlL4E2MdSbC2n34EEUB4rcXm8S4fvZ5jCfXn7yqzHQmot5b1aPTe69M62U/DWnnFB/sp6UhPi5qp3uTcbhXc//HYD5eLflbjTOJKQmjxJiUJ0R6tR4hdyPegR5ErE010/R07OE3v6mDcTa8FLi9lPxaOkxn3FuTYUaoZcxaMV4qjvvdVJwXvjcf9fvjzATttnybz2gbO2Qq2aHYdHPkrFHQa3rT4//k2WirV9sKnBOb0gMmEQCXngqG21IiQyMHgG4xM02+6810+1ZlNOVYuZlw2GqxOO2LgawGoK6yq4WFN6EkhKmuJx1km94D3DqIedlbK4rNiZ/Z6J38XSjs1PMD7l+BkL8V0SiStgsCxkdFfUuPGy3O7A/kiqlORscQ+f0sEgMSbXGkXSskiGiWDsNQxBioPFwuNd7lK+uijUGpY+jgSHH2OzlhnBzDFX8zYeIX3zorouYJ6wtaJp4dCPFQe0waFX6m3v68Pw125D4xfeJAp7HK4Pnjc4IKqgSLUt835oUsYAvxpX52nK/EjSt3e++rw69GYBwhfRlLzyBFQGsCvujslwCApnY37MG68oDPg8k84bt7m4mLNvZQpYCQF7/1kug7tm89tCp8ujSKPHXvghXd4IXDVG3bzeWd74SFrDKXi3YzcFhCn6HGmk5a1eVz4lPSL8SZaXP1c3y4BuaBMNWOzKKGB+gEXlwUNNanSwGumyC0+O0V94B09KWC0ueymYgzBY2iTjAUA8wVy87et69ch7jAvDlw2eVzjEjvjcl5iHN8aDeV/fqhX4FalEJB5fhOTX3vs4gfTJ1cyk/+tjHaALISgGcFNG5GfWMJJZgbPGMiwjhaP1rerHqYReXJzJhSn6G1zazufTRlbu3GrQFxA8Uoh9+2ej/dmrJ4p83linZGzXfN4aGnvASxjOYNcVPTt1tDXiU0rW3RRyyzgI065ELy5CEkaUeSIspRDUI8k85ekpYttZ+q4UldXx3GJuZmCQhUig5YnZzbxpUMl3sHWrYKJYj9oJ92oYDovUcxSryNEmmx1E4ipT7mELLNbmLnrlhHTAQPLbiWlA8EMfHBo04U2hPXpb3O0k/CXUDwBAVKFH6lx4cOApRnZ8HQTPqF7ff9fxQORemN/01vXn1Umas0P53dmst4U609MfYnzmwVXkSDLagY+22eR6hNVK6QQUrXVRc/a7F6y65EGDhJMQt/uS8mEEYbLiqa+yy3tpcqvyuGUiTy4bbWy3vto5KFqXNa+RTQ8rRBjDHohr3vMkMJ3Czx6CdkCb/0ARI4bPdFdiFhyVLOyZ+RV5rTM0zBtMPgo/4QQT+GQNSO1PRvserD0AAb/qLcrxk2B5hhm0a5h/+7yT1tR0DjVLB+x4koX4G8UI8S64nJJUCXa59r+CbXPDXvjyOI08+q+RVHmXZqPw2ilegn7FrBgusYRCUgLqNjkywThIWrXibRO173IKdy05bItzjJOetzaQs8a1euXiKbrtS5aAPC0nwOg6XrQEocBKFnY/34L6bU/TSF0hoKm2IX4z4BkWfw4NRi72Mh+8qUdfr21XjFYXRiJjQBOr4qiulqk3nnH5JiUGYaqf4o8+2G9gURq93I04fJ5w2lS6CICC61hQ1f9Pcf569AaQ4diNkKA9DsnhHzza66i58jCHP2foXGq0PE2+xbZaK+HYti6Aq9HHTvfSG5D75J0aH2lOhRhNzGfP086Rf+4PZTcaOXBLyaHdL3DpBntRbrb0JCHCmd75GKSjlZYZbCC977PTT2Pr4iHPDRUMiO7aA2+VR4js2MoE0rm6T3KvEmTMqkCwKfCTIZIhxIpSQIbi5Kin+V+Q3aTm1nLduRcCmAREjxOJl25tTPNZur5dc9yU4fQ/qVOCbt/OTUL9hff/hXphpkayIUdNT2wgE14KH1uoHmcYBUBO1ewVXgbhpb2E+stD/xV8hNEQuAf/Yiqo4iyJKc8xOtjkM2DW4EMLf6BOjSR/FgmTUyXILsh1RGSyP6MoDyOQLCFP163i3RJg48GjvNpPr9oXh0zh3+zuu857RlJ4HilLjEPn54fHkxabMa3vrfdHALCWFy4xPbIEQ7u3ViFr9dEUCElwPAoly9ylsEc2OmgPl7XF+Iw21cqERuM10jR60OlsvStGoaKHCgB02GhLyANo/C90m3+ci7wezAnOPcrFi9DpiZgpThMsVXF+YdIWo+/FZ/YAyMCBiUdUqfU8CdFlJ5fPx7zeSMw/crpOySX08GWBzoBqXyQ/aHSUySff3xM2XImvvkO0Ybe93Y0Yt8z1IiJKl57+6JvzPgcUooy9N9bwbBQ9C4WMoKrvIjqb51xvJgpbAGwKZ2A76GRYhRd64al43q0pnoanjegY2FBI0u/IBUnCJWzx35B1qUdidY1RFh6xGTwHKNs+MS/fG7Xq2aA4OwL54zeBhaRJXO4r9fnpX0DizBzfRt/bkKuVvpIctgM0xGqbUZob7JWhrHot3yMjneheJK1l/GUl+VpcJu9MoWcnQqDNDWG6ympZ9UuEjbfK5yzQlfVP1DWZGSluFxtNs4wKZRY379NHTmtvn2r3psvOMWVURNhqvr97NZvv/1A08nI/cEL+8J222V++vlDqoO/CmQ65AQTLA8QuHrFevooY0GYLa0f7NoK7mDhRWCpdJujMmp01PiArIMpYHDYClKqGdd3+3rR4rUowb5gKYFRNXzF8jnQVvjUqI5THDDVGhSn99hFSxFWDw3yhseO+2BBLFRoHeu9LmCRth4nHqOYjDZnnvm9OGyI+qKxCKO4MUq6u+GUEnRaHN5mDnBai4Vn9mZZpNv6eyv3SmRoKq3I5io0pEXOMies3MxbtAegH0SltSUQse3r/8i5+fSxPqgEeDG6a6uRkcJc78b7P/TtaSaklE4EC9q8+ElaqSdQdxY7LMgkrwEBcGMl8Grd4PnQniyyLxuXBk/yE2zo8wC5Hjx2rD5AHTsnx8cbEJ/t/jETaSJGYRVj4/tRpkZl6MDfcxhtjKfdzS3RcpnHSx5x6FWZZ2Y3UnIBWHpc4wdAd2cfYZktcKu2gYds+GlGDjNWxP0NrDcIcMHGs0ZLkSFlGNcinGfGcbBhiAPyktao17WMRIhKGkIOwk8Nl7K/QmEQNqgRyESe4hJt/OZUQZUNqt1V0TIQDCS2tJelr2g1Yn0WUrblNyG0neoJYXups91ojHmVwzSQvKy8DvPUPYQXm+sdEq4L44MSvQN73J1xOmiKnE7o0IQC/YQXwK4cFDi0/u57SozzxcA/6ljyV8zvtQ1zBWlpwaj53G59Kp/qKkfFBxAxS8Cm3A4UQtcAOx2U+T/778cZclvFuqB7gzs+RZMyC+Mn1H91NWxvGsEyoPo13optEwZrXjxGhq2ZGPUOxNh8IOsGkdAJWNdkIN23pPRp/QxvEj/RetRz58ZacFerLS4woR2cRTAfX+a1wdMAKmjVlTusnG9WkXYtB7S31lQAc8RWAvGmn2OZMM+oRcQv27n1sNGeo+q9NlfQQGZmxHsILAC9/eKdCrIn5wan6zcsG4in5OK1CQ2DjdAZnM9wS0B0UCY0I/9jWWVxMnkxsvsuwVy9BPWhVpwT4vDlA84jTmUf0K/WiYJA99sxaUTG9GbOGZwLEL6gQOhpY5dmQcfVpufU0r1IvuI6dUDn2pwV6ZJ6U36e5mAO3QLTYVRP//2xTA8xzCufMoBI28HM3tTPJHzI5QaIKLFteC7BpJMdCWazsQOaifbNhlPOnjv8psNujOmksE85UOOGNylcV+HBcu+5JRFwhwd74Ef6QczGtv/frSaVvuMScDDw7ys+ZHB+UrvvgMR5OvjQ8Boh5a6NHRYHMibCJK7ZgTiSuq3tFXZvRebkqMa/zyfPZUodUurJ6BsFheUli8kM+IS/8CjZFELo+nHXx4RS+nE9wCMAM4YVnxKgI6YbzI3HZvQtyHIrqtOpBGSF1gtiMWw65GIyAcOUoMbodeivtVULL4JN7qXvHhkrPDPYwCiJWHs97Mdpf5g0GQOujfDMxb0L/3oo8GOLwQteX+ysHJHsQldcfbvVeqvojJZ3MfiWhal5aXdkViaZG6VT0NDT9Lq8dDNwsAkD5Db3Q5Gy9QJd6HD/qxrkcDoEQru7aUWPVJF4RBEF199Xaj5g6gMZ44tyWehiS8sHwYGF0pnF93mIfxLSmQnUkV+jhRrfi03j+VBSaaBJ8TCoMPuSEQ8COoAgaH0hj46R2rrL6v6gXOcct6iQTKBLFVFw7JGZWGM48JqUpbajZCGn5//chANeqJ6UlbORh7d2ozKsQ2P8Wd8wAvqLHztQKpd1s3ytIZOnPj5sui8CYrxsDDzZh0WDKQLFhz+QqatoQx/nbkcmeM03/6dCGLMWfAI7x07K/CNPngWjyVjk1r1/nWfcpxTbd67gNvE6XK1ngtelBBGf26FINRTwLh2F3zZvoHVEGgTwJRQQFbZLuhMtcpFy6eeq3WNkNgqTqV7YQf4S8f3CYlTrUbd42Ct+MOIFh+HXGlcN3u0WqgZkuXmYujqSM7fgYg4su7dfRXUbepb05+saxfkq7qv2YavCVDxMGSWgBo+DP4lc0QdRtPc0niVevCK9HfFLgEpBzgPTLkoZhILB1mUQr7UdOJ02a7frOs+7oFHruC03alVjDRHH7qzbzQzma6sx1xoxhdbD+vEaqdiTbQPqgCwCm+jcxiEqHyHrNQrrj+1xT60VSxbBSyJTSoQE1tg3ltQyXFMEW7qdwsEvcfrYOQ+o4yrPrYQuPu41yZcN2c2D9SJ2QLSFpf9JTPNytqBU6pVUKjaQdQfpkbyuJi5SVL0MbNnBDtla+UkmyhBv4f5IIYBUUIPw+cci6/VhUz+Om9rFR3WZSHnSSSqxXbaPblqyh0zOhVtEKkerIaCBUj/rdiUitY42u3OAS/dw+nKfBflyiSHqdClL6eRleVUbjJw673cjDtyRJbPqNfpnD4RXg2YyjXiwPhla9TLBHLmJUVyFyNNy3bZaRYWzOMedu3Pbl7YIcv0fuvxiSGyo/n1rcvUznVxQoyV2sCorLTzaYtYFxaEvelj19LFOgV2emcOYYNFbxhuMBXIPdo49vp7fj6EjFyGtBsjgow9LnhXof5qnEXttACjPgLPkFGhXbMk45cLuYrBgU4r0AY4yRSTTXlA6M9d8FUj7Nk7Y3WJXvjhYi+hT3guNhxlryPrA3HOcGAx1GNg8uuoQXVGXIyCaGAgreuDtaCJBk8ivSWksWZbqtvBu9QzMMceT7+xB5tnacZ7+jY06O9yq2l0OGNh3H75P3aK7NdjLi9UocUvmmtkHQrQuQvQLWvH1KfIs4YXlGyF5xiLE3X4uqGDixyJDiZ8nhDQ103883moSMik6jCDW8GxcO6RHxrOWbCQGvDeYTStXtIBQjOOgUM6yo2ndMG/KppOt8eb9Gqi+6m7msmlOSVo4ZW6l1tKAXS71KljVfu6eTNVxaRFCKNNHug0aUhrRBahK0dU6v1iR7f7Gm/oW/xrlfrAry4Ys+a7aeFUGCfsMNdTFaryLXP95cSVdN/KohnFhLKsqs7eAr5dE2W24mGL6m9gsQZLp5v4LWX7YgTVczapTOe00KdkFC3apLOuVecYLFdA9QKfjnrjiM2w3XWWCGVhjXVQYztjTGqBRZrpn59eLFEkmwrVaOSdOqEIo/KZnz0UAF3ahgcJ0UwJ607/C23etbmsHG1yjpi5LmxRUZf88Bkp474gRDG9PudRageKb4Pp5rRA7g2wyF8kr5PdIpwhrPH+Cv1t+ZfaFSsruZRi3NVHj27T8aRAUqMdiKueLNG5Lj7qNfhvfIFyZydisBKbVTnQo6StVSns7SPceiQy9Til1SZhgDmshkwoJafNMOPc4D5BEiVmK6oH1Jj/7oSwbm2UG67g5xYhwH2uycHw+u0cYhzednSJjVB1TQDoDbzxWmJRJSdfnK+uGKpLpin05oolwSE1qA7b3lIrudQ3j1yBMfYD58PoJ7iHaCteL/o5M4NGOeNZhbvdPQakkAK6EhPc8Q9mJpDPJ2NSzcNnXeyla7oB46FSLQ9x/1/c5WLFSX/+WfACAKDiHAlY5Pf0tDyFmsDIGsnHyeR92DD1JuKYamwFc++lNB/XHK2pW7bD55XUZ2NmY16nxrLUPyLi6k4uZ8MBWNYmlImtYOiZe73FLNLiqE0FMSDfO2GGe+V5uvECyTMq3JWbF6xd4cVkGLkZpvdalENryhdEVRP966FTT19H/7/+GTpTQ733hcXAagauQMyNqpYtaGAlXC0rArtIpys73dwPYWc/nrtkgGhRSyO2TVf2PozlXU1YUV2rCAp65MZmaulsWH/cwxSMPyj79qcstdKf5J7UDUbnl+67UXcee+DVPUEpx+pTiWbS9oUgBg2qZsE6kRhf2EdMhb5rbihnT4l1YV2cU22M1p6iYOfFYdWTFCrz4LBT61U5ZzGFcuq3TJb/4ZudJCSEAnr14asJDHTM91fKV+6u338W6/41A84qBRd7F3twgmMtBXp12iiDNxSFVq43UgOdxiX3wC+wYNmLfLwAFs8q93trbQ1KnBAZUxL9147fY8vo3PEeZBQuXHgs05zWDeDhqezptZ2DFofAFyA9oyZXmwrkdUY/SqJew2KHAGdMkkXYea2Na6oW8TZesbhv0ySuiP/n+6fjN+Lk+461OP1PqcBWCABywUVevr8rgas0xGDJvE+qpUSUVy3Fp9f7Qj+jKbbflpX3iL9SOju2LA1ld0MyEiVuK8vTIXr4SKk0ZPCiXnbDLe25KWLffvGJgKupVQ22Pek0AONSML1jbDzFRCHq6QrETCpg82PWOBfoPVxJYZj6PYHE3DXq/qHbvDLeDiv5FwVabXR8YmImh+bgVEPgR26Z21xCbNbukiLSjxz24qcVhZ3KDnVdVyVx7xGFixAegGcEMOPTTQxdT+n5gndMEshhJBz3XcN+gamE12EkC6ouj341xYKBo9w1GjTf3Xwkow31u4F/Ve0Pi+hraxBUhnoQsw97zzCXamfZgYXukiuhXIHgC1XNm6j8pmOynwIsrtVFU5ABLMM59Qw0YulMJQuOPVy6m55O83Yq9E4zr/nxUFjnSdHEYUvRM+fpaiFwb++Cr59cGDTpDaeKQliCiwP1dh4HZGljdxY4PYTyXdv0pkqvZt5mlbXrNRKMPXJx6DBU76Tpt9EOnTUSxWBaEMkhhvtFLpznhlAfAAfW505xd+x0eUFDifnyF8hwvybvRM4wQhzAj3g9mYJa4dQ+FZjs/6JZ6nxmRQZc3jEe78KXUUmlig4ncEGFaLM28DVb7lvg9HUKapyQrTW9JmpprsFvuzMZ8rXLPP9Ns8YD/ax4dY6jchCgpwfjf364iOFaJ5Qovc9GxhxyyOyM4x2TH6uZf4SaAPGTDCMaO1WNunFSeLGzREwSjtCKFx912+DEJig9
`pragma protect end_data_block
`pragma protect digest_block
9b4a68405790b55296a4241942f890c45bd2a0bb5204ede5b867d5f6c3c31b3f
`pragma protect end_digest_block
`pragma protect end_protected
