`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
3Lm02tkwmCliPQO9fTNdVw65y8GxYajSts0f5/qhxqxBzLtjwcnREpRgykAwGRqse6FidtSF4TMDSs+x2y+ZqiSGymCnc7FSOAHZQthpI9vTDWGM+58UZlMepaCcH0ED35WJb4PmxzrRzmdNy1JvuacSJ/hgB1SHrpi1Q9TQpODPRL5fx9Akm5PID9bDmGWQg3CWCUw5dJLrZ8X/bL9mJ9a1uAs77b3kj6wP9olCjNfTQQUUk1D1X36vlHFsTjQ2P0qBdx1/FVYpCXSaaNzxyNOCXLsV5RZP+dJd79+9F8e1bk5upvlpAFHjBw8pxNbJopUxRc2RRkziumdo6rTnUxnZDf8VZsCGHDI0XauO3rM/f11myinsUc6CSEMH4IHwk9gClMdSWRB/2ShG+e8PmdWM7qWyNIKaWX28VtSPcNq+buABFfYRCAUjSjH8STTruqVYtzKqUpsoN8ZhId8bW3CLqgxGHNUzgYj1J08iTGmr1Ukv8BoIpIgG49MtKoafIsR3DiFHhF80tCTVHJSJJWCY7aAh1YW56FKvhTIARap74XbZksFzmhbbcTSrkYJdks4U5iBvJMkMdmj/WKO9PQXIPymiWRhsqRUmLXlQtnI1FtZ4dDvJ6nmBDveNFc5RirDcg3BNy/vMZrVCeAEhYRCDH1ypJd8EjNs+fzhnV51uJv6syuZuxIwhgAEpuYpfEYtAvNiY2fNp2+bZyyGaxuagEo9w8uZOsfb0RSdcWZ4dLnw/1PQvArqSf25CdP4CZjr6xP1LAXLOAAuFIGTXQ57FNdsSi0GJtchFuc0GYHk/yuhCnIje8DCk80mIlOY26od4qENDgRprl4suHM9d2Yok6yBOiBMiUxFvNZoDhX0Kn9owIjzvQy+lVVCUFz+aESx0dP5oh1pJbJA3LYTIehjIL7P8TlRB83Kpcf9nHzQXTxYfLqt0Wtw+owF5HZVy/dW2mV0FAKp2TC7iBeCoD9pqQyrgWgqdmveztNTWg/iLhRhbmJ8JvKUe5rc7id7g0dgm/bIk1BO61Tjfm3I0HY5UWl5Ed+o8Bo4LXbyUwN+GY4kaFpVFOtN9Dmu/YbuzAA0SGOLmf+elRVp75Uzgz+cBpEXIfdrKp7VVlkcSGMNXlUlqCj8NS56Rke7GF2uxwWa/wVBojMHyPU/ZZEfTTQocI6P78sWUm0F844FxpK9ELE1iuSSr60vsjyGKrKIevmwBNPfqdBxPBA/TzZO/nR8m4kekfMO6CQacjzwC6qF3l5B+MyTd6VHnD4n51zO9As/AeiHboiA8zIubtGt7xI0evZUiKMSCuuW8Stl7fD8BGh7U/vTWu7PFGIs1NjnuDkuHAzROH9nXaCnE5KeIZ38uVpq/fsZj+TJrLFIu4JAPj43yqaEH9xCcdvaLBG+3VFd8/4VAgPgkvUdugc5RItmWIOJ9Lbpe8SgV8ifMlrOF67qLrlA2VMYsazYLP+gU+oqpIpaok7t/SK/aRwF8YkxVSPTNGK1oMFF7V5Qy6nRKd1To+abWChCOA5B5av4RK+AaVTSgKZ8iBPNoDhTPuL/+UQSmbq6HlAcwLag3QV+GVp4sMWxXkwjS8OEcb5fhdlisHCEI/IQndtLYPeCYikx4zQJVnvFB/2tRYLp37QnNPFcuIume9qDBljkl4AIl8WGNIRpHQ0HSBr+Z5ThbSP7dpyjkGVSr3iox/xE60qNgECpIufhQNQmxEcVhzwvG7Js2GVBc+JhVAB5QSuxQor8TeVkxB7hR1dbrW0PSfRB8Gs8k+eSVH8FWUskwbauAm6ZKw4KRwZO8fSl4i4uUZ9GJzGe7FbSHspFaI2YtbqUgozTjq0EGKSVv8Y9zAot9cW6lxajVZdxzcpzf4eD/wNNF4KK/GKr9Bq2xfUN9RDrMs0r+gTHWMupoZRpeWUwYlIC/0oZymor28ALsz6WICCAGl0HnuWFLFl4apl/TabiV8ceKWnY9l+M5R6gLyb5/di1/NoqW9sxUUM/YLvyoD6UrDZaOi0l2scggoyk7T/HaYCpa6gDtxYvqqUiDqQuv7ojbU/Ho02OhNwhY3+hHB5c9ymPzUNyuUZrtP5vYbYWjKG0hmBNk5hdHZ8GdT49mgdcMZlwwX7+CpyZJ70lXu8ibDMpEWuPgtv+gG1E4wtLGkvnS4tQIGMd6fp1dcVLM+o+BwK6RsuKAJziJ81Q5RQeBr5LplXGKDDLKqhxd+KEBZpnEoPSd13sH49M3Jy373FWcCqgDl3knWDLI1gLsE8CrAvNDHMmrhbkiVuGnUu4v9wp9MMljuSi0XHs0/Z2rIOoXGhjPmY7eprl49mli6ryLhf+bdPRnBTw6PKlPDfEoBhTRRhHG2biUai3341bxFRfO3Sr1xxxKK6+50Sb+yi6y1yi4vyZppfRQn81L2YNptNwec7vORqQ3VXc8Zh2gQ8ORU/UZa2QVKbymMKA9/NhMtVoQ9sgVr//xWW2rm0XIB7IEf/ggn5D645dNSQU7t27vukTB4evMl8qeU/PumyEzUo24fjyTpSZJeMSr4CYX4W1TkC5CVkjSh65gA+GndIFyNH1PP0ZlWqn0NK+79FqyAAZG6UKxvJcyxinB8doC+rsbug4itpp8Ay+rPsD4KzHMrhZRIr87YVyGoCpcrCX42TEXiUAhZVV4Wj60Cyv7tPGvUmtDZm2WGXsm+x0DAVLKE0pmPsygPUUuarrhvJNxq/+y5ngBlxwBoFjUGC9XSF8P4qSsCRZXHpB1oTue3bv0DsPo9V/8CaHvmr67VFSLGpsqGff9fOZiei+qPP7tpAvm37f97jF8UwZTF5yD4IfrQadje+3rrbCYWu7o/3DBKhe50iZribc4d8Wxg/lT1AIHjUSX02DKkg1wqbE6xqk51L5R7P+OxGlC40eEJU0v0RJkip/02Mm07kGS+wggLTIvgbi4gMRxLTqXsy7WNEIrpS0Gc6FKWZ1uM1u6Xf2LQBZV3t5aS0G6e2VU9rV06FXRwki9LKvBlBSTpN5hRO1P4EvJ+BQpAGsxGE4jWeG01Srnb9DJX1hkdl8dr+qUebzxO6x6om9TLaaAznDaerI2nhnRhdDNhDh7tJtvzcGTgqlPtR3Rw3od0EIbhzv0WjSFKCkuiO3Yb40XvSPpD6VHY2aFjesa9OH0m8/iaTqrfkYAF64pWBodtk8y+zArgWRd6PruaRjsaItl7dXrv6EQzvhLtCkgRvXOk+U2JaoyjNieAhqfr3XDF6QUoP4snWeNoIKUeaiVUanXmvvEWZGOCp/j1xbBUpv/7CPkbpZ5yAf4Xsv2Jr9h3V6jFY8oTOQiHINQJDrqaw2qoI7bonweqxzRWtu1ii2UuOEYzihR6JIEHXyqxp3W17kgcUQuox0d7N9yF4oNosWDEqtwAsLvaWise3NOn/tfvmpYTMNyzgF9Wybuypj5EWfPc9Q+eMR3SlqDopuruFuBNI5TtFZoy39dZj38hD3a/+L5sqhSd8XtsktGRrTV98kHbXeNAsXmIGNNd79YgNV5MVcBTHO4O4Vn1KoFA2rLD8yUD3THqHzKLefTI7TwZ2ROAdv/i5lG9yH33ipMtxLge2LTExYjrWcaAoRODCgj7Ui94Ujt5P8yL2kZBmQlhQJoLseQFrvwNPAa1eCTyMgjrjBw14UNZu0myWWoYowj0zVRaxp1U3rXs6BR+v54HFytwHhchp/IXDYD/l/HXxapAockysNursjFC3OduTWACV64RnX8YEhaIFzORThMtvvaopPIE++/PlrmbisTUNezptHX08tixyJLgnSegzeeq1cDL2JbgDNofr4POntOhftSubNV3HtMzFEjr8Wc7GlUFvZELLCo9Wfc1rf8cMtjNGiuPc66uooQepvJfMSvM7BugDdhi5jCG//bq1+E+S+W7eym68QHKI+JHZdLmFUU96YOztkUjbJ561/4Pq2Cg/TsIs9rJF77pV1rp8K523fA21IeI/7G2+6WVAXu+19DgPfDu9kiqFvyV7+T4JNMtQWK/3JkfVQO7j184LTC1xMX+prNHLeLeg+aALjvKlTOmoZ2BeArQxR1rMu/syxH6pzG4RbhyarPSpBzvmhOQmFue9rkqMDXY1hqI8V2ujDlqB9FT/d90W57Kh8voIGb+SiNEyyPJH5P2brB4FFwbCkEaziN0kYEMPDYGW1YSvBuFpLztbHhUGPZsmjY/VMeIbeE8LuuYDrHKwphVK09Ik5AAZxqCEYboduRQN6MME7aY0W0Jg9lXiJChy9BW0O6BON9oPLGcpQynw6vz1pvZLUVq9qH2JruJmeefNm8vXY2IzbYjJ+wFn1r4jgwZSWxqnr31H8dmRNE5BODUBnGwVwW2K0/gMtDzY6Mns4ZcfHkR3t4csSnDZAKgcYOm+PnLYXfRbE6G7nfvRn1U2M5brfiEHNfT3Ct5NShDR508nZDaPXe3Xs43DhC0VlChE8ij6PlPCC4S/tB9QkTvisOGtXaKk4d2ky4pm35e1Y76R+Yr1XUpQNdkxvKkIHxqEPg49jyf499TY+Kp427my6RiIDrU0z/IORgFhQgExsnTubKLMisoOhF0Q4/RpN4IWxd6OA8A3tCq7SuYeEA3fmlUezk2z6Pzep9JhxdlEwaM+EKuO2N3tXMyJpj/cfJkV0XV3HPq7rct5dq44R3qOF9ZZKRUfv675ShofHsXYMxlvwMnPRKSmlFGCsq5XbjI568WlnkNp8PX8wLeCseNPXSzmNBKnKgomqZXRBcMzRnkgZli1GmvDezF0IHFckxt6V/3nG8gXbxzRaygSA5uRRNXdDBRa+N7VXHOhOEjPbAaBjzE7oki1ym2SP6GSkDHjZo8LTwLqYOwKuv8ML0ERjzKR4F9rpTvjN9WAbjObxmksNbTAL2HWRp+B8w8+lgs6tqO5ZsmwgJpGF8QJJ8/Eh1vM+Z7zrybQfP8uYwTytMHMpFR6uM+ItXlozUJGV7F8VK9ACCr1MUdwUYNDsw/+ZT2nSsOcTpSQXktqMhgJYUpw8f1MTrq4Za38ipvmyLnAOdWb3EgY1DTGsZW1c1gogeUd/0wAWt5497OJFQuWpG/IGIGIODCyHR8VCIfFc0cqYMOTfZvT5ybowd5Y7SCg+qyzd/qCQYWZfOHwGElBsqH6GAyRGNSfAmIXSeVUEly3EysGrX/Lm+xSlbYiJYbqsx9hFOcLCAuX4SXdOYggQDWTvlar4uv4lg50/ia4ZX3IPHEO7M0OhCVWyNRiHCJBEyOEglyhNF5k5FzmrL495fVTfKb6pAmnYpk+vedZ41mBQBcfHwu7ZIX0LXSnkgjWhrYPX9YA2020ENd2OeDReRdnguGrFHLoZoNGLfH4G6J4cZzi4whs2KJaj5cD224VRkf3D0vTZqWy3Onm/P8vj2ZjWazuGnueqbnxmk6ukZpCW7/ki8XkOTvNFWxoMj28U8/AuyxgmfhK+Aja81q1rCqWAVPJ6dCwiEGtVqlSCf7r/jRtDfzFRiwcmshsHvPrs3JZBPEppB2GoC8IqxQf0j1h3M68RW/Xw6Al/UpZ4DBr7ujJ/dQpoEoXsqRzFItUyDo+HNOLzrMIqa9boSs36MIgsY7OKAFZOKqxGvDA4QEaqF4KFJJ7BmylQqLGcca0SG8nbyAp3lhnHEP25004AYM9tLsdBoiw6MLFsLvHribGLZL6ZlDvSBi56IJka2jW0OJJ+u+qZhzZAFLuVvpUnNOcbN45KPKNhlJS8NX2prjcYfian22ee4lL7T0KaN9g3oTiwgqqKCVfcMW8vFg9NUJ6fSVye15VyQvXCGkjuAXWArQ/RgOeiduGhbHEG5kWkD3c+ds1N20sPoYdhnQ1m6NM1JVgyjK+MM9mv9Ee5QBC+SB1exeWu9nzwfxORazZoUKfBZk4/FFByUv+5u1CA9Ccp1skewMwqcL28cFY5JOzrDFhl0/46zM7SiZ+DlC6q1ooDhJK4Pkv0H2glC1VerEDXWouP3BkMBFWdhNHTeI49odJbWJ5kAxsrC29ZKCrE/ZBAqPr5P3XcBJFuSfeHfo4I+6BsH1z0WNC9TffBdwUHW4jaM5YBvdqY0pNcUyMhQqouJO9EWr+owsnXYvOV6Vi2tVMlIV0ZiMkPGW0JN/K+PgIJqz8G0d5z6UfJu/Q0HM0T7ioSW2maIrBl3GZSz4ylpSwvcW1QA3ZHOFsuOtwROxQ/QPI/V30N7bcvSHCuYQ8JMU/JejRb779Tgc6ypJuyJugLVBISbyNg/nFzXBL4jqMr0AV9+Hp2f9nVb2yEIEBNB1p59GB0sLMT5M5iFhU4vQRe+l9OresBWrh9LKZ8NaLAFETRrrTp4/UNyiWGqK19Hcq/Ew8cSQ9mkUCohRUAdWhBA8LchZKOHCPIRU3RZ1ma2ymF2NAme/LKTamsA42H0b1nL5/OJe6GWNPRqgeS3R9C2acPD2L3sieH0pXaJH3Mr4uS9rEEyKPpBdIFUJrS0wqeuM/lT5qkNf/SzI7dnijAtMlMUmlOSodwQc37hwcowtILxg5lvH1NrdSdAShAdztEbCxu9XVWcJiW5B/f7olCHZBhrOyB4DwlH3WHWPeDcCi+QambEGf/ENt33Z1OefV8YSMRxFxE1Um34+cbvx7p+dwfUo8dzQs337+il4zXAorCjwPPPTEgAvqOqwCxwZTKudGbvK8CELpJSXSKCHEtx7cc9IjrndySjLHGZPBs8LcpNfrDE0LTpLJ57D45+nlmgZgxhkxjEw6p1BsqCGFT3hfzt/1Q54Kb2S2xRJ7dihoF3GcjU8g0Ef7k4xRBVK6H6E1bqb9JoHLJ4AN58Pu9AjS4ZkiJCbVq4tczg61yCaARPxrwQvLL+eEfwZNezeyvmGaiHk5dsFgRFsjKHWxlehEQFAeDL9tA+EoZ+KTFuF/7AGE0LLCxh8qi/J6LfLSamI9vQbyhOQFuLJNj6OS+qNi+k/Sl8gYf0NwE82xF9RwAe1iBh1IaqZ/Qku7NI+nNjQm/gQohQMRY4bHVJ/929Uu+QdrNerKli1l3f7FBpiQUowcQHAzkCqM6NQU643tI6tE7vi+Q16pUnSZfgoRwR0OeBGRVEOKP7lAWI2RB4mtA0jTQCypC4VQ1qsmNfINadOCcC15L6FNRvqPDgbc/hEoNPV9/O325ppv+yyNcBKWObk5WPglpPeRNVH0H+MtAlFn/a26LaU4uiQ5QSa664pTmoJNGdRdwLXG8lDnbDVuI2cjT9xjmEySe4buslfUSzcf44TqF9pr8an4WCJcSrXxmUoY+lqPNP6+InTmVXBXgXq321gieLE+NUQ15cY2d4kZy+lLRcShsvcCDlscsk11MjFwhTmxk+vtQMaw3O4JgrbL6M1+3jCs7qeSweGFOjSfoytevZJWAq8txI68NeiPtAxaTXzg9nT85jHzXPQx9xYBqKUvXNKbrptbLltR3tpPi1I0sez4ADYobjRla05fCCr4ncVa8zo/AO953F7U7Kq2zWElIvvf/U7HNWGCb9L4nrWHMmV0uPpPSG9noYdkTLAKmnbosHzC18uhgJHJmQqDv/BwJZbLWuyTXj7OOqbXgvjsWU1AdxP6HU4ZqCfqygBH7Z3lMVAusr0rBiSPjcIKLr0jxdlxMuDI4AdDcIeh/d+C/+7Z/p3t87YAw4NIAHTjEAUV39l+sYCucmNg3otvd3S6Kukr88LgHfSQetTAftgfT9UU0VwfBlQwqAyKoReBRhkFTvx194fcMvbDaQo5k1WGeI0onEpmvZSB461EqCHU2oWy73X9/1ptgdcFv2/LKUkE4SKXBuTMTkoOECPp4oYu66D1YSrcTxmI364k87YYdnPABTXcSb5S8rIRRdFlNuydsPUCU/hAEbkF9G0pImPAGg70HQ+N8M4Zd1SU2I11jcWFknLLAng+E9IjHfQnrCIZXeUP2tHiwa/QCHgrNzB/J10WYbGcE4FXeS9aUWHjnWgsVaSlHvgNuN5j9NjaDr8Fy0wfijV3CDU2Jd0o7smmBh0kEZIvB0UaukZ1X2PqxON2Ul2WcZFCORpdfvByupYye7noZIYTQFzf4X5IDu9RkWQNgO1jjgZ29ArDAdjZheFLjG4eeMOYOAN9ZC40rEDYcXHbm622/VvPIZzbaxUBWauriJXhBvhTfUfsvOsJe35dSUvkx3vsXhampvPP5yNrB/1xoy/RJziyLKX6nl4aejAihxsZvjVIAbzF1Xr1AJTfNVgUW/2IVcOD+dYYRqJpjyc5aOArUSd4oDjoWt4ENe+sjPDvuKCLoNVfroQlXHo0c+J3VhN8qUam0UOouJq79o0ZTKIszrt2Bf8qle+1DHo4BIJrWJ9/YzwBmy2O0dS0gu1Q5WbyoWZ6cOaESLzrqPy2Y8x0tUMhPiBPXTNred1/1jMyJ0GINs81pocbSoUU0oW6na+Q9S+hgnSOe6wRy6OLI9B1Welsj4W+BmWiS2fN2IOVnbibo/VqU5KH7fh8V1yTTNZb042QRaPxKfzwF7yptrt0jZZtcv/2TatK4secY3PHzwSeF+nZTNCsxAC/nLVDBQuMnnb/8Sn6oj5/4suGFWg03vYzTvp7drvsZvwe0FF/+0piPpe+EaxzULKZV/+oT491fAtzshfiRwKGhyv99apTYjtxT9OC/D/Es/YiSI9dyLyUUKadrc/xxEdrOUA/RXuV+MSI6JqDbjDaQO4UHjYRTdWCs9eeL4MkibNCVRgBhwaDXYhIByowqxporwXg+Jvupf68fV0lAVRMcT7uU8VTv+/si6QmosHBrDc1Q2t7Nkt1r72QCIRrmVIai73P/O1s8yt8G5iLPlBIXCGm3UbL/d8qQJmah91K+V148wHonEtsnz8/2nC0jm/7ByIVCBK2jJRZkGPis2rFpeJd+6YobYhmfDsVeQIrqx76oGfwcX2RrnkgX+cOHsqjL7AE1SkYOuKdBVqupIApcB0F3vtlOAxnLM3GjTZiTK4Uyqq4zNrRQZohj6RTBqfTWyqVXuuBMI4FM0NNy3CvHkLY0VVwfApt6WJy+kVdcTkKpNlVgLyD/TdTeFC5QF8QjGWGbVv4nZus9aQdnHmJvz4U1IDexqh0mbDXIo40gT5gBhkzYzSzHhXQ1lXS0sp0eWiR6Ag5LCt+2MnTpz/nB1LBWlzZ7HMHVZqUq/lMWOzVhup7REsCvyTXmJnxecvs4h8eXGKnlqYZJ/ujZFREb+HKAhZBhKMReRCm0c/KKzg6S31eOwNt7D9+41X8SGWeMN5i2J0WpZB6hd4I4eVrMp6XBAXVtbGiAR4XrRMbPoj91DhhpaQyfvo6j2FxxCKSnX9m722+T1OB1xHwzNpmqO7KXRkhuT6UdKewWao5s2wFeC5O5qtghunucyTZHzK3bj2nBePhNY0Frm9MAzk6F895X7eZa7SOeeuIcUS5H6NkrKEXb1q00Ih54HD55XWyT5yvpq3AAY20oJ4K+2FiofZAxURxP2B38qvZTFGM200tN9OcdP9hNN0IaLIwjxzrty83goCfWycSOUGOBxpructJO4Ae8FOJSWH8wueuU8ZMiZqhVezlWQsOPQSwfM/TvFWRMIUbhnUmyyjfaHqnBp3ACQiLX9sHbPD3+cD24tDgMhoKsF11+1bgTs0YMSZfiiM8gkIymKhSGF5RKWfptRQWjO9lBHQFR6sxwuidTNnmKC+Pt9oRLAHWmA4OVD4kMovUXW8/JLwOg9MlwdQo4vvznqe0otd8Pex4E8nb2A2BujLd7Ay1qxtV6FMVb8+ssskzWbwGfp5KmUZgy5+SA3xaB014Ne1KMKTAyjl2fIg3Q/ROmrQasz5/1fSQj/Q8pNr1lF+QuWf/n9ymX7rVRklkv3xtLCX2f6h8NbXXzOdwe75tXOoULMGz4VRLdj5MrcAiwazuMfgQSq0cDl50cdcQv1xmVZ/4i1eEwFiirPvjwf+ixYvCqMCsyXfHmBvGCKDtLX5M3dSdemyzyA0FzfBpq1HdYFBIt0+HnT4phBYrkSdBteRs9uFC6mXCFq7PWRNNAucWMndg9t0rZejTvnN9XZ6MHKiFMboqO6KGZacUzf44RLhZGuE6SmiDI1fkKDHI1Xtdzvk37yMPvLPF5XUhH7syKzxb1fRHIWe6seu8JJgpRsTfziIMYW0pyhKGEVQSepTAEWLgFDe3zspbxKUsTFjzHEpb11wQ6Hm4gqJUgtdVk/HHl5Dr6k4xr3ow/V1t1ujQpEaPnlyaPO1FBCqj+MJT/lsfqQ4vQKdKe9FYkcZEyPHVHr/gMdERmnaPf4OA7xNSfgFNRPkxgav0UbLEjZtpJYanmA3LB7kD88kIHXQHrLVHAWCFQ46axEwULnYV6qW1/fE6PlS7E7ODMnWGvvnvnBJuz54bqiKlu/nvwJ9AbFZsHr0ZMGrvZnP502hcvGiBFsbCd5gWg0M1jpK1FMp3cPWVlnqU+OivU7+gVEjVZ3wg2TeFrGqh1/hP/HysuMm8jUpMmMPmAIfR1SdvDlV5Bha6pENNYbCbNfL3kb4FZMJ4NhfzTWNMeuvtwZ+XuwesQ+AVTg7/t+xbGso7nDbqmx5Q9qOhKSI+k56IgaTsr9tO47t6lNT89ZlHXmBHtQG2l2zaAt9OTjaN7E0nEDGcw66gLx+uBtm9/M5cPc9uHG7hlyGFEeTsgT7h3WHSmeh895aFpdHI5lQ4tpPe8zCm1qzJbdJpmENm5itjTEq2uor0NMvGDVSw9FmwA8qoesxEuwa/Hhjw/bnOIfR4AmHCX++XYHQ70tpyoH8sYsuzO7CeQSLZ5iZtfjIJWn0hhY1Ix8ornMb1bj+LI8wU2I5XAOXFSeTcKdz2S2bvg1wKiAu9RqVW+N+1qejW8PrEZkeMEfDAEBVT7P5G+drECObhLBeH8Kw2Qt3BzObHQ/0+G3LRiuI02XorvadOOS9GO3xSVntIp3oyonSIfDbkN4QZZhm8Bypcemm3jt8eSbnykPLtJJcVOE/EUTJjqyHpFItNQiCwpDtce73S7ch72CSK42bPbe2BJW+mCCJ8a5NhdJAI3fH92bJfLWMG7F2ko05u7QQFxvy7qJFo/xoZi4wibjJIFnrCHQU7GxgzESPXuExgpwLCTfw01muaCzEl1Wqo7QdOWvAqRbU6dp57rUxSQn+L+0wIEVCvjRgJOie1KuyDu7NLbFeAocupzJsF5KjroCvCNBN4U8GM42H+krSEVnhzt1fHq7FQGbUSYu2d8KwdJ6xdMlxroDRa5TxM7DisxkMLiXYBLYtzncjvuq97Nq/w2MMDMNm0xrYaQZMLPIaNMweUhsMM4jqQBzGujVG4P9h58NOQ2X0OIEL+MNwj30/9Iu/h81Fah8qR8v7X3AIJRveANQ001UmyB7EOG7gPaeHBUtfuEIms3gKV7CrNHdiKoTLc2mHLHZp95etG+K5fw52HwZX3W8fn3QgdkkN9LSxGY56IGlgd3ZR4QnkOYuQGJPI2VfqfqhMzo6R8pHpwGpv2+x4B6lI69PEykAzDKhEOMyaLzBGnKfYCM8WqNXVDxI2NG6Z0Sc1yNiUmFbw8ypkLleaMqywGLiPN1aaoa6ZRFDlVTmQgCmFW27HQB+7Gx9pwqRacy8wUltzxtZqCCYUf7xIShxkoThxJwDPQD8MPCdZT7ntWamBFgQ+y+BoZaOsrwmdpJ2Pjqg43uWSobrZwyU9+5C8Gb32tNRvEIdhmQUGBcO1/wN3gQZidWQ63jdsrL8Gm79wqkiMnC0gj9U3WFaFSlBhJAhn90g4DMUcZnrrcXBJwiwemJFOVkUFCKJtsfsOhRqCfNkoA75f8+6L2Ldl5BioIL0zBufAFnZTrazLtBioLRmJpQoght6mEgLMsGQ26epkscu9dsyZZF0lepobjI9zz48l8VTZwTLQvlkLaLasM1nx5H5lIVhJVdS+joeByNNin1H82JRPE9jCjfTd5d6BDAOpiqkBvTc/cfP5u7PJN7l/CjsxoKtb93bU7rMnbneNAV58Gd0DIChTsm6GuMDP+yDxz+Z8ZF0DDCobY9eybwZZEOj0LYcDod63gp1Z6RXpgQqudhixtqpLCQNIr3yr/Cj7PpJlUykUuAvd//0nKerClybJAdCh3pCQMcn886noNN6Pkk3OpjB2wehHyT3HLrApDeX0OiFxNf0INUrka14umNHcsrc/KNdrya9LV1wApSXQG5hyyLg/+Hgab0SU0xoSiGi0+O0fz3iui6iXsdVBm2bnja0WTCKRQH/fYCkN5FSoCgdFSczvQfxU8nyUcnm9cvf/scdQuotH6dHf6Tf68+Mk3sARci/f39YIFz/YdQNNMN1M9IEDplSAFOTfh3yfHWhr0LSOPNfbWIK+Ii2HZJY1MPIyPjRcrlr2RWK5lchz4MRtINSCF95STLlnumOpOgDccR/RphHhr7Ej8rO4ko3N9g3xNoM6wtaXpWhZyFXakS1eIJRmfGKtg9q3DPp0yCG2608tc1PhulMr4fr2qbWbjVGE8JVxMw47+GjMLx6UkJkDozQGFKmOZ/uK4sQEXrRcTbbHep3wc63J3XVAhRTKet3EhekSWmhbSc20DDofZgRgIqP/Qw6ywsZby3W077HfAPyCw3++iSRKBZzkKuggmsWifdBd1p7Xxkcwpit+7J1oH82J5zen3m+ZvOaffcL9yb8grRWvqMJE4lYhiYWpGb65jYPb/m3LgM8GAFT9HaCLhl1gqDfosjxqP1doc+UmoA5NnWRmwi2+8w/6ktEVfIrrFSdzF+BTuaxwtqQYdm+MXU0QJ1/JW3PEToxYKatYqDQgPbV6tTMNLiC4IRTJP5/Jra9BU1kNgxCs4B0Wx2Vs+WQ2F5FozeQa4hF/g67Wmt7/rXmdUOo2WdqWt3+j7Z00IY=
`pragma protect end_data_block
`pragma protect digest_block
e0ae31d3785a50fd96cdf2f50ad9e15b0da6f423caaa6c78dc4d076ea819aec3
`pragma protect end_digest_block
`pragma protect end_protected
