`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
Vo9WwmOI8B2ifBxuAKuvATzsIXcoExogIwfjVSd4uuOdfRT3XmWU3gxAwe+0eTfCMACJb4f9fzLzkf2t7nAM7x8lXcbhwnILSIeleZeyEnF3Wgu6hEVph6JsBmJ96HQDHQ/1Ad0wfKiqwf6Lk47+gASoH7rW0lcjT7owOEQUp5IRCtBa1F0gvbt9XpRyiQCEe5mMg7QLPLtRl+GmGgK2CbHrLRXPWUR3EGUymJ/Y7m0ExcELQS7yqr7HtZG0LlqIX7IhHYkgZaVxN6OnBwI8vZORwvb86ie58ALw/L/wfYbDSyEsKTgs5k6KMl/uNHiyK24D3raky+Z0iek2g2ZMhBkRaujF4DbefFzUm+eFiPsHRuA6h5oXdZ5HloEexqIrFSEirgRGKtpd7uQVV+0IBbnHRo/VgxA+WU1HKHtsjvPFqkm2u1k1Ks7Cbf7gJG7R2veU8KFW8oMt9el1NQdImFeukiZI7O5IdF0BYX/Ta/xuUbWDN+W6gb8gtp4mHFqa1GeqcYWXQaPKt2hcoo37/tcN4rEKAcqfreDy7RKa7XnERKGpLE0UVF0Hyh7Oh0Im8gJ/0+Q5HNb8DHMj6Pdhyl998D5xl2MWTtLU0wVFiZJ7zoiHrGyaA+3oJzeHUPkAjrZJCfXQoDbxh3dq5PLacyonre7L9P8DmG1WTu1vGV2HbTdtjOw8OFEqP0tEY8kgSv/SfEfItVd/7A0ccU0sxgVviaIJjJ25x3mMxYvkuIuxwNwU8Y0Hl9aDTq1mE8TupJ1wUA2d/ifvfWcsSalSq5clGxQedDynsZZKSQ5R3hJdAgZAQEtaxYQcuyKcgttHWbefHESoG1NYF/7BW5vuHk9nvZB3kScCePEYlJpoKy8/8+91FcJQLIsm16bYq4IG0c8J32YWtUSSfnUe/q4NivlL0wkBJ4ICQHRruteDg0qa/a8W7jtdEmfHMLnWSE3Z4dCq28f0vUX+3njXCBLTKVEtJ3L/xaZuuaEoKwyCXElDeEMnEsEBubhS1NAx2m9jAYzGVAqTJP/7zPTuJ6wH2Bm1JOmY3W+0LsdtBZ4q7ToB3ce2E4YOmbKXMxI+Mt3fo2iJz0YlTMXyV+Zxapx+fmFh2efi85vHLJEjQkRgso+0kqBndGPcHefyaaWHc3cwbhPDEHv1WXhC2OmPZgFLaCtfCWNWnJw6Ahn5LjNylB8TywgILPZmrpJykhm3Sxb1qjqDAkhSzDT7gCFvmmyLn7eXban/lwFxXPeVc4lMIf7yki3fv21ie/DZ8Jspq2HnmOO9YZ9Lq75YASSnP5fXiOHkge/8nyc9F4PRJCnJcSc5Rj5m8ZvG2RfFWpqJNQKjPxDzDNAEcz6OmJPL1WpDfeBiPOvNySbdi+xRpj1ohlqqJ9DeubCSMUwq7WBS9c31VcR066jwdTX6cBMrT9Ndsum5636PKV3vkiN50vsMzuYDXkvwoS+iIBf7VkZ8xh6qJdpM8Ks43B4nquJOWkS2ah+45k0hdP/ZOwAtbMPjssxoSJhmJSNrLyb+sAmXO49vPe+JecuRhsXcGolZO4U7AuoA6PDDjYJqrz9kA0eCnudKH6QnmATEBvNwYjs7NDZ0K8L+aVl7yQrmsxpKIaXDXsoHZWARDi/0VtjhKWBHVrPt7+6olaNdiEe9AAyXXeEIaFnBCyYkqONmATyRj1JYh55SZROpe6viUNN8YID6qt6nGCs3h77RDzSl4Tm76ZPYEO8yBH4CDDi1NmNG1oY6hNleg9OSU3VoDzkKOE+eGcF3ec6k/KT+h7ZnGMpxsaDiBL1VF+8QaThKL5yoM12AZhSa701axrB49mNbJjOGFGsV+GXL7qSDZRf0FtKlHItN6mODbdy0FsFewIErVwrOnTFNgvGcScCV4KaAC1mDNq8rYr1mGJdudHigd7nxs2vLWKo9HyJSGkIWBJWYumhqDs7Uix/llCeEpBRbn3hKKRjg9FFEwSDdLWbQbtle6qlZAx80X0TjLrDD8am0xfbz/V1iZeZWyLIIiz5KcqMjW5/dDySTAcAPco2rZcLGmusGR+GSY9+euKjvaTRI2CkfRPkPD/57DIRu/G5FrFu+De283RXq4R8KMDEzHfORp/z8QCr41LgZd/uh6sOpj5TQGTU+ui/H54yW0dIXPFwfZ/8ldbih6LkNrLnoZKVquIpdQF82E16J9iPqCDyy7KBIA6Afx13Ywmo44JZ7ya+hJg49d8a2SqhvXmYrxNf5ETT1uqeWCz0cGK9Mlm7blEa1yIjchroC0ELhq63pYt81zteNBcSWoRt3AD1xg1F74O4k7o6ktFYnfg8T7miS8XLZWZHqZjkIQBLN6vyxAo+LnMDMd76VjZHZFJkJH0F/MKhqsU0MyospTwcDg+ZvKXehwYTclR2VhGMsNBiM0hBWJ295o6px8WJId78qMhJanRXtBrc6calkf1Jbiw80Ldh7i2t2hksDNVl4h78NPWiE87AMbF7lcIMCXpCV5/PPVgWgzIHUuI5gJVI+OWL8USta05ygb4+AcUosBrSjCmD75rop3SfsVCETPJm71g6cJPpx2IhVgFeC78AKMNG9wbx/sO2UI4tXVaa71UuHLFEtDam2lzey/oaupAD3RgmnztNZFTZvZzlJBKb2GZX+8LW5KdD+E2SOE/ij3cSj9Njdu3vYOG/phZHjm7nDzVViR+fyAbhInDk7JU/NdFqLQWy6UEwmDCOySM/WooSLuClyBED7eM5KppJqDZ4XXJGHJHOnNAf19+yUSQmZfXcVTPfnzB9Ji+2r+Z2aD8F5POV+L60QdIjrWIJgiwKXQAiJaMWnRXDaW9l+t08xEuSTXJBfNtnJGJvrxx3dso1slPYxJMrqVtULiL/apclYM0XMVke0q+4oUf6cTmbdaYZUvH1ePrzqcMyYobttFsbX6VIukiuX6vkdTGtQ+1a0V0nVvao7lbkAyBOLLp+2j2vEbxOQFDOJqDJRXtu0cM6w38Yl7qdvPgNDADTtcYDH1yIb/r9a6rsNy93xh/Jy6Y+xZf/Yb14EzPmzcEX77U0pHDTB6dfTsi//99rdKjNOG3YCFdqGK3WUQe6H4jDELe+70TfSByVVhAkBB5kwS9XsRc+989FqAXtqOaWJz+wst30Tp9+kOjkapaSe5XAIhH++gkiAgOnY2kaDwr6/qVFH+ijgmnjy62Mq66VHRUkiyfSlNC3Q5meIX7lGzETr+D1VjpuEV603au5vp+oP3KxVbFNIz9RnXH9FfPqkuM34shsVvZyb/qBPmHnEhkKaS6FBE9VCWddAS7aVyG2VdjvXfrXwqaZ2ZVaIKXHqnKcq5wwWOaE0QCH2NamgjH8uo/CDE1HGdgfCgKc/B7kKH5CrzTtb8/NZxa5XwWb1TZRN4Rqf20uWhZLUrX3Y0+KqJrepcvx6fxB7zeFArr/LzzCIQlbyRz2vyuxwv8XcixafBCE1hSB2bMpNi3aN6jcnz7hr0PIfcNi9U7Jr5/CM4mypk/25OozJ4jwy8YA34ZaNUzSWnYkhq4mdfik9l/tNmrEVFeg9NtQnefvOxK+0iqicv7VbW8dwKTr9wJvUoUBp0uNO9vZaDJvuRTeRDoYuxNDTfQQwqZByFcP7yFWPcF+TG+k1OKyX9OGL3pjx2GyqzIyTKneXIyHDny/9srrX2vPChAE5pV5G31UfPBt1xOu2soMVVpIXKIpROlVGlTs+0tTTRP3nChbBuyFfCZOLqVGBi4DjljCUTCsLDNkp1c7VGdk62rLDKkCDQOS/6eu3B1geR9xX14TC8bO5JM40qYOQQLVZWdSgZNlkZzhv7rnFpUPgxJkCzbCPCTNCtRF0FcuI3Y7hmtEIbF61PDLeVsTX7ZkQ7Hbywok0nmaHvvpRVrbltn+QECjukm9Puza2gIP9YlwY93cJ711S/bZV9/k0zgmLtJedlYkO55nLtq3RJyE1vSCp+8ef1ZeFvv2czYTQ3vPWWkbXVWDL1QzKiEU7tHQW+ulOSUhrdonxDFiTwy2M41FQXqih0a7m9QDNEuVQxdOwXbWpcgFI8lPH9j+V4mS6pKPJCNcpzpEzKQRj2gvOYHwTE7OPkcREkAp+UbF+Cp2WCI9L4n9wxTJhsQQXTZ//urxiPk5FFFGtXmWVtyyeieniveWNvm0TTI0W8Grru3rzfvWYeBvKyZTrFzOVzx/MiBofrCttj+TRAUDdTW88J/42QvBuRRvl9M2gswT54gY8TgMfj7Hd+qT+LdXxfdgSlmJ++GLwTocKvhaPKWjAZSa5e294xcWvVXIBtdm4RMtGYTuideXCOKlyp44kRFfUfz+NtbcCwmN/TrqagptX81LF5kvrtPvjsBqHqS1zszMoRgkZe7iAiBn2BhXslijhPhKyvfnTDeV22JNtKVd9gwLJknisSGzcRNlYGCGzKlITkB1eFrwCRnD+Es89WTizuIt+SN8+0ehCMsmGKb07K/3Z+bxWYMcUIjWIgN8lLElZO6Oti4IY4sLMrL0XHDLQz0mOTGPlzjria1lPA/WYz5q50Tdn0QK76jDtV4AN++0kebIi1Rl2WkTUnAZdRSJ5fE46YXGeyRXNtHgjf2CxnvstI4AHPZ5ybz+Dlavc0obk6IDO11DUo+G9LAHDd5UF9BQsm2Nyc5Ly34LN3UPQIlJAo60HS5mKagj1VphOR8fboZMA5+U4sXg6basF/LhIJJZSBfkAdKD/b1S7H5NhQIw4210OVsH1Fb/7Vmgw7/4kolxvk1zFFDdy3Q1alIFlbkbZJSDhoy+09MD24Ei2I8QTyenT5PVewpu9Yr7cu6fnHBoa4atxXzr0XT1CrrBuN3IKkYnnxWvW+e8HpwXOrZHXrlZIyLhMv9Se7oGnK3amzlQmfVxboWra8hZf8JCupCcfhoqoTFZfk6ZjJtONrhcJaq4Lw1bpdXllBjN3j4+zK7OpjgK7NyHh7JzXK3TBSJGezYMHY6PzAZYm+BBNKGLbE3ztNm+PZX6txno3tiGaGoggd+inE1nVWUMW0a1QsYt0VzFRCNBiPRqYtK61Zrv/DNYyvDt1XWwcnuYsOvzF6CdIft+ooOVPlCVx8avywiAYfHtJUJLysOMlx6KKsz7bXuuA3W3JCNL7aMypt8Y+pe7S4QI0/MkbUexYOzpJrokbz7uJaHgk5uHlyUcrcvhsRbIKcGMlX+b0QhzCu9+JRyEx3OiuTlA8hhVghNHgK9rP7e2QtBDq2AHWDfO15KXNIKPMJHBMs4dCO8X4HkTs75m6HUi5vjZS2RW8TyfaUNp4DSHqX99eoJcNQ+UciuApciwuvtfjPJVpUDEmyhEhePYu87qpZgEctzF92PocSqBoPmGwIj3433ZqMk2IYTYo2rjv39GMa6RI47cbBAnIjBQnCfYgiLZiumISyh296knd+bPvtchJ/FsUddZADM0NI+D2SzYHMp6u3YMgDCqSbmVH7SXrYSfNCkIleRhDFPniKQ+8oX2l00E2X0zmAK5ByAN2JlOTevp3pEoOSusZ43yp19OHVM+5CEVOcSBz3Wbhyi1ZLcVI3CJjCsgF9Ru9EjFNvp6GqtBMuLNwdMwbdz3JtkTHJYkRVilD+4WaejXkOwnPzQ4AptF+VNq3f0JCVIJ2Bed67JRtgqw2P/zjgAbPwfKaMeLxBjF3sx0DMHTTT21HsZU7aVa4rF+wGQYj3jNKP3uDdTpdhs1PK3Yxu19GoJcxPl0BqV0DxnZ+RA+OkKYyjUNRMS7KaGVaUiLFdStM5Yhg6/sFDD0SjIcEA+gRTgvkR/X+Z9ngQavmrsfA5Vga9EKnaOEz3ci2TjrZgC6oJLzAg/OGkNOLOYk9jH9fO0viGtBdiK92X5W8no1hsogC7NlDdBkKqdzCDqFdUSzxtsR43438xssmqrrECrhjMJATCfEMYkFscGNfgVf6yd2lcgTvDUgUTzgLy0h6Jrv/EU5LWkpJ3thVXE/3HkmOCVUZPF4Or9G9QBdkhFx6vn9tu/A5E0t1EJjdCYW30pqJAo+OJj3BgdvdUhjCw24Rdhw2fmoXUOlBP12smKVb3/ESR+2FUtGXvHIBBnIx2JaWYNyf75HkHaX2XSO6iuAb+M/3zV7EYlo+R0LSYdjm1rZdV6AIaLIzzWXx3Jhw9l4OBwi0L/oR+/6OBp3BTzzKmCfoXl2v9odejEasrf++NjW1LpVjh9+Zm7UrabJIKQxJ1AILEkcBEZrC3n1X/bw5of/KuBZUsd3nQUqpHzL5exEYshzjqLH3e8IrZqXuZU5LXFmvgK2ibF9+Ds06hIzfQMiOTZPC6k6MM/SXYv0uwxYtx1mN90okAsRD9S85Cv5FSInrOxSetvyjXWQbcBXMwuO3/HFX3WSOfh03kchT8D+2YmxySeSG/6GRdA+KXhYDN701p+Y8+0UOtGk+Qd/0bFtONsM/KUUGbeNv5Wp1O13F307utGYWzzTf05ln4qLMj5FNHsCo95+Mhg5vOqWmClxHs2DVeqEyv7aWNZlfZwMlruu/vqwEGfwmT2CI0nY5lS5HgEScrzpIGMR7hbs8l6AWEwbyRDKs644idONmbfAMLiG5EhSXQcOkTwd3LGifziem4RU/Te2QCmKRDaWExrXOvXAt8CGyuQgIqNIkiKAiYPzGhbwGGHYJugK9b/QmClRV74I/iKLmNLufzsQ0O4b3eUEv9vVEF8IuNimIq1LOZwTYPaRknix7ChJCHzu/y4o8Ht7nGv01Qs1RvkiylfNYO9E1ApFTqbvYUw==
`pragma protect end_data_block
`pragma protect digest_block
a74fd60148becc28e48b5d342b7752ead9a1fcf606f8fe1a192d2f66b4b71703
`pragma protect end_digest_block
`pragma protect end_protected
