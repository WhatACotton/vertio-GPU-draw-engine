`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
MYHcJ1+1tzeukL2dvSE9Uz4QYLoY0jA14qK1dHgLS+lWbv2Sa14T5n7VnZI+7GGc+b3JV/bN4Ly353IUKq7inu0Fs0xXA2UjfKmaLpCKKW4lvrh+TexagWnrVXTGtFAFRHYgWr6OJ43/+oxYksrU9f5v3XQ7cd+9Tj1QDeCj9fCe/1CEw/sru5+xQkLgXVuyuJEJ68tdEpcQo7UhXrWtdAyXZ8foaEJ0aPZG3iYs6RsAe2hIY8drjv0GU2erxOBAKlqRwstkaJpc8gzQJKNlCrfrOxWFdWC96xKTBIDwgDGmpgA1BnUn2TK4USiMtsV4vOz46/gi5A8H7r8XnHyJKbjSjoVKez//zKnkdfAvDBtmQcbgEZSGvVohISBaF5YDK6aMM+vvxy+c9wb8BSq1k3RpVQby4l734wEWyN0BSKjcuVjvqEjnicOaCQ18hn/hWxtbAEnVOD9X+WMszMX5zXDfT7J9zcRzxN2y2AlvXO2NizoZIpi8QV1zKyB5+gWypFU2O7bkCqfildyLWUABTb4eC2LGUje4rXphv3R8haQTGJbJy5jfLNV4eQpsL2lf9SIO4GzUhnvvTBG8mXImwy+NwwHN/zrgel/ibHg7Ep3AADI3sDhyGnyFaJBpRYowqnHF0QGa1DCgTFkBWHMejYWE49JyimG8yWa/Jq+dL7OzkmSee8/M3eKE0oE0CGi2RWyVmWyZXYdeQ12yv3KP2rRC2PDXHlRJLF8kbI89Ag4S7ihqaGVFaNXPSprcEaKx3o2Qzgrc/EE8jBuAq0LcQnxdQ6Dknl9+K6ttOOqPJvenMpMQNi/HCZ1U7JOujpGcn/dhTsvL696vIdqRiJ6lVMEIpY21Oe4U/Xx2mKOOPFvniJ5tx/hr80HXr6R9muigcMlGE4SSIjLnGn4Abl1beCpCaWdtkq1ER6XoKvQ5Yh0oTYpFiV4m8UnUQaY92Tnua5h2PEZNOYsG4x1JBvm34TQ3G7YkEVpnKwge1j876GG1AxSMz2wFYFSuHal8ULZ7W8fGtiSKD4U3IwMrbKcJeM8d7fyOh7NDOqzzUrArYdEfDDNZR2RywdLzXffID45a3VM7aqO3DVCYiDQ3OpKrAjQsGVXv+m1JHQF5XMhs7QYVaoWKoRbnhzmUjmrsouWeY68FH2n4u6ou6G2CC8/Rd3Boq1uDxyLNw2orA6jwB12ZJybtUJABCo6fjEuIvyvTz14NaIhlDJM5iIvsZilRDePISrSctHCPz42IWYU3C6DhMiixiBry52RPQgW2sTJ+ABixBM3aXtuxncANJwa+TDjwqqObGIBqR991JTCqDuuouK+CkN82HusOydywvvd3KbaXkkCVZX5qn5+4Wyuy98NGvLIzJAHsWkiDNaGR1pQC7GyNii1u2om0iCpwDOJOKiNaJto8KGcJsACg0cjAVy5olsq/zr4zWp8NdQzOapB1vQvMAOg8g/csAgriqNUA0x1NiFxiw8Lkfrysd5tavvYsej/G2kaNrrbTqseAM9FGRLTM2/0NUoXUwRKdYq+DuRMVSgdfr2u0N8PjtpL9M/d7Bo/I0ZomGqYAAs44AVZX0AiDMv7qgITrLdsnEE4NWbiZKv4FftODDOly03ENlesptcvySpXJrOQcEL5f/0BsN0b7rGlZqUDfsqBAJJkzRftoifUBan7jEh7KqmVRq5n4vuXIb5b6oiRGZFW9cTOWu+DxdgLz0jCDg0pmmPZEJzVSTHTm3RxodBH4+AbTHUwXBYsLodV2mKMlV6ZxEHN6RDWlmrVpcEoaLUghfutzNSotO2vqJwiYZZeUNwlHYg==
`pragma protect end_data_block
`pragma protect digest_block
a232b6bf0fc0ba18b3e73ebe0d08835a446d77af7995cf072a3b2a6aaa957cb4
`pragma protect end_digest_block
`pragma protect end_protected
