`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
GJXHwXv8kQ0oTyTddgGq2cQMpZ1Pc4/EKDWWZuEvBLg1gl/Ln0IYOOLeQmy4EFS+EGLs2J+s/oJJc34Ivr1eP7eSgns/zJPwwfzZMKmas7gt/C5EeySFItBEc92ER+9WjpwjTG8QkUCevUmV3CDStIioxSZ/OLDLTA4BKdzkdzTX5sqbll0Fn9gAqoob0DnAWOHjBuF70EFrZvNzIeKqGsr7pkklmhwvaq1a2ckuBPrz7FsjDN7GumSb7b8aIG7M4CtczFvaEz6Tt5iCD6/yX7tBFof/sfFaDKyoF8mf0izu4NDaA+7+khA+q6B2XjgDk5yWpynCCgq398OoM+k2CTk3/ZX2jK5d7Mx9iIjH17JE0Z9Dye1OsxVGTiZvIcdzLVAnbJElkfFQ9H8yGtgIsC0eeniD2KUgc/TgiKTx9eQYAjOZ9lU+GDwGUsi84KH22eL+09xnp6FrlcnZ2PWTb6uVAmzm/fQOluAMCct6nt4fiUgAxeAdwZpNQsfQnemWL8afy+NDgR8qgqFbjvTnf/ipVALCI5AMp3khyo3R1DuVibW7rCWP/Bd64YRIXUlQYsK2GG2I4lK9/MX/bLX9qz2XrWJHWZ5kswTBJ2ZzqXwU50/XSqMBvehmpqlGSDiWITDjiLNYdzTihwzikOwd3O44q4QXVfCf5d9bWzV9DSZWkGOlulxa9+qPbwC7eeOrlheZC+f/JrnRcDClb7+VhK2IEK3NpHv++9zZhnEA99zXASGM9KAWB9S1WLTGhRseBCsijnhAzuaBB5YXGlApgrJEEnsaipOrHBNiRCslrglYAQp0FH3vmR17dD3bquLxHaLCrzQsvmD4mkkWTEtkcPyZMVLIoHkBgvOZ3vYAByNxGoXdNuilqg4uf4VLuDe6b7k/JIS5GDP5G+O0feoq6FoeUBbbMwBKmL+F0Ww5tFTiKKoiO7eMuidjuvJ2GTom6KkPpsWymaKMxdZrQSZ5Tb8N0vkrLhF2TcfmwiQ2w+v8E6SHNVlUE1Z0jbFL57yRVWLACTDzWPl/ZabsO72Gqw3911H1e3RAMMKXlPoL9UF16jsNTwaL2sdgYoZfTIm3vNmI+0DdCJbG30hH8AHu5CNlRV9pMd6Z8vn59D9pxJqOatIbejo37iC6KgJZqLn/ynryfSmSfcIJ9nKhExmxguaheY3pOi6vtLNlrbR4gyG/TFGRoMqK5V8L9IrLBUwIZKM924sdBmQynMkolUFRhDJ/EgsfIP3iR31hOwxGFpn4qWKc1eymfC9nLL6jmOXkX+Fs7ANoZvX2UI01U2pnSmX1yzsHWa9l9LsPcEfpFMfFdzNz7O1+ytfVqDDvbosQTuT27/hAzeY6/S75JuZjmgZRc6FeCYBq/bJP3f6OUwf7++gmgeVk6gn5Ppg+7GNkcKy3+uAkuL4qGF6J9l8FcABCuYtVdXysOvfC1kPAKqV8EmfzIwuD0RNrN0TG6MeUFzwUctnkKikXGycTrMFymMS1O0ZK9uybUTvec3V2gIs2NBAXD+oFTiZQztM6U0nZIi1vdu6hed5Z5NQ7gdTloK5DixQl6/tIhe8wJY+IZO+dcNqnRBI430JThSgNuy1rdZol+utqy7wDSIq3vr+K0FXE8tt8BdOhb/GCp4O20ZyO/r/NK48hLTGIi+cPZWRxH7yF6xNGvo8myFSMZhV4VF73ZqOFSMHEvtY0SJCuyLx6iUkYSYeEmD6jV4jONzL/Qb3Smy/7gphh0shAPOtqu6IA+8oYO+RKeePNH8cyjk7VZ6pdKSOu1pllKl0ez03ZjH9T6hhIQCBPxK+3qtNylaBR5FvLydzz5HRQRCERNn1ooqPsiEpOOzYFeEDSd5Yyqx70epfLpfFMPWFoSqxolCwJ8r3vp1ymmm3Nimp+T2sCeQ7eYutiaVZPKVZYUdR9H0jhxC6ownkBqu0c1vPouXcx4YGXfBy8GmGKWib9PXXseVF2rtHdCO7Qsb5HhELRMTyjIulx3jm5de6ISHL8mdC1tPIjws6dSyCyHX0IfrTEjHI6Tx9gStSS9QFQTKe5b1/agEar8ShU1SaKlTiIVrLn8hpW+PvtiYNGC2lXhr/awCArjLcd5bbrtB+xCwB2B+jFTEyoipiiBfccPmRpsohi/aN5gqtuSD11Ma6lrAr7FGNdHAyL7HSD0XWx4wuaBlxwkc+ga/sOmuJAzsydFAFHL2Lqu0CmfsVC437euFzub30zWsAWEjBGPn0S1Fh4hKLBvuxsgd6jLrL6PR+wD+PKyU3KRduwiOCqjodxKVRIkHBykZTlUgCdMALo7zJysxm+gcJi174CF0E5SCd3GtkIJdBOCe6vh215iBbso2/IvWAwjEcWOsvMMJt5f69Bd89jJuT+ayP2LqNSBHhTyr0Rayx5HI2Mh+c3x+27yFENubR4WK1jJm8NB7gWoUWnAQR2EY9o0WpEVjNqXzTl3NtNt7WWxFI7nM/t+TwriGR+B0k4WB2WE6MMHA5ShNmBeCSyqmP7tFWAAGjGsUdNA+FBP7e1228rwro0MNbqhg5QMxY0Hwdu+bdg+lbjH+p3FQqmvyhoxq65uBaoTd44za3+kMKftHmeo/spUsxowXnkTrWe/C7HKZvynV3XqDfLaT676JBN49n5hwjri/UerwVsqvtrrT556hoBqCPBgavGbxM+vci5EI9COCwIE+QwKKJ/u4573TaZRb8B763huwLvTiiIool1rYmfgv/fjQajtem0HczSBU/o50V49SwRN8MVP+iZgMcc39VXZROWQQ5IcL1WTRiER7/hvwW0CNQgPWNgPVqbB9almgp2MCsESqvCfDOKX2DdXPBEpQU4tgusLyc/u5p+m44Hyp3lRt8dlO2zyOz25GcoKZEHuU+T5j704m/BjjdeAB59ko9fR/RS0qxcsMZnlK4cDCIqDAEhV6CAUZYA/YsSJkyWJFBqEA7pWj1X7NDFf9Qzbiixjb2b9Kln/745D+UPNo53TBQMZx9Uz0T0ZpJzH0eTOme+wxgNod2wUqOUsgdD82swNGLJBOeevZcuXu1GHpyv7J9ngd9DF3ZnuKAD03GjFpfBTNC7sIyQT2J8E0tvpMias3TXujBwBj7tkrZ4bR/COsKVyV1Ur1gWo0DyWtMZ6D57j+j8tQkEsT/OqDAu32ubk1P7TQAywReTD7fk7nu61MRhq/APLBHsDVEdFry/KOLoxhPN5rVcUbGX2uFcGoK9u58CPJ0uXyCdIwcfqCeEgaJRu3qDZgKYhmaDkPNJzx+AjzCEwKvajC6lOk1yRxnurR5qPqIJv1kfNXCN6JJkaMzyPephR/ck0yvyB+fYH2Kce8NXxSclmulFYGIPMUYyxIlVpmhwEgLVdkmuxHTlj6LhK8JtR8LOgjSInBGVtLNdkI8bSCPywk1S0AcqDs070iQ+a9lz0XUBBZaOawTYVUQvJbQzS/VZCgRfkMzEXwk5DPBdnhsjeYjOxjK4H5O4myih2yzw7Jv1zdfd3ri02t4CHGgZKkgB3f5zGYUW+tEZpkYSZAm8gAbfez1/1dZBJ9WZWjSA1BXG1yVr7aZfK2NhrkxnYdaw0DY1YWXhySJ6EZpVxdPdKWPH9g2bfZwVxlJToizCgDjIRh0iRNA7vT+6S01Wi5S/TxsPy4XPVL8/gXVQSyHwin1UKlugDRe024wzPmX6FFJaQwOcaIPQeUhRrXJ8qiJqM4UhS4fdWl2KMe98NOlOxGW2uHADlVu4AX7I5FKteYqlijKzNrqr+Piv03MLB05k468E9u7BH59yL4e873d975EOVHD3iuaeIMtpTqWl4GsA8yJJzWnzmTuwCxEr4HiJGFsoRFY6tzYyRsChDqh8fFxeq1zpB8rk81/E7rvUI+rmlqQ7H1iLPi1YuTYDTgogcsZrDz2y1AIqdaFu8rR6ulOt56bv2gPPhKwab223clqe2xCPmLsCIwW7qYzHE917GLGcjh5RfUkmDWFn8KhEtXUdsGMC5X9p/C+fvUDEgYZGFoIy5hmDFd/AtexL3oAq04gkK+legnx7qsc8ecySrRZUhNXx8l9qiECqEwOhfE9dKmYsJbQMySvxNRZ44Mxxab2kT7g7Jix2gfbrzmM4VwmT5UlYtGYY6dnBZyWsCtcGKsJN70syagrBBfayH8vlGC+X64FArtxlnTGBNM5Cws1/ccWaf2/HEL1H2wwojEh11hVjaRL7OD+RgJ5GKkLD7ISB2u86D/YfHXI3hEXxa8axJwEFiTyx2kOWTNx0dRYPD1jha3Wg69X1rRQ7CIRH13j60lkI1goL+MYgwXF8ik3YQCP1WRJsT+XGgwgTAmjitsxnaJIL7PEN8D4GzNMSxnuaFGJSWaIOb2nGTFC9097DcRocRmvNtEuxkiCmS1xwnCua/ZWRKJz7W5t1EQs/5SU5a/vaynMGGmNHyZr74UITSSL/6mYcC2GrqyqzGCLEjIdrMKDrYW4FI18ij2WTvlrJXlfr80eaxxLNr43myCFGEz6AnEefvB/9z1zrhJtYeIeTh/CjedhQA6mvD2nozz6sMsgWHW7NJ+xtP1FK1xe8nMR5SWzISoRbHh/RB7OcPZrE9aeQdkzlcuq+AYwXAg3H8EPDk3C5CjNICkzlLzxO6qQiA2ewLkztfrjerX2LnpV7drxySKGZS0NpO8nhIhbfUOc37jhXt6V2xAJNYFWlCKW/bUNAXh4j78sPk8t6Nt9INQigKQiwoyuh8x6IUueLaW2RuGWV1dwQRNdOwHsd2oRCVrkepfBUWPtubr7wVyeWeIX5K91NWg1itKLXR00YE3ZFXkVvT6sad+Hj340sLhX/c2tfyHegh+pVBwyoTMeuIS/V7Nl6wd7iujfCAmLp1APcDot6zmWLUgi2VYDWIfxYXHqZFo+oiXWdNqpoOJ14vE+mroyeCtLUVWHjZscxK16gQJml8k0ZiiuQdRTip7qCsPVPoE5ti9WUmogm9DS48ACtnQ2hjoiT6yCYo5cBqCjCm1D6FTxZsnWrxMyHcWiHllbnhBz0yDr53P28gq5SrMm+3CSKkagal/qMuKqsKfoo76Yf1Zf3nys3BnFTICYlk5Y2fBIUgyrCpT+vJH5b9/+l0kgJSvpqu2PI7XCRzkBWBTnE77QQkyFVEAstZoCPrZxe3IZFodysPTP1e+XRrbpLH5JaZm8u7JaB/eXgQa/qAPwZBtnjO76nNpjeNcNvRLkgq48oHywdo/Gty0/6Vv9ANHnnTmJ23UExd4M1pkZ4QWDOFTRbY29TfQ22z9DGv8uuM1b3MDkvTKU7kzUCgVDB7SeA8d4lV6zPcdGvNH8u+CAoneUh/4eahZPldKl7zO5+G3uU1LcXf3ZTKBHkwtraC3CvvZ5qcM+jqrNqs0KPnCNFxUvftCUlNZh9+JD0czcMWiqFSS1tmIi3Y57grM/V8aLFP9Xw0NQPGL4cUxDlDZcJQs4NjZp4CyFB0FXQhdYkxycpbl0opvhXOeskhrrt1BdneP8wR68PYufgJC7PbZ92FETni0FtN4PqEEHBdk5KnzLaIgo4kMOo0L5WFZio7seAmwNjQ3XaWbkA4h7jUA0MZGlQinfElknyRiA9Go40WoG9q8nmWgneRINtBCMIKNuHBZC2dxAJ5JJEDeLotfFvs/y68xM08mGtgdJkdEPyWeK8bIRMsOo1SjY7sAkWnbTkSLdOPpKxNpcd0Pat/U2RW29q44W0iR7O5z8OkSfqknrHAu6F349P1fXaNbjGHsODXtLqVp5oTnmTsUBXr8FKMjJW5xXwdBFpDYNC4YoCBGEALsw8ELoAuj2JFEp+XX/ob9O95dJbWnIrpQUDKZYKUGlJqSooNbZPKXkq3OCCpkoKli+CMprR64WWH0yp7/pUo3ucs9OJgou52Juk6CDmnupPzqcuIpC8Fm4IxIps21g1Vcnxcd+YN5DWm8HIsAiV5Efs3K/kceBf1KUq9BhtVMxTTFKV4bF+Uu2ltatPx64jbkLffyKX/gGQUn/q5otxcv0y5zGBE0oQN+VBMA5CIsx09DzEKlEAcoD3ZwTprUAilUM9Kh1cHJOpLS65qbDRVOZV11TF3NdW2dwiiEnEDvRVbedj9DKw6SjUeu+dXMFAzavlCKYmPkzNi+BHNkl48IuKjaTSrL29QRHd0Vchwb0rbYOb93Q3Xli+2eca7XL3VGpb0TvehviumrPFdi77t61L2VquwV+WjrOIe+OmGRdAgrHwv83nbaGeltS+qmSbGr5eyiLpvN06z9dEoE0l0OxQb8oX1bSyrLLczEAGlUbeHqrLr1PFsc49NkLOiNW0DWVnrpkP/e6S3k5ZLxJXRCWJr2soDDWurn21gR73LzSIFmdyjy1nx0cqmLwBuBJyXw5zH4c7xG28tFin6QeCOiP62uBhiOZJT5vDdJ90wEEYJ2SsVQHP6VKuI3rL2ZGNtSFtzptlkriGBkCpc0QoQ9O+Ey3n1LYUGk4OM7fhPzXD9AclzfZrw6a97U4X2+Wi3l82hRXOm0c2GKOFJKELysY4xtnvEhG+YEg2y5WNEXU7LPJITUdxKeOM1h+euX0nRRZjVTCPFGkDWXg4JyKe3oOfBXpRqpE4qA74agmLsFEDFDEe1P2AZ/oU8lMfceoaT4m3H+YEb34yUi6gKu1VqzYau9jbihjLDf2Va5YvW/DSAVVC6dvX40CJWDakSDPup28aO+eoIhSBsXTbwynI4Bu8Y97imKVMXRqvX/N+Ox+ZAFlxD8Gwii+QG1OHeTkm+dijIKoknWtAs8CH/qq1lj+uRLVr3ETZyuQUARDQmlD5qVm91nl5dCm1AXFJdrDQ+xDFAhRH90PGacpLLwIxnCtbB0fBy+5+iI78vX+MtXK8YA93eXxi8tfX+BSItN4CPkmL5/jDi77UGAHdLJ+IVl9cTPQsRVKQvJiQYgTNdxv2JGhhTjvSyE8HputSjS9Tcv85xEO+OzrByqK597xGQ0z5Fzh6RfwvHbljOzzzIvG7upEPa2SZX1G8svppxs+e6f0swtX7gqQ12HPxWw/ptUtMwsdKEJ9bmJr+DsePV5l6tnZ9gL5AbTapniyJ4kIaBrbULs3IF9dqx6J1jVcUINclQH+p+vvamvzD5Z0ANHT3R14a+oh6oxrlQnVNAwjMeMfiYExR2pRHhwLRuE4AVNSmo9RzoynifRx576cZ9pnuFQDDp3eBKUaCWC/lZpSV0n2q260nvvFAqZnteIw4rZrlmiv0XYSeAEpqFA6QRtUi0KLpNgJdPvKJzQwXUgnTu+lGtUbP9eCyenrFQ6CDMMSvI9xjMiZ1GRJSD6Jxceb3HQhCw+scUVxK98WZybRil6VevUvxg5s14q+8EiJdHyUXVYlugx9H76fqrJUHTzMnsADoWFBjn2Pe/ScquRSVL29RohXWJlFCLh6PKBCBXtJSsSxV18faWow9Coub32rPjDFtuOPwF4QZ7fUiAYCelIvw5rwrsguW3E43zP8FF5IescjqsvaxprkhESfdz3JoAhzhcG+HVtTETZIeztt0FmTtsmwH8uU8tOgMqoywoYIL5+Zt5J6FzL8+eGUBWzxn4OlCQkVXsLkjEB0vcL9YB3BKczVMxHar+gDvH4zlfTVabTErwQxpXngbs9sQ7gg/5KilNXmSB3eeM5Nw/nXjdcw03fLSbHpk7ChW5GMBNh8eJatI+z0sHjuzD9UTNdDA7eh7hj/e7YpF97hlnlLFqkVQNUP85JjJbKasPuATz5clP7KFSrXdhvQk339EdJ6FWqSWyIahwab+AzwmJV8V2/rNhM5nd6w6mwybSxW5y3xwsVSejy3/Y1MBqitsixAVRXa/kARsHt8QZuw8C2SO0T9nI9F/7j3Cy0Mue1w92TxrDOZGQY1fWNE4qzUIaiK1Ocr3F9l6G3XGOOHM0DMowWDYmsLFQQN/Ea4R/4kjR4AgQegxeJ/3BcS1igEimtwFZWgTQXiWi0L+xtqQYrzkvS4QyAHz3UJULuviSeiQv0XWz6iXicHFAFgwqgqLiagse/s99M6pkw4jBIBUeXF3dK1aG0ZhcMFgLc2186dxVw2ZCir3BHeyvCZ22oTNsJz+G2x8Z8w4W5BzOsfomzTFW7p7twIH4tMWWGc+u/R4SntTs35bVbvg7lP13c6c8Rnrrkf2/u1T+ipEejXk4VoGy0bVJel/BXGXPlRMiKhYIku/E3oJAuN+nJAMB6Fdv4B7MBdVqZkOhZdZFn6DeWLHZdKbwBG/ukxWoI7UAsyI209w0NsyvNc9ue1fTWYRieKdPJacUt3Vc4syKOf2nnqP94BkeeIYo27/nRF795GgLuXPncIdU4xSinnZEXSCEVURUODojJxeBjB4HiN4zOMOAuSRcEiEIivKqkp7QSA0yWMyLzlwJp++uGIpv9LAkQI8xmWPu1jqXsOrzn2kcdq5Lf3ICZsc3ofIWgfHA6haPJmv6snUXVMoeYKp5TFkeFCj9966OrhhP9YGEiai3qZNe+ldf4P65S8VybZyQqIip6HaVJcR/VPBsuhgHQf3OKqHByD8Lp0OwYYiph3Md3sPIKyQXaR3R3+w/AheDmPcyM9uyrd/CkN4+IMI64WLNPNaPWvMvV1J99lji7xwMTaUr7rH/mJCZXe8KW0mrxw8aHkvb5U1mhbrkxhQVZDcGU7lfbKzEw+pZFP/6cTkKOpJBlwGCSqE92RmtWcmwS+SePpi6L+6IyNuz4Is/F7Xo/GDjYqW2AQcHaivSUytBNdKKT2mSj0Y/4By6PTXcpBcHgUzI1T/ThpAyYNW6Uwihey0QVEc11J3tNkIw4DS72BPWhXMOCnS8EHeW/vfp9guqdvq0z1eM62usgUWFJPfNWrVC86Z7s0A/hmfrLSF1pa/G5wSrvQ6WDqQypsngKM3+Wa2RaTnHZRBs+FxIDOh3GXZLyeSiBFeP4pjR1yGfyJkZwsxbLCucQunGqZ+F5Qz0SEPVcL3OdDQ9+1SUenh7b4D13g8EYX7JPn3WR0rZirU7RerOb6Msfv8L62IzZ9RZVrGyhSQeW17+E16LQCJ7UL4Onnw8bFSGFRZSSkz2OpmIT2Y8OayaaO2/cf6SVaZdrySZ1O4WZlzwBL//y5TmWMBGBrIAuieyFVICjSKOmoxOzYMxFjSgXzYEMNdFcTvd9CpoYJ4IFtz8sM9zEtQzuS7LfAV2alzfQ7UvhOa8em7lHi28j0al56rNuC+qcAIlL4jGqYKZi59CQBRPvpHYvVRUhT2JzM8ILFXUNFJf1mQvGvAoOtg2GFAttgj6Ymg2lC9J5tkLwEAD2ZazmtTwk1Yd5tpmfLGGuvw8aX9g92TvMARjTR1yijYHfZVO1P1iBIL+NOs35tDjb16EceYGuC9p57kwqzNLDYmVZ0VWgGzzaliGDcSHdDKM4Z1JzcWVZVmxplRakPM3W4+eVsqMEVH7q0Bf1gSKqwcKhxnm8u8H7pzmgLYMs4wtA98W332fNG45GptmZhaJB67NI6mJQck0UsA1LfBVWKxbBjOecPsNjifjpRKVJhwfGcdeEkkVM9f33Gt/ximM05BUn44kQx7BOcreb7bk9TxG/BWhfpH4eB2OHg8fq0PSseyVblKo31zTLtAxlgdj8nC6WrXT7BwW4S8meMvGqbE+o1U+tFs9vlqM10yte9plH1xAdHUiJVsbqjkLv4DmQKYuhceaKpH81Wj+EoscriZOUG8TtHvFjfP1xMX0FqcxVkqFRCvysFCXLl8uab0AtGyTeLKQ5XgM86CNB+gjnAXOee/HO6FzqMXyckgjsW1aUZ/H4He2Bb944OOn1iylopFsN565sE9Xo4t/MM7R8IjbT7U71Q+7Ak7eahzPxY3zc1z2mlIpjhahGWk2Gzizq3FZ7eMhN+0qpFW6l5OO3i8yBIf59auOTNzsnIgmYWKwX5cXdORsDxaSXdjricKZ309VlsQUvMX5GknOuzILKPjX5JuF4vLk7hvda6xKz/fSMJAPww=
`pragma protect end_data_block
`pragma protect digest_block
083de30fb2290beeb48aaf61da2944ab844dac0e05f42b85b41cfe01e57882ef
`pragma protect end_digest_block
`pragma protect end_protected
