`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
bU0UTbNECeAbUy1YHNZHL3Ku7q+1SF9sCJqO26snpkZ4u45QAGMxcm1ftbe92vNwuQlRWWX2LszkTZU2e7bTvtVtbzgeGYWVuTaOn0CawqP27dUIB5aO82k5WUi9hc3PsuJQo2PWkPUwMM9SmlObGZPP5c3zSvJ84Yqm7izEGYOA/OYd8oFywLyVbVhQh0pxGiLrk/g5xv/tevCkx8ke3H3sU4oETP6jIG810BlCpLrc1JvWkTFSwLOEl4LH6hKsOu2sq49csgb8Hu6Ux7n+iWKJU7RsMqVybzPx+pKD3/KOx/pS9IgsjYrXCMN2l1EQOdKQrue4FO3/8fqTW2R+2uT4UkJP2fqqH/9IAzP4AGyJoYNW2uOYEMkXqZw2eMYOWWjnp96HRyw77U6ichLvoDi2kMmLzBgQ4VdwaSDNaeN1vVH62G3T1f9ymBcwCT3JjO95O1d2YWvEYcdbtm0RdgmZkOfix7t7JbvVUCnWUEmZembg6kzv2hs+SBYX8WnO+BBOLYQsbEADkedj+OkUnhiiJerKsfUX4OwxxwbDaarGfL6G4NZ8MEiaWzmWnt/7IdlvNiDN/SX7K/dpYzxnM4+expVlr2Og+gdBgzA2i+RX5l/w8eXowA2e8Pw39nsLERnw8kuH89TKL09T38VcMzj11qd1uMaAyyLCQdzFOpscDi7k8gABgta1Kxuubc2yKYGUYWP94slA5W81kLgWPx7OvpfwR5+SPBK+thm/WFBq7CdTy5D+XhJ6gTelBRq9geXIo7Fzwb3xnuCbO4/A5UMfvVNjdPsDmLzaok0yomuqZdQPAaWtsW7wIv5dpUutX/QFjer/zFyZqNzdjAy7Ct8vWEIEAC87AMPb7oCwaXek+fojV+b9TlQq0/2GyAlJP1CNHHua9AGsb1dOVSeS611ouax3sJSNxWurvseLarDEszE9NHp+X5EfC5gGN2BEitpRbklXoTsXDgGW/9PpKpAT0O5OsCwbI8McxxTt8Y0N2JPggfUGxtMoHJltmgQToaE6tPvk6OPQQ5Najc+AV/DPm1s6H7DIO6GhYpHdL3IPxBsdTa/25QutxCJ0EKNq+3mUq+jEjpM3iZrF/vqmYyJQ9xBxdzUAm6aQhNZB4PMyVxSLmKQY7OaXrx0qChUjfTtK1BESJXz4FLN6DEGPijO542ZhrxX9KVJNhaiaUQXFjYYp+/pwHOD+if4O+XhEF0zmCQCIcAv6DL+h4QWVYm3XOHd+1mIuLt0TdDWqFv9gmQyVQl3xsWEsbptkiS8ZEpV5GPgTxc5ppLYloZqfMSfa1RMKilGf6B2gXXj0s/2InyDx3ixIIz499tJgMTjbshqEhwgbD5tXHsVa74fO7k0kXp6tDJHWoD0OTcF/Ov8wiFhczKVwzWACn/gBwDiZSYsmTH/qVLe0fpQf3NX3CTZzSwppRxbgxT1XePFWH6H2F6YCP+M7Oin/tvIvKBDLP0m8Zs3F9U4pJVvgxKXU8XeH4aeVr08ktSkV/E/ByNPwZOLKy+lHTQl44m3M3Ci2kYfbFR46wjZYXrvPlPxCzT2ZctGIq3V+yawfHLjHDVulk2Tx8EjjqRjnRE1Ot+lmPY2KKaNq6kmnf3FwY5I9+yV+OlMragw1X6HSOuscjQHzktDNywqmqqIR/8DkrV0vAorVan5BBqLRTD2i7lg1+Ewppe2143NoA8LrSzLYSwsuBWy6YyPmfe6HXDdWj/plfIMYRmi35v5KygFkVVWRU80BMfV/7/nbwO1CuwK194LVgpMBMp/c5SEHGtbZGw+t47/cFtRo3dQ2uX9ab2qh5+Eh68rXptiqCymL4F9RltYOxS2E8linh86GZUkB1faJJVp/SNP9NcHhAIiMH1f2xxv8yQwAZoVM4Hlf+KyICzd5pM/cqrn1oMhbcgzrUFaSRzpo1hM0FzSe/i5e7fVO9B0kwCJ8A2qj14ABjg5j3sq/tBfw8hld1SK9WdmszwVlvsyJJ4lwhS4RHXZTuCJ+kN2t8N16QR9qLGf3dI9P3lAPBjCs+ZsyUtVlgu3ZSTQarADu/047Fn8J6mjlizO+3jlDdLhK0bqKLOZ8xRz0d/hk0L5hPQFWkexr3t1G/G/+lD1UYoftYPrEBYVrfRhao5TiEjv+oYwaEjBQUAA+Br/aUK1QUaLfQ8UBOBaOE78C5fHobFP53fcUiyTXpteMKucEjA8K2+msNcZyPesH4EkEKfYGFqBuNmgJSHVd+whp+vmvy9gTQtokeCriHMKWiwFmiEFNQH5jd0JSlsV6oak6AtQhnBAI487kmtUEz3B3z59Kdgq/2/Ekdy+9cAulMPBY7jIzXJW7H0Q/DkHulqTrVCnYJW8IxQfhi32EOfYIhNJ3Y/I6tOVCpcaOvUD6G15PBcXoKQN5cxqPHzDZtzJPN4bUg7ebzwpi5rUP3aIQpvC+EQQjehQjf0/vdURLb6cOARwL4Tm9369qEpZRG2ZtXzOqqLzGt24MtTVBZbuIJiXZNwWVHZ1VCWkb1ops7z4vubbtSd346Pp+JNa0UkUpErv+kNUFPr9lTxl9Qci9xr2YB7LtJQtTyCJ1jqdM+jR8o10/FW5QZFWRxB41uLfXDQNhCtQKtBHA4GglGAIAir66rZd8QYjUaFf5GXM78qUIAVCHirw+esQpHx0ybtbG2hWFUwm7cwKbchbwYTB0DYibE/jPemb+AsCO3WbFOiJFr7Ih7VYBem3w1yHnZDx9iq7URvTlEWiJFpF0sqR9PM120w6zD6sXZ5KVxYlL4ujwjvphFIaoWaVcWBDcOY7Igp3gFD4S3v6al+cPJAcAJumBzrNZhpDIm4r1Sie53KwoqFQE3w+o0xNzjKTrqAE+BPo+LVO2P1faCiw62DaP5T5nkXG2ytJEEqCgtoiYJiR/MRvi4o8ucFEyIpUl3lMcrJOKV3q+zIYf78hqRyYof1idNyMGicEE+uf6/18Pyb3Q5uL9M060gfcCa5mP7sLBda2RonX7FbgiKEUz1bbw/G/55vC4tMRxd1GDhTonYBqHT7t4oUoLlfoDl8xG106YIsiLRLoi/jhbANCWrQAZsDl67rPw3ilAAzFd7j7FegryhLSnBlgsfdbwZR7zlOlmjOFcH3dwAGCLKpopY12WES8j6LyuFs/MMWrpU9zSnAEAzeLb9sDjAxzPteCH6Xmgi1JYLFtvfZguNLtvmMV462+veQbD8Ggbz9oPNTeqSYJ8jVzGw60RikFt5t+g6cYVS7Y4P25o61VEDlfjIiRn+sMFn5J2xiAUD6MqHqZ7jxNZipgg3s1/fKgRPSXTvD2QxoEQTD8EwXZEF51fV43iLTtzg4zb0gjMOrL96Jx93MBPnABaad6cd1xDyo2oA560kMdwnoyTaJoW28o4gflUOY64d66elYoBk3CPN/5fNMOuDkUT0t4dG2JLF4iJt2u9DnpftW59Euz8Zn+rdZDLX9rtWrBectm0ADmPj7KZQlczwebEdlrVUY1VVWWhqx5wunA7eJ97YAugtVfpdCu9cwqJmFttGLM2ECqheFAI56afPz9lJBhS4KxUeuRpsH0rB+Z+PydtO1bg7VrCFRrIF8i7MeDyHoy/FatzCAvnob/D630QeQo/6590AIyRgUqJGIjSZNEL9A1NwYRo1UdszwFYccyBUEuq79EJC3Nskfn0j4oHRTYjj6iXyAMQuUgdUSjymlhanQ7tTdR1AleyG2UJoW+OpAaqdJeIJA+swd8YFvIKlzT4IqfGyxolJWTw5wR6+U0QtYy+QLLgvrkmIf6kUiqZ96AG8037d41cMZwTL/L2Rd/dYIq3ROUc67jScijtj5LHgz7d0X9OzAPIaR4cDHKubRASYYnvZiG47ow6rBDT0bQCO76f3dp7qoTD62yKRHK40klyYdrX3dUHcrgkzCjsAD3Fz6Tau5kjwttLJRRwvKZvxHuys4JGs9kJTW5HB9FTASqEcKZxIjreVpFHsvCTCtOJUWCqB+RjMfYUmqGmMcXYYytQENIrfcNuIHAsg3qwkSPGCue3Lp8wKa/X4boXBQ1WxQYuYTsZNhv5BRsWVq2c66MtlGd7g00sGLlNkgV4tj0Q+0MlAfGnmuei5yzFl47T6bv+tlEc9aD9vsBkcNoC9yTjKRRHteiHIb2Hy0xHSZLKnqA5fyC8njyPCKmbBvk3LarfUmGbOfZeLjmcVrEmXBYo25Rm6qQWwY/0e2J0SGp3Mt8i67GtzEAIu8sBeM4KnIfIRRFBxxnqLH4GsBbD9yXNB+twepWmD/0LsL9aFJoqu4Gv39NTcXAIaaU8GQ12nerNRHVqqOvx1nSeXsPtw3E0MqMaEIv10p1+sCVX/FlrgDrProMveXuVYw5M25I9hgiEdjITkrHwBxbLxAXAQuLlglIUcIxDejUu1lIcUFk7jBKvFY3aZ/4thXRfJgiSxBIwbI+rMrU0lQ+4Q7FTB1te5xn4GucRNp3h5M+Rh3Rm1ql+xmE9Pckgobk9WBYM3ujyoYu9iLUNCbILQgWrc0dyMPOdX/yD1Dz3idHqAytQG5pXRBuTJTPlCIwjLdoVkTSTuJnzP18SEBBGv6HAVpMF0Ub54YzMVxCHbFGUtJPqewX2WaudsZbOzEHpnJDrAOTj16/jEc6XPgBGzvD9uYrxcRGKlU0kqX8OxBAa7+qvDWfZ34yQwYoVz9aFEBkdF2WZAFdjk55iw7RdX8jF+CQ8pxSOioPt78Yxpxpkh3kOY4ByiGaBHJmecsJG7kB4EAg5MrzBjlGXXK8B8jX+csF+FR9hAfbRZhh0OAxQXW+YM4phn2IaAtwumYQ99ymM+/+h8EEEMYBXoohe33hSMEqOx0nUOO3sUQtJ9ppavHbD5soeCDZYqkQSdpFR5o6NcZVA3mdCGa2zvJuSbf5jJUIlfQmnkhhgqKNmNr9pmZ3Ikut00IFbKrOjs2iws3hfcfdWa2vXWBWYoGZLEaunkSP5HzPN9OBOoD7hPYXHAAaSMhPl+ETpriMPEwQlvYD05zGpOCb1RBGdrMg0Scs5W3P9/WzHbX1CiSrjrryEyn1FBiFc7Gum4e/oFElLTNQyhv0BewVKW5baaxlTTBHkdi6k/P67DyGRUqJKMWobcND5+56h0h0lKOXyVzuY5s7208oVhiDd92poRe0b4kIWJnNlb0vQyMV3L8GLQuFdO9kmr133DkDn5rxCMK2MjrMNbG9f4Kr9zLOtFrVnLhdOnSuadKPlggebAiAXdZVh8y3v+YvJ4bMfiR7qeTIMEQRdZsH8MQKDj1L5mfFu4rmHJ2kxzydKEzUzsa7A3LwuJkvvTCMENF8MG6Jh31zBdtklodTB/ABP1zvgy/vQNsN8w08jaTQo0QSEJOY8KBLIr/l7HYbPUhEVa1BmCuad1+L4DejDEqYZAcDGHgogfcqUBlZS4PhRVaEfJ6Iy1x+eBMLIJ7V81nTZOsxgeAKDxWkBZgq1UqJPtbegPRjFoBteX1WW+ZrnGgVdRzhLHDkXjvE1N8jjiwNQQQ9Y/Co91frVgamY5ZCgxiMzI2wCwyE+Lh6g//5dapSX2HL4GGdNGk/Aq0FsP/3hgvq9mSNyYPlZoNGNKg+LxfA9DfbOJ8REgN7JlPJ1G0fBRFqgcH55HWhTfbgxd/a7yZVQ9XgRAuM6yoHAJy8oRV/38umEg/Cee6LmahJKHrBPnK+gDznQB2OptinteoofAJhQOUN6RHDfcoGDAEj4qNc0qQ4OqWMbjbekPEAqmI5+/zUtdm+q4u0RbU1IrsGdrgD5ddVdJvQxRwTOwV+2Zmqa16u5H6RrqFZB0Qi9n1WWLkxejq4UeuP0EVCv5oeRImG21kLW2JE8L0CL8mqgpcHDShZnZ9vmEuENyOjSHbn9CDtZj67ArBGCt0KCYSIfbqDpJQ6e/QzluBeafo5P7MlbuFAq7jqBVkGFW5fcT3U5Pp2MMbmlndHMNQjml6yxKcfMai9yYSr5Xgan9nnHqnDffSPKfYQ1zbv5GZ/R7aKhjLCRmHQ+NSbk+EeDHeqsLgWOYlehTXkoTbWRPjNm8+BoZ3EGRTXUYpq3HC1u8mSKuh4o6QrKdWAeaQ9DpApVA/xE9JdACDx/hklZq8bQ0R8Novszp6QprvbtJ9hTEPP2OT/zab6IRHyrh2FubqFAg8XuH2NY4VqKzCjnatOwsEvk15Ofcx6+l4J2I0UP2PoZZSCGtV8yGBLPU8Mv4IY2B32yk6hZPCHG4FBOjtcm7fLyPDORxOf6FGU0YS16L75Syc0sj3nrHVCSeizAkaapLzo29B1qFu610HM/3sh1209fbaFgHd6CTEh6BcXdQflr/zihVF+hUlyOFeEwpqlLKlOdWHbj3IQp5HsIy+h/0Q9EuqABJsNJQFPIIufwUwzYFzA/royMT1jzzsybnqwTacF9d8ROD06pLmyGkMFPAPZVo/8bnY+weHZksM2GFVeQ5aIQ80q7unw9Axzv892MJr0NNN+zklD85AmJDQo23fzcPzeoF1CSbBQQZIy3abgbvQ15cVTWXBaRxnUfuPvfY1w02nuZ/CoWUxWDAx1W/obexOKSyUCrsLzZiyDCpA7ykyXoOpxwnVo/mnHVITl84EWhfwzGGxwXKPJwr/t3fD8Vl3IE4l9c96nBSk6HbXV5+LWLUKXJBbZk1r83iIVfn41yAfUZUWx8hfIyjf/LeQg5R24bRaewKVCQHbGxdqYLSoKvkPmBhP7XVsQJn3mmm3as+vFTydt0aYLaKeQPPHzk7z5VrLP0RAHtDHRSkvhu70asuNSqp19MdUO5nb3Ch6b4tcA1J9FJSsL5Xfm6sXQGExpAlZDUoICvHzCjcQ9RkdKC2tQveb2azTlC/JiiCTCCxB3EHanF5Np1DpBdHAix4PUW6hmB01s+gRWFM+NpJ50fIxChEp3fOKA1SPd4DEvMjslRzk5CD+9jdr9PKJ2b/slObkD73mQY0ifz7gdYvDZOtAtrdfrGgo0xFn9fJv490OllpZ8UkD7auAaUvg85CjKRTRos7KMVYKJMuniY9pRc5B9luVtX2954fCUCGfHF1yGa7GcWxXxzbW6rbdCY++XPmT/c1bjxeb2r6hU+E1D9/grv5BqprbcDGBYwdJJ6o1mgTDd7xz5j0XQNhu0yMf+y9lwPVVKDl3eb5qAAzbEppxGXEQLWct4sWUgN3A6uoieR8N40iBFjkNDABKHOCXWSJSwBkVTLUCzXIUnzN2/TgaUKQ2VCKZrMzZVIPhsm4PIHEtRemZ6Ai2UG7Gi5gvLesqSHcMdbf9WnTUyZ3OcpHtqTJAJpUmjqvI3vvUI3sT165jJf5aSQI4foFi8IX4z7m6kBGaFZP77LNqLT4SOq758u/T/eXUZ1YJAPgQJz/irXbOooE7F0RNi9AIC/xue0GlYoXNq4qe14+7cFu3Ac+MLZIYqIg1Kcqgaqu+3Ul1WcTWpiv17ZcyEtstrhM5VPvrZqdXDA7EFYyX5Y0mI2yyLOOrVbHk8XxTRIE1WmDRH5WPCoiPiY6SctnPQY9jKU0+2rMdCCyGKA9rEykKyCgP37qrmj2HT9Me8Byy0aS8mSBpUU958X/zx0PKDpsGFc+t0RstC+MLGKBVQmYjJgDFeVFdodwY0JKQpLLc9NnYei+7a2dY9ho4eb/VAfed48D57WSW13iCTBGKAuK7mUf4WzW+QEx1BDojH018Va99KCcD3AuPX3XP3qRgMnUvbTSq62BrybXohhCgnL/8gkCB6BV/dNaLgV8qduNitN/NgjMx/vRUfIxPruDMxaxwLKrIrHsgJD7b8S9/nIGYeRYOu+5kIWrL/XnSeGVDxgfipAxYHru2Aerm+ACGTgG0kbzJ/aVHOBT6SiMbUSbLwJ173eMp54Ahde1UoaQQI5k8z262pNr1I45nBepyh6TZ1XUcnONAxtkg6bHpwwnayrzDe9TRqiJ252CMReLkHn+06i8IEeZ6Ohu+b38b3aVPQlDV/Kbt122e6eEwJhvscQcnISTilmRBn9V2D+u/8nwFz9YWtav/4S4AyadPl1LNPQ1xqd22TK9VD6JdF1Zt4BiXxr8JLyfPHrCnX/CHtrSKfCrqzVU7+kwrJK8QRQ8HutS4q2CTKyQJ/KkRfRDj5mt+c3aUOn/Y0LqgivxGtf1GAJsTeVKf6y8mFRmFKb0VLBv8KlotBNUcFiTr0RNJkiTJxv0muPk2x3LFFprt4tYTiqEKQ5C298yzdjBi2wBumkPPlpbVgdgdyx/ZwX0k8nARH/pxMiVIUZys0IKjjAWxn/BNUJyhRztV+C8IyqAs/oTWMLP4p4FuRzGpPveuUGW2i8DeYvQ31xZKeA2AkdcRvrEvbzBaEgukbJp6JyJYylun4Wd61432SGouFLIF4zikiQDGstIv2spbHzG5mxOJ1B0RiPTGiQTyzE4Fb+7ycU1R7YSXVaMyPKCWAK4WdMClm3V0rXOXw2PUUFuGtiIxETRI/ENgyB6YkzPUz2Tg589ZIJqemNP40gRsTkBjGiqlTJ07q+gbZ1IsFBiKAVdkgQgjywq3SypIUIr1pCOAKcgQtZG2fZVOd0RO192Lxv1QHHSkMS+zj0Rx47DQADBirk0aKR1xTh2ILnehkrDcmGxewFwLLJwqVl1wcuUX98d+SrD+9A55b/41l/HShPkxmMpnV4e+7O9ZOkJ/t1XFRirObwrfbIwlC73ahnTuEg+xSIxRNBehicmlWqCH7By7IvCuCC/SBihzzJC1YD0dpNK0MVsyWAZfvgre50aJUOU930otVpfcGh9eML4VJccfYGZeX9Bmd+clh7yVPMrX+De7PWMe670gOZFY0rFEYLO36lTOAc5XphnSxTDH27Ebvdii+MEfws/5Y8r07LmT+w1gtFhJIsr9R/eZ+sIt8UX39mT7H72RYLTwovV1sg5zQMMEneXsNdjhfhHCLd7LmWanNubrcul/KhjhfOFTwarOfGwrczk8n2H+bSUj9eh9o81drJxx/QATfIBH28NR0VzQ9tMyDmaM3g4z5pen25PDaHRWSWk2rfCAz1pBJba9fxTOVuG5Czkj1GtfKNKUDCfeTFODN27f01doU3DVvbmRTsLO6EbqKQYblgBFEbdKpAOO+43CmFvZCznNInL+klrnjBq8KVPDfTb8O07TdPY5WCTeurSMSsBOjOA4OfuePI0b9J5og8W78KI4V5uMHXKIFHEKKDWmL9/dtCHzm2+cDSmKslqSUhDeFYSQ3Wr9OF4RybpcjuvMpbgqPl5hYdQiYzbbkvie/uETBWt1fu0q6Uhm5IlS5GmrHEDjkGTMZ4ko7NQ0mIM8FwhQJOMo5LCmyK0Xl31y2uooYQwAgXVX+agmlRAg2S6gR7oJp2WaA71cqkgzrfQUHfpsm6SaHJ3oFy9qqe8+U9g8PrNiXclIUcbyVQNaErVCdKqfoEjQ1zqFn/Htqpqh3guwgfyNtRcEmJ8TRbGy2DcDWHEfjLnce0vxLt8mnYs6yxsmio0GABuMeBf5j8EM1G4r/3FHa1NP7CxoQy7wg85BuGypogv/oCRZL7EwOZv2TD4PsMNhzsWH1tgUtVqRI+TzvD67+HeRsmHEiTUen4/5m35E9BcNeZd8g5BrjeO1JOkjMKOH5xHtZtRiodzmbTljUFBYJcrgMnrSNKIgiM14m6koU6VY4PweOtedecHH4tXni5nVFgZ8E40U7knySxQpgPHtaM5DsYfZ1QSO9ZiN1jfwTMXu8uqHg/8rI1qKLajtJrdOvFXPusvCRt+6OPDNWbTPKWSJ0v5x+Jpv3kEJPSOWp73XXuAl0Nc06FglVLOS7rGryiX5HkdKuGDPX7uxrOl85ZnN3mLZBlWxtwPQT9WXboLF92yHawTNMXYv57hkIWa6Dn6mzlb+zSP6EgGI1KthPt6GkRD24jkux5oT9EHFwZFpNC92YWDy9On9oBWFfsKzd7ZlsQdaWgMqwAKh3/443P+F4NcoxTaqJOhUvgccE6ZN1KeVKaa7XkxxKdMtxWwuYP9uMhvX/Q2U47apfR9iYsRMtyXJTeUB7oWI/HScclwqLNIRMfhbO/N7PTMjyrpJ7k5/lo/YIrY/6Tq9zK/gv2M8y9WOz/oo2rKJBQOh6GHi0FBGYlIJbeyD6jNuU8ag6JbV+wRqJs2PeREY7M61LZB8rRG0NnnYdA7yLGO8/lIplLNy/nGTpON7j2BXzy8IWZou3wk5Ae4l4OWKyxvtmr2NwbWoV0Z4EEi2UDvhsNccpFy6+kIEmfOFwEITld5FngvsEyN/Rsuw8PaSc0FUnUn4s9SEV/E8w6ELtFwH+KIFDGs7R32IvvT/61LayDFGb9HVtw+Vo19mh+t0CiglQsXCII+7oTWj9qmCGsbbTQC0pSQtM3XMSSpQ7JdKlTa6Gpmiw1z7jKzYBd3gXI6Viid9g90FoT5vugplyAAnQ8zRY3NxT8V6MG7lGvlf6pBtM31kzGvt3p8rvckQN585IJ7qm7RZS6xwEjoNlYy6Ncz+xxrKjsHJvgzV88s+lIxQ1iQoVLFF6F64NQryE6fgUU2IM4iMlWhT1F9IGBFKjlypHcJa8EPjAyZp8Tgo+8yCrd+9/CsfdmPw6NYWZmFWLSE7zDKL9Wdie7BCG8dsk9ACM9h7EeK/T8DaA2iEZ7i6L8+EGEtxWbcJl5C0P1Bulp+wT20Y5A38I8kKKcggmwxVRY+TRPiL4oRTmsNaDCeO89W5ZinOSi3tuAZ1Pou9afHbDUgE0eVLnKL55PpN0jIT16Tffy3/ws2wIBYmQGdIRjElFFEHFqJPH+6IvQp3x6gZpVCvKxbw7ZnnZKKT/UOjftw2mrrA/gqvOaswtuYSTJgggL3WB0/JNY4Lv/IwUbokldmOEPpXRNPdDSwbMMx9qNoCeeU/Qsm+MKqupy/yBjO3wTDjPhU/fGLJyZ5HImnWJGn2/xDjtM4RLOCURHyxol9Faba3BTWZbUfbGLWAIEhwRerEDI1AialHtH20BHFcCq/kIN3Z9XQy72j8Bqe2cCytI5kZ9qPyccGgzVqqEZfc/73y3ltlXwpiZVHCweqdsB0D/pvLXrmdqFMrWcPZIwaPQJKjOUciL92PE+d49t4luoBQlU+SlcwoyOMcADzxm25OD2nJoYsm+QwW0MMxUwhrqMvL4tlOEF0csQngeGkTxLkFCGL5z1WZGUJE7cnp8bfUGUfTH9xcUgK1vDvEm9KKOYtif4MoYrIL0fBXYIsSga0fWGaeHzvjwjy8Q6TDf0b3WsvYuL6f2C29pf5/Byqo9Bk6XJ3puK5Zwj6Rf2VIrWiPH60qrLKyBBiblGEzMR+rtOU93NoEKWqOc5rrop8q3ZV15z/TB5RimCfnhaijT09ecFdGgI0xE0k1z53XztdelxuifqrEVBKhusCsusNyzqwap0KPwintqGPSb/d35QBq0NfkjLHHz37S86tcWMeYnzuDzT4Y/gckqHr3lbm2qM1yNwboZ6yRACp3w+F9bd+HBqVeQI7jqJbtPp+J47es25zX+RA5OV7NdNYFiKW8AIWAWi4Tpt/jiqn5/dm3Ng6I0v3GeVVZUdsZuYTm+JoJWuPylj81GnPNllp18hwVbkXv4MlD4190BkXGNcJRB+e3KlnHNSRV3/ch9F+HFebepDH4uMZVIn800bfKr+I+6j5C6Wwyw2Fh/GlERZBcwHYpR3ZoBJS7xq1mZRH4EZxW239obUiZ0lk1IThoRw5guYr/rne/UXIywksNS+Z/rCxL2CUjFeIYjzkb9/Ob2uFmgozJqYSGglqec3EtiM7ju+mw8OfvoOugaigwtUgAY0PFxapO5IIjKi3ni4IDR5my8I9/IVecB/ZNoGvGXtKACucxuneKbjVNH38Af/vWRni8lnQFcPqYICUyKbKeGw+pg31bsTCYCaVX7RrulfFlgPZcbVJTKSrpqD8M8C6NfPBDXzmRrzrvyqreyWUAGFB1iN6lfAebI5sBNFU1h+Nd4mIKOvxHvPhfLGc9fJrXnWEiyRBeCxjsKi6oQrImLaF0iMANKNPStJD/lqPUaOW99ihb+BqFQqgqxm8ipO43Qdy0iaobS+1iD3zeEfpb2syANd0/9XyuL0XuPlSp6ZgRiF+0aCwG9NOOjLNowZ0GCDf4Fq7LYBe57KVO6CK8sjHmwrsfqovqWN+FMT9ypZ/epKF1xX83pzuXOaNu8wffbPEi3j2FJSJ14ehUnu0E4YvpTR/kgZANv36l8I/IgOg7fCiDJs2HFfHyfCITpTZnDDtuDW3/Y8FS9K4+8krug5tiIiTUvA5JKnaA22IqWchFiW25n13hADFmY84GB/0pOxPT0uI3OxlySJ5my/72vJPTFNdE9wKhm/Jy/ZEKOSrNO60ivHMnR7o2xYnqe4Q+Luw6+M0TnUhl8fynqCoB5DivBPsvoKF1DV3IUAh4er0Gii/4935xKhnbESWfDOx7MYj8Kq4PBQTPP5ocXct8pmWwc0mNem2sF/NAuz5dTeln0PilUqnD35MatdvsQMnDJhfHrWk+EX9Q3NrFRKw6WQHgkBUh4AB/P7zVQLMitjvGjts957KJNUbnpwZAhuVujLfso2/9SGZRfAvjxTxUVlF0WPNJ1/EIx42Lg36GYhB7LOww9wxbz4ciIs57abPvwSYaUvPNbqEQk+JlisO6X9iA6BAKRbl9WXqYdWynf1KgPDMafemEX2BN4qvjyJnhUYbA9h0a2mSUWAKVzbYaCCalvE1WOuBY81ISNDAimvIGokzbWigIUvLEUuq7rBunSbsDoMwntkVW7/4KTatdolrS+1T0j+z8xmZe85QphS4NZ1LjZWJq5uYNqFfGdMGucQgm0pSbk+psH/ncOQyTTJHo+0a5B4zFOlLZvcZfWtznojGBg2a7whg1ycgllK4DiXpdwY5zYPV9r51bpdJBOonHghV2Z7ihSj7q2Kb9yqPOfuxLRo7AcwkV4iimYLVWLIQvRPt6Nc4nzZjt72jG4PPH1mGsIf8o/fpeWAx1G4vv+762Y4Wqk7IWWmb+DYQsedwGBaPGoDFCUS7WkYSnjmmrsbMQ/rFwd4N2JfTce26SOHSeZpHkyv8BDNULZqAZD12ERWlwf5FKu6WGddXZfiXxM5OFGE6OYpXN+p6Sq7QiMC3srckijol1e29iojldCNCtXMEFOQqLE6HI3ZrXZ41Xamyok6m+d7TX1aQ/nKS22sbNTQs8JrBh49Psk7S1vaYyIkpH/iMenakamYtCdo8rLx2Rn5WhwPgtH/JU/dVJAv9BqtTNWjCuOUzwy4dPtSgzIbKTL9iZ7lo/hlzVQLgCZtf+WuVhUJzPLLyxSgMVGTxro/maUnEroEftQMOCKik8NvGi1zHVfyhGIh0B2+N+yee49WJPbx9q29ocWkS7if/yVDQZtV0ZUcwhDwxyvT6y1aPxJKRtx3yxozNQuOchrZnytdpKP0zuw1Y0RSLCaqgww/PjKGdEjibFKT43V9PJsm8Q4IXmTpYkdkqFEcQ80lnOGi1QFdPn7HACpsm2FD3t7pd8SaePhEPoeYr6AJ6ZZYNFnpOZSJSHZD77TQb/msjRyi0luUdbcBydq1a5wBUtuD8BsYMXuAvpdgNDflJIpdTWCRW2lCpHaiQ9rR+gC3C6uXSINAcRa6Ys1TecvSikC+0OwRR5sHtZmtG72aJbCe9HfkYlhQdxZT9fkDmMXHQLXR275A99q1xcIJiimVALsDvvalBpFnwhDnY3K0vJAT/lTMCT57wd71aikS8tPFOM09gsZ9iwk3CnAifUKRNblszq8qtmzb2MDmZTMystoUOeW/BRdxNyyKmWqlTMRDOs8T2UFsdIal7zbTbZ3RXUuuwEMJTjqV+3hz7reD7zYSyLhly1Og6nNu3csm13bh96wWto/8yAanjsTZGRCe2oA5g3sCfr9wabSG4lAjFQdAkghl3ETA/nj0ccYhdcdhAsjIzmv869/GAKndzdpwDl+QVczUx+ugkxVE9CM2M+9N2QN8tZTPaz7vt7FKat/HU1T/rdzxNXeq57MgHvHbSWeJDow4uDTzyWFttoUY13jUzciZjzZzTZ72yGffTCoBlfg5QBEJ62ujUl18UKWP6octYByA0TOfhHQK10qt/jKPDFlmC273NaPFH2ym0vRw2P+Nf1lvuAJ/vjZrNqJAYkNMCiWAon+j2Qjpn3ZLjnjuFIn0EW+NuifehDM4Ycatjv3CYeCAQtugrHxRugbZr8WhuLUUkOHWaQlO/AdwSF+K1SrwM1QHeOpHN1TR/7EfJe7S6ZHA8WloPV+f11wZ1Ltu+P37LcSf5eSAs6MYB70IU9Xjq5xFpJc7OkJIEZmBY6+Emr7/lCL8N/W/pjg0EWld0KJI882o6jfAob7/7au9yYdadZsxsYfkCDWe6Vvo+0vD2ZDyZKshGW3DeKQKRycbCSf49qPxgYkqUX4oW33OZCfAQbyLELYt1izyy0/zzik4IqHzipvX8TCv+vStesDTKugUnQNFzSTwtlNRGIFEGZJ12eaipDCrzHbmgxckwf1lh2ain8NkyZfpmGamS4OiS7duvig3ZTEOz4E9g3peYuCLcCXLfBK5PrRabuZwck0T68sOND4Ro44asKiTUtvjsH45Ms5mf0WfzCDvFi4oLLo2E8YwjWjFGffhPf8hMaXLQQfszMvz7uqwEN5enItcX/G8qSeQIqvarq7oz1ebzD8zZ+WZuxKUX0OK+Qy2p77liGzwyL1wMcEfEAmbs5axjjXWJQ7+06HbUfsxns1ib/kzhT93TTkldS407rb6ND5VoU4GGr1BqJ/dXxDPRJ9IfBn71yAMBldG69ALrUsy3CYvh5tNaZLRlel2pyI1xULkilHr7DxvbXC6Wvx4GcBVHSrQcPGHgzay3Ey7zgNIYnqdPool100jgIxgSOXNQ0FP043nTNTvAmXLl1msqUNSWFGaNJJUhMpxvi9Ew91BUQHYYQ8bbigZnlcOhWY6ePrEJ6sqs/kSnIXwrcLQHpBzGD6yRhB1+fNfPKYKM2UQ8GgK4C8UpHLx8dg6Xli7CdFFX4afXSZywCd0otqmxBjoPVTBj7btP0lpdgDioHV3Unc2qSJa9igGYvsrUDnHNMbL7gHhxwlmyn5Eth06haN8dFm+NGhynhAqnfGsBLpnP3oE/heeWHQrqShtbD8NAu8G4ZvB54+Bjnn3Z3Ajg+rB2f+k3Xp7dD6CbVBgaHKROBWYoNXvMkvOUKhQcZP93Wf4L7jD9RpWpXRufceMsB6IoKcSFt4h06ET2XMyM0tjUhBsufnZI/cv/2gYj/V5gBplK5eNlxOl7kVgJ6E3M4kzAbQNpv4qpy5/BDnFfCfoCCbCJfyMyfc9tQEWN+QeYB2s7zaZsv1PAfDiK+kaKs0Anl2H1qT6niQnIYzkVu67RPIgzS26OCbXV9Mt2j8RQHUmZtDU7s03NiisloXlvzoAqWw61aTAhG8rV/w//oaZsotzINa6gJTSpWf77Ip6jFOX9q+iEtneKSM5AJZpiVFK+HTSlLzi8g5AYVmZQAM4pQR2Ln7cuRF5pfhp/5jamZL5WRG+eUpqkgy60fPsn3H7bqrOkze6CN0sA/K8RQDZfiGD8FYXnHo+h0OGQzRrk9CpyodYw7qgiu2I9B1BndktN006xX+xr1ecCeu93xZDkl0kOq/f9J2GYEarTjV7q0xGWaXiWOMUoT+Js1q06YbsIiBgnbDxPVTRWivKods8NfeiF9vSkcKOaWivmsiGhrFjjIv1Wva7hJbZ3V20l6MvsTnj4LNx/Ito0vVzNXumIInSSAtxEY5b/cY2Lvwq0CyL3mG2oWBy2w4mmjdrGAJSWVqa26I3mATC55m0K/krjufA1rIJtvSUCDU2tsYGNV94qmK/0T3Ro2rBFHnh9gsWNacdHIS0bSBJIQUPTnRHLT3uf256HhPj74EYAmlRH41d3pk=
`pragma protect end_data_block
`pragma protect digest_block
c58075ab50ac770aa3c9f0aeda40e7b848d6253c4c726e5161158d9d630bc725
`pragma protect end_digest_block
`pragma protect end_protected
