`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
nf6ee+/U0G3A6CuD4VXYuCXGdfBswUHP8dyY4YwPZSAuJKPhZ4ynQrYhyRBFUU4aUd3MAEIfkqSCMRlLN/a5dWWoaNUpgeUba7y7FJ4BzxDu0488+8Ny0HiHw19mLp4TxaSxLigtmRFAxTMEyNjyOdpHGrxSn4hR1Nw9hxg0GqEul1yknts+CKmyb8ZEOq9ZLLYGNyTqPHX3/8XS8T90Ly3u/OCS4s3OpWOSTdzOtVfMkBDYzRBSfJnZ8LBGm2UOdAz7GL35GPZHEkYJLweEEqtlEIh0w+SEYxjnSACFYgFglmcqqbC8Yzy85KkRuzwhzmBw9H85RqyrdlPIJosy5ywjYnaoSJ1gERSTZ4aJtAl+Zu/Klf58f3oBcurGC8QRIQT159E+0q/sZ3aPSHgWrxDp2KuYK9mT/pKe87j6+KARU62bm07rKT0pMPS+8BNPz1raRAuFZDn65OdKejE3xkh9chn0i+6hYuyorRWeFHbDItmnEnvAH3qgBwrG0+K0sKjchXGNWnOwbftfAOeWeZ5pRLJ0v8gPinSoqfwPcX7WfQfEXGh6p1ZR5S3odWUFjUL38dVrlW2xywehxPNUGI1Bfcnuewx7MwubgLo04TZrPay4jZSjQII3lXPGAonlWIIrOVDmLlG7QwCO/lXTfCDx+UORIGW474dLWRAu0czxAhvnvFD01EjE7nCcKl/LLsNKroO/N0cIoFTUWBe8HaYP8gKpuglnDVuQV4eUt6e+ol2GPBphcLb60iHgJGhI+fTzkOKPqF7P/4o5Jpumr4a29HNmcFgSdX8v5TjiukMzMcnlItnUOkCdzzvDdUzpuZKXpLw37THJoqprHGm+8yQxmFLfV3/4T1ZqGA+pGk2aQDbw5P3GFzszs2+8ac9edmsyn+tI/v5zEnawW8nAR/iRnOYkhWsudb3VATDqEpdfRI8iPX4ZUUhCANc1dNZhys59JKQjAm3BD3754CXgJ9sow6uGE2nEWRai5x7lkxnEWVzy0CG84v0p0FXjlaCqmZIABE64lqww6qdWoLw78KwWsyCy2ZpgWpZ3CcO4IQx9u3HBim6ZNaEbstd2Z5R/jVNz1SCO8Y3Z/XRv13YQzQ/PGE2eL5BPE/imHAh7hSJAbTLl6z9dQfNuhLxBRr2zc+e3LE0GjwYQRtQxvdei8Rjab2p/oGrpNowsKY/EBpnSywl85e7BrMaAVdbHJ3q1zMga3v/MtfT8+pMMzsw7IRNM2+3sgcBLE+Wxsp2799zSLBE+Cgzc8wKWj6GFWrvQyCc0irqKLGiT9yVrcm0ZZOIqrPjwSF2s6HSbvR6okGwloWCR3ISKDWbAEZjtndBRU61eKP7rCxgooo/nDqG/6oijuhrv4r3IA+KlWZ6gTFTptRfJfUL7vyowaD6kKYTGivGB6fYfy3EU6t657qW7zzZ8qKANgYnTAHiue9bmaNrh7W5kihNQnM7Ei2lZmUdNS4pp1tbA/VPm5wT88o+yV/jwEfsrOn55qpTzVsjRmZGxIRjnH02hiYrV9WX30asLz0V07maQIoWsCeRNC2abo0cDjFZh8xaVOAHkFOMEqd78HEW9af6Om3A1le8+dYHwG5EWIYoyi/gHcvDj9b75pcQU9KA2T6NrDDsjr8DycdrGovnfH5pbMBfsRFVAh+Ruc+G0SOcWDCFF07z88NJVxV1QYiIPGq41EOibBy75ITlXOVAcjNNaYoTGjRtaj7NTQeQB8ZldX/IqTZcIIVsDaHWRsE+6+MgDeqO1jujCK9tGpo6h8ZMlPbjtW7fqILlGEZMaWSg63SuVlwMPJl0djkPAoKjxMfSF1NU6CSR73DoCfkuqoYVflHQSEBR0eTYx5D9sqat0CMWNb4OXt+tivg5iXHl0RFWRhsVlDQbCF7D/UhEwfqR8dwnjIryVvQ9vzrsCHxyRmF1cYpurhh6GTahZhRq7gQ+zAL1XyPl9yeHO7fSBYFnRgk13IQtY5i75JbLkE1XlOnDWiNbYGz7Q9yT/jDlhfv6+pvg5eLVn9t09VxCek3bOD3qJZDG7XoAirlhqYQeLmwIDetyW4pT7vn2Z+a5SyQkZBREejkzKDY8OrU4PbMbMiTm2CareWQTsLzEHsHwmappJszFwR8L17+a+pn3ZkoMY9cYzXW5ccON2+dpePTxQqD9204x7f/7PC5TKbH7hbtfTe12qutevJ+Z65ifkETFIV8Uu9MNjdyXuunyBCojztL6XC6VHMUNXK+8pNGSagNHm5sM5elpBNDBgqXvFez6qUUAZpWbKDy9YspaltH8STK1GpQLxLa7kqmJOCJvi1KpYUfSSBdrlrCKUi2YCA/6z3/KnlkVoiBUYCLYj53bOffMD/oNjO5/J7tQdBTP8ZnChp0Qe3uZ9xdWE99IC76E+NmLnC7dE4EEjyzBV646Us1S1UM+XOoOjf17AIZMcrBKOh2L4rNsxQF9EqYHozZvSIeS4iw6B1EQCxxPQAuyWPFx9tRRDozeF05Bdwq2nAHEClVlpHf5qczL7hgaNfKNNYiIWyR4EC5k8F78YHkZqv52iSKuMRExt5CkrThTvHQ4RA8UuU9F3Ta/MVkspAop7dBgtwpuhFPNPuJpJbhCMwpWk2nVhKV/9oC8iurClxzjYuNStCa0YDqjaaVvjVQxInt0vhbjKFFK3Xe3ozzWQf67zVyXDcqYGdYO7kVUjejybkV2uxynZPRT5klDcwQKZA/qWGlSM8TEAVBgcJTkdkmtMMsu/k2lJ+zllh22lZE9/zlJetZkZeAcm4M/qDLjszSDzJjWj4jzTboEm/p2u/E1aFIlpt1Vq+JYSU/P5uzLqQlvC195ISCGx6PmHQpyHT/VD+laO5UYOpv7xWESeGbBFoFZAK0slpjfg/CO94iTdxcAe9pyZNiaCwfM90GzXYx8zny9RZPyNKshVUMOMV8+Ad+VNJFroe9mPTIM9FqdkaqswhRFY+EBaXt3pPhA8Fp7Dd01CsE/9VXqiFWc0Ae6YWsyRVBnjSNeCbB0EXP1wKSaN3i2OfZywE2YThHRc+Hb3Dul9rnQx47ScOBYWQ7YMoJSboc5xnduneP8aLTLU30NKkm3xqoEh6UT2dHDZxFzMnfONwxdMn2xzS9TI//6ThvxF2IIXJfNZqlTrhUOPT7/Y1A71yHlWcjFLpcrSWklI+76n0IY6Xm9aMixBhGA/Qp3zYi7Cpii/bFyOUZ0G9hBn02y/VbI3u+q0nQnwOaCL+OJPF+RGuivjUDc9thiHSkcuRnJiE4srp5q2VbYjZbxgAh7/tkOY6s6ByA9lQRr/0rLldmtQu8Ra9u6pr52wMs+A2drkrHZEt6XWgPkOOKBSneRaBQdZl4INdBk3AHVgdk16I7bcQPBBvvRuSlUaH6K7N5qICL6NFTnr+x0yML8LL0X/IBumg98glTRx81tlopg11OKTORDc6v8rVZw17hLc9NL4ajK04hlGdIRCF8/E3biQQsQUGcxXd0ycCeY54ru9Hm1Rc8GpDXe3DxMm+OmwtOU2alfn9CgqBZxT98RN7WTn84au6LP2a7/3rhTcdQ+vCNA8FOkvQ7jnN/yK8fgXRA8siC02mrJAu/8UtG23hFGHT/4+l8j5QjntvRDpiN19Q3jZD+Sx11qiVh4cYhKOIXyHw+FaWcqZm1J7PxZB/FbKOUaenSWc1lWXNwMGL1rtBEch6CjCJCdO66Rl7T5+qGi+AFp/mPb0P6DSF5cB9lD9rfVfIsm2DDcm7Ecv6pPJY/Vg0uaT8hh51xrUmhCSQGEtDvRX22o/bWMTN8Wv/88CC0cxPJxgjXbmuKCEF03jabH2NWPAF8cMmtM28lOIzn4lPzAJij1D39iJmFSY+khQDsOxwMbiU+70hn0SvJ/MpRz1Lb469MtJZ4t6lGSUjKSVc7MWIbdMauHccTbWf7Hl1ezLRXEYMVJ3Izw2uCe/Bg/uYHaDmFsHCRA+ELhXrW2b177rGXa5NnkHiONUwFIuhJmmdrOGmu9vJbHp2kPSfh31d/wFQ24nu4AquZyO191OjFIejrxjDPNA4DijE5neR5YWt19PNiLt1xUysEThk44OymQbVKOJWFFlJhbzmYmu/T/y5zqaJu2vD7jcrLijvNOOtVrPzhlhNxx540S9Rrv0gN3icR9ld1ZhigKg1iY0bq7kwRFj0ARxK0e6jSfDjlfjV123IdTmyocvj64wL2GHyg+Hm0wA1f1IHvM8HV9B7teQEgho+q7x9NmOvuHcuK12p3gG2sCHos8psiHkGIV1d8QoJcoRaNf9J0j8uDz5FuX86iNq/Nn3FIRfXA0a5oysW3eFbAqtvLNJE44/yGJmb7bwB7CzO7PCWado6F3dmQ0K6AZi09mpgVVWU85a6UI6bZjNZd5NideNgGCzBBYBlCjeRxBFY9hGZ17uzOPKKli2/m5GUReDBNg5Z9IOQrUHBJrPxEzVIIZzDldmRIIXdo5zBoXscLlincLXcXOSLmG1MfZUb+Tw93Pd1x80PGNpzAYqcLdXgRnzn8R4UfO/0AQ2mhKy+iGKZh35NceWtMqGgx1GlKFUP373eED9lTlmDHLTmZTl1CZMd/9KJC/KdBKNtqsm2cuFZqC+QSHJWZ7IrANth6UWvWHuHyjYXT/5o2JfH3ui/erzrODOItZvXJVLRrK9WRy6IbwmRPEFCyI9IxXEHsv0povBMZPGyZNi86x94UTKpE/C9IZGn1kJ4JfAXSGU7Z31/0SUkmsgtbtGwg5XG3zqgcjY4A0yt47vVutWApvjHt+a4WadXe7+0Zpidi7K0FjNfKs5R06y9ww2Yt5heEEEzqSNl8lv0dN252fKmgIkxEQVldQOm4eUT6P03gpgSLpR6d/bIdhOuAC7dRQNEPvz+NwxHdjpqYVu/4AWLc2pMZU+hobP59l/+ZF06SEVTNuEIU1S2rOqEZAjnvpxwNVMGadsQ05Me1a5IBlJfO3DMkPM0Zaa/XOASCHN/YUVCWW0PaIcnyK70wK77ZrYVy2i5Z/eL889h1SH8n6KhuGHvhNKExiY0o6CSWZKBC62C5jWesKqpHvK5KJGRLAFPQUm0lOtWcHctkOPB+5UsQPz12tYmDvNY+dkDPsTz14tM7aFSXRBAw9CkvsDd/pG2/O0lrspixZMht0RsHOV+0g3lBJXBq8uhsi7nrY5awsvNBUyD6HpIZ9xoOB1sm6n6un+gyEgWLwJx1wvejUraCJokOyEgNxI+szFBxLd+7+rT9uSBcbnvnp0kwa5X3ZgCSR6Wo/Xqq4oF1H/WBVbnOdVCRfLpajx2KQiJf9Ti2ILLdFZ8iY+6Bj5nAn6nROMe0IH/PRk9ayb8xay404Y2+78dazgJ1kqKuikuxXp2X68pWkQTX9oJBxeTkPHE/3x2yveLy8ABxdHlaF0UsOsFX9qAi7GOx+zDEPDvzXSR6pzY8ee7zUKCrm+Y6xt+w7Uqv9tbmq3v1exR8DML7g4PJyD+NnnJpEYBDTvK9eruisJ0cKfgFt1xMvWj/wwwZKJn5EsX4H5oW/MFao90Uwy+IEiqEMUP0/kwvaYWgAMxarPDQr9dO/8uCXLnisLn0LpSllBUf9qpIjf3Dy5qB+AYusaoIHW43iHwijGzYGhVFpv7VvXmwvc4EIrYuzzIRCs+YXGuwbHEpOxw+0zHyQqDZG5LmYoCnqYi6bYNQJibJHB/gCO/GafZDV+sR7BusDXoCY0g4NU3So2FuKGJDIVRfP9zLKtpmmEaKv+WSV3/Ckpk0vqO2xSfGS4HhxiDFv5wFHpFjMXZDPUGIA9khIsA338HzugqlRghtkPqfC2Cy6/yHWMWRBtSm972jZBdCo11Z/TGoZ3mJ394kuVOO7pNq5e8OoJ6/wqnT4A0hbHZQRke61RTSYK3MPELTGKMMVSfFq65v3vMsidAGMogHrbSRFtE3UQWg0cSHBcVZKDHD1jZ6t4eigY2kuWWxo3eNlyOFtUQjNYV/g6bagnMWm/J2dp8VIf5e+4rlgXv6uL1Fk2tnIV2mbc087WPKQdthEcdPPvSS/VCvtxpeEA60CEAf8hLNnttlmc4DSJVo0DrG1+UckmpquuP8LYt3vpK25Y016tkeips950iuLnY+57METVq8HJj/SXGqwNKJZftKuWLZbz2mUKIj8sbBqulyqdXBDmUAUdpSHcmU2zfsl+jZc/UfMYNCl20RHyW8NCe9nPYOrnxdGS056symiQVbVPmQkjBFW2C+l3rnIZHTxzaoBAgpiMXkhA5BjGPL1kOuJi2pJC5/QmWstt0gAMiV6rE00AeHO/InCsF5O7WmmxEY7sY0AgiYOi8YDTDx9E5tYSHbuxv1+VKh99BBTqhmAMxbvsRgMwOMmMRR+4n771dgJDpHE1m9kIFM/qYwuUTiGaAA8ZEQHHa+4BessDOIW61NDVuXRT0hvrXBIqdn5mrtq5Irj4B1QmciJyz4IHxH6LKtqPKm84YPt3fV1pJcPSIH0MdmOFq7gB6l9atp8qaBF91UC0X1xz1uxpepmrXWErpx0gVgeHeBJPYa6XJDnWP38TC/0TDtFuVFumz3y48RDtx2B6SfT1zzOS0/XBtCJYxmW0sNdLGTBYbouElUFAm77gBZVFaIwC3+YWHcMjLBSK/8rl684I5gKntI1Fj3AhTtfzjsQnEX70HzgqBmVi7TWVfzIsfwjOJcjM+YutCmF83ub9V9C7t97/36HfYqYpF1DQ+qGAt/yEYAR86xmQfzSb4jNac7DzdbbcLf8aE2kCXgmKUdq5K4dYGXneIjRWifkSO6BX00CDBDxb3HGwIDXIIoiklBFqQhShvGKnnyeFG30QveHIheIkuHi+29doYASfg1ndI4mGV+NZ02JV5ereLvfhc0Ri8Lp8/xa/YGhZgu4NToD3olwhSCAzdHM0aLpAduVmY36fW5IPjjZzbYT67gkuwATBaASUVWdQEXqcDzb8xc2K957InM6AJibEENmqJRpdpX+oKloi/ZXFJbGriYiLJfkYiVbFaBaQyOgVXfj4b5u2SecSvqUjzIXkv+NnYTTk7g4CEEh6VOPPy6zHq1ntMUrdoM96swRl+2jDsY0VVSTpUrsi18IueuDnP0ajAWAHWrHD0+MFDAp/Mqp5/wBgbmjp/cxY6S8RF7onLAKRgwceItdSZo2Eadj27y/GcvMBg+d8WdBDohXHeh+ds10WRM6KLC6aNbPROGVKzMpa8yzA6Vog/p+Y+xJNI6ig6C4sAcb0jAnr03JbsPrn1Vs3gJu9cThpvr74AMYAsuZ4tv8lIS7BpH5o/1m7yUKZqHPyF9+6jqhpX4zMcjcB7mriTwgyaOzp0cjFnqOv83MM3ZpYYFht9TfkRfK5avnj7kD+THpNX0Mh7O96tA2OQMeDk5pGr+adah9hUKI1urWeOsW0DZEnBM9rOklz3sO1zFwbMFxVWeXj+fnP9O9t5tOi4GiXPF++9O4lwALOV1V2bGCEggptn4anaw0C3Jn829nLh1iYig56Kd12vAiFGreiiQDV2iSJYr4zDeyH1euIGMXSfE/8VMo5ljiyR/bbJQ6e1WEYcDyUs32dgImrd7pfXWcB+rToyw2IO3k+Rnx9cVZqeMGcrCAAQHcd8kll7SX6cUB+imkpYaihYQ8LEfNXR+VsiMR68X6O+ATJVfEv7/uKIEAiKBrSz9WdZ2f8jq43u0PQek90E1r7wvyKFrBE08vJdToso2jdqj5g8R7lvjiFJIN8wbTj8TDq56CQS3itNS4hD0Fg9mbNlwHSFmGJuzjnh+IaO5s6aMrf4Bc7KXqDEfkgEvDWkxdP8s1Z8wLtZQtfT8HxoHCdtrnKAlI46ae4uqJJlNNbxZ6+AueDb62Xax21liFxtVtBxZzC/npuBqt97EjGu2a3TPJd1VdUlWZJw8ejejDqXEMX2J2aTIHKfZpNxfk0XbLLl3s74rSWLoYA4EiRZyTdxKWxOJYb3hK7HLK6dC1iAXe3pmRqm1s8F6QgLDoq+T6Iw0G9/kN3fJFxbdtGa1NKU5wvJaFPG9uoxayRgE+pk0NlElYLt8VmIx9NhL7w8EkhRgizhPljxZ03caooW3hUQYqXIatMGW2gSyRih8Vmu1rALh17Y2+esoDsLkTR9npFl4YxyI2gqCVO8aF8EotShNI2R6cZUiOPkM93NtmfFMvCssa+eXdQpDywetupixhVYDJJdn9iI/tM2HtBAZWjVqmbFFfYyeFsMw5IdZfnuq6ty1RDuq/evh1i8GDyymqnKYbLnXV3z5Vw4CADDFTCslZPqWxzRwLLGzODud/FF5DAFJLoUpToZzhsQyhhxPHfT6y2z5thDGXym8A8k4RRUPvYeGKTvQktEG6TLab1w5samYPmfJWyYa2sEcZGI/vvSWJNlky4jJvLOSuryt9Y9abxKBru1D2WQ6zKaHggmc62qSBbLgPouNd9S+l+2F7LIRAaHCiQkB7m8WNpilG05HM7z40e30V/Tary6kl6+8BBElQWaF6g96plJCaAy665C0SNu1PBTwz4WERoGmNY8OdS5diJe2AY552L+qFtXQBlXp12vo2vPzgEritr8enNAWbqj6ix/kOVlUf11eQiYUlkMPIh0pcVoDkuQK5pZi81vvNi6/pRdP1s+ASZS4hCIHNcqjhjb8abL7w5BLlh8DI3TWnp+JIr0fpQUxR0SvOEp+Dfz7aJFfSLVEE/UxfPwEfY0TTbiYaoPumtgHF86QbUk5+vUwC15233OVLmWp6MWLAVj9NoIqQtXBPYFc7aGZavZDCgynVz5buCGXT2ldo1XUmgjAEWn/L6urC6xX41k29H7p6C0QIIQ0URiryZA3pxZujcAQVyz6kpmqNrRkZrfauLo594aSk6TikpgdovbP8UDDxAF2hBMdNqNJKOaoDqKrnfOs5ZXIMiH3fZ/fQb+gheDfjInAK5iao4zZ0LDsT1Td15v39RvechU0KLYC5u7kzGS75euPgKuAdqMuptZj5bXVf9otimlrN7k79vEry+r4h7yMpkvjpRLN6et+xRP1kPZCWaujnpPX1JiLPTV8e0F/TKKADeuGaJPHbzrjkrl5rc+mv5EEBonnXGUSW1UUjcZslKFeLf4TcAV7QyMBDTQTcqjWzeS+DFrJU7tFA+wQvOEOQWoipLAgr/gQyj8FOzEC3wvyi4SarhCh2ypYFUdSYWI3QlsRMcK9IvSoAhBhmGjqpeEteDz7TKkU10agazmoV3M3F7LWuV4+a8Q/iooxnhRpKMtr+mHGuYRIiQ822QZ+xW3R3WLUOssTlZZqOcb/VZtm8kvzsawppIIqL8ShHAbLKLTE4zbQa8IHE0ZPTwJ9dL4rj6CgvJJj+Pliwc2lwneIN5FcIffbHgsZHFjGq8rPCETmTnc0QaPWxR8n3Bv283+uIOUVbgrWWqEj9kZm2RMbznH05s0bgDc4YS+RhEEecWPvTGNsgjSk7vt3tE5UqtkdssKchH7UKXcGbgTGf+rxwIhjDSnBD9qH1s32HcM3gKiOE6E+t7+d+e6o9UjQ2CeN37MzJ49DoEhkhGMLTFjWdRcGPzIVbH0W04d13nOTTGPIqvFBxITP2RCeHnUuvz9de5P6Uo3YV3Scq/iCp/I6Q+l9ffDXyXN86EBJzmPpLSMO6tyfLDeKmJTJjzmqIYzFaiULYzsCLLg+bYekVoGHi3dE6z8AQ1AhfPlbfVZnjDSx9myqTtcyUq3c5RPZsQX+KMk9+oSkUKWL4/Pdom4qBlwdRfiE+oAB/vmepU9xRnjgt3AEN5t3UhcAEIRgMazRdUJPA8QDt8vo+aBEEF8DhmkTyzVDz9xjtE1SnHLR+H2z4/GWNDBUUSAz+l8bwNEeo6wzIPRlwbFJVnrdy8fvVYV60K4jA5MDSwtSCkQ9i9Ayg5rXbZlbVjIlIGSMtA1HRpmqb8qGqxbSB9TVpGMP/DYhSDSipueJ9Gqi4CMH+Ann4AjUmYdx/x3szucjxvew2xivS+w40yIB3UO2PIiTKHoFRosbMXczDiJYaUCSvcLVMsoI4IAmQqPTrMwfGx6LckYfPB19cnWcn5Ps54NKR4l64U/Bs7Bxi1kcXvu18HNMcZXFZkCBMsiw5LqAm7cTK6vxr2aPi/Yc7J7BxQZBt8dRlvB2ZO4v9IkuwfitjSv8W1VfiKbvo5dAfbmt52DqPfLWps7ZZFAnBlhIXCyGI4RV6upesTyH8Dz9tMRwrYOwb9lmIkgkwTkzs+pG9+yxm5yEYweW5q1rKpfNGnJB20qbx/YRtWrB3JpGQhjSDjb7lVZ+JekYIOTgQsMszgylFKSVwW2tdEK4/91g7nvEjCx28SUGKOZjHcnD7dMuZHOBNHF7hnxTMRRKPsPpwM52GL9Kskgw+e2PHqvMZpHoFNnAGEftyjmTx5kZDZ1qpEfGEnQqPtQhgYySABr8QATc2o/NkjeAu4C9cwiFEGNEX4HTfiTpAPKzuajYnwIBtTi5S+IncqRYaUny+X7Gh8akXCp2eRy21aUNWBXEV50jITCbJ5Zq6xQjmrqGdW2ZlZN7h+ZNKVkMSqhqBI/LXDxNWypoePvcRhJfYKgzD+zVTabseyuIvUzFxavEtZ7ctDMkXRqArkcweeMc0qJMhcfrdNiXNHO8jQxdb26m+LeaePHfiXuf0fq4KFZ7e2ZdD6UbzvGxiSKKVj0xNKqfo2s2vD+gqfirSvAmsksYog8Wuc2y+my3HaAfDOJTOfi8+eKUiFcZBSDpnJ46l5UI9Dixu0udT13Asu9666XGDXGgIi8DXwHSVWgDvvN3tZu+KTaJyQeXnxjnSWau22eB/PILSmnq0XB2uYnaCSAo6whY0EKbgyJUYJHACN/jvWCD2QScOPIcs4ycuvbToHKVTV87kONEtq646pxKSYlSf5Qc1qYWz6MPoJKeArBn81WHKjEhQFfyW8ioxQWckglpI6DREp5pl1lMsK6FvRuz5FiBaomlVc5luim5ORPRT6UCykTCJL2vkKWU4B9TAifJOh6tupyoKjhvi+WkgldyUdDBHKqdHnzJWJgDg8PMOhorOKM+J4qA1LTwVxtcZTNlDy6qK/goN7eHqNqXooV7eDevtXFSqr837Jfu7ZtMucmuLEIt+3pw+G0g1VtslRKJgWF6DyZgz8vg9+D3m7GlfHWpxcGEFTsSEhgPCg96Qc2zan5KAQott5r1rjSJPn1hPG91GZArGmwIPxLm6Z7TbjvVqo46nL+WysFjdCY22RAYohbpt4Q5Luok8Ct91As41DVvp+sgNn4BoVT1vw2XOpWUjpuvgZbsqaQM467jUxSWBoPbjfpyIxiWgiZGV8sSQHYUlWSO1/qevbh3JfrdcMbpLypzAaVsgwrRG1++ahXJA0LpREnTa+jSTKmBLYiwft3GcCmphIfizD7tOZ7EWZ64KKfuxlckXSIeexsu7MRSi7sKVDi7FOdfDgZo/VTjigksbb6xFZC9X3N0Bb1Pm8Ce9MtvYZJDI+3nNhINxyM5kl5cEnN0EU1eoEwX02k/X8DxaY5ZblsWx8sk4Wwwkgpkuu/Jf2k/kt4KldJyqWsyt0uVxSp3y6uyg8UTgMbWXhGqPpcqtyOLzatrQQYyBR5NJX3xEhVolst6UHKC5RG7GyJOoyN2E79UP1KycDVKYRDaJba4pkFndNwpzQcN9UNEqYGQ3N1lDCb3KfUuOHMQO++NoQLq5O4ZsYcPlhoanFORADAWQQpAXFqJ7vVK4cdGFlTuDz3P8pAnwoAfIAlvIu6DOBGHE5SDu9Ps8Wactx/k67lQFK1TDCiNqquL+BjPBJSNM7ONvipAeFWBH5i4Jaj7JEGWJJ8eubsJ1IKlrpq5Mpwo87ldXG6aofO5IX/dLqGh4kDGl2n7jRWoiySqydQ5CS8KbJHl8LRbBbSKlcgstNNVOQXNUiT6Z3y0q8oKNJ950ulW4vSEdAvH9Av1dSqDm8S8K4xNagF38znkQkt06AFIcDzITX/Rv1QEFJG8ni0ZYqhtXh3EhDZVdcO5p+7ADLIyLC8HrJ6QFKwUrljk/iYp5c5eQJmArudrxkh+aaiXYiEXaTF5oiZO5k2ipUpFdpE3m6z3YnTkZaErvuP9vVAVdQGI9yoE+SbjFKoqLf/6WfB5Kb44RS43dt6Gtg7IZHuJ3mXDnMKbh/4Vnj/pX+5zkBXTYdmsWuzCXRwUlAAN2JYiDKE91fOJ/ir1tEs9dLxHLrJlv28kSfELN/pYDhdZF0Dn90/cFOMzuNpg+cOoUXBJ4NNB5d9MMcTll6uR6f+ncfRpRYmCl+vl/AjGRk/DbFBPn2hoy7oFKgPKcVfgsIN4HZqUBCF3qF4KC82siZzV41zKgnL2MQn/sIJhklmM5uvIxq3WSWaIAo1cJpcOmoI+iOpmg8O5LmZk0FDdVMPPnh/PJYYahqlJn+HRM0a+B8DAjGeAJ52kepPZxslG1FMpopDfIt19NmWaOgbEr3x/D95DI//wdbLKIeDY13knpKR/NFyhlGiejBgUvTTlEwMsiLbFacAGwHzgd5GoXeuaquWnJVD/w3ncSORbyi4aTMWoxb09Kp8jQy8QS/eilFuHUp2ni17yJuQm+ivufmUfQP6CwHO/j8J63Faqjpslb0ofnEH+XBvd32oJpmE6sjrzowvFVk7OMaX5bSx0wS1Y4V+cOby70+ptYWdnCQEAzAYjjO3F2nVR88mjNqd/ozihhokyIDj8iU9EdUL7EkiRtWGc8lr589moyUqo0TBZAyEZz+73ETTb7gu/CEkKZGce2o+Vq0WcjuOW2q380/EB9QDkQaZuTSz73yYedgTzI3BO8wCPvEU+YX29lMJf2fSkTBuk2K9oYMToXS46zBMM/WLO8WwsIiXYHC5o5XTjLcQaV2u7ZIsOqdVy5TXpTz6go3dn9CiqzI1XRlorQdvRqvc1v8wITcLsco5yf3ZaO/qpANLaE/OXd5DxxPrb3IZla6OjCmL//71+bgT5BE38Pvsdln/P2ptBKlHCpdUAgnchT9BgXR1wuFOLkhoYhbpnfovSh5T+7wuLblB7W8/nzzq26hHLvuDqMCMEtR6eufZHqaFBTKr/4Omz8TEo3vv5Z+NRN+jbAX5prj0sUOupnyxAJsjKcFL9Js+S08BehSTrwvbyxxUdG6cN3Jul8pHVdLmhupjvp+NRKlzepNvVIkT+pV+QRzk8nEzXZusQ5VYWjtoc0JH8jMqmCrc29tTCphJkh05RtANEUMfVXOFr4QuPrR/aFnRJ1OWBr36naDxc9lLViYi+w9C+KiQlEX/Pd4iF9iA3uwr2yqJToWil5Z0j+qfxs7E5FiaswUAJ7cgQbTJLSfkfdZ22W5LwJNV/OXSIs/fRZzeY555qXfCVeZgMoyaO1aX8clLeGyItJ9S0GKdKZGZmwNzOfZA1s4PUHLeE9YMrwrpUjp0XnBgjfs1Fd70KhrqtilibxW79Ju0a1GheNLiENOeRiy/6+/k7YSPHSz3q7/T1/6+T0QxkklUTQ/TKJqylYfTp253QSdsmk1qqZMbe/ZdIzwgYNTWt4WuLyU0pfFiqigCLUhaPeB+TPhYfDtbYE5Xmz2Ub0xFSqjZLdP9P1dcTWC/hlf37tRZ5RW3fdBDNE882npvXOnMhxE3NgRkHXKLrGmPvUWUcuAyLALwQAOTZkhhAesxEAKvDpPnqd+5n4z4+90ItIYUzNYhIcw1BlJRjhc8iNUh08O6WY4AZJb71JzLytIJH5o/tl2Db2hk1MKMVq7H1FMr7w+ESfcp6wkjHL3k9Mh5IDe04xwGeAbmX0HbWO9rt3gCILl4xcKHR1unyqBTWIcLMo0BkJ29lmTNBibwtyRIreguGLyMHykgnMzDNoKlc1/HRr93SsT3rdcDcT3sp8ieQ24epgrnCniJhjyG4XtiXxqLt35/F8AzJ9uCJZPzT8i0x9NsQNBkQXZKs3+VSUV7i3+YoOk0fx9advIMJq1vjfjPK/Y2rcSRagFBNZyIMr8E6S6n4mt7QSAHEYiAiuSZgM29yzx0b6YhU9dJX0b/6LKgTboHGl76+UJaSACBE9jM/wF+cE78DCeL+96aQARVJ9cTvPX/n5BcDNDUXpOHBfj8fZRO5NA5liwIMDW2+CJHQH+tkRd4O8j/m4R2h6q+INSbTEDgLB0Psz3+ujEha9Ec4G8hmFint27w4ekxJxIKi00o1PBnNwlj281D8noZnOsbAM3i76xfACcf6Smws8buDJB4CgoYXxnVjuudt7Sro7BzCUokJ/nO3CZQDiUzsfezjsRTr0exnG65ifuX83inS1hCmYjqcpbgZEfpmBkXt1I0boBOmiogV6PNMxPUIOjhWXK7AuFWp2sDFyU+aLZi6yaQ/caT5KqOu8Vad8uhLU9SfYbhfRptAFLbMZn57XeZpWZsIFpXLJDBKuefikZNQ5MC8VGkw9guyhUHcE7j6gbr0I+5o1izn+kn/8QsZE+jCWNAHUDsFJKyAS9coWo9w/MCsPvXXOBf9XJ07MTXow1c4lsrTnjjv26OHjyOUTNR5gKop4y6XIUuE3t/PAwfoXFwvKMjupZkn6xKcF29jJutME5l11ayw9V8zVVXKAuUT9yvjgWPlerz5fTvvWuL9KkxddhnGUcEpyLp4jQ/e70a1vDMFn4bWWC8tSnXHpvKe46J4R0ECHVNEC5ISWVX2XlYqWCFe8l0jTEYOtrPjjZ19zUwU7wDQ06q442XtH0r859CiybhESLKbhRo+C0YGI0ztgYGbd73YfTnlMfeAxEOChFIEnZpm2Q+eoigYRPCzMC5x5LLjUPULjoXarEm6ZuTikje2/kQh052juzUl/HqaMEArA5ohyB+1pVSqBLf+AHu1y7CXcjYJJ39XsQe6T2V3MLv5iUjyd9u27wwRUBdZXNkyle/XtsOB6wljHV2tZtpR4HNaGtWIURSWXmA/atNU/77Vk7R3swcmtvBALET9uO6htAKnWnxwHRvGHkzQ7QBw1byggBmkjvPBE+EmLQmexrldO+Rar/r7t3tFZUTpBivKI1KVilFXuS1ZEkavYvMmUCu8Sj9PcaxpiJ1EQ1fH1hRygZyUxcrWi+SzHTWKZRp0IjhqEFIvZavgEYdP8z5AVxr2kEcRrLn/YKhrQQxvwMAV2lkjZZPzWynGqN95NbBWnubH0g3+hg2aMGeZN+byxokY2chfpy+nQCnmQy8Fz5niAz2x2PyeIweBYRJ73fQkC0SkFP6w0De4LvWGvLW6xU2C+NVyDFkeFUQxY62s3IHFGzb8H0QHXWk72BpiISAlZu68mLLwr8D3BTX7gYvfgFTHRiNQBQ/awIJMl0Xbi2PoJPwmngnYM2fUkyb6DX0ztcvuhOK1ArmWJ6F0XaGbbh12B+CvSAr4MVQNa2Y0XNmUh+1fkPg8AkWaMtXKfjKvIALBmpaHHtuDgS1cdg06EFKGPe5Nbr4K/so3lQaJX8LfjeE8FaUbqog6v15X3D3UAwqkFRV9euPOS1H1OYKc97mBhX/qbAjUeUUXdUTqicVj6/lJNU7Memt4sQEDXm0wav9bbjUNuflePQ7sXLMaJl3aWaU9HveKKApaCDM0qWEcyTglXz+68Z7/stqEEqXzPKNki0E5nW3Hsy7CkfonIn0J8iATX8qj5WzCKT+g09HRXWWVFSjtEnvgzOmkvSawR5h0E2h8RmEo5I9+I++osIULMefUVDB5cp+UwR2Jp6uSSZCq1AlisAijeZJ6L4GD/pwFH1w8qUGXJC3SbJUH691Laqs+09ltd9Ycc3ZkdtS483UDaxu6x76TqE5s7Og7PGIiP9gDQKqTh6ZeyArlklUU84aceU4yaR/vwYjW7/2+N1qjKQS+GlgZq5thRo0wZaxWfs0BNy3YIGga05vpBOHI2IRDc3PkHfMwZ4Typ1ZTLumK6VpNuULbkPjgrBy1z93W12aJbhx/Z5kxWm+8k=
`pragma protect end_data_block
`pragma protect digest_block
2b57faef0035e9f89944cc0e0eeb4e72587dd4d2542d23ff67e60ee72b06deed
`pragma protect end_digest_block
`pragma protect end_protected
