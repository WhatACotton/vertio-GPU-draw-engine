`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
hsHg0f6yNFX+NK4MOMV6V7VOpFywectJf62zbItu7k61C5wGJAVvJPWz/5Vm/lZnkq93bQuGvgUqhJR09c8xUoxuga9V88I6+Pw5UcnQKvi64rRiWKVG9kryJJclBHpv/TzJ03Rh1bBCMaOW0BZ6eTuUC4/mVzKbrqjPQ41hZPPfBzEpCnh9adyhYxjIIwcHGqGCwG6jJn5UpkPqb6GT0+/A696CWHjkVHRHUMzxK23u75+Fw8BwD4OuvM9LsJZtBKXltwWF4ftt+nXXSs+GRc1m09NuI3+y9VSAMXMpdww4feDgnxv9BHZ7Xfy1tXTciwtsh3lSp0mtBW1+Jmy7Mx9PNglwm4P0D7pG87BrNilsDDvvatBS/IUpSc5ZwKbcL9NPSSs03XflWtzfB38TcV/de/cZASj//vEtbe1vW5uKIAoeOhITs6+NTYWsXUi/basHVabXpZ63i+UHI2E7irNTzQiDipNVymnveKJGgZYnMI6PN9pXWEhyD3BqECHhAd16YSjgelz20rucP+y9EWwkw/HAshYX3Uu62Dn0+qn5C4Aq3WM6+NJ6eLjxjSg3wSPTz7DIrsw6tx6HuZzOY375eW3dvWfNdUoXfhKw2MTZPCEu4+lQ03HXKqocNg9M0UigOY3hTns1yOnuGvkEbIgcG7FYb5Ou/TQ3BBojjEoM3y8IVLwhRBoAkGo0qVVKUan30fYd7VJLUwSrjovyGcfcyxk/oTLEgxskZ0UZJaKHnSzI25DHVTQdWY23/KRRRrj5vtF8x5yZ9vmTC5YEPqE04ZT06r9Y60TfnpsbN5/MUexctrPMATiGjsfbjd/SjJDJOF2J5GnLr7DANA0/mhJngtegXU+zP3gc8a+SI1SflP6hMyYxK3Vwq5ROn3LEERqh3UxhhRLj3C5BFocqLPLZlmfFf0rsNk7JeLWQSRAXdxdkaJ4pY2i/27XxF5BtBlB3ic4IxYBk+YDpMPJ8vO6Qzdiwm+hLwFBQbHYdBQifMq7StIfO84q07gG8zzg6n6i/yNMTqCbDKU9mp+j2JSMiKTEe+fzks92pEr9ljzamm2odLGKwsR+Rrd5TH8WYeLTDFwbPMLdGGencqvbGm6prX7LF+OGLY3mvwcPKjOLnMreY1SoOzo84NyOTffTUVKhVgo+FqDjAq/8GnDbVLMCtmVeM90RqGzlBS/Y5jJDpEDApkZ/d03bX/rm9ww40/k6rxxbTBx68XbqQMGUY61RNhArXr6/JR6fA+05kOhEXYdGwsvF4grRzrTA9/7LTqLS7cCL9pRapu5gHdZmOKfGnTlFS9zFvuokAxdekC0WxkrVmzBYUWgnsUMA8BDqMcFE7L0/0HA71dSRT2qCKkoon/HDnqaaJpwcAsIpXThYGn1MX2l7eiQAqOV8feRZuVrPxcvPRQCdHdlSRri5L8ePLpA2KtG5Oygw0UuUwVAhGDLYVRbiPyfz77SuKqfzKL5wLpYiDCPAbb2V3ooSpZD84qcr7HOCH/g253+wGZiUbMS4FIVf/VJDW6+DcM4coPFlsS2OcuZtwd41jBnI4IUS6X6E36yvE17YHrNUlookqa+M9mLaU1HX8knjT0zJwmrcqJdk799O0fxw7Iw/BrAXJS/bVgaVmb0dt02EK4Hq1fb+n38cn4vz4FulS6Sw73rSZfH0PV5cCHMzZZtEevVHWLrNHKhyoUEJe6SgQNgUPEiAt7/2L0VJQ3r+2hq7wz3nVKFIrz8XLIoj0RLyb64hVc92uOu6YHmRur0YGvI6kIy9/8Rx0wqgQuJrMseC6XiBI8InOP9MmXCEG7/aAd2EZs3L2F+rNIqmuEjL4JQ+0qsBMC5v6zmONP7ayq+hxi8oE6a9maFIH7RjoCHXxKNDvzkO7SDu5470SW5TIo7cDqwq+cx4Ci6SqygOzmFkOG3NHPAtHq9RwpgWNwnOUxZjyDMtGNkp+QISEIZm6mXUONDAAVrK8vw+/PJ/Cl2uMEN4BU1FveK01//eVg7IrD7IqMs9bA5YzsPaVDI5CnuoQ7XRRzVRGl9c1gL8+InZZo6fbzqTZnPYWOpKHvcNewUo3aEHHXfWdDc5Dugt3l5ogdNzug/PtDLbJFiwt6b52C2BPOWZ8llfhte2633PYDagAiJ4/stILKXv0aZ5AH622+UoxdsRbg/d6r4y8IR2hOPg5r9NhHa0oadsQhyDRfFEhg5fKN2EaFJxfzWx8oc8gfyPzaJGTH4ojl1ajBIjlivUdd2yEftNcmMOdhAByBZ6e7BBe0idOecJoSD3Kx5BmdlF8AsKsi2Z0H9UXffoYXhWPnsd6ABZnrqi8WxUKRwy2gpr03FDi15rFVUZ6UJlOb1CWrMRVqW65XRL4Y3S8NszhRam8GuFsU9HH3rvQDpYfiUoWQo5C38H/fpjhnhXvLzhSbDWufkNCNIw0BC4QN3TRoBsmJbCEv5WW4m86CYq82njGuQhcz+EYPw1QZ1Z2YXjtt+sZ4eyF1a5DCHD17J0v1EeEjGon7ZGtrCOwvdzYnSp9qrRX+b7DiBn4Az70sWCXxfRndNTnmipzIv70rzSKB2NRdLJqMtEm0PCMGwz/r+h41T4vMghhfk76Of6JFvks0RrtSLZpNfxNoc5t+G7OflgdN6aR/AtiGvv9K0f4rQ4AvtZWqIiBoH5mRZEs8cLQc+JCHz/wf48Gp0/JXyf8OQ6QtvYE6fefhwpGgTNYVM/yKwgWwHNRBPCxTBvU2to7u9MBG7Tj+VA6ZRtJ+2ZGlAtmfiaEjYu426fAnHZdyrMrSEgN4Ovj/CzUHgK7fpHIUWLevWJP/Xdl8pSCNrR/c0k2sLsjEjSfwdI+I3/bepytN2ZPz1YXIduR9nKDJB/tD7z1xrCVUfgW14r3zYMzrcMdiU4U6heQHCRxy2JvQuI+/q4w3ypLCwrX3lFw25UGOjH1f6Vyucnr6lS59IQJ6aYcPW/uhl4/1VkXQNuKeMma5YHnlNdrvgeTArEoVI/gAQQxkhL1NdoQ9OTmtCtwg+TJlOInOEh/c59A+QUImiuuR/5t4FpmzyW716MiMYR+vNdSOuHQgNAYhtEf+kXZhHNAx80VaymTYl6vnUHTvyroI/beMPy43088iqZZTfwuD9H34bkDh8YvUkYzombSNyBQvu/16IlrGNAc4s/dUS3gBzG04CFONUyoF4eC1UgC9MCctOJSPlK4Q+96uhNTiBZ5l47CHTmlKXZpRKtlKDgFTbL02m0MfPdX9fh7l0DKWGpjk/J3Wd6crXkW5Pr1YlP0nCiTdhYi7DUDG8k8By54WnnMqwWYXDMUKEv6o+3w1vqjrtU62EbdMqAeMsyRAs4DB1gVPjIYiPpiDYhxYnC1Rpc0vTBMOnkqFjBiUbNU9n1qWbMuKyt35jn1ZGx52YcNc3TAx9BibhUlBmSahR+Y+hsq6Jr9/fZZ9i49yXQQiPWjMV8ws+gXASqD/nXXW0I4vxfigrcs8+enJfeb1ImozfSfpoc5oqi0MZK6QsHI3CEUUn3qwc6HqKtR1xupCKLLpr456PC1NruN8JdCck0u+LBBmEx99fEMjUMOiE8FJRWGwXHkuISfls9wDxKTNJ8xSYCbenwKL/Oh0eTcpEX7i1SnU/yliDzTKneVrE21cXhfBSydY8r1z1Qy178mgj8qyFz8d3u+o/zBg5yf86xl9wghJpMWxV7VOhPt7RzJeWykd/3B1pWttKRuY3PSGds8cgsJ/5uQ5n0QKR8NoIJKRG2CyulLeJHAcgPDkm40De/3SwVIMTYsrwzMQ/xwRXaai9KzhSWDLIDrMEAzQrGHPu2ssh2zHx3BsZCndJp9On7YMQxiIx7bB0u+2AczmTx2RtS6ukDYJxSmqR+PsdQfQOuWLH8mAW65XvRmz3r9yrGuCdelLwYP2M2cNJK6RDVAbc6uxo3Lk/b+Gu7LMqQ94EI3PHIxZKsqQYw7WA/HwgsVgXu1pFhyOVJWv7e5Tt6VGyI95UVmbS1hRilBH0c8I47VEiH4o6a90vNrsAO1T5OnOxdEossqvSEioiv0kCgVVBUlULPeKXFl7ouObsKihdRlma3cihYiZCQk1O9A4FBEtGV09Oj7ULM1KisX55fBkIBq2mpdyWOz96pqi/dWlbR3j5DEl/RDTtRhqo4KwoWPR+k15Yep248RahwDncpVU9wga5HP3z7GsZ1u7PPkssxGHbLgOsj4V6r21bJDhq6C3uXkm5ZtoUyvm3YLKdgf/vAZBqKumLJ/TTwJtT2U1IzKc3AoyNXO67MRgBf0mLmSqf3CKwTcVX0ZGTUt2zsKMK1N74ejHcPpIbIHsiAv1Dk69BRjGCW9N/Tw8nG4teuBdLnAZ1rc2SDlwT92xNdhhFzgtTbdHr5CtqSWI+kpXDp3maXGTGYKoq6SuMInN8zqTc8x+WpBeTv7erQU5aLclpoxovxSDmW5VAsBcPOucUFLvDFW9nY0s2RISMQf9pc2dcWgKV5EPbRNcwjBRKHLGhxfyATPn4MEwmZkxzuoRh8q1JPgWtoLMiJs0BbHQ6OsodlvziSl7tof8g5vyLUn/dlnrFOVh2kw93PRJcdOw5prxvW3qa+KXJFW5jPQH6EmSU0IuhX8m8SjID4I3OWz0NTfDkYSO2xuJ5Gu5eliLKB49mzEZUwxEOL++XlY8WDP8PAmoaPv7lQoXQvb2Bi7rVbF72ynn70BWkT9oft+9Vu1DmPNpXNGIMez/mXkGwH1513bjsuwatpQgu8OhmLbLXpLWz0M0L6ja6QKR208WdnSRTQn/BWpCj36+eNPPfuANyOyyuabpXWaAjvIVRI+AUWWJqIALXPwXvV/tfCwvopClZjSvRAKcUjEsRU/69YaiIj3pyWZzs8bgCb1SBmGiz1nPHoBJ3d63TaaM8n8PyLysemfdmoEThMEuQk5RSe+XiZxOfSs0ZLIBS5ZbE5JW3EjEuqRkoDxnZvnq/DfT1iX6C+icXGxDs4b0XMELLBJAYiNXz7bpX8K6b+RNAJBK+jcB1pHQiyvyyaL91Gkhs91PLRZ1cTy8sJqcNTkjHuKKXhO2Sd849unUcWS78N4Ipi6aRRS6YwJqFEPfXXlXFwIyyDYrNZllhIa/mb7dFsIdf6sbA+uFHn/i45PR98B7J/iFYjdLq/LtyX5xmudLB8SZmMqvKX9CGJwhzww+0iYQFy3GbSDXF7t0fcwFg0lDghuRar1qOyg9rG+Eg7vcPGWd/Vto0GgJk0aQtBVmd2rD4CIlGtzZ8Spn8gsOgNazaQbExir6rM5Bc1aSGMMY/1XaUsd1TLiYLJj8jbq27v6PdPCxOE5+xHdIp9tPPQpcIwLMjhh1r4Ii0VPCXQFkHQPwUVImuBNH4ovlBLrZHaCwTCKY7BtTIsWeRn8rjJtv4MrId6bDvedt1K4vRczKRExzOYSkkmMasDag6eqEvgj2ifH27RLwoIpp/LgEKzjmLKoY+tCQk/tF/AuvisrZqruBMMU66zQBXEs2Iz9vJLFsxCHsOu0c+TgroXaCEItvVO/PjyDFOX2u7Mg5X/fdGB7fe4RVksdaJc19oCiEwV6ZYmjyNtVyD97tRayzOUC+/cG5KotPB+0VL6O+2uEbfwVtz5Ci9a6L0u+dbqMELb4DPsJGBRQoRg1QVm9qCPtW2JRX1CYD99YWRZvkStTKWlm9YXkpZSogiGmxDCJXHpxLMpbLFfq/RiPD6F5IXUmhdC814tApVsH86EJu6BKt1EQKPr2pj6Q7eC1tOqxuz3wWW/pGWlhT92BQ3ntk+7V2guhGotF1lln+ZwUaLsEMkTe5ogUiDrp6A5Tnjy6dEgLTwW999hfayzfJCjsqIPe6tvyqYD3YTch9XmBNPkyJN0YBGj44lCpaqMjWrO+pihkJoDyaDjqn5RJo4hxX0eotwfAhVtxI/RVux9lTmt1EVmi6HeiaqBCz4une9v5mcZQe96xUxQ/F+BIPECLohFia1asdSeBGf/HdRSvE25R1VEGGbTlXotMhQSed94KN6iu8o0n7D46/O5iR5cSWhtLaZmBdNJreC0Q1Ce8/bNrKtKRx+jA8crGgRV7FvmurYApIWvIQbn8YOz9AYNkmKPRQK3d4P/L2luZ2Cvf8jGdvR1YiZBWn6Di5DwM7Vxnfk7jzgloCgyMlEhzETOiSH4IGJeiinvnbos++kEHeIlMFTi5Jjg7CXYHMbPLDQkTPIolK6Wem4SyaXafvNxnMqRI6HMw5ekvfQRT2hk9r7aOZAIwxAkrYbByeEarmUNBGsfm3SoWHUHNQtNGOlJlTfcMT5YfLzg4kyZeA0tnuwRsidah4OVFV7Wb1Mgxtcc7OdHcyppU3o//WSxy/KK/oc6Y60SQZ+6wqHx8UarC+HHWQYgjLZHbnuibD3WR7sqbY35mF6eNjP8aZFKGQVE0xaToJOOn1ifjeG3tFI2ilLTFkFjsy4cw34iCNywiq9g3P+U+WO9hOsVUmilZYH+S4hNJpFdEU2kOe0OWwTc01Q852c0OvFcJVbRXixnAa8cNCEMnQSX/euapEtN8Ycr3cTFy/HHfv+M+ZmYKTRgnkx7HkaXz/7wa1UW1O0WDs7k0zLi+/1xTvkW8nWSy0EMaYVepslrxXMbN2dnz6M2T6k7xfwfmzZV+nhG9i9uxivIXoxxjSDBG1wPrMJzod3c8ZW9gwvN0hBQOCUxabJIbTMmQhddmVJIjcCp3UkZSvwoUsh5kr7P0F1/fjomUTQgMXIClmYuzvPzIsYmWnSe9gz0uZ+tBKSXyNDECHHAqNPnSz0b9+tp44w6rT97LMTOKrzyCKbk7sZnPtS3iuCXCdi9Rr0h5TiE9wt3Xx3PatueXGWljIaNcf3WWPvKCcVufsDmvglaZgdYM1RkvCpWMRLb4DXRGTmkREHePWWIaL/ToPZUarRqJujLDd6x++bAwX0LhB0I20Ri9qBCstQZD28B20Q3KvgLSIBzpEvfI57zeiIMB62B4OJfVdWreQj7/JPeWjfXl6o0CJ4Ci+89Q0EbX1og70Jull7NCRraOUdKTc9LJgYUtA74AdU0XuTJyhA99hC5Et5IuolXqsYbYWCnlsZi7PX1U8hiy00WjSE1pw3Sa6W9FBYeq/JKXzoWybaYXO7Vq44UKpX47WZ1mO+KxQ4BGNCSZ0cDEjOPayZ1KMBOsP40iEVtdNgpys4ySEEbG/YLBh4d93L3gjSMX0joVApC94rquXvwWK69ichOgGrWLGtsfickO2BmZly5ryAlFVeSLWZ6GjDp7QS4OMpQ1HoP54OpQL5wuyIIMHjDI1OlSI+VJMxuAIpJ/5DAn/Xja4NLeq01m2JgNv4XZN+iPj9KTQ3Rxocfst1tA7xzpRrIjqo4yhcxe8JGQBDGOJbJN1BrYSnLn8DGwCoKoGzRQ0cO1rTKPZDwXuV/lHMJVLyFmvgk8wUaR2UPS3Mrmwx5kU6VIJ5Ky01skUqBcVlfKHi1Ay/WYB3gg/+q/AniW4gTTdlNBX1g1eiiv84FFU8DB5aMN052p5f5zLUcIGQ2AO3X/pvU06IsOa6CXJL6fGRFR5/B+fHq9tgh5BJ0v8zO68zRtoemTCzTOB2garv0RKNMKBbDl+wlvO/qQiQcIGqimcks72DEipQbQSrhU5GTFEnwe3Dx8LMGs0X0YCceUCOX9uc4vdXap0ZzpOV95kZSDQmGAxlNGFZx58ToCU66NiwlSi/cAxTYfWAUQjUGHrXPA/Xh1a6myn+RiWFALWSbW311Qxvncyq2ka+KuRBOk9IqBrGP+v3xejjAIP+kSHH6oLexy6BmcujIM+hWyZzYJMf8CnNKWN7eezCTzmyxzjvMCkGB3n7whhNud6BnQPUoEmKuPYeeg3rEpSXxE2rewQqJrbt5cNDlELbw7WVOKlNxQcEMx18kYG9fLdgtUMkOaZC/EGKlZ9uVi/CFPQPSo1/dPcWA43QtAPU6oxiNDcCKl8lvnJQC54LYGfz4e/AhY0KD1Qg3wsSQfgkeeyWsdqxrlBnkJ1KQCcfSBaarXHBhSE1NDjE9fAjVD8NeupTk/8vDpBRLNR4qi9S+Prj0SiYtBl4XFessQnVniOsKiMagAz24qpq/0azxbE1Etvuiofm8UTwVJbTPR6ANqxXMG5md2WBgv/r9lQHBtqW910i4Rn6v+BjNQI70w9KUuiyt+tZGnOcSc6vuyD6f1MPSa9rF3TsKsS93sz/wQnY1bG+D2sFBVNO03jw6/Rwauj66tWyixo6XUMY8q3R5pTQymZ3OVg+zj0zXOxK4shqlz7ZBW5AyYIAB/qpmjYq2xOvodaThsfnl/+zFH2xfzFpN3nnJh6PklU8Y/YGSxJJilxF+1GCMDV/FUwdp53zPdYLlIG5bUOD/owvcesEnReWAUaQ9YYNXAZfslgbtOyruQX6ybatnfVNTROVAuRB/sABigHFwkOtq4nK6V5toJvPWH/0hDNAK10J6amfZJ924rQE+KqWNf3WkK1dsJA2YUm3hG25fsidVDpAl7j2TXuvud5RgqkbDd29dTEcXIJT1unjkBUli4RigrCxPnCJjXVPAL8+dypTKg0IfgeofO77i7NytQl0h0lhE0Ib4HGhNGMx7d2AdkEpJbgUOJpNIyXRP/4VBkCq9/l34Lrsf0MJHIW6TzPiqWE51VC7Pn/Ve7DSE9bnuGUsbVj9upWyeFog6JEDF5Wtur0X7QE2LGYPrgSAr9i/yzahsk7Jk3RECWQRX5sJL4QohUSW+pq0UpDghq0BAL7kSB+c969cGejWAHUu4ljDuJLaq91SgmbKWtPQ0UlcYV5rCeHhfBaFQpgEtR9vkXQZeH6NM+5P9pWGqyRrRTr3FhbeFNZZJ8IjAryoEXYVJ9HScnz/h+wxyIHJIB0hxTDCq75fTressx37ZhHOai3N9jzbmBnZnGLI4hr175hJfPlf3CjFj2QgNYqelzpjcYi9qPs7udEgXYTORN+Dz3AycVi1NOwW9N3Vobngasx4xLNdNona1lBEJQETvc43u4klQ5ap816zzqAUfv/6iQhphr9PJYBaRdM/x/Z2tQiWv30cgxl3sE9FoWVoJ3G/U0fAq3W2DUi492UENXZHnlptC/+wTXBA8mXGruDbZXX2lx5DLS3xs4ty9pNw8cOAo+ko88g+TvgPq7OTBMwpnBh8xjs6Zo6rCNYNKDYpc12jXy2TlyQIqKaglBnVaZEmGAKPBrJ87ZlU4kS6AS2eB/Zk7Mra2qRQhItJfzsAFgXzQagxf9Ex2Z46wr/byGbZfF6MmRoCZYcGLT3HRB9+MeJHrFh5TFnlL9JWCDDUYZwcJIYvxMK94tt3YyYvMI+rhO61YbC+30m5RqMl8iU6m/h+23MPaLcOVOM/mmXVv7gYLD/XMAimF6f1RSmgmdFQ1+9TfWWSFTPHLFujoRMGtgzz4oZJHIG8rFXXACSW3/i1My/PStBQ0ewYMJNfqJXwj6N6A3vjUCS3MGcQiwIjQvgSVy1pyfjZ728h91/iXouIxWrNjWKMIv/9EhjETdX50zHILf27HXteA2REoyaslsOONlUu3lWSQJaAtOgUZgutVxg+v9Rs3Z7kbgkfoiPu4hLgPwr6tmAJICSlvkhXAmCPQ2470TZXOQNxt8pDgBnBQOxK37bzfm3/nwoS9weR1D+XreIRwZrp3zwlZFfIbwefun3QPyog63j0K4qGnP093Ttbz78S8YFIJKgv1LJoBuf8P9NALmT+jitY3oDOJ/h9/xhtJA9w2+eQLtAZKyeAEzNk8PbOJmme2cIWv24MoC1L1ajREyQ6zHrOL/J1z+Ld0qeLy4e265Nqt9Tbf5s8O5BSVct0uJGjlBpHweeDtGO4EuSkpD+qh9XQFA/ym/WOjn9GSLLj87+MtmQhLvheRI7EFaPMXAr0AgV+QHmMF7jF9pAv8Tq8/1ex+fXEKKzxr7tCoJnPP3b1JJxhz/7mfzKtPfJSPOgRP1FdCTKZ8GUgfpBFsSyrEH7BSL7xsQmrZGquW8wv3ktnK5wwFq1Vgf58OtQaEelbIrlBvZdD03dRLw15hNirSsetAtpAoRnyonQHTopXzrYEm5cDFsa6KNumda5hR2Mf3iYfyfBZYe40KBJpo3SWPP/x+DpB12WjRIsB8x2SwbbLTXbo/Mbo/lR6w5mBKFDqN3WdH0Qh5nZNT+78EyAdoblZG7thG0vK2WbIjXZNmWvBzgXLf5my3cL7c1cIKr2yUn4UjNJ1L5VxTfNvggq9D5AqUDrDVthu6YgO0IeNdien0TZmH8KxghJSndyqlbBoEGee2ajNS8xp/YQZFWfYcABrFi57Ifzn8s3cPvMo3K1TYlccv4vcxBAYrFnFh/7PP7yR2+Jr4wPs9QaxUZp5vd7H+deEsh9VQRsJAsLtzGUjAqpJ39MofwP8/NOtDR+grpig50EsaF7eJ/8h9FEZ9xKZYFPcBXClNDTRpCPZSkYugNWVTDr+4VizNmJUPX606nPthnmOUSHP+IokFM3c293LuAL3RLbgXLS3ItX0/8jTZ3spooxaKHTY+0uRnPOiildIoTgieAqlNHqWxn+tQ+XoFomn97uzshnPun1PrAsOOuL+ZvdB6LbovmRlFqWTE9XewRazPjXswub7670pzDlvoO9e2bXxxsqEVqghQcU0RArbtHE1TPE9qvkVUWBNpTc+mGOUqp9LB4ZXe6oioXmV8vlr+8t/KWT4G23o2mgpcCq4zqXmZ6drfwm4KVC1bSZROHgPkXy4PxO0/Tx3YQRmBttMQ0z3i7alpHbvlLGdodkeAyEF0XoeGAW+jv0J7YRKWCMoIdTBksB+W2P9isSvF2px61svXBIA4LDQbVG5gqZgR4fOrCPmEBJuYMoHvtm3LwLvZCTRea7d1ArGKhG91+X0EXnLor21WDQqlTy/it6NtfxpjLm+HQuDkeS7Z6D6jNhyMsPOx7xpV4vYNOI6/ZE6WUCpH6gx1fEWiHcTmpOPvIg/c+eyRhoBIlSysk/R7c9+85H2po0m3fqnn1x7pF5wnhw0iHnm5NLj3P+U4Wrkkr5APJwlU5vMGZ3ZcaWf5jK4vGpC7b/HA4UKTVvteWlv6wTmBZQiRstpS+aJch9Dqllf+V/zVlx3HZf/iPoCYRH8aiUSHaNmVWvvqOEs4lVjbX21HLjMPMDDB3cG0FeXnx0raECHdHKuHL6eo0/2ORf0/+lpITv0tPZoydlZ4/6ZCGjxw867LODz1B+WY6fEC2005t03VF03OTMPNMTtEmIjYWDGALbWO/isk9R6Jk9YE68YQ3kpi6axTcJarkyzfDY+4Vn1nEdxXZtL27d0P3BPxDK7jWSF14S6h/E3EXyX4C1BhYSq0RspxB3k2n1qe9S4poGaAfY6zDATYZQ/ea7Q94cmSGufqukJNzgRcCswJfb9j+a6xt49Lndu4TEB6+5VOK/matB4Kdh/XNnXwGSboov9FGtD/Z4jQ4VEuX097ue7TgSuceVr3JFgCYXFWhG6HzBWX2sluZobIhP6vKLLEb5hWeVGunpu/HtAb1eB2XaFQ0AvGTG5iWCedu7IUfFHDUHPOgv+zTPLKCdbQ6S0fS5OdpzQ4RhYEVWQB1R4PZY79XX++cu4rFVEtJr0cZvkyioderblOmXcJ4ZCo8Ikz2tsr/4yEgzhWoWc0OQeP2vvc2VGoFSag0dEUcAnPjSZvUtC2CTTFwmR9nnRwWnN66jQ0DqZnh4FjpBtZFZrQFyBMit1v1v+sBXIAPyzWhBJEtKcYKV88osil6HkIiv0MK/SrBiejSSluxqwaDpPY+Fd+VLzqSCz7nyNW3piITcpdg4Pdy78kPDncTXgc4ojzCd3ATouRPl8fmS0Noz4wz7CeYV9GvHZ4i6Qq2jlk4N6U82zWVjaIlod3B8rX5E3aw6x7xHddKztGXeJp7494kQXGnqkoUypH9a4OqUqV0N6jEgtnWGNTT9G9MhJwVaz03MAKSGaUR4VmaKbx37pbIOPSOlp8HqM84FSSkgBRLc1RWBIp2ub0z4z08LauQzu809QV26tOOvILqBj6DZyUcSdOzBUFIBrE6UDoM1QvbHxSq3jMOWKOd5hapJZEI69krG4SDxtJB552jcscETqebBq1BH6UQR4qOQnMI8GR0p4t1IG7IyJMsPv7tNRPSd+0OaE3qJPvhHrg1ARP0/phwI+ua/YhbpXi3169EoHZcDI9X2GUH87uQJVsXwvWDxQAZ9b28QekTSSQKSx+FbnGTdmVQFPcS4pKp67RX4qIpveCetNcNso1Ef0oOZW151NqhN7Lnr65OMAeuePEKK3txqbfvC7tGyBfWR0Kr20bmHC4kMO6D6hgWyais6BolToB+F/UenfogXcCCsFlr6LSikorboPdlhqTsaY+91MxWlefdYble+9hb6RPqLWzMxX5a2nkNN5hHI1ox3JxVO2aqmBLabUautG0DId/iwZ6U3Embxxj9Ed/C6vxIfVFhD9IqV6hwiSRfa32j0gCKlWqhQBmbjpb/7+s3o6i9AYjfeU/A9RMzUo+CUm6z+3vZYK6WJQMhlL9YlrhDPA/2jDx1T0VwJoDcMdbHU3KhEfBK9PDjbpwHFTYLFLtBlPw/mLPRliIj0tiX88xevXr5Y+DCeBE/TZe2A4NO8qXq9sIgI3r/kP1RqTEcckU7rQcfbSZZNSNVwPvLRbG/psP4RHIxVlmETUe03XDDq0QRBvCkwMwE6mdne+H5vxIF0Fqe235x+UqpKUE2nUdgQ6vs/psc3dcbwjauJYPt2b+YDWuMVWwoyI04gm3Qc7wc3EGFMkyaWxc0gI+6pyrZbsKkTrs366b04wjrDxFdM4BVxL33UqOt3tKr/I1RxRv2crLzQ44ZE9V2jaYlVQVzqlpglkgkx6duI8LHoJzNi8jABCMKy5dAH3BwEw3JlK+iHayHVUbHsGoXNut1/DoQzn2HeYWYx0ogrEQ6PBRaJesP5F9wXeXvugmkJP5c52FPktAMhEfFlZKatVYKRkbF5/8N2Fcy8Dz6aKknveXC7dsQJB6PnGHyzj0snP01K9Fw8XBUVqyPVDjnLe0FYF8rjaSukg9V8MK1rTm1bZ30emb+rxFweqj4jDgv9UW1r/McvikFWt+fWnv3tI3ydOkntMPHnK8WnVan0mdE5OSk4x1RCoW8ndDSl2QTqFZgYn89hSVPKqKqzwZ2hA1XkJxaoHAEpgZ2nqqYkEHZAzo0HwwZgjeoSqjlA5ZGYVNSNKyuHuNBMLwkoKk+gG71MA2slUUPAJJZ7CacdUopC5mai0t7fCtW5DzcX096mX4M/JI4NZVA2DVsyuK1w1eWIcA5a6KGRl0Xm7zrMkxrYQEhVcd1RPjJPpSShMqiP2+jwoldIeP9W36P619O7i/GP45H6XjfZEHeD8CvyzgjfoJGOHmcXVvun8ZVnKuo77DALrKUFpBoqM5IUb10J6d518CVawP4/lssReAZ8plFjJiBaZnbWuDfs0U0hAonqAUT3mapKA/NRWxvazlPpMEQZZRVpz/e4unWwx/ywO5ltjetDIadb+J0hlVJzeIDcbkhngtGM0Mr4hTDqdsVyM76oRAzs4F9LETGqK+eqfhV5pXbu5MMBlsSqwPH16M1fpwUkeyo7oNoqwFmoP2HpyY5lx6WrYKHvjFRqSeXzVW4aLyRPVCzXu8xEQB4GQrOpQUXvgLkvMa1DihvD6Icn86u/ulCJFl6T80pngQowl6+hx2qfEyrYO77R06jybHKsMeaV7etvtnqW4jNwgJfjKYNt7ecr/Uw1v7USh4zQus6r1Kbw8NexTXIEZsbnjF8XimTyIRt76dmb1i5Kc7DeI/FdHNgUaDutG+CaMKY5UEPXup9/XP5PXSe3Cbk7aW4Q2YjfkRESwwqH8eR6IAVLsrsmJuaHmgKEfIUr9/GLylnX+7GDEouYcyzbXeZ6E3C0VYWUrCoy2odAWpHRunvMYZRwGGKznQeazxgmb0yKGvHtK7cWAU7dxYUGpcgUYkfafIVE7/wJY2pQyszsPJWe4y0PUPBW0TBMh2C6z8biSJBJ+fqF/WqxhNMkstCyIABX9rrCA47dr8n+7lAy0/AsDbsMSb5yQVwGTpADywC9Ro+pw4meOS3xwk+a54n8Dfg+zLE7FGVpZitV3b8HH5/8FLdmEPwGN3+hduYa7ox/74B6v/JbAwzLeFx4R9+37e744QiJswC41SGF5A1KTJhRhjrCa1x5YM1Lne8dnR67Q10uXbLkjdilRjKY14aupK51xw1APD1GHSdeovsRz6mWZXdlJ7Ks0lC0SrUidJ/rpyXSTa2APRitUo5pWAGZyYNn40vU6WuFlJ66Bu0fHjycJ8FewozRmYyJE8gZBeuvyyl7C7KKcG2tMc6Wzb4PCJc9uRwWzb84GrSGblE1/uA2T/COX8wcvKny6awdFYsRU7xOq2zvZJN8ts80e92vMGGIiHXYN9TALqIuXhGAjsx+z892/WhStVWYcRuSBJQGQtDwguKvapmiu6cXQZLn6J6KUVJT1OO7tY9VuHow7vFgJktMMVqNZkdEHctrUSV0FT+X5O0414ckv79SBXoQnd555xrX6U2g0AZDjXo3Z6cf4h20eaBNUzGIqKuYVP7paUz5QBIZx5kjO+/do2eRNKl+u9JcZ8pCRNz5x+3jXqLlQpb280nnGpzi31mpvLs8Jw1+fa4mXKrDMACvnvQiKxXx3wGwavCuhqMpM/NM/6FgKHZ67D5UDD2ODhs04GBGJrxB40L+jc4GD/YhffBaoVFrXw2WNssRx2D5rhNRU6gGdqlyPcofNZpsGzUPYeMcgevhj6J6BEDvxDdPOtgf+8dOF2GAObKw8cbYaXoakRP0B7R3Ae/uuaal3++2RRSSW2gFYevWNIjSKvyIYKmRewHTg3c0SHJssdeSJfPDooBW1zE0QfRAdhcxKBzx719m/Zsg9CyTsPODEYLDgtJ2ktZ1csUf5xyNUOnFopLCIdENNBn3aTBN2U0tYc1MN1gX9YkFcTnCmzhro0IX419oTSTIh9FK74okM6bhrWPeTNoTvlJK+jQBlcJUeBqKEej8kRFkVvidWHXDTrdm8QpgjW/EXzQYbA+5inS+6snYIqNpnoMf8U73OmONNzsVc134Wn8jf9AWVlwnmqiWXaLkIxnSg==
`pragma protect end_data_block
`pragma protect digest_block
5834dd2f969c0b416d5824f3434ec06697a8553e721782b3da9748579b0b6b31
`pragma protect end_digest_block
`pragma protect end_protected
