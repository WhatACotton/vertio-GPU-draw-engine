`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
ZcDCCHIlFlAZ35+ekJ1BwaC4fDsEva2KdQaB9kCeO41cd46qWCIdQZrZr/rIobglQFX/cHWBJoIjFQ3bVJXu6ZqyGGN8DpAslPiiRCKwHwndxxeVlHLY29J2wd6BQZZOCKftrV+PDMMmklNOh9zDYKeRTdysvwzlzT/z/axlI+Li24kuVAR4Q25txiSGrAkk/DyZLjEoWC2vMi3PK6yXEVYuYPQa1fU0UwbCd/fhKQ4irCnSwQ993hupmUOBgc0O2htz0OGi8AV5XbscmetRQTUHSfXGQEF8dZ63/K13glD5SbDIA5pXhW7OARERVxagtzMRt81Or0cFA4YdNMDTOzDjcOYgs8fUWJCnc+RBhz6lxzNyIfoRI0DxreGS6rAysNQZrwhNUcncloLNIE3YqJPlCba917eHKd63gJoTlyujH/QIrzbZJrOQtbOUGMlWjWYG6YaSthc9a9+A0/Y7E2lhFaCTRrS+kuVFjvwnwO+TwPEpaNOailj1GgiubghwWBXdlitPWpOhX7/xq0m85qe2gNSOtCZuWc+viNpWG6BULWe8K4LuANOEGXKbX6iWPrXkVdixYXE+ywnvsjm2WTVuj+lobQZ1nuix2KY18SmnOwW6GIZw8mJNz/5sLMSPwXQgN9MpXdSBVpc397G1LWaiabCLHuhLoF3rfWfm0HuFWfy7ksuWP8JMAg6L2KRQa2c4tA9wNDHzBVnn7XQqFFdDFn1yQk5Pnf0n2nzD8I6U06H6omtHGJGgi6H82HSN5bWaNbNq5UqkwehN1DVJys35//oPpVV6n44U6Hxs7ZeU3XYXd3eRegIlBPfDi4xveRgNnVg3B+sZDWiM2Xg0KtngNcXANSjbCS5r0EmBo7umwZXlbxTmNPez46jwgKRrD/sZJwLsCU+xt0QQe9UVxJbHxIc/vR8YL3Lp78k3aRXbc2RFwc9vp+EWPfJdXLJq4ZOh4VPZM2F7bB+tgI/XVRh/7PYusqTHhhBKdxbxvjjUJZd8zp3wIr8nSs3E1BB8mvdsx9drEelqZLXsQ7IdXeblKh1OaDL3PNJdLYyTeAA4lFGBO2f43G1/T4LwU69GsAV9gFmFDYXQPRoFHOXop92Mqbc/QrzoTQBhzG4m9fGbjE4SlaKrWGMNrymAMayIq8CuEBfp3/nU6OTuTXuISZ55mk/Nv7UkDKAL8viTDHlCsrd6zpnXrf5CeAgY381EjxXXumdWVNn0z51msqAoGWpHs6ZbrTUth/evo9EESSw83L4ZRT8+OM+RsQTkpcUY4BCX2CRxm3/9XSMTxtTTu+KCMPpU0KPQaJCQNM37Ck5RmrLiokOGeJA6bLKE3120oOBtWny4nyr5Am7Z/mT+WxBBC5SOLIGDiEG5gmb7QbbhqirjLBdBpiDpipQX9A6ruVy8ocCkiJnWaJlQ6GMMJzQO5UJh1TuM7/nllpxlt/XxHvggkIuLQO3UQI28DFr/tT6PZp8W0fgk8nFUe7LNUm1/0GsHL5euL3iXD8M512/a/QksFDzuh5AoAzhB7THqXDgDFqVfBwo5FpVbqXC3fixedUTAjAWS87UONoguJ5n5+xjdFeCeQ0gLZaR1cYBly/bbra2nOR9ndRRSO/MjtnxEKpaIrBocC65uTk1eE7tv8WEEWE3cdXsrXk7qTKPOu7sKzLOgsrDLZNBqEaR2JyAifuCBUMyiQepxOWwMu2DVdFAfHszznX+Pmw19Bm84lagELmaddusjYrSu+47AhtwTIRxx+9JyD3RVYz+cb2hXmf6Bwkto0JpYFpydD2p1QsoHGrFxdNKI5gLxQCGjGXuGEjWXc0IVSvsbNkbYtkh2Kpd2a9vaVXNDHLE5AsBmFaY1lZWoMEWkwvm7LOHE9ywRhHB4Re8vpj5H99MEo0op79q+IKiP72+QEGJhhFSlaMoXdMuLyNrpP2A3c5+RagnYSCWEKc8xpamw5kflkW3xjTqWcAibgD3/1EKSphUORyt17LfqOkoWkGux+dbo2xBrXFhoOpV02J4pz27WJFnXADqytemEv76yjIX/u0OfTWk9pRQyC+v74973WTaCCQ/B9/+tY21tcgDw/sLpg+k7+a6+PHAmHSeJOaVYCZw5s30fdQpThZt57GXT75HpQvdHqhGZw6jDb8Ebrncgzw6EsIQSxvTEhsOserX8Aq0/l4AiL72FBz36Q9rx6IfL8ASb+62eQXN6jy9CdHOjj7u0cWH8o6PLesLxS/tD+nFZbU3rXE+6tY1x17gFtVO6zVuJtMDbM8kEv/tSJEC7oQCe4wJJGImWxwYr+UEx7GHYvVHs+CwKJ1ay8YQ/JbO2uJ0+pNv96qsGcZdQh5d96qhzakezXThO/YEMi3XyEopyI+qeVpssiOraK1sK9ohw0rPXNogiP9ihm7MAoYiJ82CvVPx+OEpW2z5xrA6Uj03SeeD45uWSQczFAHIqDdatuBqCwMgjWtwSDxeqSsfZ9OnMranLXBA0+SYaNbO77g2hJUMqZTaA1Ui1a2GCCglqAcHoUPBOwz/cL7MOJ5fWFqInocABATKnPSA6WP7kcI1gPrA/OQcc04cBOKvd2h88goBbRjLC7kyu1Lq6PmBSzHEbXaFYelh8ZcqJwa2S3vUhqGe6fjCmY3SU2YcOEto9xN0O59gFweIB+nNa3TC0VpZvE8hkjMLDUqXhS0DRYZDo/ytW2/ypRvYfn1EpX3L35mwi1f5aZnS6qJixz/D7RxtYVAIQv9PLkT0vJ2p7z/D+SH4cNoXBvriLuLQ9D1tiSsowTjrK14SpTM8aue6UL5eqMzssuIgsfWAhCb/LgIW/PxbDnGhh4ZOCfmSW7Qs1c/3dZHFL/HwZDjB+JK9HnV9+r6PAPPmsnwMqLBxwOoS2MMPEvgNTzPM8QvriUKt+qfL1/OVkNdGOCYgys/TrRqS2ljTA8VkZUk0RKJWdN+63yIa6DWD64Mde0phgcQ4VldV4/d7ZwxI2AYwI9Y2oEMICRWnbP+JgZS9xu9W5oKn+6VzNwpkh3mkbAgLNPQvXAywCsRIbv1+gH5TC70WS7P8nMWyyTauqSYFdCIhRPyZ5kMN2Mj3UdRo7L2ipvp3ePBw1Ik1ffOqAuMV8IhWWuyzIr2VeX9F567kXu+3T/9kJcKJ7KXi6U0UlPc6nmwhSGeT8yZpS/8DT63Z0IgdNpIvPlIB+yvwdGbkjE+yeK/gLF3zhXfCFX6arZxkpyZlc2NXZpLOmZGKspJ4RikNNlNBjMR/0pcMrYGSYDT+0c9eEeoouI8oM/wyMR7Y91lDvfGPIaW37l2cJsA2tmJnVXdbGwIIX6conUDsgyW0qwNra+qqLKbNtTJcNkMmwlRE3Ul+KRir4+zUHNwqaUN2vAkHPuTfI4AJm6LjnzO8mPW/qZ0dOeDu0V6rZN8VddIDUzA8AeqywCisYOy5SefS+3gDxrQ0Cj79SuogjtVsPWHsmrjlrvBNxPClfR3AEqAZxU+EI65ngp9UxmhF7ExgivCk=
`pragma protect end_data_block
`pragma protect digest_block
766956f6b078d75ce96176a4404c852b0f3b4e157f809552befb3ce5d9d53ad1
`pragma protect end_digest_block
`pragma protect end_protected
