`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
/j33ptlPz7JSqb5oCy5my1vFLE6JtB+T7F0yK5HPVI2a5H6xB0+LezD/g00mZo5hzKzV6mD9Z7VHppSCOa6uOhTdNjDJxRFczViDhe4vAs3Szmv0Gh39D+JbaNcQ84345v59SAnvL/yhmTebK5aufu3/+EYebyoRcJvW/nYLyEK7vM/DJzYvxGx0UJuf85zYCa9v7JdHx628MlboVkocYh3NLNcPWkI9DWqE3Yqib8AeD8qc38ZRhtw2yA5RJXXbdhlCGveszUeDVyCY+21gvZDiQJLm2WvxQ6shnTcp3sDab9tjWFR+/61ZaB1G/F9qI/ru0onJRT/Oo0Vu0SfWuO8pt0VEaA7c2ArS3WCgUIFDG+inPTaMruYgtV39XMJhk6tHPCKp6Gd+J4H/UrrMqQJw46jQgUJwR9maq6n2ePetGCyai8LgofMPfq3eB+WDMbOV95C7yWPN8+KSYRXVEnv+xOd0JcB9sqiuFNrSFCiA7/6lXXwcmLvrBLTB/oRZTgl45B+1Cw1JFrop+ZJets6HHnCwLlb17TrN3nxxqjHfV9u4ggFZCPhyJtFQutqOsSa3jYw1efiS9YctodYsiVZ4lkfS3CfBKS9Blw9mNpJO65MFELC6naOS9NaDoCcenU/MGW68TLIzXtMuAccduWWLXVi4pvWqUXl9E4QNEbrioDYJ8xG/dDRW2yk5GhtJSa+EWf9r8G+5ZtktqBX8kXcoX2vVBD8uoVhlF1Qjz9UAlDklP9nOGERHvKTZird67jnwvSpm6Vndw0CGAqR9moa0BFRKG32XaSseDsZZ5MraUAXuJHChJtKGoLs1gOnLyvNNUsgIf6A+ZdTUB5k2OlDm2oHr5Yj06Y4BYIaDosCNcK7vCvpd53XkmtqThqH+/fN5s7UEkRadDcuUO2llIYxZj0XTPCrLyyitrmBe8xOxH4MkfxuZqfrptF2PfQaF2WLyRePyNpu6gQ6+hcebh8GXGN2j0hL8AKQwERQRyjRLhKtRXTYm+7Na1482+N28KNOW6lD8bkC4yGwxh4AI9AAmVYD2BO+HWAnGSAiZIhLnk8SSvZApqzGrgOGpigUwGOJGc+nt0v4weNDM2G9TwqN25ir4yk2P1Kw+O7aAnTYjqBimyYJeLliX6rTH7o4FzwMViwhlXx1dri2xN0gAEuxAFdhQ8cr2f88R6dE/0HGe5AezRDC4YWMacSeC5cmF8r24I7oqvYUHl+v3ip7xC0qj6o/gbaOE+cfV6xXfrVoUDhrBnMrCJAAeCzwtAzVxsCnYaFkeRQ6UlYTyPeONGY8Z+bRGD6MA1nJIyzrZHhMEIZGIgaBmYtmgYVjrb5vXreRzn8YGOLgEXVqyih19oEqp1mmbbS81wwk2Yenp1eunBLwdkZgI9q+7sgDpZz/jmeWGiEPeVDcXtFEs5dbwoqVKMkh/juTpe1vKfh9EXgNPl3P+cVx0TCP8lNsRcia844BOM2jWU8w7Pdsq5HbSIcrnVvHq+ENbtJUNxrPb6mowflYIqysQZ+QZxfDSkLqAP2Ek8Rl10DS2/VfruLSOMJOZkPK6yJjBMnO1DO8Eu/dGo1XTkLddUWV/U6uPWBospuCJXKpYdhMr3Kn50RLE2lGLvJp3vsUAWs0W47tWMJFN47NCJusIcXFguAyd0zF9gNQSdkT9KPxoVxX9M9Jq8A3jvom/dgHBD6aaA9pL9WYdq4btpdEG6pMq5pV6UVl2ewIbdr0vN523+SzeNzbGQYrRWerS42oNszu10AP5hwEAS4R5453NN/eDRnautyyocY+waLVtxbRy+LnCrP3T+P90pa30kd80pfcEAPikxJZEzi0h89sgEXVTLyVGaTH5CPDPh/sD1A+KtAx1wKkzaBArncYsyu/6gy93pqJDuyo6GcOKdWH9UQiSOyq7uVUxRGWh8nyAIMObVKgDh37RaZI+PsA4DKzxYR9r6zH3HeubwwdkTK16/SIvrH7B4NXTqMA/aqTvidE20A9y9l7UAWZWK1/Yf06tSVaX67Cq2aprtuMFrpWlYUEtd97VvuSaj8Ww9CdeE+t3i0rd2DOjzXY1kkv6y375ZFtCsLpMB6mJwbCkV99XQdBfhiL3J0BR1GOw+GxPUWRQxyci03cR1f3vD5zelO/utJT7yR3VNqkeQCJLsf0bIpPoXY6/2B3syrg39R3fiTNfKcnA5sC+32rvniTWBS216kciHXMlOr9D1cZRJWn8Z0u5GOePn3S1ukhCMdMcaXsgvREpmX7wBwCpW+zMuTyAWGMiAtNGI12UdObmfGFCcLJMCljUdIcbEpqnV2Iz7RO897/7dFQwqD/dNd8mNsxITSbA4SQvt56SGo2fdza5sa7e6ofmm643qTiA58XGgnVtEkFeFSuln38pxMf5l8MBH/fZlivzg2ec86N6jNNV2kcRPBZRRAdTBgHDpAFDqMX6Kr6HeQ5/Q5oTeASynLa6LBHWBSGb4QkUxVIC8RjKK07nBpk46mZ5uGhj43M1lb3Yfon6cD75CaZD8vZTuBS0Htfoy1gkVA8jx2Pz809UpDcgBCs6KRulekoeDgbBO3JqVrKfYIMHtPlbqV8lg/ISai9jTVlG27XfRujVn/3Fs27gXOjDGBVBSyyc142GloxtoHioShM/dQeXLf6xrGC9i+whde/FH8i0IcjqE71is7auzBW5Yj+j3d2HH3nsL5mx1d/vPU3YETS+PRFD6c4+mbj4j3NCI7C9kvNIyIRII1gxDG7aidWvCY6qxdZrqkrjdb3BKx9LULtNiWoSRMxxpmSBQ3b4oAR2H7PihVHYBUYLKOnYxxiIiSgRG14OVWKetlsAXZdw7hfbRx0IFcu+QftVEP1nfDlJ5Yl2390h6PfRo3h9WomtkxqRIl+bB3VnC8DxCuRavdqZ07ggi3kNUgSuiP6QSQ4z3y50Dswun6oY9xxvGKhVU1sLsHxHWHSeRhu2NEAQH0rFFPim0fvBIp8+wB/mK4gziT3RVw7SLPZI6pHDkLM7Hx9UonYWlrkkpBZachFzi8fghA8ihO2kxphaGwk1LIDzVgEx+ok1FsJk0zfcph97hn/JYakJ/Ru0/PDCjC6geYAqpdxcvQ3JX7iv2ZDStUsoW+W5EduH78pi4HcPmcvjMilrSs1lWibnJ7gshGrjrARHUi60EbnKLCga2OHbCgpnr+zRAhhRGaaW5fC+AJX4op+Iy8YUtxUJekQNSxtodzHBXDvyyWNPOaHn5/vM35Rp9rPsXeReT3cWF4MD2qlaXTXucsf6uRwYLor9mQz8K652depOLg7yPAvTeSXD2Xg9B5wRxPBsadlhcaXYt6HHk56yWlMAdz5kq5xN5J5IDEjQN6OOMub8tRbWziTsr5w5fHvupMRilZzlnXD+EMAkyMlDgAMmcE9WRq9hdb7oT5PpbnpW0//gg8DX7YtL7yNrs2a2NfOLLf93SqjPqiePFxL9MKVQ0Gy2z72QZ1l2nZ4wjHLlQILAYRlhBB74Spetfy46O8wN1iAHcv5e+rZZDvjs59g7h3+jlZrhKVB7r7IMovTg2eB9n8jiZxk6m/YS8trgdva7EBaz3J9tAjBp4lSIy92qLWHP8q9n/CXzLyOvaPNxaiauTgEJTAg+FWQb5Uq1UaA1TRD11j+JIS9o/dIFpSorBrPtO7heWIOVTA3L4ZM+QyQ5uyQ9tm6qjMwRFbJ/31bRPl5pDUoMUiFFDk1FZuP0pPbVSEHNsFSlv6mvQH6Gtt15Y2gwBJOxzlhHxGVcY4uJxw+isNl7bIucfjeJ1AqrfiU//Rho/q92J1h6yaV5xX3eWkfmEgnwABtdttyttq3mSvYqQ+ORYfNSi66nMjy3Fy6Lqqtsdg85fW9T46AfJjhqGYPg9r4dB1+U/Dp+d7AVws6hJ84sNKVGiw2X/PZDw8+HiXysA6W+v6HNgsmmfcgFahUznNghnQN0c4BkcQuAZXRH7L15L0Tyicwz9LFJ+u8akiV9r6RQFBPLVKJ+n3Lo5wyuCrJK6nZM+fluXi2DQ3VhGo6GAXsAvtx+vSuUnlHpSBwnjOW8ncJ0G3Fb7jNu64kBgVneQZBuOqhSBdhRILVnqrSp+29pTfhrUa6SiR8x0VQjWkak432d8rnwrgZHk53PmvhuX+yvCDF7Np65B56uIlcTsrPpEk285MlsC8VgpL1a4L3Hr2K805v8IWPHVU3eTIDVkid6oE50MMsON2lFXgNzHH2dvVD0m8DpALGEPfTLCKtE0i0wyTM2HEMaboKQ5Ad2mmxfGC3vNqaE8mcfyXAEt2vFwYu0qdEIaRJQ8Eav+m2LQbZPihbtjbCLlz+6Ojpju7/G+mz30bK6+JuQ+EwtHAI1N/dGIIIjHSB0LAGCGLIPxpmFKjUSIJwgEH6cghpa+KI9dyoVGLBO53mJuRaXw2qPIQGzDlE8hWrT7sdkE8qwWLtpuioKFjHtc8fOll18tBtR4f8FaWW0+PR7KfE03ARKub8Ze5EK+Ke5XQUMs6c4zQhOSaf6FoJImq44hmA8022heDvp61i7zPhAC0vbGRhUoGw9Ufo5eGOLAwc2BEFTeoiV8gwO33sMMEoIGBrqCGR7dhXuVght1AjNpfS4DvfLfr0f1FJsWUxkfgTL1PLPNjHEz2kX1UzV5pTOIFTUpyQcxcfrqul9GFXorXTdJd0wsf9yUPPGmkvXKR5e8wJWmzsQgAwttTHZCUEWae1tg8fEvecpIijnvOFqOGsjT9W5MteqFnEBjMbmPDXnVyUBWu5aAlKh1OpRDD+ASW2hXoyFmxPeUrbmxCtdxJG0FH9gWWxjtqOoqFsZvYPk4SgKrdb/6PvejSQGkq0TL1xI3/Nd+Qcw5B31lm3OdawzhOP6Q25glrUslXI3osk1ClhGLsMRSANvx7wQmCeylK2Sqmz+KJ/YpX+bu5suR3sSTjXQqvkObkMM/a9rL9YiQmc787YILRkhF0Z7Kq51XV/mD7nYbq81YELYkCCm+/5OdUW7BGRVxPx9VKSMOHXDi3uldG1rcVyYUP6li+ZxPsE5WK1meuwkdgvd4V1ATU2F8u5zibY80tyd94XEZFC11QEJI0EW0BXqboUgyZbGGNNufHiPr/YGVyy0Z9FkcssD0W8O9TZwL004esee0VPnxp+6lomYLrjeNSk6K/Y421j/Hj7CtS13OZ+udsrVduVA+jd9s0bw0H3pvA4MVXYtEK7zizpRDJ5Iy1LmAvvZrOFQmwwkrQb2K/dnY3dqAOjNXlKSnQ2MC6cO2HuYlre5gPbOVkesBzMfqbkm5W/HcGiYLqniUjnVFdgIzHo3nXAMQd97I49nDOWFxwVv4WzyVwUg2W7sE2sG2ydEPlI5T+KsZvOnMuDuDPadSw49C2ntH38h4Z63iis7FNNhIXHTQuE/AeJ9JZ+no336P87W+Ks8x10Tvxj7YroQavbdjG97spyp4kgJHRmftj0K6cs3uBSSlYEoa53Pjin9MdOgGbH1twhs9HAoJ8AVETxn+PQcIu8foTCFLLC/cDVZ9cnFoyt6YWQoLxh9WLGOS3yFcJxFJ9QoNsE2HkeRKavgYz3J4z/fLQeJDN7320BaCJZ+2MHRdG5aaluQ/oz7X9l4wTNsU+k0HqKrAATZsZ69HfPt9EDRLKi3VeZRqqV3jPr8HU1USvHR4ud568/ef6cbYN09L8nPv0h827PU4yICicqwhuk0dNuRq4QF7RWLZD4SLHQnGhaXzOanrhkuZQrvqeDDyf91W0y+pvjGzZJpRQat7834kqXO2UdBoFnFYfZ1dKKc4QKeUsV01RlX1s96wZ9an4sT/3M3jM3r++NJUJaZ+WByXqKhoy35RAnzhQObGPx8mRqPjnY8w5GZwn8weGHqX6WcQ33UDWCiSyHe4QQeJRVu6nVCAFGp5eiAciWkhgHEZmPP77Bx0ZcDXjxOC7F4rbHq7t/HesZw7ScBNyJbUjW6CvSR36bE0fZF67SxwnPf5G4SkLcDxhvxtwAN2ToPXZgeq4rfn+tbB36UXr1Yg+29YjDnQKDe9Fj85IlAZ61S8qoYPwRkl+C4g2QmK5Vbtd4YDsRaDS5pG37D+fc+WtrVT1uKkzW1lFBT+zr6g3ivN5RsLA3yXMcxqKFH/Ggxsm07l3YvIo8LTbBbwrIYN3sQUIjQPzxQEuUoPe0WS9EWsCsUlCZenubM0ydJmvcRnxSIAHi+YBlOIbZYu+Qlmohn1W4y1qI0ttf2fSdHchK50PKsLUR/GYXiXehnvJxvfJxBShBwjVVjRobCqIlhmSojeG2pNrWHDyar8t+oFGxjRIG8q70jMMEwkYPLw4bVnXn5DY7cE1f7M8BD/AvOaCc8/S1Cl57ad8xTlGzTPocWC9Z+RIz/sU0ZQqpxEdiZT1E4LUGMyp9/BG+YppWuiuBHMxRd3Y/g0m7TG1QhY2A0i2h4g1GXF0hv5z404IxdFIFpmC/1bpEF7LGLSp4sANdkd435LL9KytviZKF3o9qDT96gmXd7FYOyL9wNX9NHT0FIPs1cD7N1LwtuotNmBJmgnGwWUiT0Q+53OKBsJHOKFVWmN3keSkgxqRKAlkpULXrSyfsINckPd89wPFfl3Q4R0n7qH+NsnlTUgoVPjimeMcy8bniJofeQQYZFWiK3KIlz033rdey7/kbQIZdFJtKDaiPrvqgpJ1Q5j6vFv1SSPM/dw33PlPcyRFRiNhZXiydkRg44dU1cxkmzLasf65DRYTJC7l08wAr9sna3X5nuNFlXUpMwdb23ppuHhiTzwpsljU1UiJkRZ+YGvTOIhthVChmt87yf7RDdXLAZuo86IlDXywYQZIsgfQXwbDbR02hU6tf0X1Lj5IHDDaHN3bf+0ItEm+OctORESTab3SlY4Y6OG/tM8PRu6T6GupxMzTk18V5OO/yqUOLkZzbYIK+eSjHaoCik4AUQxNFlPBa5c+veSZY1QFVPao/aauPG7ziMQXOoTe1FJA1ylu3XXYvFYlP9qmMg5rBiXybD3wA8f/Veb9YDWUw1vBansv8gXvaRMKG8ywXWKiX2tAyU2dY7wFmkrnCqOPYuVpwlWGf5VG9dj3jc8WecIh7KdG7ueoxgud1sVAX0eWAw/qVHbKWhr3/sa4ZrwNGYW/SyP+cPurpoCCyQUEgI1qgV8JZg87bodq1TlRjzpcumSDG1M4FV+nckpjG+r/Kfs7TqDFe4S0Q0OSFazsleTykwzZ4gef0v4dGXPbho/nZiizssn13M8RzHxbiYLdhYhzfOGNFK7wFrmBbEGk/oR2Z97/nyDi8eM4iMfYq6V1RRNeP/bD8zG/k3fYB+/5wJjjMpkBzpfn+Gucv6/WlFpTvel2Wuxjz36quGCXApp3ITrkXgu79Jv6RJtPfg5Gcsymqyg60LMOnYPL2n0Y1ed/XBlshKJusVdrOVoqbiJX947rDQqx4me72L2xunaWzsLSUFwJJ45gKzjJVWrdWNyPJlxlFRBMIxU3stKG/jcsDQeo/NuDw26jGCrchomytS6mceVS6Ls++csGQc0y8uWQehaFSjxRhc7yhj3Zg/wy+zO8JAOaWarvsROrEJMerQxMPtwL6ENGF9rSgQNHq2aa0Vjh7FuQ3uPIgjWLWE7LcM5RDo21jdfMNC58iuoX6ZzaVhwn8P0QW/qwnz8axWcXvhDcmiJB03NbSDtiR18BvZ2BPosmGB4NAmpzEi4ehrCThAEYEF35EltnLysIgkWWOvCXK+QHe2oG1VOEsXh/35Y4/hBHw78uR/m9qZKahrDbGMfrp1vD4yOIwkkpcN8tfVAfnMZJWL4DGG+gtqgCiiMvZmzV8bpQoxNkPurwg6ecg/iWlQKdzwox6Pr96Fr6Vv3aZmloMhJ/Z/FEAwAsAAZ1LHWE4zPdog0AedaDcWc58IaV/D4OS9olreJSg33DV9BOhEnYqnEbxRJKLM1C060wTiDtoGMd+ycC5Pt9r5CVS40v6+FAdbqJ4VJsoYMZ7Vk55Yr/Kh7llro7PYT2JSiD6DMRVJ2eky3QxD847B675HfB+HBoxJm9XuuzjhVXSUlOLRTW0waD8k5WSIeMq93umqYmL4tLL/4brSjY6iPBT0ZBNh8L25Z3L0nre4Jzim9hUWgSvYnKW2s5EBHTHbJUDu4A0VNTVyBMpSVZjHTk8UQ5K/ZHpY/uinXLui3QWaptuh0FpFLe5ubkjtp6nw2GLsF8GLKeq/I1qpQhWdDCN33UEjtf8Ojp6cu5ubOkDtbFrYvzlg3nGH/y6C61y1cRLaVjHk8tjuR4x8iroC7csxzKbYuWRuL40+/owMotFPaUjYh71CaOd9DaNTQFsVeY048+ulLGXVYzgFzxvLx+hCq/9Yi6geMac4V+sGhoKEy2kIH3I2VVjO+2OxcWPF4BTrR3pPalgg7uYJC6TFXihAbOQrOAvMH7xMt1evkMcrDwxAV5EI3T/1hd1l0I2GHSmiIj3bS6Fi+2tv9d1EtK7TH+zIJeo8kvkH6f0tGR+D2YCxNVlYmh67DHeRjVj8OSwOSXSejf2khh26Zmx8zc36eHqWfS5EBbO159z8rkbN+V24heiipAx7uvZEgO7FIN7ECxnZvLqpQ4Xl7g25xAon4UWQFA2sE1jFD+C0esPTyXXbq+xl2/R1YqiUFQLXQ82ziiF1KqGKv+uxlHvjOw7bxHY9pQnWrqKw/IgDv1iRRJCsYA4ps4v4sFZNK5TdSj3dLf6UKzz9GkujP1sftC8NvPhNAGuqdh7+SxXUokc9RKRvT+H2D3R7llbLm3v8DQSNjxKzNQTXatyUhyqGDYwcUHvIf/HVheoZ2uuGNZg1mljpvS74e/jFUU84qs2W1ZkAb7bRKt7rVfiiQffwjhPhyHZJd8UTq9jkDarijqi7Pw4xvDA7+PuUVlghnqgu23L2pyrGbOk50xvfD/6ZfBHgy++zaa5JTSo6trZ8z0H/E/A3+murTuEF/OPln/jhgBEVMa1usqwvqD1iO+hJGbVIOVxgKKMcygPqqzFWxLx+AXNbNeawaENOmDVxod5kEmtY+ejifbsYhJVmn2csyZKxKUrlyOZ0xVToqQ7gee2aVhXZDVlPgaLSrNkbRXguej1rQAbcE6cUDwle0CBrkjZSUdf6cF10FlXwAnkpqr9g78kVbE4eleV703eYML/uYK4NlDeSjn0+OSVAj6f7BlP91Y5CTyLgQz5lojsCoWmhXe3r+GxDqfsU0nFytdk9susb900ufvz6DPh74qvm2OYz2fkUYDuJSWEg4j5leL3piPvcbLYKYZIuGrAcJz/47COqsErnh8RZTkcPEaCDMPJLkyXWGjjzynDFHW0tIVpqq/eU/a6FS3Omy1Bivc+M8OqWcC2YwL/M51Z8w7Pz0b1J06K1xmR9vYjmsHyCithO4EuQUgUnXUID6tU/8Xtn3MBbdIP+iQtqLVC4YDRB9QXpZSW2nljsQQb1ZGP0OjmiJsmPvG+ikAMI0ZwyvjwqUnnPzGeFNej4vC/5sSHzkIov7mX36BqdwL/eFdMcP1Gl+9chJWRU4w/Bfm1qinnAy1dP48YadodN9RCFOHM7vyt7TxEHmM11e/Etfhak63pnuRwT3z7i9nO2Chk+kQ7t0SdBkRloBv0F5ENhGVK4DV1pMc62y0foBnmzCN/Z0k0l1ms+nHYXH/tpcUdFnEOB+wuSU6hCYb7Wik2YZRDt7A3J+8btheRP9sTHb1UJixb75VqPsM4TcwLTW0ZH+IpX/FQjimmsj/848axjy2dgZbKpv1X3DKCZjPUG8DPj8itjO8SmaZ7ssJqxWBvwFBUBDDbvcFLV0KBHbSOvke0FbJx/OSKenqEMEAoZzlp1ud66LkGLkXm/E0ndxsbpEmcp3pLo4cRC/tAuT1r0tTYGKRM2tAOzC1soyUKX8koNyDwApGmWuqle6VXusDB54tgMmKQ1PfHa2jG9SyCGCLT5UsY+WSRPAseycYA/XhUlot6cUONIyHnfn5w719U5aD+MCrIGKNBa45RmOY0O3XVqmuwttHXXzWNCWy4qRLj/iYIc2D/+JWOdXHTQhG5sqqtuSNLD0aEVvz0+jYYHo6vusFqBaRZUeEfMqUXSkOXQbgr+TyHjMWNGEpXlTcbKXIg+aMuqgG6E7zNSXfi5KW+zWL/HUGCOVFP18/OmhRF3T1v6df9uDkFTF5hkHQTmzKEurr/vzjek9basRJToEp9Z1zRSGQ+XkU19iq6RsQmGrbSVUjgOl7U+BNrXAdSSY4Wy6O/nB2nOQcwnX03Ghh3WRsKSoYp5X8ZHunftXCcXQdCimcBNFGIvzK2wLsxwvuSYLbe/SXcvDNYydV8QnWIrOyPfbKp8puTap37gGqucgp4qabKDnoSyC63JZZuV58fyzqGSjq1X76fpBgbpTxRPzCbyuHVJK3GZpoCCNcQEEebgc9Ix4NHdsd21QfL+KMqu/Y5k4hnHaoMIMyHX60GzxFjzUaOVeETvByATBgoB3jJqn647igQfe7yiicMZ+E0Nuh9ZFnQm50PQTDDBC4p1TXR5YNA+w00AHS0ugXbfF04KqOzFnxjF83cQU2BkyEG3VBfgHHb/rZjeIbLE/ys0Qp2GD9pKp2RkcjzK9rXuZkhBBNkCC6Nb3zjObTSWHivpQGnch69Qk/NSfkdPMM9ogHxWs4cF80U8rQki8YockbLTNzn6kOuL+auvqNQy8x4XHE6NCHnTPWnqK4O4d2XoeNE1u9PgoUjN3hzh4ZhPrDfYMTf7JW4HzMgN09a3wZD9VrYw6EkKojkDxwyAVqP9cHJ2wjyPXD5fJqElRZx2qgPUG5SHP1sCz211saRfLlxh4hSduhXIJz4wUOhulUyP3cXVbwGYjAiUqOeP7eXV9zkCeTrF73v/aK0vhbBNljgY3b2Ka0vaYMKS9V/ZD4ePOzRbRzOcJqaxu+2jOeq7P/LxczvMY5LzTnRpkCakpWYhSrQHjudGe5ONfO0+dACSLKDYq4/kgxH4+Of6A2Tgz1SfSNXzbZB0EHQoaBuH59+PytmtWi70XV+cFqd9tx1/NNIweRcNbqQGHinpquenl+k2MKrUk0CjElmCn3ZgDIVGttq49jDftFJfPoB0+dVvq9MZDT8Cpkbn5oFJLqiYcjjlYy2PWAxi8uRE3soCqzHyvCUT5/Edd9NDiSBk3e97F/NlF5t/VkV1TcVZVwxVA2Co4ICfs06Kc9TRmRLyPoublnnwX3fV/MIRC+5OX4aHRhM9pPeqpw7U1OokVC85yiPErbzp2ljp2iVWEI6OOkhg2muVmMyn2ZMRlCsZ1WQwviOYJ9S1AaxlGyfnRCjT3TEW4OQC2rnKghOfe9J8k7RBlIzrXvZUVHbQ7320MYyL3qofgH9jaWyD5idi0s6CJn0DDfSq76FcAGMx0EOc++cd8/VQ9wPVFIpbNrhUGP43K/tB63lELZALCNYfiJbjAH4UGw2pJZl69CdJAFARgdKHUZEiJuURha5f1S1Ln6l+SpbjKTg4S9JmkIOS183RUlzpKSfSe0ir7fo9ZK+NAmybpfKtsXTfcQGJoQZ7LxSj3Gbr64r9j7yoHbyDntf6j9UZrJfd5/p3BC9bQ80KtOYA6x1rgzOaXwmjylrAsYggG103fRdXMRC1I3aW8Bw5GSfS36KwrZFEhdYvHLSgF5rCjZMP5k+UEu/C9CK523b9n7iP8O+s4bGfuQp2OEnvip6KB8+KCtXzKr6IAHlH9f2EUjIltYk/q/zlmVnvy17gdE/B8IUwG4EFe/vAIz8Eb0BTV1tvtjL/SIDlN3D96/xFS85sP4b33MVuqIxeqR+q2x9nokZQOuWSlOJX0fxvMy0Gv/fbMmsiQlvhByIV4GJl54Ui2UWhUQDsDFQVMEDlAm13trC2kO8i6MfOg7eUD0/IOnnEz3LmyziAoiWKVZehSlLWH8/ebV+omonJcXclzBXnk41g/8kBnY7aD8CBVNpvW7WcM7YLQRHKF8UnCVCLMBm7ECG+WpHKce66AvwaPVBFw/LpvifnEIv9NdBSaLWpXIJxn5V1znwH1+HxfbAxPD9QO8MOxcTpiX42a7XFl/2ZSJ7VI50zsJHWyd/GhuyTz9hk73zvH3yxol8OBS4L5e1gadko7wkeuq+TpSmLqECRaGaz6hC29pMVn9Kgm9uBqSxto+n0stfxFufZgaexR7JoG5EDmNYye5aBa+vGci04YENRhoLQOP43ITYKRlGzsauhDiYVBbyhbtVlqqVOsHbqBENSExbOSxhOjBVJe0rlCvgEHT2Fbe2pTY2vggJXOQ4A8t5GCfBw0lgcMfV0xQWmz82k6B6W9C/KLpmEiwFDxcBOz9OkUisOd/2JENmqfor0erAtDxTwmHWhjUvu2No4NwbZ4C43N8RzZgC6zK4ZAPsyPNtnGGUxj2iGkw3FrFa1X3vEw2oFgSUjk+ibQQvDjBJiJZL0pRNhvT1RwfsSOnn+kLH6Vk9dDzTyLDVyy4p7ZzFr7Nv9pHxWQWuuTowCvUBHBvXUkpB23O2nXiQqTc0tMDpX86pqHzmPWcSAhYhqTEZHLkSjLzq0TBX/er0uyhEqfcWmL8oA9CTpIDC7UKgJmHkqFWrXHyScOlVfMzUec6fQLYlhygDsw7NOSYJC7/ZfN8ti+Wzul2mP7QsOUcUhoVFbqjFWexj6glN1FwjIXKh68/6gM4w6TN7LYGmcWj03VSDj/NOfNDx6aS3UEGF4pYJ1c/Ed+IVOf+03t9ysvP6SUhSuKVMtinOQedSa2nhNZsDlGhiB96b3eWKUMIRkj485xkj+5jdLOGdXQlqYaf/zqJIhbXmh/76O+K6dKnTJPfUCo6OW96LQNt5gd0hlUnHazbvWbFt6cHwvnzQDjcnFSuPX5m8rFNWAJIKMs5E9DUCLiwL6ICflpkSy9jwArpuWZvgPn+BxcGh+QRHwfXlPpmx7g0sYWVPUufpZmhN3ydPg7rXSd0dtSuWi6BTCFazSDzBzbs5ZhWogZl8PTeFxZq+1EwZ8puFfe5qO3qAeFsF7tvoTlWQC9Yj2XAKCRfpenC5GIEmJoQqkSARZk9cQTh83eUo/jDgClkdrHHrMURvOAUE1IJoODKGtqbzSZ8pepiraK2T9w2ZF/n3TjhuUSbcdmmCcfuczhh/jImnxuR9i7Wb4T3duHtD55WHH6YAyOvvCYQ8/Dbchsd8ym4HbDfkIT/QYX0EG2znW1JyHUnkOp5wLtTgHlT8Y9T4bYdKUVMBI5a2HDFOot3hVwi2Dq6xI9gyPO4ByPLcvFUfQtWIeF115Z1InUWeqQOFDFJjNU0X9Uj9+PIsEot8pzE5Z0sOapgfJe0YqxOlpd/KLfaHvd5x7i0CSwomEVrSU5EXKeDPvSet/7bRulK5iBc4E82sA87HDm6DH8Hzw/v43kGZsm2k4G0EX7KdItEcT7MMDyGlsKE8gzL8xnQHVWmMnNas9SkViCpLwFKn0ka0NwMHCz9BlkWRE10lCf6+ZTikqJWFCFFoUyTlB7Mm7f/ObzOadXSZfUN6Lt+NW0uY+ARDgQi1xGEYcOu4/gZ7x6jApVuQIGv3I8W3WLrUvA6MQnTNmzM1SLrAQI+cozYJAkYw5hflfYaE+qe1FV7rs4N6FgMUfLj2/sUTSSqUTuX5L+6VJM+EP4CcCNEXFwYRnB4TtHEISmuDmg7kFqGYyVNBOCAWrhHhatjO/9aJ5exwWDxBqAiMihdQPK8Wn7C9ae0yzfDXEHYHc56CtEyjsfNTNCw7SAn5v6GgXkQYz+fTE7we9Ao/Oe06dpxtPfqqp9Bu7UUEodti1/Yk6cCeyYp+meU25jx4NGWCms62PAAU0JtloCLHLhsLB4YTHTaYaAwPnD2E7waX8EmcuJADV4o7nfZscYj18yv7GvvtDS5Qyslh+TJW8whtzdg22cwhWaQam19uwxaa68g8Ysn2VjDKPuSpZSYNfTeMYzQSzRTTdqxOyM8yEYPqjV227WD+PbQVlQ+0ny398ebmLwjZmwDl9lWptHsz5sIf5oKT2IMiztysUMBEsdHvI20/v9l8w/tlMf8B8U2Mfw84n2RrMAAH/mKda4akZ5UXGzDvNIxOvy1/2xk1CecnT7Fek7ps5lhQTeUeh7grBZNW/Lk098P7RtD2U1QXZ6ACdo8Ec4ixhxC5wsaz0ng+sGPzKK4FkIMPgeIzBFiBXXIHVYlKJACywan/4txgxZ/yNrPiGFhyNHzOJaCqu7KwLNqJCKe2zjg0XGzuMOhJWcb0k4BJSrqlzC8bIibeaE8Lbu8D486YRXNdyXc4Q3G5yt/uIkt6biKIIQG3jaY8sobuzhbDuL+5fIfebC3O3qBSe/iTUcdCA0AOZ5MRirChEuVExxBVSu3ngFXofpmBUyYi1QrMWAK0jOt0zxatYy3FSm6hjmdujGc4Bu1zsicKfH5rIip0v7eMWBtgS3wjIs7AvSO15qLk7O6Bh0j4MrNyz7i4/wLquA20uZZBWRC2K8xNlT1DuOgFtkCkOMxdy/UVZTh2yWtG4s1TRQpv5DPZge6aoopzQ/TwosoIN+LctyTXrhJcNhjvpRDCluEulF2kfdcTTKnTexzibxGVAedZRbxb1OKkse94sNchBqAWHhI0cVHvFnTX5Qg9PaY5AHpFz6i1Yt7AjZ1n7xF3ZMVSg3hHx8323KvWs3dfR0azFAjCfCz/XP1q2I/0avYwT47JbpJX+MCl7tWSuQ476Mfxq+bb64xKrdg3xCcx/NHHKzOUCkdvcFd/AdhreJ3rApOe/m6LdwgRwsBlT6Dvu3LG1sv91GLAREja63a9mkn3loVSPLy7sfCqhTuMNvlNMF6WufDvRNlxeuU1TQkKv7ptI+1STrhT77w/95/NLvZInf6IPDfc+GrQSeV2fE2dtEZvIB2Ygq7z1PhtLTGdjgVZdPRPGaxl4IhSDYamg5Eopq137IDzudrmxPN5Ut/1srojVLnJYsXTSLNGw/x7T9sgg6U4WVCJlAHzO6fBMYxCKyiDSqFvoCPV81sJXuTsy9naCxBWuHgULFExPMsEnNCzByXqvf3kxYn35+uoVYC1sDj+4ZbYuZC0mkEuLoaqq5NsoOPg2Ls7EEPk6qeg5MpYgOO5XvZJq3PWmNHs2UBP44lnM8Ihxemo7Bt4b2676OL/HmJfp9Xexd27E7JeegYmszioezetD3hpKLYOkQaegoMQ1O5/0AFycOkmVxt65A91P60qoBe4kOTSk8csKUOXZ8tmCFeMA/Y1EvMa5xd3ggaLyczjM1iUFQhy6McpJR6MFRu66fmDIe2QIclTp4hVHgHDGWFz1BOEjaLXPzVjjLChGYzNT8ZBV/INBo5XYG4HsJ39oLOQAbdMLG5HjUkWxsHwM4iDeaqgs7QDT9oo/sR+JAWrG++HAG6lZ/DSCfCJnk7Af4yfFcovA0pSF+BOfIqTIyZI4yaNXcIUdCM4H2ZXLvFGNo8JG6qXgf7lq5u5LOzQS+0ILkcODjga//Yt9+2l8qZlGf0QByQ86hQXMrD46/AgtQaUL0K314EReyDZnfIrio7XMLADa8yEeTxSPOaDpBP/q5WPVR1MrxD8PUXIsOIBsCrseIIaq6/rBkZEC0kYrpFfn0+l6GY6W9kUKo4gmU+2I+398BiIzl58biU1z4PnL5u4Zy9Ia0kQFiSYDpmcicSgttmS2YTtuph1ZneTaNos/THg0P6OdhhwdKX6rIF9ipPjfROfdm95+CXet6irPGxRl6f8HRMKYV6P8KwdccYkfPXaKovI3LJ2tuMqXMyaWjk5fdF8vvKZ3uKAPw1v49pTdXpSmwm7tSRCUd0VUCaKnm6X8aSBk3ZJ0hyYoAXIaWuPBxpDuo0tSh+Thq9Vs+ZKHqNd2BAbGU9GDBOvlfW+k8eVcGBblQq6lNeLobANAQ5gSjOBVHwRz+itw7+Bi/spQjrh8VznZq8n2doU1Ar8=
`pragma protect end_data_block
`pragma protect digest_block
2370f4a1468ba0d087a7c652b68d7eccc30590411fd3c67c2eeb4389173c5c46
`pragma protect end_digest_block
`pragma protect end_protected
