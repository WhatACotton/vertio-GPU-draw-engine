`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
2IrDmpEVHxE4rHPguN9ZAUhwSgFZ7BU6wqVqzPldRkDdVmb0XxEG8MSAZUqLjqmixA2BhkKZ57nSS0yLz/3CGRlxsYIou9zcVXkAdm+sYsGK9iAa6qOkuQmwr0OwJPz37NzuNa+ffZuF35pLw+JV9TrMze4R/V/9NR3fLfBIFnymGPal9dzNabhVwLOm5N7+aA75/6tpkTvW4nLhuKt7BgRisooxHVqS7537zSoggCLMn2fReA6DD82hzE/oOaDB4BHirgjyKjbLiBzeNqERPM24MH7QKacVKVICYHHZA1+sUQiITjTfHN2ceN89wbT7j7MhQabyjP5b8CWnbFtxXhyZyijtQUNbWJpWrZyVa0mAf1OEKwVTlAQHBQ2rYyZl6BU2HFKa/5yG0hwLBUmGVdEZd9H3A/XbusrDuhcMMA84snpWjQveFx8wOxCY4OUMbpIC6E96OWvSvA1bA/SMfGb4AXhF9oxZGW06P/YMGlqI1CIrqzHXnO7e8j6XHPS4iQUkuFsCeVeG3uEo+r8PIXRMALMxBhLKTE3OktXkyBAhK3psFacLDiKWf8VMt+dARchW+Gr0VpOTbQEbSNklJW570cuLOI6MOk158NURj0Ku7+GOdlNtVl50LMkuG32gOVLOLXFE1tVRoQ1jcqEX5SrrbJ385COo+OcRacRk981bHmbAr9cqZIlRC100lE3YrS+LHQaZJLpc2nHVsxEgE4utLeyt8bQlIuy++N/OQOeFNCrDKVxBp26K8knKlSpu2/leqn9Tz6AgLgq3XREBZGgbxMoyujRpFNWWfsnU2O8Vm42s2Sc9B8ira1RSEr5iAxEe4QmGNAcQjHPMPQm6fgHxuvp8TO6GS0YQL3KLRn1hh6PbvWua12EiXKcy7Lb5fVUfAoHUFup4igNQJO9Qqh//ZyhdEV+77NkoP/1QHBSYhbMQqadiFQa+iT4tYPcR2584O+yVABj2G6pSj9i4jnYV/2xAucR50Bx2oh2kMzlhoQbzz4260gYQa8Hnc2aw0WLoj7ntC5g21JZDljQqo5Kb/Rja5ThMORQu3HWxJhfjdzhSfjpFymIaMSjA+srp+QrYuj0UMGIC7ywMufm7OxPqEE1YsKbxrZQN09bcGqTI3tJYjpgU95a306Gk5YUVfkh29OYO/uN1glcVbv3OImMar1TYE+4k1GEw0L4pIXzYVy2MQPe11LRUahb4nGT3zSeTN066jFAUqGCFho6G8SXP/UBEicMcqS7Js6u1gUFW3Qt6pTLf8CTn1ZQj8tu4EwQe0mrtGS+PRtR24X4S3vKrE0VLQBHwSjMbhvjxdLTuws5Ya+UpQqZIM7S0fgToQteQqFMr7aKNZQAxjgKJkczlQweQhIIr+6FX/d8oBYhcrZMySIkrm6RRQ2r3CGwu6BFBRGdAr2W23YahAfqdndBuqJOk9u067rpn2Gs7uyBHUeJrGXvxmG+II5QZHtSFtawIu1I1QwKLgik+0EjfTQWjjs/jQhiN6w+qGIgsqT4Y+5LUOdnhAaim5G2jNC/HXL8YuDGZCcD+Jcyj6U7wgXN4kenhgKWTRRydwayEUFSQuoc2pBi+pGBI62BOFLnTIv2oar6IYoDyWWdI5lExHJNCEbvDDiQmvcaT7Jv7sFERs8b/hyvAqbdnR6E/L3DHtciICyJmu8KNz2adx+a9T8wRecwTyAxSi8X8KypZ65AKlHgsprUBfJrYOb1W3wm7lQAlVsm1p/E9traHF1tQ2dUm6ZeNzYi+CMm68tqXks8Cj4WasNkGz7ebCGZb3oyoxflO5SNrKNOAf0IRlqCT+w==
`pragma protect end_data_block
`pragma protect digest_block
64464727f907406916ad3242be98a785f9b615f47b37e19d1b3da8767d36d8b1
`pragma protect end_digest_block
`pragma protect end_protected
