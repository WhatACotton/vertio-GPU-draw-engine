`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
s4556xDMYAfCtexbdkdETRbopiFEb2tH8FBXQcDHsZgAbb78+xjNhdmeIEAvL6GZIko+ZTz5pQtE8NUhQmJPVtANHlFPOryGuEUIxTj+gDVdcKpXeMSXcw/qWq66teVZQ0L0Y6SqFtKDELuSelTURFSRkj4eXziJXaYlqDIzFkT6u3+2iMgT3R3wZUxm9S9GnbBsYgVsaSe+Y7QkHG+u1WTTe0wans6VKu3mufPg2wqg9d4+qn2wa6RhVKEUHaeShnHZ79pYlMwzB8RIzGoWGhzQ0ONWdeG17YN0YsHo3KsfnQypxBg5K5+DLXrpSV/f4oFtiH2HraAgl6wtIiC3+gW1mhfo0eyeMy7dmzu3No5vL3woKTFvr//6hqqAb1pfx6enY5m6hiF73RxUg9tq9uBYPSWZ00u802j2L6Q61P6o5ABw2mu7TfCfr9T/PmystQK/9QPiaL54mv9huGhd/qooMkhAOzYVZ8Vq3qUNeZ7L+4rPqovvtZ2Mr4wFAQmvY7QiGbTOXJa/inl9lu4N1yiw6wEof1Sh69OCYWFJojKy/aQwbXba15JZA27z1WmNrFPCB/qNs0L0097nfTPSL1mtql3JvNX/Jxg3aXnTNvDbg9CudDOI8wu0Vf3RHOgDuMR6hS1PoVrDKy/IUeqe1hhg2KGS5UNc8AtTQKH2Fpvm9k40o018AzDMswmpbIq8pQ1LkA269+j9PlEIqxGiuoGkcu8yhguiCThj0hsNGDFTrIjgNG8AV1wuXVxRASnEQs4Yryw0LvHG77hFNh9fZjXAPZa2DL/sAmC5FLDp5JKyyYruwx5hBtMOn3jD227HWpts+8g5lQgDCgrbmnkzsgGVUKM+XsphT9RdhXtPvlfXdYY8HPmitX2OIvrEpYmwjm8wJbJe3PBQmeWjenbb6pkhCbd4UIzZOzjFHHqCm4I7x1bCmZEzQFPcm39oDsXf1/Zil4Hcyb3WWT2bHNgg2vhKeN7NNR+ou7+uTRAC/Cf3y8HTcCp7XsawCfHGYAKfmHQ2YGdsVggHWW8k1jf0PBv0m5zWhkRz4SlaReS72k8Fpr7DeTSo8WMEySNGxCsWAVOs9VirjRutB2rMffsmpV+v4avCPNijpwaeSOq7KyUlqn5ffEBvMbkVguIbQOQY6k/xmENGntMKWHdGWSVYJa3B66OE1QyVo/OS0NKxmZ8fM9ZqQYkkMLwH6nQknkxBZhWqVKLKa4BQFjEJkJhjWOeK5ZbG5qtRW8H1zH87UvJSp9q5Ga50paJz5Aq0zYiLDIXWUFk1nItqYOA8xzlyEyeyOo4JBTnA4kNkB1/uRyv1qMUZyYTmqb3gvsCYk3EAyQ6wmvJjXclhmwnxAwD6YNTVZ1sHpj+RSfxElBjGcogTBLYmHxotw/50PeLbdxMu2HZb7QXReByDJNoq7tFqQYdoKrQC1pDLRHt5AhPzmh7n5aH7eCclq+k7NKPeSi/1wa8jWP0ktbpphk/UoMU9M+g5pSl1HHtf5G9wE2FkjnQ8eHjnHGEmuFVZq3iWYECJcrT5ZiK0e7/yF7CFM0s1WN61YSTrk5rUj6G5+jY0g766dsejD1tHl4LRQCihwjNikOaaRGSlNYXOorqv0PAikvMmPxfWl9fJ4OpbvPgJ8wrFvfETx1GY9OfXFHDbcd2eo/l7E/Q2JPX0eWi7MPWGZyr4vxvA5Vg5YPTwqEfuAuOYfZxm/YHQlt1z2ziD1Ec6WZtsZ0G+o+4ZpzZH2lGxs7SMHSV9CNilv/mkkkhhYrdabhe0xEyukdCFIN1PsL1kn3yrs+X4Gr2bmKohN/fSZUJcNpVBYJ0CU+3K2DoOZRgqJ6g1TPPUav7lcgkW3LXm/Fnu6ajYlmcsMT31JKx/YsOXbSuUTWfV6eyYjgJTuPEHKRtIsKQLAhhXeYBNgOmIrk4yUs5s9J1hz2oFhEO5NkWhknPrbItNSflwncPWVZmQ7X1/6nDWXLxTZiLSFrl6LIJmXwFDGPybvKoAcsU+FPoCqcJrUTl0z3ypHNNJOBbsJeJJ9Rn91JyZ4lbJankugnCRhsLznLvWzfsikr/kVBeAsOT/0zSmUz/N+uVAv0Dq0DqSalMRcr9mVbll00QxrpzhSSK8DTVmP25z5sy6NN80hXzcHe/0Cjgrgu2UG7pU+2gLbr3r2B4b0jEJyAUOZ2PL9S2dauHvgSMKI1A29auPYCu8mt8/GiqHQAFTnl0fV3hOWojnWG310k6Da5M09yIzUzkxDk1FAn9ZUXltLbJjb0TO5dqy8PpuF35WiqRoze0nvzoeBdofWhX9nrEM8IqcgC7h93P4bhqp5GupIHrpER/KD34dQL8KGgCO09H0n++24xayaeC1SP4m/GmeNhz0+z0d9zgiGjlT9K6zDTR71twISodkG0kw9GdRY2p2/QqRZjfWbNGdN0fqWl0cfyZLI0noss2MWNbW530jI6/7uLDRl9ZewXXu7BylXgUfiv1frw6AuRez1Kph5Jy/nhiYtv65wble1KgRr+iHThvsnuQdWRk/suSfHPkf4PkYw1nCstIwolCGB4PnTnIOG+biwnqksHA3152em72jxJAjBtFerUP24QU9Jve6hUkkuMyTssHUTxue/7Pa5acHJ9mMdwp9r3WOET+28v5LYTFa546VKghK2FRyr4V3OxR8FooFhuvJbcqv86csBYYSVW6eZIzsWQ8t1folefXPdE14KW8wRzPl73me+PSk23tNsUi51C2oXApsGVf1rjc/M0Jq1G1iOuzsn9CNL6QIKUK21ZwABz16eyhAV7qiTnwwIQ/2h4uEosn1UKev/aPC68PnIHCOUrh/qDfWPRavK3wR1j6jCF3W8rSTJS5tdcVH6fpbEFUBMq2WaEHx+P0kIbSTmiiWdrHsgRYes6ehrupatNuQ0qtETTRSug/TM1GOSWKQ/YehQfhKo6lMr/XNF/TZvCCfRIF3CpPkIKGOmUXM2sJfN88SKxskiB/+m+v5jEkPbm/dnFNzMTLUt10tRVm3/oddoaMZyLJay6bGX6By5EdefjITz/Jh7VKgGHO+znOGdSyjZdeAacOGeDKrBsIsyJszsof81tX7w2ZG0tBsDL1FQmnNUJQpSI2SsuT7qgpPdagngVRvqHJGwSfiz8SyZnXeaWcDoeJ9tYUMI9HiCDy3FAADYzs6GaX1oWLHtuEdyLB55g1iGGu18FPjI0pkx20OfXL4WxA4Dfos/y+XNOcKQQFyOVpj2lnLnyIE45f5+s6QXj/r15TqKE7gye8NljFEn3mv0jkKOueqDzjgJEmb6E0BrBZOj1EZ+Pv4Ea9KS49DXwC5lx2JPNchbvbmLRLtda+kD647xK3+6Xl4oLqD+TPop/vl5L1tP4QK6T6TPpGDl58ssKkP4Y57kC/xXNd+p7WXVRNyO1LptVEWWPPaBToQgZHpFOlH/ommZ92KCIrINvziEzDcaCi5OpVKtRKJJGfzao2PM6C4TNcX9qg57sBI1eS4iUAghTqZ/S6iWeT+rLtmJkD1Uqli2vZW+sYkRwuul50r4dREeQdVY3Zfg03Qqc1tLX5kb7GNQ1VBIlF2v9HbgVGAWIuLe6n/jwFnJ2RPhzx9ScmqQlb3uWwxi0JGMVp0K+ZYCnAha+QUlcSIDgeYwgNF54+Jsg8R4QnNq9LYm/y+B0u4tsCWAGY4FatuUVFKh6Boo+0/r8Dt8jnDC4Jvea8KOxHv+XtCkXPfsQBw+eo3K8JpsUDq2xHKFvfbtVc1T4f2Cnsg2afW65wj+vltkVsyogIljn5o27cocy10ZZGKmp0R4PVoIILUDg39VWCfr2aNKuVMTFtWEHWJqGudQTdOse2Q0q0up+L73PnH5B6/lkU4EPOJIrWr9F4yAK73te2E/CwtLdgC9zj9EpQ2TylXodrHh4uvCaddYcBOPv0530rWZ+mOuMcvVrc9KFt3lfbGEEngfTdwI3PmRJfSZf2RW0JoKt7AbUx7KCh5bNVof3pYmgwJFa/jbSaEjrgwL3c5VSzj4pBN2G+TYZINxwI87SVFnsxoe/y5TSEQJsHUVho4fx/USNmTy2c3I3UbGyQff6QMURo2nrmUpGZGNGi6b9VtwCWf6581IPSLbajntqhS4RSr6FwmkaySAWdxBx6N/2IPaWmH5lygCTVQzQiT5MQDlVV2fAfdQyzSPU78TXNrx1t4JO9H7Rwnzo3gkbUnm03FTyeSz+BIfP7wjtCdDO43/l41a4dri9ySMrRYmWomCk/GydR3vMpOyEsTR0Xd1QPIPkzbq29sw72tkWwdn4QqqZ9oc8jAMI3mIkG8nYA8SuTu+8saRWnzeTX+gVSJ2ruu2hdWGRBUrPV0rKj/k1+F+oFrEpyFNXjE2en4MrjkFLeFyVWrpkpmTCz2embW/c83rgTwcBlKM7/Vzr0fY04iAzhBmRjJUHSW+1o2XerVl95o821pEvUouNH807B9YB/AUwT4FJC/boeweCDdXv9AIxI+Eky2nXEtvd/snuyq75IwTuYbZE3gxczIJ6BJLVS7JBVPpJxCTZcKSMv9EWYDLgnFwfueM4SwSbndNtgEdpIfxKZRHWmtuPY5WFSJb4iMAjxW56/Nv6xTJLLdqP2htcnUa4vG4PDwz3E6LEGEFrM2jw6jC91f8a2Pexw+D/yTAMWbdlo5tIEflHC7QfonQeWSI0PRlSPfM01bd7gVnyOSsfv+q2HMalS6pxbY0kySVn9RXbe9KgjoAIAa2jgEiw+IyAHhJOlBnbyszEwbXo9UG4pX8KwMx9rGxFWfNTb1zHAmyeJcN63ljbOZepFg/VV5Xe++VluXpJpK5zA545iPQpz/uhfvg2jifQe73Kf0I9nauQfdPe0+clvn4fnX622plauUvONGekqrJnuU/bpXQlV7ywerf0ogseFkc+4YFdd/VnA19qVxXAnqta062HGLvmYiP08dk5UU/yDSpeDZYUAHkSJdaXc08QprSL5UqJxi8RhtUEYxIFjde3wmlpNX33muTxZxfT9yiHzPor/bS6cEq4OE4f0/WcfFx1h+QQhaFQH6oiIHturKKIQ/+f37zeNQM+Pq16knOP4u56ajoH3yaNvFKa7iEyeuhvDRvpiy2XoUD1REOiiBQdLWgDs+vtYZWWOReaAAsLWhv9B7xP4UHPhRRSjME5xyt4aYL3IuSZHCpgUn1OYPKOEI1kG0EdVrdpQAfw3NQQtccYHnRq7G45T9Sfrk+8dNynPBDt96IOMFPhBEsAzIZHM8OI+J0JZs5w2hJsqQSRqhf3L3tCSGVV0Bi4CQmx1rFj3KI8IySFADJhgGWo44DsCREUV1zs9qQds4BGyLaLnfqxCEx+T0D/AXqcc8RMKKTwrjYGDYxiBCJUemf6n1APssmMsxCfYyi/PB3dYaQ49xJ82/4DbZ2HyBTV+o9bnNiG5tSd/MuDJo1uR6aIVEgdi9bh2hxBNEEx6OLUjSJ/Sy9m6FU72zL8nuM8gFNPLfRgsXO0qyCLoAKF1YbQB+Qt6UXjvUwQWQ09fHRmz33H0Syy14KTsRL4Qq5th+F9roOcbhrPPEwFuezjM35mnBhUvlf8BkT1anS+fNYnrm72HLDfOzqmEteP1f4dXoChJVbSNFGRKjB2O41zaCrxBpSAR4H7NUJyexPRagoFnV0uoLpWj0+0iiW9F8mcHdP+MoFZ/MLI/xl4ZbrJvVA3zhTMkdI8471ZO4V5+Cssb8LyZhIjz9X+bc6B4nYzHu/0ceFLzf79zpMclETCu49DPTRixPrJQYizMEIqHOxT7fgAXQ18HJzDa4lc0RtKzU55EmX93oqvrCTwx6ZHuF8f5Q/lRKv0Oa6SmpVroRKZzSBW9XSabwHbFuvu2l8unSllP5hs/KW3xf+XG8J1e6OFqL1cg4ZA+DePv0J3G8Ff6qHR+6RNMdls4uC6wy3CQ7KQl+sTZrtclNMai4eHiD6qPAZnZjoeuAHvGnV5pZrRr8L5M6oCAz29HEqNf/8Xceabi5NFKNUCHDwSjFCbA/xUv+YOHrMM+D4AjVuMrF1SsTLuuOz9qULyi9AzuKTifm2KCGylOttb19QHJtTaethkjxOrZmIxS5QZSeLMcnfuHvo6D9bI1bBZN0aW0O9fgJj4agJuDerjfawyWD0TF55o9P+YgsG0wHzEKuE/KE0jdtujbzfrfrj5hzmanLCxdDuMc+YVmEFNfNyIMJHcDOGUgpCGfOuQALURrFNIvfTdQ2nkLChLv+KGgo/Du7jNjbmkvN27QeOo4SJfZ8EaQ2heu8oR5KfpMMZZ3RRgi7qwyMw4zBSrOey+z2mvv63FVAC/mEcyCfzl2DntaXZjhhCjAfqdZcmu9ewkkhaxUt7aEWVrsdRO47eiNJFfaSjo3mZjA65MXXXAMl1UB0fObS9FARG2ULEspsTivo7cuBh4KUNyYQbVbX5BKccUJrTapvKaN92CKr6oy5wD0MdBMO212gIwHadzhLXc+B/jh89mvKk1qEIbQt8hUMhjACdFONan643IVRkSaGNViab/uqzcfF5Z3FI9j1Gv3GX/W+gq7GMj3Z+2Y2b3aZTHBoTvphPV3OAkJwsuDHGaUS+De7w82WAXvPfC67lRLSzZK4TXIRWAuzg4w5p8dKDcHnIrpUpFhdvG6Ddlw368OCvz+FK+aEPi1QowP564oseQAaHzoT7OFVTLHX1gZCmN2NvZdwHS+liOh+e2UUFTJn4wWfDhvkg882bhkQ6GqRgMY+PQm3I3WYdpLZAsrpY4s9aiMFDWPwDS+yUpvcAdbYw1RGDQD7lAONPWxSOBlnx0mLLajV4ocU7Kd9W7zhbY+ySGH6zfeyd28+OLPTJMEeZqww5GDF8BsACk4ZFSATVhqL9lGMFeaq/YsWGC1NruPc59cIoX3Kz3zhzelJ2FKYRfJ1k++FiOe/AOQKCxBCmKJjjA1j+6HxXIcUVFyLyk7SMxkSf77eYMjr5+7VYt4UO/h2NFg15RZZ+7wFMznyMhTX6Kvgdkaiyg6B97czIa7E5b+5qGRQmwn0JLS6UMT2TXcH8pNOxhRrev/Qnbfne1c+kGPScfv9mKgodEeux9J+bCL47vAcrd9v9/GRt7nvqlziC+1ek+9opzBQhb3XpdhJI7QOHzHuLWlMPyFsKOIOyal9EhmoqlXRkQ88Cs9iRDRqwLFjAf7df8SfPLuVI2krEsqOV2OZSZI5nL2vVkpBiQugsVEKo0spHWQq+on2Uo/s9IeUVfLZFFZWI60cOIhK/xu2yo7/PxkJuO75i6qbwJiuSewxZTN8rNZk/6DA38+7fukQY++UEX5doQHtCZSsZG1zmx9hfaUGcRQD/7vnYGwbtJrprnmvcb3KKCsmZ3JLeyxpQPZyD3uHD8nliLaJ63Re/E+S7Qbb8k3AojKEyMP9PifvxctwCp8GgNer70SUpro2zn1n0K6ZCKOSSlHZwx23AXOMtXdJFOxekqgCh0Tb5wDbn45e0CHsQepVpS1yqT+YuUggPxcf27BlrpceNBPcW9mMzcTrj9bayB/Ba6RFcfkaEqlrTR4lacOqcdJWOUPEAouzbQ8EmpjRj3AiZzWIwpdlKDdqlfGtTF4hfREmcsw2GhHd7QdhLQxSO7jXwxMbsfTUZ5RAECJwwpbeOpPjpCt9Dd+eweFSmSffo3KRU1hmjvTneQjHylEjA3E4QnCY7fxighi0Egf0Dplax+n+MgzWgzyithwFcxYk80IVk/shSA91U6r+url6C/7FCdfUKjyvTCvNpuvWf2aZN+IQicNVO0AXVsxRLyBG3xnhXa8YJU3vZMkK9fCh2tQFceQHf98aLQj4lP4nbeNXabF6tqSMktzA58gij+P42NKV7t7KI5pPBu2EwUTOOQf65+PaXQCrIq0CHiIhPgZfA86ggROEnUAWsSJ6Y+VQ69FBdExnZHcyiYsybX03sbk9f3fj+63dv2n3mvOz2SP3RulW+VClsce4Q6blX9aOLeCIwg6tuU6UMIklzW5TFwgmN0Q6BHOyI41qaxpSzYGYgdtUOm1yLj4KxucaWweGlMmn2cVh6r/QKdXp4itVwuEXZCUPoaqNR7C1Emkyhee9prBSwvwgZ2fF6FzYIwt8yBcfgjc7RZ7sWK9EYLsTqr2YlRHhSI/FhPUfqb1pFNqd0mWn4+y0rYKdDvm45uzKMWIOAgwTyqU21Z7DVtYlErFqPGDNUtmGqHCA0Pe0ftuuHqNjoz/SXtdZoxNjoOwG0K14aZd6VYivga9NZgh7zeMMTTmD9oiUAKykd4fq+CygSMZREWYRMoU5Lh5mK6ZjrOcLpvPR2zkd+7cQUvnWZK8WqYleD1mqvfAynczDyjjfqIvY5FGqoYoaEnhWAtuEGNk0qxJPPiM3jnQNNL/BkvNRm+yZVvEUzod6vJu3lSC2o0aAUQNpOQN6ygq0hE2i4PbQ04imVGgD80wqyoXeFCeeamLngwQicdCLPI4g0IpTippv9Pq1r14u4ifvZN4/gSO5RrSS1ylDj9wHVD/cjWP0uHK24hZSEG3oK4bbwkV7UZN5NB6RdZYFDI24RbP2ja7Dc5MhziPSfawOxMX9C9DaCC2sJdIdx5Dink0quPhOphUidz7D5zrj/qbYVymh3Qgb0KSRBLRcJgJF3LsU691stvxXqxTqcQhs8nkJrgG8MRFKBZVEzvEgwsm6VJKCd8ldIWZXCFoPdELMFnu5lzlG6aBJY+ZrrN9RlKYD28mid/y0JgA8DlseBCQvSk82qKVcXDJn8fQ8l76XDv0tjBhOTx8nqMDeiDIze4MQAdMzZFq/pi59ah1DnHjaReb+PoFWJx1YbQXZnrQ1AyBvGi8WOvLtVNIZ8QasXgFqefGgAOeCvxYHCxHi9UbXAoU85rdX2gZpe/C+rvCDzxejWYTuBjYsaACL7/+u9/two2JSrjNHYLre5GYiawdA2MpLLt4g8nu8zyyEGln8uyhLmoDOhkze2s5LjLk3dShu5yBHYyDvUFZuxf3X2mK+8Pbdn3bBaDy5ok2Ay7Fa+7x6PtbtA/PXsBK8b2l9mxt/tQHa/xvBSX9dd+bHCtcynZ8yQ+x7UnoLa3c4p9reL1K7jplyh0vjK7BwzGzYy9FuaBW0ra5HpHKhPo3YOh+sLvDReEsXsO7U54XgdqDdvBpAmOQ80djdG6sLZKUIhWBJ+fEv1tZlt8L19SrfCe/finZvJK3z8uz5dxUVlVwyTBPmtA8reCY6htNDWe2XCddopcMG8rfC6dMcrn1IEXiK4FmP9paGAmuT3XJWaQ/P3/GsoNCKFtMIkHHHi+biyOC4gmMjVs3It7L3CkUvz2Cx9LgKJg0GvRsXsQykzQaa0yxAY4aUNXuGPk0QQwcwioC5A+xTVixkZXPw2kxCjBGMFlpjgJZe0VFyDp2HqEihTeQR7BP+z2kZeSGa04y3svIWnRih/OTf0/qx9Jlqfk/gPLkdWrCvs1AZeQY3gCOzZ4V53myrOph45Rpa5W1xz/GfWHTnvPI6a877XNPRGA/P8X9rW+QXp6MgXAmbxgYXt1vP2agUCiBt9w2NOB8XL/9xGJBIjx73xomlBmbUn3JXX60lZVUwjLRwfVLgfmskTdS3t52yoh+x+ffBxwXHnSOjCtrHXCaHG6C4T2JglUPmz2yP7XO6LBFvbH4bPLqHYNe72tU3Ncq5yXUZ+n8OG+9JA5gS/WXcSNcOhBs6P2e2RwE6+Yrp7USoYqOb5jvL9tVq0RrmbG0uNeNhxZ7hVTap+B37aSZCNyd46SDavR3x+5PT6XJ66Dqem5gmfW1Y9LLozIQh7msdkpdnkArVr3A/yEqr5iADXQ+nTCoetH7pFseEkca/QHU9RSvyvHUtIkbmEZbi7Rvy8pgJ0MppksbSq7d+4ZMdAj/Ay/eLxGOo/R7TXIktcnh9ab6o+u+ZODSpBArAWd25lIQt6Hib95R+/DOl02ANkkyHfcVN/HjUwQZrZy0ycGNfmlh5J5eS8S569T04nWb7wCcEL4Va5KIFYxZn5SZze89l3ie+oAu/hmHepgYSHujEhynqhQvA8W3+W7jWVnk2cC7zPOLAr5m1Snas7weup8DYA+Orw80tgta7V0cz53k2pckCrbAX9rEmjVHzMmoWKamJa6fRt31nvzR73NXkES8Fu6zugTNq2Nqiz/1KJgAHXbBlHugcwCoTEvaFpnzmD1jvct1a6cUoYQxNlxmwHmD8NG1K5tuwHnW2yK9kSiS5GEIsiEFQOAB5xEdfkE6TSWJIqNOod8nQuCE3OrRHu3+n5UiXi2O46Uu/PELT+eQQcuq1AmUbE2je9VqXieUvJwMCkbsiX6ieHZl3LAh6KbLqYgbvPn8fq8a6pqfHM0jcsa3hfto4SiWannGqOrgPf/VK9Jn+Mh2uy3f1XfeBN2aHZ25VJfG1UNV1Usg5v6v1WWeWsmg8LsEKt4NM0D67xnq8ocFDsNVsiANsp/asLtkgXYpMSVojAbBixN+6biNDr6ANQuuGA2ZzdMuJzN3S28pQa1vlOm0BbGES9DU7ULZpGpK7IzyCovEN/9U0jvCETg6QI5OWl3rqChqSp0Q2REZaha1OjnqinSHxoW/xI+ImMQ+lcxSjQo+YEO47bo6/mvoILevbt3Mtyi3oO0bsucnEnw2Do0V0x5f3/cZIxyyMKjssQ3uK5hk8LlDq7Dmyf5/ryyA5hfm1omKvlo194e2K4AqO64QmHJHfj/LQ5SOCGiMq8qxZ/K/Tnk8OeOKE9HX0Vh8XS36M+3Wpi33X/Dyh/CRKLzFsrhH+y4D8/1XM05G1yDaFatJSNKhkFaFsjmZidGVo4i5crG39AYoSMKfrZMIx4YAUvLGvyOlDPRt4fxHp1iPvuonifpNDcOmzGDBXAR+p3gDn4NzDjvTBI3o43SrlaGe60ISkq2bwa3XiW0h04wD2i6vPOjJWgt73egVLo2Ap65HD1A5NPLmOAwRilmibOrnQSU5bt4/n1fFWdR5cbtMAtKehRl1LMcq5IhlXfkZsfabaDv89pLANFp2EG682dPPFiNUbayMCczQElWsagnH8vfyrd7ABdy2RznhP4JdvHfpPO4pI26IvpOYPPJxPen8FjrdbQKxNpd58wIyBuKX+t7cdCMb1NMJpUl3naqAq1MrIydi9pZuN5BUSkV5+4d0QXUUjzl39y1A2gYWp6EIwaycsRYUd/ig5LpFn0q8e3kGbb3cSIN7JKQmFFcihRmf3PmyKTimw6yQcX4WfxHHmsy2ejy2SHQcx5kcpt7VJdrweQA3bqMSrerv3+LzVdyOqanloqIMWfLKkEAXQmrTb+nCwyPMazA9DXh/cc1Xyxsax+f5wCUx7cvmZhNYbPySfUtTQypYRQn7EuUPb2+oX5LIUWoFe+E+AjkGQtraRH5uHw/1Y1o0GrbbBQLVjshUTYoNDNj9e+vQavK7P24lCWX76FP/Ah/QCkNYdzpv/rxuaT0TMdZoC1gmtAyqfEgk+qjIR2ox53UMxtafQG0f12WTVNhEeIFj9zcUqOBSX5d0kLhJaXXLxqPFA9dP6NvLumDT9Go9VuuNiK0biyNYhXmOEx7QN4iNsuriaP2QuXYC1TXfXGwYhoCk47mfACB9Ih7cX2HdSKf6J2Wl6+WoC+4L8cgBDyX8FGC4a/ciiRN58PEjsOd46EVqJHMDPaGjesgzv9of6cgqszEynxjWJYiYJF+ZsUz65riWmTnLYRj+MwDcXrGHYfHFP3n48R+aWVig573bs0ZbQtqh1+Z+clwv5LkNoPx/aKqLGBPcSaTHBD5SojpjjaoIuWWkt02aKJkHYJPXAFivtF3sghZoBG4CtrAgGvvFLZtz8I5r2HwxhfIw8b8Y4a0quaxQLasXlG04DcJJZGbWVsTn2v81mAs8SqhNhkj4h1e68UfXcwSFEgAgPeugmk0QBJx71v1TD+3Zsy5DsTcnjbpes1fs/q9k5E6Oc7LBKxCQhBq/zE6FPxjLtfm6cgqOUb6Bols40PkJGbSAAJdqBSqPB/nl14FdeUoJEZoT4FaYErCcN7LB/Xo9zKHbhTEliv8gtn2FLdh+5MUFjLpkiFGFLYzWqv5yHahXxsqzLB8rmDVi+kIsKUdPb/yTRliWFTsa/QuYihoCCVbNUukqY1gYyMeFwLRw8JEsws3OgXUu15sCsw6K+OmsBLeEosut/+zvYWxNGN/DJI0LrXtCQ2pXD1tlYXMUr4KKY369DCJxt3Gkn94HjUbtji5sS+uAF6ce8kElbsOvcVYnU/l13KxM0AWLiwFIdL1sqMHonur86ESqbZ0DOrhhfn5pd6JawyEIOW5N/IAT8GYZkKwJSFZwudx6bglOglCeJmv8EkZlSsCE4CB6r+4q1akmIPjIl1cNUoPwmLOc+Ohb38AEM/6P0EqAkrjT719V1bzhy4uu5YDqOnu6k2w4ntokKofRbFhcQN16MigAaSEz/8AC8V1N3s1ejHC2pVRpwxH+f5GSkh7vwKBnMHYSTwcmqLlUlxk0tKEY3T6fVhyv2EQ+CnB+XY01DWq9w8AKy8Cd6x/kXxRx0BI/5cF3EGpJbW8JDczuotdYrJtfEf+f+zq2h9hVc0IssoUs7Vod5e2mbnwjAEcuzROKe0hOqJ4m35gjf6fdTIMtsvVoaN6Hb3hbw9brAcEFjt+6hyXqdcmtDFeIgDQDXfSutj7nJP8f9EuTusA94uvXExfFxRDF7VEppmR4Fv056FU9uC7pdhP5mMdHlGt7gbcHn+0To9Qgai1DrEyvc6EH7lqB9kxUTeEbf0rPIk6+690kkj2FcO93dcQiAYSmlJOFQyUhyN/N40XIYMLP/tuNYjEbvlBIPhoT3oAkjfqhmVr3kvwa/cGaF/3e7e25w08JluVipO4mcbW4HvD2pJgY2zbpEC7bZag8KaKuhIvaHfV1UY8LyVLDrIH5a2YOdW55Ne5/ZkoEIWeb9fEETL7lGLec1W8oRNEvIGbUv2wAhk52xCXO5JTObgB+i9w24c/8jBoSkVCKBt83pnSNDS8iLD+iyzEBqIPz8+vv3E1mR8fEKkUOCzlgS0IonrWd2XhPoF5uyRMflU2+J+z5wQDk37NqUJr8k1FUO+FiVPp6D32i/YL/XOHH7+qe+gWYJYVJ4gQO4/F6617Q2Cdp3NRYRNyJWSG3Ert73ZjabdgKUNtRp1ZwWX5bZ+X6dm4MpUDa/jzIkRe5mNluTUEvE6WkiL8Hv84ymqp9d8CdWv3DSyfaz2bGQ5cSlmQohV0htvWBU10U5MarPVS1nXO3xGZw2kp/chcy73X1ll3nfU0pRUSH7oFP3lseCopMQ2gRn8rwgwWSs23zt1LXbZdhQ6ItjnNjqEaFHRmpzw2NLKPjG2lvt4ohmy35PbSzYk1BLbek5DE0L/Q7eUjaqNYSPgXdXwpV1T2iFUUyYgp03ZYuuxTHw5RREAN2apaMKimKwvq0RhtlI4iRgyO+cVnIfl08ySNIW4mFvAvtcfQWUTOA2fZf/J1qzCOjgB64ijxD/yLN2stQFevrWzzcykrXtPYTMBbuP0vVmGrvC/73hmcmW2nCe/QE7EuPfja5Iz9diIRN8l/FMzPV9kh+UyYQ+kdQjQmAIGJbAeqIcJyksU2iThbu9jmdx8LvnoHx6fmjmNfqs2LDI6UQNBfvEYbUO08e9GujPTbX+mosBpAF/VmJkTQkBHorJjyXEFgSjbtXnjEZeNoe5LXmjSp4HefTn38whv/w8xn54h50y+1L58QLiLLyPZQLOLoFonm+ecL2pYJDLN0E9eSDYKO6dv3V+rPKA2ATTaiX7aUxnP7UDuRHUaWykEFuT5RFL/Q/kqbyulsuHw7f20iuoCpv0PUD+3iNygOd7DZWxuKfZRdMuIlk5ek8/iRqt1MWktUZ/Q4utC6w0Sl1SHqPZrFP9sJ4w2MhoL72vc0j+4JGusoIcgeCzKLwQxXfPMfj2FQWD/LWagRD6GZE7qbR/RqanWcVe2P4/06kiNlefMfzYwNJnd37STEg54YlGAVQE3oDZoE6Cl/UEI6beDtYy1YufXSr9DWVeSDBM/JwlvrN3YY0UhUKP5tgoUcb5AhPPjbwSzzyYVOUBbqt6rMAsB/QVj/1FfIBMvheJNFt5OU6C+BmiE/4wMUa1ES5ni32yPV8MM19+CJBtmuO1AaRlERU+tmmFhhI1tPaUNAHmXggpZp/a/R1nDa0eg2CUecdXWuIo42SfOrb4MZlERGKhcZQcs5g78xEAJderERFq8iYqPeLUXgCWcGsPPIUlU6V/NGQPmyrCUdmvoc+9Q+cXYfMngnpLdBSoeiD/DONVdhMa0FjzKbTd0rGZLqLE+HGM8t1rb2HtocmT336y6kSqaZ7G71pdZ0LD/TKPh51IzDMEilnCq9LlLLW3FnXHbi5V+HYds4O1ZvseJAilA5JOAsjJsqmt0GYNtLfKQYUQZZV9rQJjOU/zw8dD7o5erqSOi+QvrsvozPz4+RGYR0BtaKkjwX8RcMnDOpjxOgUZJwk5/2I/2EvDuN4/cBAAb4cN4OmC1XcAcDW285tMzyJsn55ipgWTyv8ZY31wr/wnpB8mTtaTAJGz31X8vUlRHQqe6wUNRToCCmEC8FAirMwwuhn7bb8y/WkD0+MpZTIMp8YDgZWAUm6WSMu4+Cb4o0e7xoM2koZCFzxbM4xTaaVBt/pRk+0eRLKJ4YFHyCMmYPzhYGX3fLXduHq546CB8ibuLr0j70WDfRGDReDzIb7SjUm4/kuJjGpox86qgh/mtbsalbTrfSw2OjlqPWQp8Ca6PEYm0AFiNLGkFpAK4eUxtQAGoo/4okTVv447qqsGcb+GlTxGhGt6HnAiTdDJeR4NUxmp8iO31XSKcdqG85SQWwroCgZTzunbqX+jIMnn6uf6OfbNlqY0c7RWbDVfEmW/h1S9CrGezNXkAsRgSiyhpEHX1au/BKebfAVb6rpQewQPJX2DdVi3xJhyt/6/8MEtp8GKtVgbrDiyN9LVL39OcwitC4/fRH9XTs9TTJgn0Ojp7/CpakLq+waHIciMQTKZjTmO3bBVA41T59CAugt9RcEVpbZuv+e47Xa7+ky0myI8hi5XGiDx6AO/heat0QgNywJ+Ev/ojxctEJ8hL2ZmKHpbBx2AcHYDki3zWtEn47xEZCbifK15Ah/QYxw9G5LLnNvEmUjGFoYb2mX49Q8NelZpeTPrhTXSR35wC12NfcYvfwoGkSKbYCShLbAOWoaZukDMs4IyhHilI6z/ND0lVIygMT3tDW8v1r5iatgWOCgkK4fFznS58PcHQNr868EAmF8yZPAZiva5nXv1as76Zz3p3I9qH6UrOBc3WzsfP4+2Lw/bWZ2T4O+4XQbG1isoeXLWscF0WKYMxydZa9hBCeW6xVmzL2bbp/UeIDnl00cPDudNJFo3tKdiYLuDy4XdbvJEV3DlZuJyh6ZSZaxRgVJyYvU6UOYqFT3OPgiXwKewckVZ2wBt5/6vSplpJ5AdxTj14DC43lrAlpEXnfT7UKzib2YLOgbzODDXuFfrGIHqYk/H9QW8xKalsnQ8NHIzTbCnRz1EBISdLG/Q2S1x9+T6wmZAW5LRAfS6ND+w6FBDHKfH5Dcvi5dInzOLE+Y2iL40oRe4xWHFLRMMDy2EZJEVhbldRCFZFWPUotuLHlnJzPRU6cYvwUnn3MXpKqBmzSc79wiXG9wnv2+9CJKXLMKu1eLlsG+ZYax8zJGjKNzI/fT8Ip8q1d8dwNN068b3GKCWe6oo6QLQTQilC+LNPWy5tvbsDm01WDNQ2bB97XSLxMt+8BIB5tYZ1dA9MbkqYjBT2myALafYeBq8fEUBF8kTqQQljT/RyvKYy/2JlQbQP9fuyKHu6K+9FNWeFSbfMqrtDAiN86VyolDP56UVhcXG44mf74PWr52C+oWrozsbJieotm2ctnl/BvJTrf6Eu1c29O1TuwX8j2axSSQHRmwEsvOFHEW4BpWLL1+4o165ic88nzDiM90utwh26kP3++xGzEN5Vhi97c7fYs8Bd7oZH9+KHFaAP3qyN8qDy35HmFKMTwvaDb4+oa85k6feFSMqQ4qrN/0A4XVe4ZEsiJKuZ4dh3lIU52DHoMgVZxE+cJlL6ikutkTK5Y0ZG5Phl3lawhd/r2uxx6WUtX2FkYZf5Qt8elEtR4h0Nwmq+g1yCiPpwkjWLqf1t7P+Duvyxg+6a08r0n/pE+Qs0afibVAtmRURWwXR9lIf/iIntdZBeQN1D2j7wKP294ZK8XuVaQhqEdnq5KKwRV8kVpWeA8vervTaxG6t7hJmtQj0hx08yh5uwcv+mJwxbLnWgN+6dkP9W/1zBezRoR6x36VdXPUxNKfq0SJQJfQs8QuTwthJxxPpOvDeGEp2uhKUV1NNf8n0U8dJ15+iMexGLdcvsaH0B2kudHjewjTfNmpXycgJ0PeKDlCNTGWUHib3pJY5DDojgtJ7F7hpmZyOPD6W6cVplhDeK3smTj3gdho3xPxfa3nLHk5FoeN40A3myCyBfxqPQk3pmoyLE6eWUxqkg9EOZrKCB5dBgxzQ6TAFVYcfX5PlTbZsIPF4ESc0kUSfqOoYXVC/VL/G3ocXmDW21kMDMZB72LPt4z126ymw8LIqtH5letw6zSO5r8opupvJr6RSjbNoTp2pxINrvEDrBpVFsZknk2xZvtEM2Q/Prjoksciig6mtd5dLHVSdaUV65oEWlfVWWaV1NZI1daoFbU4jQ57ivTNxsuwGG1GhzR4WLz8I80b3qGBKi8TvpG8p0YAmWSnlX2FqGO4sGOuAy2GC/ExzQw1dpUvxt3iI0unQxV+3/G28RBcAKI/hBAGbK0IPMeL3/otZnTncVcScZbRu7aSrjj3120451Ap7zZ9YnTgvYdfcXtKwIUkezptxHWBVEvGewUQm5N/zmj02x693KKe02QlNfehel+SpmaiEVe12h5txWKIlv/wBL0FVlAsB3DVQU3mgwzTEh+Z4/Epl44e4Hjds2wdeiP66M1fD5NdrqtCbDpRqPESPf4u421oSNg2DRJ/HUxUEzjJp16x8D1zjbMLPEs/GbLNSe4QDAyBRnVuj4qfH/rULaE2rKkNt40tpb9GzEI+gJYw3jgtZ1TJaB6pwmmnNr6meA4iEINmEvHMQpErhUNmIeTfd9oqpaM9TdVzZu3MP5EtB1pREVFcIHJYLNxC3RgDa0A285YdY+onY+Wob9H8c/S+LY6EY93IYpm3FDs2jtbpuRFt6r5N8usShhqaAWIjUnaxqIFMnPivz4MitmbiTlK11a0olLQwggZorGxoaD9PVv1A80buJ7+uUtr4zdGxWAn5YolfhrTSHEdKehjhxOpnOGzhGZBU9jBV9DahiLY2v0OQSqTXHHlA1e4zbd55LgNt5LBgayqKEqi4SaezmnNOvn7t1UTn7yUywau74sFNzjsNlVr0t9i3+rtDiTZHEPQfPk+8NB/eHo1Gwv6rAlxYFYvl2PQCGuG67f0w11yjHNQJI69SDX6hb3oQATmMJJgaxjOfd+qWITGMLHiUWpRdDMirOH0EwGuGltc4v9gIjs1eimMBjqstW8zIWWFA7ARmTdoe2RLycDEDBn5Q+o8dB3sD/hNid6oZcefxIcVm9Kc1R548wLA2Ly5+2z2anzAxJh8vh8hMYLRLYRVQPYrx6QbHip24rfx1swmEclM5gH0FDeMgXvu9Tl1uJevPIeyl6rpZen2pZ0NqpOprE4lZ9SU+ORxV7Mzftt+0OA89dwVKvEE/SbBrjxfj5re8NPi4LSofrxr90MeuOH/WNTquxM2nhcrST3JSYrPq1+StpCahmjMLIHRLegL+GVyNE7XhPLgBfEMWzTDJ0su53jBNXOdA0LFGKmE+RBoz7JSaEvkoItFT4dQsCscPlaFEM+O2ovHJk9qbETIpY5QEzccAk2GJqCqIO0JD2ly0wQ7K4t7f6ht9V8lvYb2Wde9ejt+YdmbdKVfsr6AUHKybaCU80VxCaSZS6LR0Ed/Ahl0qB7KXyTy8If4sLqXgxvTgJIxvUUMHQ9vQBKaNMiJv6iNZcRq4dGAJIjDxd0Wzv1L+CUrOu9oYgimp55sYT/Z9sDK/CSoOKjUJ9XqbYBjKN2zyqgcPfwPAKk6u94n0B0silyMWlAzBSMrngDtoyDP3G2PYD4vP8Ru3APEdtb8xnHj/PysC94TXITeoQGmy3opExrQATDWtNHbxiPH7jM41Y132ZwKdJXZJ1uifQ6Ml+XOK8z/KbAR3Y8NtvfjrW7/EL+9PisxTbkOJbP0kjS7pPznIPy3FQXhZMyoTsL8wrxB2RIM348RYN629eVEJ5xjoNj8VoruqD5iGZRJAvsg4E5OsKeZ3kqUYNoTdqwaG9Mv/gvQDRTTKGALb4kRRvXFDb9RFPLs042UkRRdSXbg7fsYYXI1h9g+FGRHuQ+DPesk6P0B1048a6nAMa/f7HP2BfUHQLDEkZ+Dctz812IA1v+I/c0J9+k1EUZJZkLDF25VKZHr2dSLmtb4TQqIVcvI2oQV9SpbjRLWpoUhUCJ/QypZb6he0DOHfo7BvBUGN7NVFJ5Fg3n2+LTlm6aGzHAqRc+DvW0mGudAIaLQHfeGzfl3zJ5ow9MqG8/ZYdWvzp1Bc9Fg/pURgh5CTm/4RoGeR8Gal97mrwy3wwVn1A4g2WPh4QnBENCzYK1LQLqhQwUZRuEqQgZPbRLFY1ZLtPrpZE6ng09fuMKB75CbXxqF34JBDoM3Ga7udfqxIis+R+LsgDoaFS0EHO68ytK1g6StDKRNcSR21O+RQUEd91cT4lqWcQ+fJCBNCbskUg95G4xur9rky4RNv3Fk3Tlbqru94QyLLKAo9H2SlA5dbem7kDCZ5KQjbQ9d1xJDFYdGHyq5iGNCqc3N8HThI+v7OAGNF3jahpzBbScag6P+ZXHvZjlirOOeJOfGMTN0hUKSfn6RntQCjyiGpbXTizM4HzF+2TkTwHkbFVOImNFduzFi9FVEkS3ciqxdivf9sJfYA+iLi8YO+I93a34bCaFVb9pp8VQQKuaBz8MVVuu71qT3jKipg2UjCsF//z3NEXBp48kZU9x7S5SrgseYTuGuo+XLibJmXh9HTZ7fOOb/unXop1IfUag/TKkLidRrkIScAn/X85LprafPLTG3zsklyI0k5Zk6zCTWAzl3szTyDt5SwwD5aMdQH56+AOnVPeeKzWMDNKL8Fc2KRkr0yTQizLpEVlqEEloDMb1xPqfHTBh2iHFYHROCMcweeYTS78/8Qmdh76od/Sg/odNNJuet2/djqOzkB4KEJcV6ThDPkqKp8CNHCiBKhpAuBPstC7lYI6hpuP56WmN9p5wUQsgFmXazMmG2zPX6dAhZ5KrMbR7BgcUD+MS1DrMJeiYUqTVAc5mSYF8NT/OvCFHqgsN0jKPVVwEpDZ5Z7JK/CUCUz8hc6SjLY+P1YqVWJV2TjVVgEIMMy0Y46ZRmYnfVvNgcgTVSabs/l0cxlrIxoGJqyN18dGdL8fMgWpjVL82+OLOjsA2bgRuCFjej6DTwmQnjXj+wSTaaX+6FMXAzzxCqhnsiLXPoMPA45iLPxmQy+ebPfr/Vl/j30dM8KI3HyJHj3kpv6NPTHRqzXDRJQYQYlZjKRnUPTC55Z2Tgaffi92fvV8AmtlediskLxGgM9D/ouPWB9Rax+LfYm7Uj+Xa7ongQg3LA1vZzufHBZuP6WsmzEXe+kMAQfLvcuW9OMQCX1fc/jkxVhuzLBslWIL/Xjvr8mbNUciWsYbOkqeQy/C5aE5fPS1zllXVBtmcIv0FD7oIAly5gn4E6xX3QVRjXuG0PXoywuVJth2xrGEN22M2etxIP7KzNVzb3gwAkBkr2fDM1vckZWRDvrt/g8LslEk9QK/dp3zRnrCUpE107wTZ4F1IPdlHrBdBbn1CSu0gjpW/oG1BXPsuJobxDDFRYt8sNDQVTTfYgQ3o7iwgnQIDJPAQ6AsL+MzxBTnp+hAg70eINDCOg5VJ4LtNN4WDTLshbqMUrOrUuBSpyLzKXySpbwxi84eSLo+CTkz6FJx6B+XAHWgTBdM29EZqphRZQUlnP9loN2NTeOR09iBsB9/OZBckuZHdlk4o8MNQ9EGKH0Fb3l0+p1ebb/i/cU70ExJU2kIbJIZkPEPibPpBoXYKVYt0TFVc+ZrloI4VwMuFuEp2mVLy9iqZf8cautrn6CmjLVcs4GKUHdMIaXkFUmmcilOLSvrJyuktgR/+YdksVCHYNV3ml46PW/7kEf4EqWtAQWDOExKsrFoJAdE4CKqkjvFmsIiQ4HP8CeJErbQx84TBA2waRw+qRe2ftv5+V0v6cw4VryyFpFzMO5hQ+s1BLN9sVTgx+rYlUCEVc+/ZswS39R9kEu7bUv3OldwOBNYCNO2a1hl3D/V9BFqYqFexJI2naitHa2X1wTi9dTz+tGS0rH9tGN783G8jyyiz0agbDcbVxKEGegQqC1mdy8dI5LEle1u3nkXOGURTlGfGz5rTJJyfcKE+ZgX1C94J1wRZtVlGuDudwQkRUpOo/s7jusyjxjR7INnM5NbQf3cgTaw115xWOmJl2K9XKWfDfdp8yTjZArjkIdLtAW3dtk39e8EX/0M39w=
`pragma protect end_data_block
`pragma protect digest_block
72a5d8149d4b148c58710b7dc1d6f6eaf1961f546b404411b47f936c3e66bf54
`pragma protect end_digest_block
`pragma protect end_protected
