`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
4kNd3CW8eS7kE6oze+g3MZNVt0frmV5EWLLexO6uEKdUYWgykdcBfYeEiLVyiOo13wCn0qwmoRjnZOFPwhXYN4oPcotYxiMhetDuNTCXfo0F4BAuNQ410zMcagZ6YZcbx3F8cnnIeZytTbTXcb/dI8HwqCOZkORDVwrWjlpnbpv96jM0WLlVpW/SQc/5A32c72iXXo+UW/EzypfzcH+lmUFMOi3VjTwxBQ+u3rGc6Fj5Yic8odBEcCQRBVs8FoGll4eKcC7t/MDYinA5Mhv3PyjmpCwbamFTUimmlt6I4eU+Jlx0rtDCBe1I8RbqEQVEPhnGUFJQB4tqMzdfa3DUk2LR3lMT1tFUbFvL6/gLnqrNkOX2GLclf955h1o4C0zYNMaSizE/KRyai3QvQgldHrCpULF3sVQEElIGVjfaYqUnGK2Qt6Lci9aVtvFlmWtuCFLah+FBMag57PeB7X7CZgmDDu+fHe9FHHlchERJ4ayNXiLdcjVHLrUZjpNveJCCi3Vn2573eSx1pcbNoUAJgvxaZ5HBuBff6AfVZZexNq4gIU1OOR9jOdfeFPVIVsxeGhXbZEjD7vBh8nrJlE85CVGIjZMBSxUa/YfV0TNIqGF5W2k1pTYMq51dQToaexryVHFIO+tr3RAMVtfNjD6J++sHD+35WSJa4g01SZhM2kcVcU1GcEo9IyKTmj6T3T902zeOK8r1h3ZvrMs+FsIjqXdmkNgITyvVgq/BypHX2VDHZL9pJRbTgMI4fheoi7KMMEGB3VOREP+GXpzEp4e7Z6JT4jmmVyE7dbBRBWUJ4BhDYqokdZhBARkjmuqzURZ+XvS8Z+6Xj/llsjCla/OX5LRUhlH1iqoc9bCK7v8diOa1SP0Xyc+CXZmXUCd3uwyCg4PQx7PzFmr35Kw6ZdtaUM9P4ZCYkaqwUNtUyanZMbz23IXxGA/Jnbi/UpJWDDGQwDNrYiLiulG2LmYGbfOhictDO43pFWFI0329Mio7w2GTn0Y+dO2pjYsclNFQuc2MW5RxzxtYRFvOriOiMhSqj04mdEpQI+mZVXCftmEmTTfKfByK9idP8jJIXtGeZKwrhOyrzc9x1oAIz3POygF2EVHILtLvDXNQ3N3LbD++E7+u9B1fPCt81ZQyu4qR9z8Fw//5/De0WYwBujWqPMFMUTOjEJ/iX67LzYYLVCm7fqENq2G8IgOIDH/tucqyUfht+jQer0VwZbh7mfIMbi3ATsjfuPlWwqt8+ZBLCXyMZjnBK6HIKY5HHmGfDoIanVvisHdmXXLlp+I9OKWZZYTy9+j5Coe+Jiw6ot9vRiqIXG9H8YQMgqaoz6rjBl90qLbPjR/mJIWre1Kca7lrLlg4z27SqgugkQITEI5cGbeGAYOtIYemhTdQuy8zjtuOJWvJhNST0xlV7KF7tjoMrXaUKeBsrthmMMRWiwZsAgOcTSKhIbPftwbbh+CIczpPPPXv/wH4nNVdpSNRpou7tBCUByMZDija3QJYy2gp/muT5e+ok38AcoseWMVjOljQIQ595vvsE0n4CGR1LjhnlH64C6etsaeuTZAi1S4nsd8vPE+N48ASfvdEs6Rz5YEcPHkNtxcLtpk0IdqXN8zx3IU7uJOVmfogp5dqh7Gu/eHqKh/Qam3lcNWMqOdDSwWSUKriat4vGYoz58dZcpL6MdKYqlkHXFcB/AG+/qsrRvvNDyMykNfm1vw7pSe5mp5BSs42LiKMUJZ4N2nuO5ctHbwN0Gc7zoSx0e0v9pe3yQ3RQavlZHWjQBEwq8BwV0yAgiK45aHGOzQzG9RG7sXXfpKT9g8UN2apyv6lD1lEwHc6fIPBiAQQTY6Gq+78sPTVOCaLUP7rq+MrCotKOnHnKINDMVhNfHk74mgSVgS9IiqBswNp7V2ujCT57c6Sts53vrpQlMDFzGeo0RI8pWoje21rK8eO0cGbztUQKJvHfu105Slsp/mMI7dnT2oAcn2lIvx5xVX8DSprHkPN2o0aipsvOunyWlYJRaoMRZkMIdS/OA1QXE+zJReLI9gl2iX0lzTOqh8vcKD5sVBoI9YuKTb2kU+cHIiglRqOhd47KzZubtCrCiTLLe2CisOEnl0gkJUBsAgOYcHHxpi544HhUfrfrrE9vGK5vBs8+pt5h7vaKm0ZjJAGwsSrv/ATNfSXrV9H7ncHthkkaxIrBtQZBEFwJzYS1rSb6cZw0U8CAh2JGu+DmT2+PUekIKxORMfTmlCJZdR5CToY3ILZsyxePf78KyG+Ut/GMAofD8IqkBppsIaawz2o6Um6FJoWQGm+eAZUdporZ0a4b0aA7oCV4X9Po2s/+HhAnEltVIQKN2unH7x+9Zd3dm2/uJP/gudTiGF7bs0TZKcqgkTmbr0nY+4d7fl60H1CyrGjakGgdvfjwo09P4QQZYRgW6683N/TYBrh/T/cS40Io0W6KMYJPBWAnODH4etk3U0AvECAA4xfPCQUg32m1j67RzTeCXl1jPkWzD7QQeURS5AOle+TJpdTysizttepfHRKfYPWSu7XU9parEUAjfUBMZjR6PEm48+JglcqFbeST0fUZ+qHX98xf2LIGmPQ57wgUsEjMmkGNLn+TRIl3o/Nn8/S8kcR9ENvBLKJTBzJLtOlw3azsqvcoBSZqTChSYBWn/MkokDaNtBqU1oA0DWB4owy1PSFGqn3gOah1+/2+tIzM+TqTgvHmAs18Z13CKM0U5jpezrdl4B/ZAvYdyPRcS+ZB93d3s5/A/tTWHnl+OmBYaRvT1x1zSPp+NvidPu26OoHMjgJ3jU7//MgPgGPt8IHe3MtcBT/7kaV6sbDJgtYWjsxBYaT2n8MaNUTa1yLcd4eLh8vunl6SCSl3Lgw/5e+molkkZFXw2cZ9z6yf6TvYVUkikMJv3ubVzIoDdK6aCrjv+8fScXdagPR3AmtiG74rCrmgwIlYd5isZgVpBvvjRnF+V8UXsc3D+KWC7tCG+CZQFbXDN6AsuEK6jySnbDkUnjMfGWE62PL+pRqWeWeHmpjLxskE8uRmmCTMprd3jWw6hOPbH9xxibseW6ILTBYiOuroG6irrWXqmVsFahNLhWqJEyG9iRqlbWra+bXy07CAdCVvfRY1JPLv+squoQ50CdEctMCj6hvldoT1gswjO9qD+nPB9GHyhU8o2oogKHupaNpqZR57mTPGPHTRhxka6TKaD0y6T61Hr9pMRI5JHdQCSjX2KT1x/7FrQh4vySdShhLoEaO1IbCTb8Aw4ZT9BX+u+O0u1KEZooMMs2TZl6zno247BP8QJTAidqsLCfM5lUZ3L3sOIBjUozkaDrwHK84mdW3eGSjSxxNNGYrkxENmyIT+NpkeVhIn392yfYMdI5ETTWO7UuG3PdTNZlD8+1sSxl5PMWzvKIUV84q8m/VdRPBi787MpzAWRTcNAVspxlUqsmwjBiBvi1TRDknIXFVHdrZlJWLdO0SlUMUm52H64vKEaxFfqKiEE4jmr89wd3MON77ouV7lYWr80bclH854WbMEM0U51NM/RtMv83HHsQ8Z60vVHP2nOLn+Ho0iirGQsVTgtZr/IjNgI9dhjvaCwlukf+nH8elTJWbnJhgr8V2uxlYq2EP4Ip4s4vuzWv9pJ0D92G5HD+pd/EF/PBA5umGSHuhAeDeLcKraVhAWHXVcoGNu9UPyxkrQe5gODTxG5bZwfeMCwvJXkBKwE9cgb4AJN1AxuGk0t9KqOrN/SvX2Z85xYvthaUG97dG+tRuO87KHpBb7MEk+TFhz7ZwR2M5LZ52kqMGFeQhPY8ZdYhLgtAy7ShRj1Dsd4tnDuk6BKAKC/RIIIQXwYvZddujywB+chqkxXWChUpUVu1O6M3we7h9f/KoB9BFrcQ8ULsXvA9+p71b/+VukHST1Fg0mF8W9zS6F06XFZjbDJyvdK205sUetJ4VqQUiR0qdIDSlkri3RQAvVNoyBJY3geUXp0fWos3eHJrPboCfkYqpD/nISCgv8Yp9TdweaFyeTewZDZ8SVCVeuIxG0GMMbtqxYGUCzZVLeVFz36w39f+sRmfQbgCQamj0On2U0E9EnLOWMHigzgay+lr1v0VvRTO0/x5yUnJ0gEjmMHHOKPal1EwDNRatSDMlyAYWLF18a3HWSVurxJVat8ozzAN+GaWzHY76AEnNcsADNZHLot7Hw90bHJto9YX/nB8Sby1lxK3H/40xXG9HUgcnez7mWPqZ+CUrHnA0CMErH9+rABBAHFhJysbvuBjg9WaEVR9s6WHwre0GC2tSAG/OzEKMGpcQS2houon2DYcJzYDoxLSQaypXeFL+9ujb/PTEXXpYnIQfcc+z4r8k9SoXbDnMFjdKAWlaPCUGoyItxWvxwWkKPmHb0XpbkVZw/nm/MhTdJAoURIJOXi1+nCyEB7yo2US5TnZ7nRnyZhako8lrdjUyxsfykzO9wVwOrqylOC1VLN3+m9K10WrfZhzenhO1BuVzcolM7NnGrJmyz5zINdV2rznt0dNIzmoxUiZJ7cKJHIct+mqwQi3hVZ2wAlWcpDfuNn5bxGm0b/HDKOCoQEKtCDmrsM3G6FhodVcltFXmPC9sWsUXmjDPpT2l0yb9BQ/rqkPCeZmsaLa84IdEZ+vPcalqiSMCPfcDn6JgpQFd6lC0cBGwsq/zwiv/7J1H4RZjq1RkmVJT0J8jHznEHXeQwH6+VJmeA8jKs7ML5J7za5y5LvcjIMLDGi8TmURUH7dK1FB04VCOk2MRk4ZnrTD7oH+9pEEC4CdTXL9Glh7CdIgUvB4NrpKdChO8rQTNFzIZKl0Lac3o9FYWROuTj/jlMd02lg/QiFIiToQw2cTukw2A68ORHLe8/J8uwMfIT7rplNv1Ln1+FB+Msgg7ntTUdGTVNqKRIRCXEVARSQ14I2nK2LC9hB4vOnVjJ8dn8GZeGf6xUcUoQBCC3YlpSH6+80BT9lr8aQM5Jv2zjFqxFkDjRdmhRi3FeuEo07UCzOOYf2yTyF+mZcETTdmIyEjcBz0cjR3SwX7gdzm2v2ZxKLLtTG0o7GEjD8CJH093A6vYdSAaKclG4CWntldH4pCSAJqVWeQH7DMP2EY3fxlotH6jhLZwqdeVy8wzvUFHdM5588IL3sY5iO3Qhpx9AuXa0i/3CMytwwqKlo2THUFScwuCCiBkfzhNaSFAwiiWQDdlKtKU4sHwATPFNK7rYAz0S21taLqrLldOkcfT3OG5jFdU1rTUdyy1UNg7rTEQ/HH7d4u6upzk6rWdtQBFjpdAX8vXks81+uo5qbQhPWvbl37vpwvtucFDNI6Mr2QLE3ssOGLAG8C2e2fgvIDY7lo/bdAmH7mzxq+9HXV1mZzMxytayx7sTUBLQG1/ej6AoQSUfgRuX2ukmRMWXIxlwUaxSE+wF7fngs8aH/HH8jeLPx3noys2D0mBwJlmjFjS5h8cS5+zTCQqR9DuMQ6maelrHtOSoZsX8lgOmn7t58LUx91geNvJhIZVZlVkDeRcNfa2TGyqCjWb3j70WLTnf+pfOBZAk+bdp/MAtTMGA8OYwumeb9X4t9XNwQcXdVwE0JuxMEnjyglG/VaH/PKcA5tKGclP6pVEiCCpFL/zFcOA2FRcbEMZ3TAqRmwkLlvxZ90RsyxQkmrWErH2IdxeJPeUSZr52D+etc8SwDFtfh1xMgmBcnImNbImdX5+0TVLyVuOa02CMButYjRx/gG+ONPDE5avAucDRlfcNAG6WgyG4aX8FTvTyWypdb9ZxoDqSkZNOP/UkJbaObO3ICfn4e5y3PluQuuf0l1mzhGdwSLaq8NlAYTkr5kjX/j3xG5TOHtZVYsoI+pw5kyr69jQ54Md7XG3xp/4O1CmLzSk+raviIXpPMBDSh9v2XtqqkjqOUeJiC5z5NMAU6X8tjTENNSM0trngMHRIzO3gDyIsd4wtq3kuwaVFfXEWRV4KSUZ0PdPH5Rlqd+7O5n0o6whBbeyQkZXA8SfY1JHKy/i03DkwYQN7Z696MkrMLk5a5uRwHDGT2ixvsKa3Gt1vvnMVC3jt5MIT2pU2HuAVkIcnTfonSt4lewbN2557VBdRF1AL7K+VQmaPbVSvabSlYwzdLd5xg44kStTd2hi+UN33Gy6Jd87E6Y+CbxRo8qIwsU2mUjtPH4HLFqWABb6xJ6mn6JNjbNrIVWbp7UlC4u8cIFjgm3s5szOPX4yx4CC6S8K4fy7q5y9GJ5UxzfpG3kRDmifpn0zuwPfwuwyBUPqoZe51nNnCox1jPJGDyg2KjZLAiWsOY8YCYdSKZVj43Or/dgu5cSwHy/7jKXvFxDndX/R2jiG3ye+Ka9F4gPOrysjO7O6/DhsR3RNJ6xD1NUAGzdBL0G96yVb8UnWvX8RkMiv6vwvycED91ir5AdeIaqpVq5Ey8OIsLAqBsSRcFqpVeNgO7MfQRd7O7u5esRb4xwPfrUHkYl5cMET3xRD1kpM5JtTnf4M2skjorkBF8PG/HZHvBuXlDR8mNBAtIojcGgSC11YcewnMqQSSUggvWYlrOkKEJLNRYTQUnoBNOiW6+ppBRNvmK+zAIK7sY4wtRtxtFv3XkH5x4kcSyUohAy/SQZa45r91FpFqsziNTTwBJ8dBJVbZg1qNShWZvb6clxetetoU+2LBmlcBXQadTmEhW7XZYj4f0CPFYkWJqL7RIxyQuVYbL/27Tt77GFfDzjKhNGnZgvMtJAxKY1dr3olzwq7AikrQYwTKByv8E4N4c6yRxZARYlUc2M6mBi3El6+nxX66+3JkUFMwUPgykuZ2ub/kbhJfF5sLp1czl4KWZap2dvLxU2Yx/5Yr8kG/o/B4eSTtvLiS3PpppFITohvFuQsMlI6PVxJH5EzFOpe2lfwYVYHhZQe9slJbN0RCU/1JXnF0iLH3BCRGeVu8o2XU/lDgsMztskZT0XCEeSjJADmWPJDx4ry4lhT7P6w2wtpzNTmvkyvgLfcWEmLthdUQUYj9syYX8rIY3KpQNfnxuVT/qZ6rtN6tMDT9YUZ9Dwm+8IUqfjAJPdb+ma/70lO42KiY2MgcplARVY+4LodT1QH3GoqNN4MUwbdkieeniEBh7tfFTlO+bnBg5TYQmu03NEKNXX/oBvcUnWcKT6uT6nyht1CNWhObTO+ZMCINbiJCPnfOyAcztPCwKpo3unoUGnG+V27RPkwzSbxY+uCdI/YaP1RuobIWlN4QZD0Uczp6zjVVL1niNdW9QBxmGZLQHPY+Xx6iRFWwuiMkcntkox/DZAXBRJu2+5FOzVH/YrOIx+T10D9c/IGEbt+zArdcxZkrBH9Ghw9ZTpgbOA8cBgqfuRJqIfQvV/k3G+ziwVVOHWhVXAgkIqJcpCv7zWaYIurz6WVq+CCJTKJT+vs4LwUpEaruuRyyKB/BvVl3RnBUZRHXcYV/yxVlQUBLuO1aGsFnqTKOl/AindnXWznNiAi/ax1D7jgJkgUnTlJb086vjQ05OF35bALROKcEyrYuTK/DuOhdJZvZ6w+dGeAYvTwuQrWr5CPe7xpLm9fNuYhlMVQ5YFkQhnsBnE96wE0YFyDs/VJR5BMBHmsD+ywPjBudRTMKm0pQJkjCA1KBcitBwlRC7THFAIujS7MziKmRtBOYXfRoARL3SYwsiLXR8tAeucOLS0T0UbdN0YHi3/x0tYasHJ39MCH5HYpQsFWbl7jNzV1Cn/WTSwWFaeu958MNkCq23Pfkq+gZWETCQDqpjhIHdsoLnqRbia3hNYIAX5MlbyRaGUMjEp2IUv76iO8OFdG+WoVtqNsqwG73lIyLmIY+ursCFI7PH18kqlif6i8nRmM2dPXEUmynofH0uP3T/Stpa5kN+GsRd+I50lQT4iX2bSSexfT2776GF+8Q2YQSJscF95gql8SagJ+SqLGz1kQvJVHF1tUT7juIxBWl8/AOiNbAKd2H8IIDJPvMTQ731QHInCQ8D68jymOQNbL0BYswIxdkHevts9rfaUAYP2e9bUMP+Jah0K5uMYNaaRul6KttMD4yt+iQOCxbt25faegnEmJT3VMfkXrVXIOHFpj5uMzDpl6lU0a8oSjcA4HOL3tjiQk2l8AMLUl6nMS9SBofrzbH2cB492KRWeOd0Vd9cvjAog8S4t3is9iGqfe0UIoWL/2yUfL24e4dQpPnP8dDqmA8tkN6srJKDmAyy4sIsUIVIrzwsoGADFQo4HgB3n2gW9sy1JnKYGbP3I+nL+5o5gqRWPdH7oS5gtkzjBRhKhCevPrgwp/R6ulbjeSDFA3UHMKDxv6H0SNm6rRTQ7dUz8SsYGBoGs7wmdRAiqvCBdsrDtVtb5dC7GnRKGSK3Sm/xIVp/yACb0CzNuw7LqW69eoZ6fF9rUdChv/d5vtHZ1VRqOmgsDbl7PKkXN0TH71YmMvMgv19m8f2LM9FvpXuU8n+NWNKus+Imtu/FYxBKmsR/E9IcnE1Fi0V+K8FxMvM98kjBomPm1MtCcPrhWrthDQ+Iqr4T9800kFG4q6EQ0SID0eypbluD2hvXpzDwYWuVAURQp+pkrtdwoCR05FEUdyby/m5KOV4GyNdCzZRJm3NFF2Kl2WUaU6GHwrbvwZoX/aKrXFFNiqLCKNo/jsSZkLcmUny8v6CPOD6EOgCuHRJLmhCFZ/+D/rtumVT0xfEduZ6NLx0tUZt0GPhS9Fh2y0FHcbGNex7WA87amC+9rEl+8xvArvFYYIBq8eF5JPLoJ9tJMGers8cz/MFxb0wiqettLxx4zYHugUqEyR7oOKS1J/Wfa2rm7mShEKZFwRK3181eZek2lkdsOlUjgBmu8YJD47Wq1gUinVmGru7KMNWcSfuAHt1GGt1VZNp66NYtD0xsTm/H/ZW05rEpwe/BrHwuGjYe3OSJGphIJFM7Uph+uVDLOFwVNqYiFOe26Dgwj9wJUT2wgm5l3K3gpAXn5ACwlrFlp8Bvk+2Zzuje2jHmTWc6/98ArLICavLC/AoY94Ok7svaeflbvnlZi0Ot18y9YMlAV1Ui9mEQK1y8DVSAb9yQy69lriqctZPKmeVfncZPutRzgkQnm7dHmJ8q/70er/aZgwWIN13fxqPyhT2bLFrdCi4Tlt8Tw3tatkBOGycs5krfarLmj3NrMMogYNtkG7TLO1yyUoglY5oa0vmNxqzP9rf5dTn/TZ/2BkHwr1mzM4kUMu67aLEvIyTYKRshM74mOIJatCuDAT4znxx/eQE18sRR0phlzRmVKn2+laAlw6V74TqqByd4ndSzJ7FBNuRRf9jZ4yfjRkh1pwFXsGxh7sHq+BtPzdA2QKtoe66pKH12ZIZhftjVR6D+PWqbltWjr+tImbL000aBNBcjoV2OmcQ71MWBoWIO+WtDl/JBgriC5gOyL5GmUwdiFreDsx585UQjy0W0Qf7cx8Xb6wRRmWyFxFARojjETc+DNE4aLpjfLc3iejYvcWfcY6rP3l7TfE/XdlSgGUCHzVp75Ut4uBFGuo7A45/EgRW8CLsLJHeGdB3SgrNLavu6bJbLMU7438gETCF2YGtg3R4tBfWV4siKchZZUMpre8ORurcUoBhDRCRGPu4w3eCMzhUhqCvpjtYtH8Q5+as5Oo437Wq3tCSXUfX7OM6WkTi+rv2bhGxNlaNzdQKvli3lEGzDIQ0QNHuhslqFwFneefXNnsLDNgg6SDKOt2WJQJK4ptheJVm30lvqIeIDeVBBfn/9Ya3C6yyVfGbyERmDGhYw9SJTOM78yDAr4yrLAjFWSDZF2iYdoeXAQ2Ca7diSoxnqkPuKS573Hf1v7xopte//A3MbDfpAJ2nsxniBeKVH9vO15ZHupyseUDWbXvpiJMVv4v9kuNRBTGVgAMizqFHP+AbnefLejqbATcJpfaWrZYOF7Smw5f83C39aGTtKeIqX1asUlhsZCaZuwUwrbz6nvBMd6m+lfyZf4h/86F7OVjV8I3WLy/CPy1cEQuZPMgjRhHk4UgakAWv4PXJrtuwBDHpDcEp1Dqu1q9e+bUMwr5YUgIMnUMv89Z8cfLV83SCegIc8H4wF3BKR4Xxcsa8sJ0V+aILN+id/JV5aN7hpH4QYueGmp6+UCxTB3c9v6+Zorly5Vhcdz6ntn6pH/JSOYSHLX/Fk2p/kcA4ZQ2hUaf4SVrMoyPNHf/jtwKPiXsaTRzLSCwN5Sb9R7JbxfnddT9TsG6ScLQBqkVdru+bdgM9+grDskjEuQV3eOplbUaj1c5NMu7EkMvWcZEvhFh8FRufDfN2UD4yIWwHZzjzri2z8chKO+QnQWFX4gHGRwcfFQ3XE05wvKnb3p48FEMGrkqhIzTwJ5bs6Pd8ah1u0K3K45LGWN77Zn7GSHbRRjkCCsjpTFx3yRk+SwfrekomIirl1x2m6vfHNCP7byJh7y1ucXCYLFLKLQGs1u3zqM1CbiRqWwkqgTDf6BZ5w0eUcpFwId8u8NmqD0OB/mL7wCF7ucPb2sem5sGaPXxiLUnn/KUfH7jIrPPzohTZLdi0l1gMHO3h08wGy9E7UXx/kayWV7URFF1iCY29Rt6LfFeITq3jxgpTaeHpLo7SGvCF1QyteM+CzV4FBtVkPXOedJeP/SL1F6bD82w1Qks1iRDdktCcfQGgAx5FWgONJCX58wGFm6tk7DaGaXRzaEIy0LVRXETyoZkEn1M8meHMmks1In/PjtvXftlsaSoX3l+RcJbawLkPpRL19PWiUQz2jTbySHSGZ26Xay18ieyJl8TxLvbTA5eCd4PZBG/T81GqEFgkRogN5QSb1aAlDSh16PoWoh//E+aAgDReG0pdHknieUMSnItrSRU/VCMqDTNh+A1XxjVS8PnYfAB1PiiFJevtvnr5BS9jW3w8OI5ODSv8sYSeUPSFjbTxJ5VmDDllpTvYJweODRinZwyCZJoRlLfo7bRB+JW3//2sJT/XZ2nvUDQ3Ug/6a6FtXTeYW1yBVoIo3erX1Blxr2kJEUuMemYprfsXq/BH6RJumgHzuVFa8iU/oqhL/EGjHrCYXp+FHpO135Zm0ma6d6Ov3TmFOa5DLGPk+7fFrC7ug6RNFSkRxh3i6tZ0++7A28tuDJGlQ9m87iqFKv994OD/s9iHmHWYuHWdbaoxYo0va0DMi2G5sEhJ0kk/AiKz8jJI412MHbE/ORZbv40JT8l61j0GdI38my671KPVSjB+/WuNgNFH9ODoAqE1taRuRbH/+R6O3poBY/dwqk0KOEiamqW5AKT2j0lOu58yxd4Rg9as25Xv31HizSbUXDO5gFKyOhv6Y3kwb5YA+B8/lx7Jg/a1XGU5dzQuz8Dvc54ERNi70dH6ONXaeme4cIX2hudyYLeBLXzsAZZhubngekXO5UW3t1iTiDgqMs0w6toUqbq2nEG7Jo7gJPkwOXGsLyMaLChTeyCWvNZ6BkwvhBJ6EKMuKAljxOC+rqFKH9czcnLQoqW8Y7Evcpdy+PyN7JWoS7ALlNMN+cngOLF42sWF7i/84AwLhKpmzD2xkaXpLLY7lnCMPBMKZXFmwOW3Xx7uWKxvjFrUGK1ImXNDFLYnW5f6JlQ46ISSHUNC1YAVQcaXrEQLPGx6NGi7/h86Qtc0WR2yf8MumizgATA81LmYTjb1DQ49Yx8hLDEZ2bOUhFjkKHMezcDs/eSQUlYAk5brURYMIHkMr6GvzlGpPsON1+Kiz8qGymcLOed71mAEqxO8E15pT3G65ByTU1wKJ+rk9dAapxnoAoTn7L+0nh0J9CbGwb21NqpPnUcE+u8IIcyT1cCCvFma4PIvDldvGOdunwhaNS11u4uaQ3Ily0d/Rfvtf1jYdCzHiZgOTjDqQZDTyqlUwY6RgHr8V9VdnrFi6Ca5ZFy0kJZ4ZI6J9G8iOnq5hSWzUYtvU0uVwowtlTdCCPI09xZxqwFeo/8CtbB5SJ97zLDA+xoPthzdy6sPqNJRGDX5vNoNLkNLrggoQp1FwtWwE0Qi5yit+055n0f5/Wb4AW+Hahe2cn2RMWsZ/TqUv7v4eyYHCcBCZUkV4E2KGjpN0HgXoiT5SLMTqZX25XiQdNos8is2QKaN20xj4+eU5Hyl6JiSV4PS24DtILBk7kF4wG9ljqmK6zsQpzW4nTuHbm9r4fv2XyttwcixOCtG0c5zFH+yFCTWVuqlY7Y3+DQ/451hm/zHPb6tHXSdtsOQ2X4vS3S2QuX23E+HABktGhXVk4bEUP5hEWiJFCWzZKV3On7Conc21pFCUOuo7U87fkbb3jWFJu3+66mCnf+WqNsrJq+1cBm/Bk5GzxCvad4uku7MvQV0qevDDkE7edSw5s0wbUF6S3Z3sEDlszLw794cqJVsqC1dw1LqgKIR0GPxw3Kp0L0m1h7RCVadLZ2DNWKBU3/weD5VqFqvMnQUgQuuU2JCX17xnI6fjg2ruzwcndKw2zyOgtcZOFOjQ9gg030kqZKlxrhzMWYP3EMAXhohxrsO6Gyna/4Myrnb9OU9bq3rF74TfB6ZnRXMp+T/xhvW6T7Ojs43RZ+54PjVP/gz7xMhoSWJYST6l6Et+Jvd8FAKGN/EDWPBdMFEROR9xEY9a9+mtf9UZqi6MBnsrba+XQnrbvQ3gB6YNQtpcv/g/IkjoNR358UGHcaSvmTaJLEZK+QkdYYf9fZ1X2elwxIUmsIrmPp9quU/ebwIrkYfl4TtNAJom+Mv2EvYYckZEj35rfkynBVD6Y9VO0QwHEi9Iz/Q1+chDrhm9YJKcw0/GultvakNobItautrJw5X+aZ9c6DL9uZK8uO+0twOyjzGFvEXBEpJP67D0/+EuNsPFmRuvd83OtMBqKrcPemTUaweS/OVwtDHl1V6UUIiIzAfS2Zy2Ehju2RGNvevQyuZZA2XgYxF7SvpsVMtN+c3HBNd5nZ8wKh9rUvUA82pnKFpJhs2BVBa+RzJn/wk1pegiP77BVs9JMPcxk450VEsEO/w3qRddGsZBk0FGgAjUl6mo1PAYApdsz6rgnpPkWxYChxO84xk8YietjVWrZmCgcOFkrQle01RLXCLR/h6FeSg5fdavaWRcmgnfbSn2jvkL6r+WyEWzLwL13UigXmooY1VWf6KyW+5xBeevg791C54xPZADEkqTx9cOu/aQ10F8qCf8OmapXNH7+cqov1vjuhrDSo47vIY66nDAydGgDXd5KBL8b7I894DS4yV4LBUDUVpKHt/5L2EZFQQUx1vMB8Ksm+P8TgaH+ow4sUEZUcL9Y0UtnHZS7KEhu40hHR+1vE+mBIpvXquCI5t26Mf1QsDO6Bdf2LkzTucLRtSKUAgMd7kIPZUTb6ApW6PBFjPDKvNUVjNlo9FX+rGaTW3/uubvOwLmjKhrKQCa5U+ULXBtkciZ/+qQ1UyqCmSffPJJVo26+9GJgHZCpeq3dQiRB1KNLnmR0Dl1KjT7SHgXqG5byaHGiqn99qE2NEydsBtFMneMj5+HLfFJHKtWpD6byZ0orKYmlFVgNnJK0Bx+HJMwGa+simC+sFTY2xGn6p6FT9KtmgkOnR3NbrN3syPzaP1fog1J+F0B8/CmPSDyujms4/FsRWToSb3g1yYglrZna6J75Ae7utRlaOr8nHCp3C+hVOGdb1wJN+kyIHgmNiG6raCTDy8CDJL6JArbPKqrORP62GkBC6VHeWtNth75NYXQng9iLzvFFJgyTpH8l9S9//3GzPR7ZnRYrggeGqFrpx61yVU5+Dc1k+h5PgFwHdLgOKxYDJk4FDAqG4E7+P1Nb1GrLZ4/YA1aMWHWqyVkk9LWleFblNMCsHNaCF0Hp+QSaa/l+6xTbBfb4lM41j5O/l/ZJ6DJdm+tDzaBYQ4fKpg9t34FvhNkweLpoOFi4th469SbO4yjJVVL/Wb10YMyiJhHemIR6XVrgrZ1aY8VKZHqtlrrBl/rvg20UIzZqWQQPXwx186h2hiNtU22n8MzBTicvzxnB/8kB2Dr8ciCDodEYDps4R1YCLtKVefGYcyLuoAJeFGmm97cjNWZ1qq98/Fe33iQ8Yc8MpOIz0junWw1yLFimDL7DaulhupFL7VpAvsbf70Vxe5prt84gsGr4K1QGx17RjPbjefbgpzAe42rQAfL1CJtVngEl/d//nVeTVEninekdSwu+AfUAdUV8iWfvc3YHZraRNrBFZYYBDWfhePmmxbof2EeD7CUcAIVs6Ks/tuzr6xCQa1+Jno7by5aF+WRIIaHW9O2o+q9CEngfKqHNzMk9x5kCD85sFXLl7/Tk2U4Kk+vVkWdVCZnr2d3hqJwYO+EJ2Mumy8qxjAN4PSZocpM5z97+aw1wLZdfnv4u/hX3afi0qYv7YTcZ/F/XZjtv+MtyTYON5DFGgP6ItLsU6Ku9AMXphJ6SKNlB8lxfT+7b/qjlCqcFGPFaaGnmmau40yy4EjgZzzhjeXLOLxyPxnJthXAJtIj9n6e5hLNWnMLIjhrBJTdH90pdbdLWKo5cYqz7tOVA7mqe6qDDZunJiHDbMHPsMOrxk4qp7uf/ZWpALutCrO72LFPeogeYyBuKLdJvv8qA30ddw8tWo6ZbdPI+SCP+obmYTA2uPSNrGMkc3YUjUIj7Z2j1XMINw9XeJXkQXcMOKpkgdRYGZ+6m5g93fBbjWA0lH9cEJA8Xjlzpk8qjSEyKuUf2fLgg5cTGJgCzxfjSPdhODgIah6VOSaqF8fwXKKiXsd8tRrAPfT/jU3WIyglrHwyy8KLLeFMGeHc4Pabl7VKs8NM8oZq5qKtRKlFiXRELXqsNJ1cZPsYEMFF9JMhIEnZE8QStdP8Q85FmGf3oI++BaxbQJkzP3U6iZpHO1OzDxsL7UzIMrYcuNjQr43qY7R6rQ+cPeVtIi1ZQDQ83w/fy8HABCg1KrNGSBgsQt4Il2HosmETLZfxVixyNTglNtu+MJCIh1pXQLuxkpcXp/eng9BVDt2/Bsxue1oPCHdqxCBoV4qGdOao5QVGoHD03ILprNIotCjkNGOKnX/gB7s8xr2Pm6NLR+TITnJTPKLGxneG+AghhohNgfOUCLkUSBGlbRdZmscONy/byetb6Y7ybXHbGu2QEdzOiWkaXzjX0atdHfboB5cllc3cMvVDMJ0Z7k/9Bb849yQckn/3gP9AmIpRrYqM+EGMeYi4RETIVV4QRz7wGz+v82r9Z9+rltH1Dbx3DEMbdTGZkCNz+sBMv85XeFKSfe+yoBrZ+lrxplNWwDVRBuo5zrKxPfBGu7rFBkJoF71WtcHH2x+qPW4+rbMth/NNk1VZ3x5qMD+r9UwUo/QTrG39PrjzqoxfrphCsAFgFNFUgNO4ocvQC0Zv3TjyIij9ntx9PUSko2MRxYLmI+nomQiFo2M7USw+j+lkaaSCtMO/hZhyS5epqLk6LQt63hOxPwuXD8jE6/wxLA7+IwmyezP5T3hbLT2KUXK3nPF/1eL3I3IGsWmxGfBmgH5KkgSZXRzhl/M1fEh+vy4pBhrGpp9Xr3L+cYeoGUcH9VJgZ16alm7m5i/YCuy68ysR9CYcNshSp72Hg5HYY4bLUHLU8SSoWCO3xhv7h15vjHA7RZe1A4QCCaoUfMQqh3GrodjK95+jw7XWQ3i8B927l4pIbS0RzMuC29f+rxWjOTy6o71TacopDqAEhNXpH4bs/dpfVx2PYBB1W0dn/nU/gZx1h3276SQskuT4vv43WG5uEwXTru+9C1rUq6Ocv9bed4MEqIVKFr2KJyR0VZW02AUIbcgcdoeibuoaVry2/bHkFMp8XkwXVNUjOIHnvUTZvDmJUm/4TQ370w9OdIymnmZfaswf8zSxJQYvm9MkgtmejRQ1TFPQt/3TM/2gUjkPma3c19omYIcvInJg3L4jJKnImktCzqS6AthcA0G7qyo6TyIFKsdG4hK+FqLh4H4gsCqublNXzihu6Mo0WG+dBbhrxvC/SdN3XaKZo40S353ODuKlfMszYP8+Y7u4MHee4uYrTYJIWSHc9zs1SbCzMM05fIEk8ToLOFQXi7fg2+MYQ5txvMVFXds9cqBQ9P2bwQefb4eYeg3kEJPdLszfcsNlHF49GTb/JOa0VFv/dRlOOnB8ngvzBpCKuWKMt5xVAuuc68XGlQSicou/UlOjHgxPx2m7ri8yxWYVN1ab1W1E9SJP+fEw8vKHRIrKb2qX2ATS0WtVM7yEnUkHscnB6hg02vLrbdcycuWMItpOBYcMCdo+EiLDZJ/i6fSlUcoMK2fFtlDjPwsqQHCSAcfqZPASn4hjmn7L320ks+IM8PhtFi/jf06XdT0u4xa7Xi/4zXJNwOUxb2RFmxPO4BEdWHX9kg1beJuQFa+sqCeX6q1XAxwNt9eurCsKoark1Yc+ct2qe9TXdfIkwQUTuS4W92LPKHxVBo/iUfyQs+NaBzJe9ECPz3J/nZyUzTWPKGwF2D0Wxi6YJqkGxgz/Fa2kbu5SfqxUMAUGGevw+W73NrcPenhk8qIaR68tVCKIr8+q05Dosbl0Jmqx412UOuKHMx8qmbZU+ANwB4S4zCtyGQ0vtn/2pfNLSAjlB34J6QyoYM80dCevRe2Vtl2KqLuunEZITAEkC8xp2bOh+FuZSh06bhi+yklerORtoz+bSMmE+bUWiNmWxUk0xHUGGcUon+WUmH1IJsmmI6fNMPWJIIL9JODJdBEBYfAFHrS/IALlzYvEd4EFdHrU8X9v9RMraNcSaVjUvCNteKDnJ9xs/OAwNJErPIIcRt6YzXeQHjSOyZoiLllSHDxPCowivvR7NbDKPNbye6dpTRdcmSAuc8RSYVHUq5xSOB1ftNp988+z7VUDhheW8aYkMzm0QKof7GQhExgYUBg0PIOKZSM59dZsUvktF+IDw+dNmVr/IOA2rjOIh+dCy6lpic287ZCOGW0SMsoXTctCYuovz1rFDejfosMs7HmvYZuddD0egqsmOyeJZuZuDdwKUloAwzLcFFDHAZMQP0ATkD7vAl8xDsnyDCy1TtYVdgtSye3sIVNHOwG6noeJrbkj67/Fo7fyopPJwPEwdXyZQLatHXRAl2R2khEmogLlvgbjvSFqTh3nJOTI3Okgk0B47HkLLTQQJiSaml+SEWbxrVo+oS9DhdqDReLr1i8uU53hrv2UpJwcJNXGRAVfrAHU3CzeBWPoxCwsobcu4toxreo+3G/bE8BGwK8QGUXLNC3Ywnw/7WA/inHIxCz1HxqeDdJXgRt9JV7CHC4fkgzEsTIayvSQ7+y40FOpjugzt/3/FVQqj3gdQva4/SPNDYbsP8w/xvrkSjZGRSA0fjxUYLFUqFeezQT0RdKMKFTJ5C8BsXutFj17Xrj2f/Z01slL5Ueg5HGiZrIGuIN6GTToXvuitkUwEw9T24fQiU2l91vbcjWTG0nWBFf8u5dCHmI7UK+qYt6xkqT50njNAv31vTzutDpwnpNwg+vWmU9Pf4i1mEcSsKu1Sa0hG1w17C7lm6YgfOswhuCoBVOzOFpZXRCitURdanP3F+wJRZscghbzpWJ12CctXo899VeaGTAUjaoeJfwkD5eX0STH5i7TSHYAHYuh0/d/2xOUWge9hZDupMnIqZAEkjibKVmUVaKJUUYZUmY0iRoRATMywCHnMmZSbyxx2jFRUp8e01jZmp6oJfH8gc0zrUQbkAiwvFOPtLEzPr19+1omAGc4DOVeonsdZ3r/TY/PCD1RDx9vMvxjkF1NLRrTqcOHYrLjzK4gZI9XLe6Nd62SETHRh+5FFJCHwVwXB73X84R976uEjwreyG5I4c7Hzxtn3SQYN7LgLJXRVSkAKsvk72+l/mfwyI27KJBQwy+9bqaViwD9OCwRnjz2qv/CxdvQeG/itYo3SxlKXojoloW9yQYON3F3QJ80gphepQ8Fj0bJUJPqK4i0f3sdDa9Ia7iW+ZCSRK3h+b0+SYDTzwMMuqri4G/FTCDF8dlIDSKEp4EkiAbFoYBxl1GZHQ+jHIkYWIolnYq4VwEuovH9gs48B1qZWmZt07DbWA6gyt+JoYLRS0IDeDk67ylYpb/gHM2NFFpXYm1duN4TaSX1Ec+46tcQnP22giCn7X1tM9sKUVUm6MAeJFouitDiHp3okso88L99jK4I7rN2vSL/ot7hysIYx7QbOcCByq8wD0o8/0oZlt6oUzccfxEb59IJo2ltUcprnwH0saGcNRhBEcq+1iaLidNmPG6veiRtsQhEBYLsugjjgFkKBDSvBS8bPNR7F50Crfifim4AdmdiwoLEftPZT7GcRui5ILluOrv/m8YciGO5zW1diD8NfF4PodCFMX+tyqbQtrup/ch47nfHwow/Bd376dwQvVlpD+TBQyjJAlWzLblSwdLsRlB7jFGDW5edXnD1YHhQhoYD55Yb0jA/Pyq5HcsEHbrPC82bIVaOoSjna7P75tQPShCUIb8VI49tzNvSHN110aUNP3hhnbEXQoJubx+HCJLwj5PJE6zvsw2DEwuyS7JnEYu22o2/8sJT8ecjpfsWviDrtUJqT8DDhfhxgJY9xBIde8bHUx+Okahv8lH6Fm381pQHr6DbkE2bCznhpygrd7a8jI5WTqRjPGW/nih5F2R2ewmTf1rBXF0g56FdYhXrPNsiyTDDRQNEEkA5ue23517E0Tf00CeIK9L0JZBNilHz/PK61bhyEF/TLcdlvhSsss0Eb4lCMs0HJtXLIm/0piIb6YbmNN7xXXNqzK1fMBqP6jh8ELksL8OuLJYvSRwwhu4ghZuifkgy5NNWCtts7wi1GC1jg2NHwjy4APEIvzyR3EchVd6UpnCh1F3E7Tx5ujcyDHIh/fk2KHaiCDiExmI22m8UdW97aqHx3afkLBxLdiDsjvJ8aWnjDjjpzwc0H539kEFCkDtrvueI4RwyDL8k2mJN+5Sfa0xiV7N6hCEBqOMEGrcJnIfkBpAXRcQx9L3lXkE7sffjuVy9It9PR35SuSiBIbJ5XFgOP6XBsZ7L3vf9Btx8GyaZ17d6G43XaV/Xh5W4FkkyDyT2fkaZF0Nx5uKBKXJoKE2zR7EPNFFZLIiNe5eQQS9gSAKZM6HI/EA5XLLlhd4i0uIb7dHk1Y+EOgOddbTtqiDvDOaCIl6VFHMOeWkVkLC0wPNGk7iA5Crice2GYrhWM110ba98r3WfDcIk18dsVionG+D1OcPSZWPpqbW8Sh6YLYIKHETlLDKd5ce43hgetwS2fZa0NepqRkiDyC+5viky2t7LlpRGwJqxlPEc9VPXJzQr+b0J9RaQiATQVZdn106FlTNuBOToHvwPoP9UnSy3QwLDPtBMmbjWo3sl53mA+onPVOnPb5XQMRIPDrYrcH7azGpytpOIt+VDmNCZijv6SKKgzecxgegggwSksSOdmMTl/jSlhWg1KCL7kinsTklNcgKNPnwEPZW/GumvtWQpbdwjFqNzHsA4swtn2acE4oj8MvS1V8+cAxF3lpHCWpE8o3tvfPC6Ksq1CEAr7TCvFdMNqdEspNlK7LWXqsN4tTKSk9xpPMOB7ps9gLp+KOScBbLuLZmD4UdHk+BDFERjMwfqwJTMz30AeQBC4RGYqe1+OrJHY7q5LlBLRX3OC4HqKMVDzm7msezVJbtPmC68R1EUMZ4h9mith717YLiWl4fmPij3ebau9CvtZ9WR01gVq4BIXgRE6Bbv6+xaxR1EsEwB1y6xBRVWlKuTGnxRVOnKM80o2TzD6NQHWB5ICVVHFNeQzZLiTR/50Tfq5+WBw72d0Pv/tvuCVhMf0Tzcznqyu6LfXpUPBB1B+G0vsFEstt0O5XneAKlqjI2dOEfs9ZCtzMSQ11N6MuWm9yqWsiHEdGoAr3o021eGGlhQBT4ZolWBcTBUN47PA5JlSDzQNvUyZO1EJ6RD0rK0t60YEGK/lIn1aoAHmYOU2K9P5p41lo/ep9Y/1oP3z+SuWnd/4aE5OP6qIL8nCkd387xAuE4GirG3eA4eHFv9svvJEem9oaXplNvdnAaRzwTw36WU8ZjuyjdCPTJxC1LkhjWDV5F8It2x7buNK8tmx+sjryNzuTxUe4W7U3w6C5ruWm9Lq74b8T1qwnmKS62V3Obk8zVUrqoPYXSWwGE9M49v7cS/tYpPQV9oHfT8vJ1LEW9eAe0bhM+GvshUQwek1lgY8k4vXfI/XOZGBgco9lOmVqdzQ6Z9MmnACCS0eKNezExFuLlJRTUJcIfZjLC/N2+LOMPR6XIpu6Ly2Rs/C6++250GU78xNdxFVf3fKZkXc9+it7IkQbMtsNbTe1QbGWkwYWOGXeizhViI7c/yWKYmMAnBtsbawxcztAmLoAsgn77HfrTi6sBiISlQisRmCtJwjS9mljMwnu8LugKTRCI8eEmCu7X5GibfxCCirTawqBxrjP6pbleKpMJlnA4VT3PnYkrjGjGFkCiyVtVOUvekGIiB8dH5aUWIq1oZyCh5Ef4LTToJ24pTDnDnEx3WO6077ygHeCIm2lJp137zuATk44/reMKF+9Ajegw0jRgBH2qx//SZmKpDcEnobeF6Spk2sN7bUr/OqdoVEbhAwNS1ea88UXT/X9FS340wblL5wGoORtJFaTBl75OLbpaz/y2GEpidV6MeW7H0rjfbSYeY205ohC7NKvpSDAOihZU7LZWxu+rm3wxlh6Nd90aQvYsvUboXx83rM28BAC4LEGrKdEFU1+xEGoKi5QsFxiOxpGXSMyLClZHkZgippNbPD+FX9RPYoiZ2+ATp0CwVKv80W8hpbBswBzMiyltTesDYa/0owes3G05eP0BGdDzyIxQSepXR7rLVhytnDUTew+TCe2QUtWowBs3486tzdHORGF6guQiT/jLru7WL16jMQnAyq3WjOBYccBMaTFEqwGn/ddOQGO+eaMw7sV6FdP7ojXHKl8KZgdSRu4rcHTqy6ePdeoCV9DvxPfd3afBBG2s3nI5sW+U0XEbS7VqRl9UDYYGpzzQg+pIZTSmEi91TmW1RLS4o19zmakQ+S3foTciKNH2hZqWvFjISGxqTWzZh3YD4sKtnn3lgA3rKUrFu0339LiCwy8TKouSVie018tZbwXBeqyb4di+e4y/uIgH7e7xDuMu/FJEzylrx0274In/xgZ1ZhBVZCRR6ElB+QDjDGetTXe55/g3zqLyGdq5h5e9dRBFrYvIO8SE1hUbQCEdZdRwPm6c/FYMzEEeFRe/ixHfzyOwUUtRXaSUQkKsEcjPVRW7gDIG4C+2GuAbdAj5oPV7hoAWXRfMM2B1gqGaOP/KX2k6ZuiS10iidD/lB5dxYPgQySdsahecYHPxka6mCBGfB6L5Nl5snfuF58Q+v7XcO1A/ML98IuR51JCcJeQy5j5sBovLRck3V0CjCLzZ9OtYRY+PpiteoPYq7L5Hjn41QbO2M3RjhPWCzd7GhCrPai/7XbRzMthhVh8JPjzSQaiWIjgzctNFy/anhSEUA/whH6NSQszl2lhFaAvNPyTZbxQLAcBstZpFdZvlhIxS0k6cheQimil1DZ/bHGnGjPjPQB9mb9faasZd6iAC1G/w5GloJWjp/RjxLNrDx8uINfSJekNxkXf0OP4vkj0EYpczEdCcv5NYDGtm0cnqFm6Sg7PN12z5QbNrKGkq7BNMHmWQA20DLAQDshx3ECIIzlFOLgVL6702qaqdGCX24t9OKGm2M6fMzTfaS6qgtUeEa1+sKF14MThvUlE/ZqjPklTOnObBT1kN8vQKmJ8poagVA1lL7af65TWJPLsz/upwsS+WbZPvdkNNHSf0ehInC/w3yOvMrejQzpmjmILj7wLJiuaKP/5ITexiYMTVVQVayoaLp2traw34utwUX/yDKIm2t6dEZO1DPCkmsEw8du2hqaMxCUd3Mj4BNxqOFtHXb7+CKi75QWWuN33DXXw+TEtt5LC/aEgQfxYHJ/3DIW8XodTj0TeqPKz5Azy29DlQlvg1A6i0+mf3+KpBEvontmTBxu+xC5c142zMUWqQMsoFN6KCQqB97iY40ZeXh+gdFv7bT4c0OS5HZ03+zrzJT/DsGococPnoXSVkPo++5kJ2+E9YNpEvi0Rk8hbiWM8PxeFKFc89Kl1m7ByREESMHKcWw8nFgP20i5VpA/hq1L3BbmwlDD/TULXTvfceJk+yq1pZgOGG/hduMtdcghIOvYfe4vcVvi9ysaoKeKS79L/oSnkytX7JWB/uOsWvZks+szjwuHNZdgyxIOXivvPklUB2T8E32AnfFfRUL+SM8lRkxBkIbttQTwFOlNloYUNqAYlKkWjudk74i8EPZLfZUMhsXnTNHouZtwayyX6jYt/jXjN5e7T7vdBfaHqCHdZOw21XpHEdra2nF8x+RzlZd50KSPzUIFyG31OqNF1KFp1eM/WkqvE8AFi3VE002pzK8l+iVawNlc0F1ZvRWs8h3+1lI4r+thuWPtTVMnaReZmTpzjMSxh2T0Jjcl99yYlwr+bU4d1Ts7mF81XwXxT3lk3VK7U/9r1dP6DnkT67kmquQiaOlU6tm0RGr+v5bA4eFTSFx/YzRHIyMVXKChqgzRhkl9cPBjOm6xZa5aOLxw/sitXm3xFXm66Ym16YiUid1Mu8ANouMxXmJiJiBcOCJix+qwvotzzV9ieYey8tSTnjCTMCJuN3RDtFj3kAFtJJ005zFcKMQ3tKzRuOMV0zgkQdUjr3Kj8Ufw4Bv04mtqckSrQFO6gdBdFiiWgMYNNUlIGaE/DrIQYVIz5L2HTKKgV87fQKYbZNRYqJ/dRDW19J9PxfXIHLw3TKyI1MXTq8haHUl6a6oY64fcIR9ZsIeO62c0Xv2+md0vZMbgyJ0H3Ne9h2uesxSbcA4ZfXIPck2cld9IfsT2is2oAcFh4ugDWLNt32waCUNz8Se+77cFdtlOJWBuw3xRCJlj2Der12/h2zLuk4qXf81tg7l6AXLEuikejtnGt69Yltp+Nd+LoEWlnPKM7WHwA/KqRix43y0OcXezoafo+sZMmo9YgEkWr5RmuQUwtwVbo9Z1HB9dTrILILbdtoxAD417i4hGE8gxLUV1lcQQP+K3Syl4JZ/SWGHVbx5XrCrR+tXlCk7L1votpZLeuFGyuv7WhRJMfJf1unzYXkXmDK3LSZi0NSt4JXhh7FPUxBQe794Vki/lEiMUB7UoeByrgV0Ibt2a35U2145DScR80pC5TSmtc0abxQgQ+16gfYpg1fogq72DFZw4l+CvJPsTE3AmTK4xAvTImTVbjz5KjH62wzXPpgPyJMOOhyO2iXW/ovN85kJJ1iR1Y4eZ+owBXyhqqLHDw0DuIylEW1CVffBUqlL55OW54NXYsPqL+5UpdI+mS6FOQ34OKU3Yi7bAUmwkVN5r4rSxp68F0bsB8l0ieLZIHkY5lwkFd7c+ugh65ME0Xd7ljEnYLnnbnKwSW5re9bGzVY2btQ7/MvdvpBDAWcM5QzM16v2fBwI6jbtmLeBLC89xqxe5Sk+YMFtE/s+TwdQo2ZeqIivin8+z4xm/U1I7HBncYxeyiKS82ThCkNOAlCxzEiWG1kznFnh46xd5Ro4dBL/p3bDXuafhOIJ9PKQ8uZkNSvJK/EXlDWBhZEGFAdfsj9KClQrFF0LTis3MDUbCnHjcuqar5w8ZHcc7NTBF2XrV16qfRz293piX1kPktzsIxrBOnJSL6q/LgrzAGK7jitlAZiaZcelPcHo/pJzdZu78PhbDG76hpcf45UqRRjEQz+Nfq/11TVlRAe5s/zDZTLtW6zE5BKd75TyqlhyatWpyByWAg/Wu7LNrmrkXCEriso66rZvjP5avbzuYbXsXE8a3h6qSw5jIYeTLnEib/9cDxM5g=
`pragma protect end_data_block
`pragma protect digest_block
a00092ba769f166d8373e6d61eee5d1a332dcddb40376b56272fa7183a4b08fd
`pragma protect end_digest_block
`pragma protect end_protected
