`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
wxWi56pJKoB4l2kw5PdsMBdPNgGLgx6nSAgNDASreY4cC3XiMh98hWzecNpnW1nSB+OdMfSZqbOQrgFXDPODrfPHLCfHz9Rzh7Od4Ap4i+eQFhGYTXxQeTVwFNFPRruemMXBdvHj1YJhCcLS0r75Rb0lhOQw+7H8lRG4xVdVCnQhIu2Yrf93VWJ6DcYWBCSpTy63xoWZ/7bc7CuXbSiWGHGN8eQIQzwKD/GRLkGMgWnOqjpMMtSs8T/CgFExOnDm9dKkORxldAeLpIq6lsGJBQoYiOeOPrtFgz4INVxEpWQF2MN8nXj6nY8srWpgt+Ymndrhwnq7RqsiAsREGFFF4L91J8hv5pC1uOCwrTdpIAw8z5bnRnV3ZFT0raUulg1rLtluvUnhzRVz1wHM1+BZ2/c9J5ZEXa4dla7vxklamqN+fpB+nq7PoAX54GYFgClJqc5zBiCWqp77pHJeTuqmkT9pMFUG/cvENQv4R/K9lOkU+LRU8Qcqsvl+Oes0wXUsEBAUg/e9VUFefBEXXoDC6QB2DyY30WXJWeUZNs4E83FuuxrsJvJg1I9zpX6u1HUO2VrYvPhfoa7Dauc5KEuRM4+76CFaoSsWI3NMFjOhMJ0t8Gh6RWUJcvsLmtJEZXw93DPHUShPSTEeGPseEla16iBlK0IJnhCmv7paZMOe9IZkQCSoPCcTYvwWCpQ2FrFFEdT3mYheuEKbaLjUzJyDeV2fSj2NUipiLRLZgUBqAN9YvZ4dfC6yFtPvrtkZJL739hMkT3SHF5PRD8oisjz0gQZG8PAhOciTSduEW5kUEEco7IuzMim+WxJb3D9WlRDtPMulbP9cmG5kSU4zyHnPT5sTQvrPggpcVuiyGgGLnjYG91kPlWZxQ4NkZ0rt2Vd2jei3pIDTuHwDmHeTlYfE2Wb2dfEZFZhExeuJJwMFDh2IM1C4hFSvHkPE/I+XK7wbkgUAVw0LvyT3FiPsp6OWUXnDK1HDHVRE8/xsbHmdMCHfROolrbZfy+TiISG8gre4fhhxN6lSIMgWYC+K4wuHX+9emZ57LTlskxeLANuFW4mdB6dtI8Nzwcco3I5diVxLwTUkt3mF8dgyZDPc73Ba877czZyMetxMfk0cdYWV3opmYov+z5iCmB9834hTUhj47qiCrBkdDMod6kp7hts80l546ncymApt69Lw/6buIj/LKbE/y8yr6WNYcQ7+uTbYK+tgOjlOYCFRRmdRZzR5ZW3D9Ys5Dl5ZtXNLdaeJ9g5TRHgFAarabVz/LrrpukPwVWLyKQfMnAzI6Tv614gX/XgFI2ruYKoeZ7wSKBxF/KciJWG5mZEKrP7l+E6za5bq0J0992n9foh5wqho6QU0RS3C26pzO+VW+WSXLS8Q2TssI6bnZGm8IsyKIVBl6Tvqjj4oxsjs2RIalHyvEopcF5+3zsdr9rNI0ESxm0Sxx/y4g9q6dPCk2yHP23RvE/1BPpfQN7FxQa0py0ix7s4psMUbxmoDKMtzAzjVb7bOUFZK9g577HTZ8lnNeHVwm9U980JjqXjkcgFIKn8mOewLhg9DxGMEPGagumNwbyN7PTCKEHdGIBZpXWXGgHVcp5jZwwfk3wqiJd8/E8P4qp3u1BmkC3EtamDmyBBamxQIhHT/YNggLsoInV01CMnoUm7U+aD2/Wb7Enf0qc9GGGHnTPG3wIe1Pketo8sdo/+fQXzFaRQRvrV4cggOMX9O6zi0Kx4bp4PQCjYAT2hKaAUbXbdyqIJJgDuXR78AFKupieIaL9eX2YchPbMx87jkpCmAJgRuLxkEBj2KCfe0nI9IZu5WupwdLWCP81fjWcjjE4BTrkL9Ix4Rw4HaGeWroMQykWS6Zl/ipYTTkWgTYIUtuKbtpJGPJr47O+C8byquptqTvflAgJGapGaiQ/LZrcEDJymPFWSp7ZPnHfMGjaIZeyEjkZD6vV2yAuvMxQHey9BEd+EnnuK5NzIcTUUahhyjRB3hB5lsjQu1zmavKTiWk8yGDWS2gIctMMhweGHqvjJvOnXYlOVIufyd5A8wN1MSosuccjYGWIXcF6M5RVhZI0Rb8YUWELX+Tq8P6r6F6mCsFbHprx3/Vh4J9Su3L8oJ8wedwAWHngvYeMYo0hQTcl341iC8EtAUiWMnPpanEGtDTCSwxZphvT0dTVxAYo1OYj5nDXn4EaNd1873KJC05BI3GN6deUHyzlAk5x2eNNXHn+ZQ6BGmjYPXb0ueHDqiP2t/gbEMBVwn5ax/s6DbIxDRizVMXGD1pA1+IfcWVgTyMAeqzbddJqNUbQDKWl+tlt7IOtywxPOM6e+Tf6beDp2m+3VExZHBddcSqLUCuVyqCrHyY27u8943voTESzFQTyWJXwW1SkL7UFSAzYy9HQb7pc0oNbjHCgusKLek6La52aV7hih2IBjyQ90+EGYd7HO9Ff35HefbAKehfSP3l7Kbd8g31wsbXbSy/jWNxmIkIBp1/ZBnGmzAASEhiI5pOvz7UGXM2mWYuHr142ZRGPq5WkHmPlzrtoXvCrFMiIpm60jGV10N6OssTgD+AYuE8nyDMqOD38mWb05eDjZknUwPMYYjf1cfGx7CalgKuM9uLF9Gy8DOFAf4YdNgs3dt5ADCNl/C0DP4xsXVwu77cPGSGHVjyiyRA+PcjEcinOz7/kzzxqnrFR/ruruQf3Ju1MWt6B5DMSN/4tkdNS7Yyg2P16XU6hvQvwEVR9DIa22rLs5HnwQEuOkRwQD7oUjfIeqE9/AgFuTwu14ffwxFPLSOM56ikuHrGEpA+85QNaamnlaQ3M1/vyvZhe4xxV156vZ5ARenzBbm3NybQQ7zB2ElaXYyJfI/Y3zWg9dxlOuOmCxE6s+0xQ6vwPdVjSZEIytNQZZShOyC7Z8Eja4OSWvXlPwBUucQNbzDzoGPxWqBGqVeltei8H6Tcr9Rl2+ii4J6Q0yt2RLK5YDeQM6Vm5MzolsaaO+8cc7UYbq6V9XzysIjcM4RnMzomAPe80kwDDkdAog92FrVJINqTzu2s5Nf8yVNfMXT/chVzzEV2GfN08EsOgeHslc9Z9GKbIIibuvelpOP7fDvJsNgMTxVVOTP9eKsMmzIbiYUMlr+//mC4H1IgP8qvDi/rD2ieJlWvv001ji67sNd/aeOi08J2hgJn95Vg0ZR94SmGkRy9ej3r6TnqNMXNnBWJFttAEcOzMMTES/0s1l0BJvtA4t6LVRD6QUVnkDYkldFdOfglOW0S9i0Wco5pueFuNhDOfnt3x8EZt3/WiCzWNZxQbOAsJiGnMfD8YFXur7pIUmRNGq3CmpNB1O8xQe1WjdCvmGgd1gOFIq8nb/A+smSE5UgenAc5VOHusJCUJd4swEOjHw1lqHLU4vOD2xbrzjNdAWjDJ34J7KcLjHmSGRZOU168xQMEVYaiLeYD6aF7SQQD6GhNn/ae92jYPBZwSHuWfAUc/5gcD3CfayYolqMAilePCnypEK0mxUJvkxPLC+QrSkagSYcRi2Ox93q3dAW6yCJe5SO5cjcjpUTnLibVkMkzNNWp0Bv8nfO/hWdEsu7T+D0TrSMBXGzxV9BqvDRQljpZC2QKj9u2eH5WDpJn7IzMU+dzs/wYlvgm9vBIMNnCKfY+dzMkR0/eZGE9ZWHaM7RgfAfL0a5qJbHDgJBokCmSDfnsRVqFCLDCZd0b3XNVURj+68k08IDw9lbm9rlm0W/G3B1/Op+SnayTQI1lNka3Yz+9ntkBixpNHtoA5oqGmfAGA2x9nbSEfbpPbNe3HzA5PABrEZTcoBaYjAcp2RYJ345+QQIkIgJ2n517Qy2doZNZwOGEP+c+NL2TGJQWAzQVFVRStkPAMthScx27BVTWgNOm/OK0VrBPI8wR6fGkkhzREkkgYV08Nust4T8xSYcFFO9J3vJHaJ7+MET2yLSKndqegIEsGyLrW3fBPASjnoIdF4kXOZKB4cWDxFTObgLk70D9tBfpd2MxRLn0/y3LLGDnrtyfPfq3k1Eyxby1sREma7bPBAplWnu7sooVeR7c9P2UwhbEiGhO7DjK3a/PdFZwc50yjG22jPf1Pfa/tUKeZjY5ZEY9I2KI+Oy3tK+3o5+y46CAu281QqmRxAqyJeiGPPj+CNcY8W+jZ/f+j2z3vOOXjLXP5CdObd4fcoZnrWVf8fqUQ3AvCEa/fhw8ArNv+T7eRJr3vmvWsFCr5Mdj7hkMALsnmG9MjtUDOkJSlHz3Yxk0HT4A3mMl2JTllkiJS6KkIaX3xhq0+4+HjGbLCY2lTBnDD6C9udYy9ImQdR4d3pPZ2zTDBIQaID/XlfOe6dCpCV0cjcHKBIeZd1Jg/QDrFtpscM5RDG4uqsOvIblPD6lGklfM4TLoNcCoZGcffH+IEM/KHIlh/4x+vaAbgxyvjtPDUy4zox4iHgA/SFJomSZHG5kBaJyvboL5pB2haKvdOW2JlF8HDrwQO4i7Nb36xA/j6GH1pLROeIMXlj7AB6kIUxd3+MIrrC6i7aUtkL3hKAO/PfpJ6PeyzHn6oKrihwoTT+equCDaNoAVMcry6lOmyR2gK4zFQCYN2o7G4Wrz84HH/UrzCXUR1A8KYSoJAkMIe71hlEZvglVowr4BDPkdqNXMWvf+VVBzZTtTGZJjbEQIjIeVIEibgCRWNAtJUtdTLOD7XYuWtsEMz1Cj//AGED9GmCqN0Vm/+2poapYWBoL8BSpMG0reAiaybJLwJedrfzMCT1JjWWcscQunn7RPpIUoXlPlPk6ld8UIZuCmIOC0ne/b4xgbBB2Zu72k/0EqgGYVrGQa0msXGYbBycFk9tXs5kFhF+I8hvz0NcKM1XHb2EO6VTMgT3GLeJ6Jbw+NqJHkjmMSSgH0uCwF9TunK3xkA3IFOmLn3oY4MXVSrUl+1zsmjenFgxq+dySoND1NICTsMEJFa/a5dmkYZRV0R4TEzcrL30n9e+ANbjM4MSPQMoKbKAMpwIJtSUHJ7nIzou1y/rYkcFTxuw/h4XA6eaqJPcL2Kth78Loaa5EFMhUkW+pJgskjbay6UA77t0Nvj16UHXUYt7N/QSuuVwv9Th0RezPTRIhfVpWFw5OrSii9dyUdi1ZirCAkXuq2JYMgPYpgi/r1xuja8s5nK1OURdMo46H631Zega1rPaN4orxe2ZwGalRYbr+NlLL0m5Yl18soRswc8bhZaTzT1HWroedplFSozzKccbyeonW9kwoiLQCraWMEyKVPQgBwqBosYGUgWnFPbsECElpxfkG6NVf5WLz3t+SG2CTfiHt8IfUfOcgkBuGcHw5PVSSj0q1c/G8LV/JjeXn3B1v1iTMfRruOsHRUB2n6yftPeJTyTwpF5zdNfHT28IANyF9DXurzV2qZHhfjpfaTL1D2eTKC6Fow4rA36EQtssttOwqksgCkKa7TNI/D60JBmR6DqI9HKhmiaEtjN8SduUwnSRfjMd4dpFE0YfXNZUw3zwmRJvOrP4pr8nq25R3KSfQiBMFE91nuiwfGSU0oX8LkzJHGpCoxxllQRwMtBFhHUflshc7M+DGGFihntbJXLPf1mEnPvc/K8k11wJQuz5q9UE5DW4U/AIzPbuZM6NHjw3E/5sJuesB9qqlUshB2+Edx+7D6bRJapdPuxls18T+v7MGumIBfhQ7Z1jFiagSLItm2wYqqFZnEtF9+Hw1vh1OE0Zgw4f/SP5rdufa2ATRDMdTdUyWH8gsrqXHdO2b88UhKqrAkNWc2EOTsfAnIcr2QKKXTr1jFg/VuI6EsezPKl7Cn6U3RkRrSDbILhioICEfDxtkmBzjjSec8whYKscV1gsxc5OTuktK8fIE5GDMK1Bwx0+QMiryYjQcNY70B8R7bZskRP/NLRBf+OqgG0cSjAAtTRHK2nyVx7DQ8/prWtshbnhiPPW87bxANIRoB/hsUOfYeE4WxP8gvQ9z9pC7PMnYxU299+gzpYOXsUtv3wiSXBDLCMbe1VQWbbt62LmB+xCWG+K8zRGiLaWfJWvQ3KLV2QDaef8A+ZWp+XwGneaq21vhL40/LBoT8fiuSevdpl0SQh4mYNvkNPxD51QmD7W1QD2gOskzqifsimcniC2ViHQ60eZmyqXfu17gbrUg+CZOIh55SvI4K8Fg5O4+/P5hB0SKoh991QNSn//HAp3Nulums+GdnPtPVUv9jMnHZUfGZ1hGz4u6g59yvh8ZHlAaCgf5eEIb6steQYDXR8MLVlFu6YnQx/DP2OdqFAQs/voGxc7Me0CRvN6tAcji3sVSlX89UPH4FZsOCslnYRv/qjCLwi8Zz/aLmN3rRf4HV0UtdfdRJYPuVMYpNmvRGOH29f1a1sieuEDn+mdaVBomjgDrt+i7wW6mz6OxWU4anhRIww9kAESsnrlgdC0lR4bvCrj4mNz/uvi7JtDgmXNV2jAxMQVfqyh7G+/hPRgI04cxLyIU89NHsP2hYbo6lirqTsVtFYoZ5UuVPIWH5Jl7yQnVMGyJCjuBmDc96ziX5aWro8f/MtGtFc4UrRbEiDhEiHmO5upzpDX/ae1KX4DfVMmqBRlZG1qVeqxiF5uQsfIL4gYUDZ3ldf69kXDfgtedY0YksyWh6t61ZDN1fKQvV4B+bgXbJBuJFFpgSYlR3csFnEEu0d0uSg73V+mE0Sw6unc1LptHTtb0av+ed3JctxVGi7xUJJUhJqMPWEhaFXM3Foyoh43nuRZTuPjef1LvMJTJO6GcDYNa0e5vWtLP+iJGtPQR1Yfp1+sO/nS6qRIV4kkfutzG4VCgCUPzn+1cEgQiCr4csQKR/Gq4jf9o7utW6pZ3WWKBzCrr/Zpo3bm9Rop5NxO0A6ctvR/ZN5nwKPs/OLCtEOAWE6J5+n88ND/P8ybLYoJnO5Zqe7+x+muQHQXUag4WMI4ANNxipj6ry2WFekx8+dQybkFGMQuC+ocuoQHO3dyTfBpHhLWWnWm1hVFCXNuw7kQk5Lbp5SZrV97Khc+F4gBrb5BbMZmoYxicjFf3UNgw0FaSRtPiysiDmtnV67LE3pWH/GsxCBVxr5S34rMOLMdG10cj/AtI5YtB6AmkhB47cQn5oaHVakob78gRVCuB6bTy4z0UrmdVix93DF9jowmrQX7wMYl/OasTsyZe9sFQPv3ygJ1+vM1Khh9lPlY3mFSVxNvhmF7wYyiHiOP3tVYqPgITmZGezrZOGP4xz4zOT2XopydZ+Vp+tcgdcqj+69OM1aj2Qa7FjPJ/s2YhSeBD+GjAAzsn0r6k+i9RUIRpMhvzUrljWYC5Zp3Ita6Y+bHcgmoRKj8hDVm+33M3IA8ipO8lb/nE5kowx6+H+f1gfwetiEeZHBlJSWe5u7v9paTVGl4Kl4zNiyyWZnmKK26nptUNncDFA8nA5pMPZkinkl9iA906QNJhCjXFeG2JAjj+6wHKENnU9hTie9iKeS8vF2nIYBiIKr/EF3vy8rEHxBvGGT7Ketof0i2LPDl8FEmghOXzDj42vFBNnFRQgtJ2TzAUIR6ZcheJRhCKuopwaaFPCByJaOIBLy+PTYcpy/0a1HI9/1erf+WlNxhpeqpDBrhxWRBAh6dzE5UVuiuxAp+/OsfmASqmtsrQeEd6tRYNw9SGQGbn4dnc2YqjO80FDPxcr1GKLfCuOZQr+pECc1rz+wmLEszpb8Prqnq7QDojU3VvkmEyb1/heZ9iEiHCdn3Y3OJ3q9VVnt5H7paOfJw9GaGA/eY3NtKq8V4EfBOxmzcRsgkdgXLS+MUtAfQHdHm3KKXIFcbGyyOE5SkIal8Icku6Qo+SqTuweI7U3FraCXNINYPPxrhEYEizqTTGoPaeYMIteFAHzLgIA6MPFyNm6++SN/5SLKAoYSnIpGDKu6B62V6KzN+5b3V5wEGvarDD0c07f3bqwS00Z098HP9snv36OEpjnxT3E32xJ7nyk1M4cVXRLQZiO8ieuxu1lns+ax2zqsYUJBr9IZXpTG9uW+Ef2Ie3JQiLl9qFZM/1BDswmBNnH/cfpTW3wZDjYbl2gyhWRZy88NPoyVYcTkFpx7ANZJVnEvUkikT4kvKT9unOoH/F6NmF4Knvxm3Pn7vRHaFTCCdGM924Vh8zGGs6muG4033tHGuVAmp80mT/o7rr0cZRbwPYC7MoSqJU2T5XBds8uw34Xy7A4JAHYat75LJTr9onxAlc5i0m5G2bYx6w+zX76f2AQz1l7f7k6K/GM5+IHtCEUwTH9qTW85XuLQgdyv7LuvbAPdfK5j2nH7DQQugeQVw5CPX3M7IxJVEHVjSyrCEwKMMOHojOnWg1yRa4sYql9CIMn4XbOX7ATredhl2gP41FTLujzPanwmrdzH444uLlg2gDg1nQCRs1hg/v+eWy6SlG7LQBICfqzdz5+cvHkzkSG29rKPp8P7t3tmHvYk8zW9Jh08+0WVmdRcDy2WL60AGP2R6zs8KiV9rUeAaXdUoZ1cmyr2dhiIUkVZtNrzQehD+PPKQo1WWKGhQERaEpmfFRnZSU6emme2TIwxBpyUD2EHJUtLAHo1KC6zedtnL5tpyx9heeBLBhZPoL+fO9rAtcbFxHX0KYWMgJZOkEatscn1nZ4KzhehV8sRXgld8tv9SWvjE6GG6B6cQN3R9DezxtmFUe2VjbLozWQ80WZP4i0CcAw3l1qlvk3SS7D0pGELYy85kXLD9ejh0pyhATKQYKvsV5sBEHxoZuqfJiw9XOEMADgH6E8kWONSaZH80OrmtMiCHHLEzZ9AJiYI3uE1eryKz+xf/KljRx1clfhTiDpHrKtLn+3FQCf1mPl5Fr+GS5OF8UsPAEUskfnQHUsP0d9oBdOLSXgFliW3cLyb4ajOsRKDNPppInRwihIkY70pVBdM5WwjrLO1rnOiZpJrDbwzXCM4VSRmx48E2J2yoB/dycKfxbrrJbgGwG6TUsemHy13ZSS0AVTqahIBg2gcIQ/e/tEO+LCuwPJ36qkbb8BqEWIxa7G8UbZzF6Y5HvHmjKJDjb/8Hv6Z7XavgLgIHI1rHsXCEdWlwXLGu4E965WfzwruNc4HK1Ln0OZknKwwE3h3uKfu4UvtZEubO7YcTXCJ6JiIUgREyV9jZbT5Bm9SVZ2OjvkLRMTAL88dUo+Ad8Sg+YM9mjFWzQOsjGFgle+o2ztS9FhbXgG5DD5S8N8SrCO+eof4I7WlINkN/njYnBVO4BKhJM0dhlPEaxoEcW9QMfe/v60PkPQw6vLDFl8vlHtCsjghpiA55Zs/y/JlDJJgYnEfOstxLxZxem8aA/9VVqPDpgh64PtuKpA56DYE42nBY74sCANIY1W/k8X+ZDZ3XS+PnJEhoQqigDIO79eadNYzlfh2ibG5fqm6bpazyzCy4rV82eLDEpvt/81vD7rmHGYyNYvM29rKi9XQVrawdtO+OH8LsiMxyGOhLtT115BKLL61GO+rDHZz9L9dDgwhQTJTJmPvsP5qP697+Gf6p3x4+KTevWvE2nKXTi7mx7bUrv9KYXd4Zt5bfffWtgSn9W8vFXe42tqNgektWS59M3run5uG0Eu27CYEJJUy4WwmNgWTTxfUl9OtQkwm6zuuAEF7qHVZ+IvBVMnZhDr5vL5r+e5MticJJNKtPVjm+qWr66+LhhvCvITf0MTxQL5Xz13eNndHWdtdX7dYXePtuoiVjINhfmusVJNq8UvRTDqDPYn7+RP/NSN6LEtuQRo0ag77p/Fi+mqvCvJARnWG8IhDHlPe1oUR2+J03sj2m+Q3B2pGpfXEGipKZczjGnx4hwNjHA3Rdboj0UGQ8lvDJKIYXfneViUnwySNpx6KyPxYd9g743W0skxnk3bv6V4EE9eUsaf5TEvc2iS9yz7AJdq3s+2XEHdzmEDeejHSl8IqCFfx9IW1xQfeXNFzNUM3PqkVyVmzkjcdLCwlncqV5OJcMgVGSQfSBW0nnuoQmSPaNYzTTKReNC2PGQ5e22RHojVCjuAu95mk9h4X/9FwQiBXEcguliHZzmFK2xJfgrHs7yppgqbJMRbfnp8V5dvCnB1+grbGpAZEe5YScTzIgvwOvsVmeoCwgZYhpsBMqQd9oyTDfqCiY3ZOnv6V9B2dpwFDacm3isCh/NeX0vNbePG3r4FCGQyPmV7guYuyVCq8HP3I6Ypm3DExVyAqB8BNitnFtQa3r2GulcAI3AN3mNHnwIvedJJRxi7e4IDIb5R6nW+0zsreYUVwGWRWaxIf3m1JcShlwS1upP8bOK4P9VXYZ0VGA0zxcvwh3imc/JcgXfvlBQfHgObk/8hBbt/BvlJskYkr0GS9U/ICltc/mCILdFgklrwVDJWjNfggtWETfw0vMkAMkuPLH3VEMcCYHDN+pWzgmupI8RO9EJ9RVEyQiQLUSONha55F5kSlogu3xEaJe543BA9kZIIGhPl1jhLjkMP0oNmIH97760edVQb1B54tErhujeMStDxdtWv1r8czNGvE4+eLmyBMUYGizq4OE6xGWSaPRfj/rSaq15RY/d1FeYFqgyhyrlF6G14D7WTjIoimiSA0Vv6lbbFbUq45BirOCM0DneBljKUhXbg69717cS9jOX0VQ6UVb798/ZZ/UN9UOyOZQcihNtL6ZRMH/dJJG/zAc47I/W2q84YOcX6upZUMByyXr/RrcmG6eeDO7wQygWrqHMLyCWt7YMb6lgC2L2Ze+ZBWRqfK8QyPOWnMGuqqoBP8XCByFzk0D2TY1YUoiGswZXldbSKkQsve2hLJrNQxZj5yYb+HcmtR1080tfiPmIt2nSiTEfmfDIx5slBv2bf6S7Y+ZZB0lPus+UA3zaLZsu3XsNTJaND/GDHKL2MM70EftsegD/zdeTdmbY1Ck2c11/VCe0Z4K0f5/w7TzSOuJYht4DTliMbH4aFViQTEqFjicsT2PQvB5dU53bS4Ewp45yx6TOWktowpAzC3cM5UtBpCT0ILnssBEUqR0UitV/P0duacBa/gBqmh3cN6pebFJibSr97dw80TEoIspyhzMAfkOLJcLeVvC3DzFloITc76gbZoIJIDEcuvuTY6XZg7G4Msg3BXh++uCZMP/A1l2RVnllVCgP9wb5jdjtsXmznOhKPsNjtHvrukmiCFnwETX8PR3kJUCf5A2Jp4xum1t+uS0BvVZN39ziOhEq3nBkn85PizkTVi8w1qaZb+T62RUDmbZZ0fjOJJsEfyMiYh11ktAxW1Z0DCqbb0+sC2ZZCqpq083tSNs/BYYhQba9lmQK4/+T7HdCBCOKpjD7ZPX7RnJN/kYvprA15fva3GFZ4HWvE1M2dladMIhYl1THNXD4GzujGmfsTrNG/C778Nt20bJjjoKshElp4U6GoNDt7ozyBCW8PxG6F6tAkqDm4IN4FQm+SnvGwHu1+C+VV9cxLhT+jF8y7+pJcgKaX1lknfaY08tZ12froMEz8j/HnT1XQW8zfIUAhbP2FuuCdUHd2VeC+ScISw4JmgIs1hWcAPZwtjj6OMLlXKvh55U40MDD8DIlNjsctBbFhaJgP5xsCRm4lOStxfmDesY1AmqooCtYaKmf7mGxRbKO1RY8tfyXxRdCK16qi5Paoj5cevaT0ZFOpDVPELs5YeEeE30W/pHt9mZ2GvEOoWVmRDoNiPzmw+V/UdKvS8SklM/0vb0wxuFVS3JDLIYYRRuU3rgcWwM9yB89ZO9uHVrX9hef+/xABDQf+KD6nVZidB0kXRsIhPM0ub+R95E/dy4t3JPaGOPq/+DlqkuJ4MBiGQF1Uca5R1iyMBgJ/5vIPF/dMfEyDkk5X5WWhWIFgFvP9GVbkEPo6JzuPqvACmGZYzNrgQi9/CxKnUEpi0qZY3w/3drPrC6OhMMj56S+Yzr3FkEuBvin21InOReqU0cXFD+ORHOUJyWoONCuRTOhw4YhMZvQM345BI8LlP+jj1H6XHzoH2JWgJuyftERu9JIcXinMhHWIdK2Cl/XX1A1tYYN6jgGkcUkKoYnvI5XC9IKqaNo77n2F1lm+tePkwMjsLuL668xABTRVObIVEZT4Jzn5Obsbhe/kDSkUQbqm6bFRG5howRQVtYHXE4jSP9ERPrXNT6d/xtfmD2VacLezP+7hwB5O67HG/qRZEQlilWkRw3qAmp+mOVkx2or1bLcUxZYTJWv7iDvlHraIBiFr93wluGabYLZ8hXW6qy634Z091hgjYvM4N/4kVtBhab2dGp1r7xQQGPzLYnUq25XoOReW8wLKBmnQ0wTT524fF6SCuW4ILYoXAyp5l0Tde9FWi0+RaNAtw0pynlbzUl/RgRArVaeQoDeFQVcNDA3Tl+k9WV13OSbfrYHp9b0mGMKbYqFb3qa9KgAUPTY7dThwz/Ko0wDrtm2zWop6IXBONfkOzRxPreB7yOfVbzMW++TAXFY3oksfQ9Goxmam82SsngyaapHLWSIdGd5O05B7vdS/N61oGdZBvoor8qZqvJ07ySKkZJ8p+Yl4CYWSZByVTNTsckxqNa3Dzu93XB/3z1YyedzPGUBjqSRChpD5dvLPOSzQ4fjCO78obKfUDt4e7BBLjr/+4UaiR+OH7EeDy+nHS/zLySmp7lAtMvOYwxo/BnRPg133I6D5hEbpGkkFXeMaH4QUP0jShrvY+xkU8K4Rx5Yuok3zl8tg+Qryg9BvVzyow4CBEA7r8UhaOqviatAj0Zw02mOPuEO3sxMNOwzIHkZ5ZT/g8G69fS29S6ecps3uHPWA/oehh9+AgYKa+VD0s2X22OZqv59g4p36/7qP09FQNJCyX6QKjNRs8lg82f5Hf0tRmRNKJ3jI0RUsv+2vP+jJUx/uI08VR1StR6UBrV4KJu6He7dw18HOXoo0ybGQrW5h2B9Uai/EsLte7+SxS1ElkDqb7tbwcGZOfOnHrzvcefllfFQRe0fsoXz5TsxsjwagP0gsuTe+HTSNseklBlEtGeWTWQIRKN4HbQUsumDw1YirA0zUKQssgfCSYmgKbKS+yCvoZvAVukpfS2RefmIBa8wrxx+ZE/5/ggjshNi1ImiLrYjNvKJdyQWTE1lOPu5azaeMgiS7p7YEmdg6lTvovlS8KSWK1M48Yknxbd4Nb4RJjo7b9/PzW703gY4D9TFy6VzmuHQwtvg/Z01l+I4DQYRvIQZHRSK/WykHtTtgzGYmfZ8Lz6pq59oxaFXZa2mM1lOaEXMScSKzYZraJHv+HHUNMyyu5RZwyo+CFYkDmUpzLo9pFmmTJK6s8FrpKxy3MdwZAlkXl7clEpVjov3kiPgwB6kCq54pnQO/NlcZDJehtSXoUoKHcdGQNQkuaDX3gZ7MSbD/VvwU0HUsRnwzvn10Fmjo6UPBXC5Vme5xj93+Gr3BKwzFhbkSnwJOIgHnwMeJfdsTB7rjvX/LUckapnaSR7r9XV2/IQXAMOb/O8o72NrnsBTVmNNqNzNGA3w7Sm3/l+lDRnmcIhpszUt5IO/bgO/S+tHinlTA5fLS7yTrozifYa8RErpzAKzDow5Itusg8R/+bn0mTE88tReTUV/q5MxnZlmd9pSj2bTe1d2BcpAwj2tMFuw58Y6D4cR2BjrUCbZmm2lnvq1DMMWrs/asYnTpGZadJ7Rye7SN+AlVeKdpBqJq2AxrAdrp37aFRwYXAIQtNpz9LuNAsaC3HPoclGUY3gyccdjw7Bx6TSJHwwRMp31jDlGWQBsS4W6z8Uu+iGld1PQEIJSl9ukQvcwquBkyn6f8IkBqCIFHzH4wOP681+7UQEhmQCKK4iRhIJ0Y1QDrxn8faAwgwmGzECXfOBswwa4NVPtv43vlwu0QNGZnunfKlz7MPWFmIUIJIg9q6dwLprqCUV6rFKvmf2QHHwJMiLQdyjN08zSiS4fvbpVKVq6tLIGj8NHuSIzZTucq9ThN6x0SPaM1AAE+vKgXSMkKTTwqog1YNr4t7d/xou0OMgLXWQsFbEtluO0LnZ7jY47JbHKmpDm4k0NG/GygLrRaFOPo98XKL44vI9indHzyOY3T7tjDK1LCnm7kTwbKTcVIzV6Mp9neFr47NxvZkzncIk5yGOrSA/9mwo0GKbfUy+bPdzlFehwPS4WJ0QZ8kNyg12Gu+AnEM83xXJASeqtonhug6FqKW7SwG0SINXKnwZvgTMiEOPC7OZFvneO7zCMg40ao+EY11nR+C5QEEMESwSgdwB7Zg9EioajDc+I2VXF0eIKhhLT9uHoC60LOz+pUkY+Aw8OyCFq0oZXJm75tI+bUVSVD3hizB/UdwpaDmoGrc8XGBNPCcpzzMqk55Qk6L/13evo9fJsbmqKyCdiTeB9e5SCnSma1FYitaZxPr4UGczetaj1eOUShYdnJpAyooHrvH6rbQoqkv72gXsPg72NRlkGfmmf7qSFAA6ogRBbSrOMb+41SExIP79ybFiQ5BzHC5q1SNI5oK8cXdasAGWcmKUckK6khdBoWeBIRUZJXsoFP22X9SzWG9P7EDHkGucZHvCArApHt+TBVnWMD6mnGlt4O6dHEgcjAkTI3kFIqtcjiGVh+F+YEIk3hthtDdYpinNUD/wf9dc6QXelu8VKmB3SUmTAQe22ZuBDpni3syaFw03xLg9+Lia/Xc9wWFN3j/tv1DR0mqK+Fhr/trUVf7VEOWGBtj1DWrO0MWW2Wng0gtDZGpUURuYtessJ+3unFsdxcZaqHfQW4lVOj6Gwfpk/jBYFWvF7YTBzrcC79IrpRx6kWvIH5LiPUfr3YB31sUUBukmZCWXxdKovCmZfZ90V68AScTKBtv3cufjkP11cE/n0N/KEmQ5VSjRJRyz/Nwgx7K0poCdkSoFkvIlX2jQPFQ27dSFyfmms5dbb2Sp93dKuykQvHez2ToRfPIksaVAMKvd6B7Xr/9/dtIIN8xoSXgWE3DpSM3OrUJdRC2mCUbOHvix/WF51COuaFFyFv8RWcPnUzWNsCjW2mYSsB+SJY6FWBoB0AdYU1nP0+PeHNFQGKbHwHi6PkO1w1Xikd4nq9ssOwLfwO4SKnMpO68FJ/03v0P5vRq9VT2jcm0dTzNKzgfje/DagoC+euhSstSpWmITp58hXTcdetIv9HVopptW678gDYpc5I0zKqWn3z/EbCLbtDEnEq8SzIXsSMOU/firgMrbHE/ytVVOv6W+NJYN9epsMMtkq0WMMCn9cvTgRFf3ytg0g7xcVdKnX3hO8UIj0ygrm0mxEc6V2cPIDsq6XmKxXMNTmgSg6hTQ6P/qHEXKA6b0rhEkMWTz8R+VFHgETaVZjFsC9IdOBt7y9jAVfovt8+ILp7i9J8CH6oByDogy8IxP1NqDC8/b/bMq4hoeiywGykcpRitXkrZ49sSbCoB1bSFEMgedDpzfEbZUNveoCPc6etFpyVlZ3+1waF0eRV39A84ssJw6y4JMGjI/ESGS7a2MYJwbARzlxYkNLWZBNaewvHXZIhMc4aknXP+rBh2FIVU1eBxoGhSTjTT73GbhRK9Z1NU+Xlb077CAUEookIIjmHWPXkqawj6R2+w1QZLOyPzUbVYhbJQ+VoOTrm08jb2lcmlCDr3IWEIgcdyzrfZIkujBiEd2ept9Zv0+us0vMkkLKiS+5hzJyTUCyinyivghbynA4KiBVn+8pqanB8TlFhh6LZIRbavQ8/VXcPItLE4Rfx853JijN59lB1C5iZs5lxNstjKqFPKKiw2419nOavG/Sw63rQgxfrOO/w09L/wRqUYpwoFCzDUit5ZDRVvmeGJKXsLOdCU8GwdNDYGGOEdiaSlNBuSvAh+UYib1Oc+NzHPb1uDRflBqGDsIGGAdo1ZJw8T/3fKVg1feF3MVhJf+c82dQPGTkuYFpS+xsslspX3gV0LAHTly4Xedkl1G/DQS1mZ5OXLZeZGzMQk9pgvyKpgTWvozRadSegjvnheY6jdS/mZ4qMpA4BYXI6rKzo/bnoNRjMsePtnn4UKffCTvSDCnml9g0hrGXpJxuw3vb2eJWermaRVxkrB2QV2t+wRkOdmSSymAOXqvY9NEERdpA68f5U4eD/TnVH83Noi1VMP5VBKNFk2CVZU9+VIuWWhaFTiPgloSichgdcpe8LIdiEYmNTI9+/fa/nOT8Ro2TnJ4lNvif0HZKUdVqXHx0Is+VaMwr9AmMttvxvYN2wkY2Ln+EHIpTvs89rNTg9QwlkZfXV2gJG7If05hmbh4wJEHRv8WNtpZ8PdPH2yIhX4T+28lPrG4OAVBdqHftC3/fNzwMTXAPtLDpWLPtft/6nsnzTMu0aLx+LoEiKxww5UjMreVYehaaAsvAt9VKcq4uk0C0g+2z2FKHdjJ97vSbtPI9ZHUEl8dJAyR50Tf2Q55PzvyYIXhLcE8T2USaCNmG3Cr4NobDY9DeSHa8PFX32nVzKrzKs1J3SEHEfYtRqyGd0WIAzB2+LdCeYWG35qaw+UNU8lkrYTnXzDtio27oIzHLLc3gmb8Sc0iRkvgFU2XrXvMsS+fgHBbY0ZMERQ49IVOML4RRBoSC8MWi5svE1WfN+Fi68gmSOICHeTKCuMHmO2gS3Reu6mvBbXTsC5HwJJ9Z5hSusZrfvuls1ZbN1k6I+QvixAsAjd5AeqFsf15n55jnZ7AgtDG9aTDobkCjk/7C2qG543QaSsDiTSKJsS+je3VupzdkLDafEeh5uKevOCabsqCIRlKPsL34b2+0r5nMEIRarF0gzVkIG+3V1IOIVqmro03NExgzxYgr874X+mW+DE5zgTyI44peCPZxC4GAoQ9Zc/16nDeICZT+aP9ml/xyckAjI+sT+k04a83h+F4fWhVw2ZbAViueatTQtj7x1KjomJZgKpv2Yv7R44Iwl8yQeKHyQ/fZm/IoPqm6v9P9Gw/DIg1ujzAkk6WwL1NRxeIqWQmEu8yz9K51iN0WWgcfi7v1K9+UpFKg9ZWhVWv+D+MnsLUp9XeFPTok2FJC74RgyDJTjTrGiplrhL/Dy16Gx7K1MAUgComQD+L9XVldSkbnqJa1LZXcxplO8uBVVfcUjhqgwen5Y5F/gDtXxka3DkfsyDPD1MNbY4sz+KwL1/S8vxK3iJJM7dDwcRHeHf0N2tV/JYGn6U+fv6d7/a0bjb5fff3GLd5mRaxknoqdNW9bEZ8wgmcDerjyJcSgOdC0snFnVH/rDKMyn/hsHzJGb7giyYY4d2xL69WSCVtn57DnUEo+FINM69VCQ/L2E8GFOI/v6tkeefHrqygYMfMZfSLb7PF7p2FPnANi34NUKIYKqlPdza0blUILERyx/r1P1RXb8+mT5OP4cgFEVH14V5vbO/PfQEXR7AHesxRIk9qNKA1usurpwOQ+VAwqg1PTCp0kktWdA0mSd4YUombeHqOSoo0uFAv+tPSB8nYPoznQXmQ46Z/nW2kBYtraYRfFbYqVINEpicBpS/bNjXjK+KxGAS2sOOdYSJiGRURh80R7uYaN5tXOB4BeLgaNq/VUngMFS9PyLC4nmtraUSYH65/3srmYAoKn9B6P+QAcoDPBVL6qG4JoXnnRwEAU1lEePhurw/ad1799C0tl0nIrbSxLv5sU3bz2npw4fz2w6SMxaBQwS3Dddmgywax7/On9lKlkeGKKDTykY+1FhGIx3qkm/qURP9XGy9io7v7mzlL67GGy3mPerN4Rj7liunNm33MbyhUkbFizVZkK4GcCfyIgYgsqYO1NI49c012ApsfSOxAY7SH9obXBNHAxynBqXeT0EqiZRj/Dh6U+sMMK7AfS3IV5VMV5cODo/20pr1iOf7smm2/Yg+HFmeaSVuVjwepBVXsuWewWQB0rE7HeNNASNuCDL2Pgj5vLA49HVlUA1CAzpc3TxUG+xlNXAo/O+9UaAisK3DlwwzoL9J3e4iPvnem+fxfgcZ8NnuvmbdQZcw8/liwu+HXvCwwZeHBAB9ddWpnBKTclXsRgJQCIQ1cv7MjTxSS73m0PInB9yzzW0wOAPF8oLZNR8i4SNSgpc3tWuo5JmZccs1FttaAGNaGjW3rJzaiJzIF3l1N3quS/NbVhtvqDk4SaNmwOnWCF8XZKdjDwwWWUP+02PC/eOX7HGTeTQAT2cZrKQSgBEpZUpWc3AnxBip7mWhphSb/CQhzzkzgw4Yeqaff6mYO+DGnMqvtcfOPyIff2lFUzLVTLpvbjqQghu2ffT/xMyGtvXz3I3FwAOMT27ftbXGLGxwBg+UcS3YRF/mfz0ZFADzAbIq3ZCi1OCKXUF1Q2/4WQUtoyoPg+CvRa387BAlklpzPp/ELxDRZV6IPRyepj9fbC6KuVdf35DhLKr71+ZSnGsm8Y+0XDwFrUB5L5gE1qQv8TIl0m9W//LDe6xtrLMt8tt9YYJ3pYUcsGiBfOqV/D9kbe2f3B76eUCwc/TxOeNCn9kkR9FzyoNtgztWz4UZbvfIMdIHGoVCJCqcggCaTIZd4AtuFL+1X32vLklhkm7BJ+7OCBxa8wM4b3V6CI/O5rT4l0USoqjGuqvVz/4r24Fs/7mxlhllD5iNXGVv56htjg73ethPUBps1UzF+G7ZgPoFGqphQZM/rAAr3UJEK70T6v19qa3FM0AYBcWr2WJbQM0QtRmSBAgVtDIvqXMz8v/LEmCMNCtO22OhMh8PWh/GGXeeyM4U+N7j/pi8SnnCKlncQkvAq3kPMCgDhULYSyETGEMstGrXUd24ts++IBA6+RUftJhdYIJ9sxugMm0IHhTe0Kg/Ook+BvjKa0MV0NeUDOZpQucD/Z6nxRHZT3nS3074fnS93C15US+g4nYGiA4ZJ1JDy3GZ9pxDvDefW5WiY31OxDJ9ND45icH+ZrZbuivktCKk7IYzH63WbLHB6vRoguU6qrsHEDI8hEQyMcqSCT1f8HNXvPWc36vquVqy/SfolmuU+uPcu3DlVjNMauPqZ35V5POJzGlo3WUqT/7UYKg1+9QI5f8dyQQR5COf9ZKO4ZJghM9wbX2EkoBICloTF0F3ySo+WHIV/O01k4xetup4cP7xvwJEmHmEg0zIvQi4t7oNoV+azs1/YJj9PHnAtU3GyxjAfBHcz0Wk6pq+Q4d9l742kLI9Wc1z7mTnSdJU1FawCtlkgXqYCkVnYHPM+6pyTlLqNF60KPA1yzQWjL3HeOAR8+rCi7S2hlrkz88/EMgC527fbjAZOGnB/760sdUyyi7TA+E/l3ThgsSSiV61aVI9f9o6CvZR5TznoNeUYPRFe/5h7Abnf9Z6T50OTtrKSet6y7PeWOEaaYfQWDOvWE0SI17GtM+FFauowjkFz1hcxjKPLKTS+7CmWu8TR6nFepLUEUtoHIyNErlDTL5JTirTjdRT+9c2Pvebxjcrky79Q34FdJ5qvuifEnxTQkbAVtsblYcHUwfvxjjUjJXs2ncl3wPCt/uW3mxB6kjIwOaoV6+L9sSPWS9xqB96VkVP0R6CRPWPhCMjTYXHMJVmM2WjL0caMouioDbgoyIKJaVSuno9X4wd7gVvlNPhGfxL8+55w2gTX8JXcXT+1kFzBSZoD3JVPoNTHkKHwMX3x1C6gxJn3ocZjz8uYou09SA5bat+9vTXdNuv45x7hR6VEOdsTUxByw8h2MpOeK4pPUdfnBomO+gK9RpEO6VBl++CyZqfCjhd22vlNXmYdYDynE3dnDWyc3PIttgdqKkrudkA2OcZhSVV9b+D76Y3V/PYsdCARNrL8n/W4B6yaNUpOuWDDv4z3Bv6x9l9cf5URpJGmwQkyjayGJi6ZdX6MZ9TEy9hJINoc5snaJqx10ciqceK+/XBabuq8pQAFHb5lYMkE41M+2X9Ez0FDdn9o5dMJFUFk4wsG23BcIv0pHWCLWXF8cv13Vy9JVHpo+7CKzN7FTbvjbC+qBfP+oxs7ViySv52r6QPRhq557KUkaq/DtdNIF4gx9yDW/goTo0nMotS7rv2uOnopP4E8upw1GJ+qlCm4qtifBXKMs36mlHn3jlTRmminpMsdfKlGmMXVl1sWexu6Mca9QzzRplo/iR6bbHAT1Ang5f9kii640p2KYLnR3GxdfNgk0pzxVK8x+I+6cLXUqwSkZ2XsazCnxR3mgPZutRR4QZ9JmVfNz87YpA5ZfHFM=
`pragma protect end_data_block
`pragma protect digest_block
245fa0877bfe8d258cf3c20e3e39cf9e77be2a9a97d435aba225b53864402f0b
`pragma protect end_digest_block
`pragma protect end_protected
