`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
3mZolDjIY5dg1VDfb257bMGFdkHph7VpCP7OfDfPW5bf+wzBDGGVrex0/1uNlJoH7DKGVpLb/Chr0089OBKWeGChgxwPj8iH1VpZMHtr47URiB+scoT28Ha9O0sSFemd7EK/tG/J4IE4OD1OCkdw3nB9n1I6exLFvCHS2jWpIYY8jNWf7wnHrSINeAu4S5Gfbw4mkHA9cbP4Ws/mWvs4dHYGKvxTMDiWG+JNL9nXRlENrlDZ06AiHRafwFmdrAqNvhYS+k+7D42DYLjEEKfQl9rWMobIg9PPbgC61/vY42xM+jFTznOv4+QAkuGcSA0rVwrrsfKgLoAJcDjEtARs0hZzwBILc/uLcBwRUIO35ILvt5nZ1Ihb4+cqxK2RKtnKI7UaJWsus1M5gGEU7AjS8ZVWs+05itFL13ncBwyTiE46CQ7xPkm8OIkf6fbMQ7FVruW4RR62dI7kSq4O2ncXEXg8+f6Al5pvr5yvtnNVe8Kf4UZmLXcXA24Hrxd5V2/QS/BHMssBcdWc0+1QtFL0f+73MF6eJ76ukzZf6de8svzIfOvoF2/5KcSfDFsoVBcd8ZeC5b2SgoFZU0Y+p26nz5HLrlA075SdoojhFGo2k+XDCDnWyNcUoFdaKcYwcM7QKbdxnRs77yR4ashzQu4N+1td0UoyRDv9D+2L8PhvSLi9HcnkXh1oRAZSae4KssyZU0R9d5rm4WM0ChdVnrMVMurrehLv8as/h1dueJrnnIVxZgIQd4DlTBUe4vHNpNVqSYLzlH4n7fa7Eu29GGNW4ys/c5wuBM7oamdwVfsCQA5BKiSFMUy0xKvZ59NwrztExUDcylo9/PmeWy1UgXBoaS80hismdXomlpVNG9v6Wsj2n2p5ZAyvsx7LZcXF/sG8AH3mCV7YPoCMi4rvKT7Udthiz5cg2I3v4jLo4rlofe1bPEQLXGdWcDhyjS+j+2CjiLdNpUp1CaojfPgp59yRYpegTwhPQqB4sKCH5nPxw38NixQ/ngCd4N/JHiciL0zLFSs82o1pyaL9uGeNJIKyUUO0OYfCdv9Ai05B1cmWFdd4Ww128+oXFmHBnrfdJNIK6WNW7eWXD1JgbTZKlNk5nCFobz7g07y6k7B3WrEQurKGgF/GMJRplBMdNbCOi7LivUMQZBplo2+aAWHulKY1avCKDA20YT8iE/5AN+PECvS1Gy3qMojmUfHnvnc+zdFfO/2c8+WFdON0uluyAfaRD0TggtX+MvlkojU8TyM1zs0b9fy3xqC5mVBraxdFtEhwz61uaollH+GD7AwqEmHu6czdHzlc4Ze7FMB8jHdadorLJvEV543KgX6MUaZVILzK6iUYTb8dniyIOKWIqugOrFAtF7hXqXtgw7vSU6LG8PeqcvCW/zbKGh5gp7PLT1SrWJneb6m/TdRv7vpaD5Ck/O/wOFwwpdmL6FFgZCQCnHpQfEJMySn+FgBtTQxTBAX+dpfGToLJff8SJnIcDnsE/ansidEMYeqOtdrlXaJjES7mhGEwvTlpiy7eh/U6x8vFA/EHZ0LMQv0wV8tUm9SQltGVfzxC2lnLhsDi3kQrZKUeDGvp8PwQTdR2zvAt5UBgKxYl4TiCTn4qfRogEtuVQ9rXjis8goYa1PYmowrLu93V71d46DOd1vMn6OBqHv7RTYGo31713fZndTj5P4qemymeoe69NPbHrUFM++Vzh6KHna0UNrc9OrZSDQPcYdtYfE0iaIpiAo7Ly2sK1n9ZpkKOopQb8b2Q9dOIRr1opb1y1UZzLC3xYr/wso4C0fnoZzN4RunVRw2thDjGZOF+YwLTtDgjRbfKGLKw3e96f1fUIutYqk+XrnxKH06jIHGIrOK4tTgB17RuzEkEc0XoWoOdjivxyksumlcNVRaIxMlJtPx5Pi/+YwxSpOWoWRuvzyODsqTz9BRZeV23DfT/3FslxbSm7ZoXKKNdPz1UqJw0Tz8ox/WpZcp0YU6pJGx+C8WBvw1GeVv99X2/7y8ltaLEfgSNlZqNJCnVuGJ8Nx9whgPyGe+im+H9pyKbuzEAj0aX8xXIdCH2IULT+Qe8PYUCpRr+jUITOaBRQoLHlsb+Rr6FzQyqzQlxnKGlwu7uf6YpykkvD9OtKgsqssIOoxqlzL5DgrqwNzoF23skWouKAswTRTLrXwL9aKN77YKlzqFjvEqyQ8sAfCR6yylNJnSnh8V6pKRadYkXTmmX1JMYC9iXUAVqVmhE77r6a3NdjeVI0+Qax8KIJUv+brEeMM6IHsaM4WsP6Vk5A0Fzhd+JE0oKaIbACm1LsBehg71dEHLsdEha53hW4JKuYSqeGcSOfnWZQwM86CQqMzoAsfSkHXBsTnYsHdVQEzBrEeBTSi8uN3+3FKpV5I8sPH+uS4eMwzgdSumKT+kJc4Gh3hEvbG+1/6pnZuL87AVWvo3MPjb6Y0kjdVkynuYoZL+1vXT6NBFp9iw8cpdSZAU4rugwFCdrxgmq7YTXlhwi/HnXmxCEGdixsL1rIUOi6z+vgiO+UfWoCIm31Tms6s81Ol9pAVzmo4Owfb8bzQg6AxGbpPkui+Q7DvREu8Jzei9XmEdWj67MG0zoOpI7RmNxf9ZAhzKGBnGPorRlyM93ZkcRZnk3/aOCXX2Xk68MlYgbAVCFw5W3e8jxqatR9WeDbgyIpZEwzpMs/EWoerUrx31jX71n5rtvd6ywBInANhi0olWrRkHskpR+QG+/DFvuLUPRzoNtowjpFEqpWnOlKi+nOVC9ycgrtapI0+/rRIbHZ76kO6XxUwxG5k8LhduEtz4eIBlxJYi4XA3+Ui3yWq3g9gPkxtMDhS10+0iUzPuCC31Fh+HLUQsbjsa52Srzupy1feOCkrW+YN8xowQuqbsjeyjN9eibDLBoKmnFoPMkMaZnRTLGSobtBr7TnqR1YCodBZ0jWUZJQfT6S0zdwEsJBdM32VWAUlKa0t2jAOf5LUnrKbt2QExYRe7D28mm7wBtxOASjNriCaU67CjeyrAVNvAolAuZpNKNExePKizoipMNNb96CAR49yMqtxTUAfgJHRgCegyKV6iKZEKcwXBGDJFQL1x6+wVkEQxhct/Zcy56ouw8Mn1yRSfxHwt8hdOTKA4NsedE0kcesoGhWkbXbO1yaS2c1zAJ8tW0FIDg090WC3U19GN/sb06nup6REjXZXSOMzVb5bPQ/LH3pDkn6qhjtBVoUthCcUvs/iXE9TYliwxhSSCJcNh4mnMwgpJn3rd/Cg7Ps01D7AVWKaLYF/aYmctJHcgZTsGkRXRjmv4Boacz1BDaTZyNhVykjq4l2HGkeEyilZ770BuBjOCRz6yJ/kX52ehXUQAAaHkH2ZbeHY6PX6sphL/2BhKkRPvSxNoM9M80KgnbsvuK3W2H239EygGPBp0G78If1Vm7SNvZEGSv7p0xrDB4dt1y2c4V52Pq5a3r7PfS6r3cZjNAzeoMLfJhG9JQEWMfqdCWH8KvR1CHcpMdXVavzqlOsHuA6KZUunI0Wh/G7UzIoiwFav/vuNiRDjO+gGU2rUla1qMqykF/wPfSdyer9528kr0VRZ9EbZtPqI8bBlV/2kbHBR27OtfvQ8VIQCE8A1SnaKG3/dbI0fzEzkkTHNlGUrwxFx802uyCInBw85swFyy0PWh8voZPJH7+6G6yRwALxs+/rSYTCbrIHM/WrqLPZj2Yn/Kz52JNRjtrE8ruNQ9bcJgb226YV5vn47L/0zxTOYMQdFx24veg2sjhEcH5hNJn5kMu/ItDF7A7w+SVJdzjDpQ7JkN8wg6gwY60IW+gtFN37MVKdKj7DiRMU09gUI+fuGV2k87B2Yoh+Seqz1IOmKCrS03ISzkQAAIVO1ZDTdJJCOOWgUiLPIeFrXNZsJTofsmQ8LowzXazXvEbzzbxYKoAdOpObIWgI7BODptwxdVJZv4InM/WQn60mx8IsVRtscdGU0DrzW3qMALaFzwz8fOjWaimExUoET/cE3cSsWVNr9dfOwRnx+JM54QI2i/MrMHLL+863fqmRkcWpxa4LCj9JMhG75mUGFM1wNM+hXY2gtYuFqscvEwOPsX8d+6MKBoRl5tx+OXKAdOP0DC/5Rs9PRPZI4i+hlv2+vZ2EQWZRAuZ7GBk5p6r7+uIyY2Zv58tat6WdmDIaqG4Iyel+8xHqG7QJb+8EAi6GAE8DPAMvEFLA/dhu+R+34a0S6FvCIcYd/ZL7e57vqG0MJelyafdIDQW4NU6h/uvsGrrDasRZ9e5nGO22qcDHdByPecaiTSrFXWDrvFBxER8Oi+PpKcaa20q0T1AKrzSN1AcArX/xhW0u507Cr8QaZpTAUTUogA+/BEsx/2dhqaQ0joIB48HBnlBURUup8B+G04ezjZj9aDjzhZRowaW325P0bghAg+nKqlfDjsZ5Vn+Jvw5tZbUC1utbj2NJ1c5A7hv8OqiRwaWtBG+Wjaq+ev6rpw4eSzd2ueCTSf/w3EWKuB0OkNTIXCoikR5S4Yc2hqMzvhvRtQAk1xV39JvlISurU6CQa6uOoOLV5ImW6xgbWCBc/QE10ATe/uu4mT396d4vOS1rzrAZ2v1lY9p49x0X3M8Uiqsq15USHRYTVlCvGs/Mp8pp1QgSl3+yZlwbS4bD2sXhibrwgPEKB5jJK16egWxJBFX0cboU8aEzlO4gYXpDEy4k/EHrT5RoVcq3+UakyB8TWahQ8MAkpLiOj/g5834S+TUZUZ01Wy+yHh/q1lRFL51TW1ZnzPOcFLx52Bpk9/TZZGGjHyINnPuk58ZaIoPqdUcVhuJtedBAruXUqKLW9PKy3SGdGTO4YqQC1lTswAQCf6YNvCqml1G+uIaRrIFzOazClull6ydvj2bPqGZKXsvae/kLbunjsC+yQ0XhFIOFmQivC60wsJ4s8ZSo1OVxTYlI87qgvh7DCxcKXob8YHK9Iyw4fJMK3i2wMyldRlbcOGe5TVBSNS83kUGHRKar9Gnm5vQu0g/ecz/++q3xIUoogI0J5idHJs8q1DxBWOAJO2sbGcMBahMaabxG3/6gv9wWSQP8Xml6KEKHDi3+6BJp8ZI9g7Y8eQaBkIOiPEOX2jPvoOF/yFU8Z+uapfwkeItE9STp1sukwULQtqVWbzoPBNxcVT2vZdErwF2brX2dovoZEvvPK4Fd4rFlVyxYxBElIAG80ai9wu6rMqkIpmevNGmulhgtgmJ/+rTvT8YOoPREKAqRaqaP1Z8R3xu1IRpb8OjYB3JKroR+movZJUg6O9KZsC4ZR265aZiJZ3E9YxsccJVglKGx6A0Xkpae5WyWrz7fNRfiS8jxjRDR44X4f1B/4mgwhQf/9dE8WWLOsfXxpxQG43KUSdUfDFvVfdmvoPMuWiNc+qxeVC78vmT+XniSuLEvC8l+V0vlIzltLOdIzxzXMaHGmQhbg4Q+6vetbtAkkBFEFZom0o1ZwCQKVIA6f1LRhF2rTLH3gfriorPkgGZrDMYtpjCurRrKG3dsX9OIaoc1ZSDdz1KOiK7wxD3i4hbcpgE4q2PHKuwzD0w7VapGr/opeNKxqMvw2NkEdTXhR/Ibkn0due6XX3UtsVIL/P1sooTWZf/2O9cv5T0pSdv47rGiFrudvLEFF4BZ6M4gNhAh0UUdGlaFI4bGGWARidoEfyeEAp9nYh11Ne+b3aVFP3cnEKnDrWbR9oZCpQ0VBz7ybSQ2Lu0G73+RLpDo7wubdk0InWbSdT5aejZsj0LWSaHva77JNQ+Rzfc4gX3cu4NDUMZLJdQPK+yI/oT6x14+950IXj5jFroKTDVnAZkps5TzS4A+aVzKB9ZKrV4sXYJ6I/Xg33TsTIehvwcT+mIQb5k/RUOxG26JImzzkz9DTXfIHA4LkDGECqrUVvcVuSzhEke809lJrM5Wby8cNwxV0Fd5Uhnb9km7CKO7o8CGkLZ3Yr94jhj89DEFnViN5Tuf53hGFT/wPZVHKL6aMkajj+yxy9GdMf6vFSFhh8yi0B25CjoO8a7QOL9wK/HHfKckvGR5Cgv9dI1jwVphHTu7OBx3F1fD9n8AIJlzjyWOEv5rZYdZjevSHNk/elHYLr/izGuk4xLPLlgyPqHm2RgrhZhafyZ31FNXQXZjBlGmSr8i+lqtJ9wQAiHdpk3GLIB3UfUvHc1OM5T6D2MwI45+XfVbkdpAIV5S3RzT+uBH76Ocfbs/fIP5MUEx6tN/cCd5XSwE4DEBOIS1vtsslPkKYEGZ6sY2oIvAQF2PBaD6Nw1AkPEiX2kGIsjeDjKcRcBr1oJIGfzlaSw/l98QfiZraP6BpHgrG5G4rCmNVqB9EzC5R4Xk/bjDuzd40IFIt6BNgAmrOyPKA3twJ/rSMwcWR063jA/5cMwoG5iXT9lrEtcEPohMjhDpHQo17WmAlVO+8Kw4ZwtcmClA8f8wL7FOj4gIh0LWDs5p3wl98xcsEOge+Edagj9LcT7faA2pWQUDvcxTG+u/I3IdaVcZDWNCKduHLIzZD+RnvqJipNxBQalhZUhJleOeLJhhRLCOKYyr24sIk882nZW6gMvolObmF8HduUpQumyDjySxCVMb8rRXpzFSyFea6U3pMzT3BaQqG7QZegV6/aLaZVM4mbYCx+yj7v6SQyjyXN0t5IWVCP9gBMLJjnyHWEA9/E5XhlNtQcfSz4dw+31x/2uR8AYRnEU8Wx8eO+7cl4dKTWhLj/wjR5PUQRZHT8q4oXACHhJPjFYlhcBkTzMAPzNqcKD9OXdKKWgug==
`pragma protect end_data_block
`pragma protect digest_block
89aa755a77a1d490d15bec22f3ad9b325123c6472bb5329efcc174a88ec18f4f
`pragma protect end_digest_block
`pragma protect end_protected
