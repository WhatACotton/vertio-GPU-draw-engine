`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
S+UjK5u8tL761aVfakOC6DhMCtzrHa9vLzq4e3ceSm8DPncDo5WztYI+bUuZYKUl1BIZe5kIlhGnT6jUD3Z7+9069q/+gBn/FfMkxeNCyD5bXRfeTn/4gKwZUYyIqW89tbV+sfR+yo3jxDXtEen721K64giCwAY66lDQdedX8qic9yZbY0ndUIjN5ZgEd0vLU6xCSU6sZ0gg+v53GrJvovLLWwMYbkMSKc80TYYoFs7CAMoQ7V46irT7L/6uZBQR523XQT6dkCdZmbKwjiKWZCsd8h06QQkK7V+YVV5ZxHeB5aeigoVT+cV6mwGmNIpmE9o3ywX0SzhmguXaGk2TFTIKUThYsUU/j/7xpGCvznkBrwn9Xu41f3PKg01mavjRdCyLtAIjhK3XTc/vaV3+xt72ZdodUq9x+hmebhLpIISVFbe2opMSdyCHQLQ7+XhqscQ5k/OZuWjLbpRA8oJSGg6nzQ97DWY6tuSKzVtNLPgf43VfJqody8rNl3mclx3G+xbzRtOCdmnWhG2eI4nky3uhUhXcmcfrL6qCeOfdjvQg4CbenvnZxE+/htDDgXKizMgsxPtB4JKyRZ6jHxi7EeJKPrxgqj539PajFaamsGFqC9vhie2NxHTmz9M2CVVOEuDsWB4UYheb6Ry8gyj9qvDhgpZAwnhWnbqkvykhEKY7Sze5o75gEbOaXIAnAYwAtNMok/OWG2EHmh4RKoP3azpBNNPuEpB2VwPG/qD6mdGMnZhbARTknOWfvfewtp7mrwYDVd5oSOino1N1Vng28kqg9bVev+4vBH3H1mVpNhRYJ4ya6apO7h4YqYrE1ExcYzFybzAH8Iip4BSmAiA755paqHXMOSj4ZOiw/7NJTvafL9xpBVcN/KuMDUmEHu/IQLLq/NG7BdPDCRvjvdxbWGGnmWyTVbRogx49rDZW9TnVBlJ4gAu0GJ2HPCMhE9lU5ZGkxegJyYF/Fe5JvCoFnLyhKTJyRgwsbR39SLMkT2Qr1mz8cpqgRCLNLqFqqHkB8gO/IlTXtVhRrssxwu0YsA84Ixl/wPqKN0qSKnAAmutOX4SRVeBHc8TQ4dLheCO8366ba2GK4kaO9k/njlcDBrRK2e2B9e2hwibe9My0k3hBfb2cYNWYgwtoQWDNgicyn5n5EviBpnDy+O/+YLi6UuQaMzfF6jvnU9vkK3sXI7fLJW72FcYR/F1/LxZ6Gvm/zdAi51GkZiD3xvmDur7cT11JS10+RtAm6HegrF/Uc2aKO5TsLNUf/vw7sIsBsSSPA3/ZR4QcSyieElNvBeEr+kUzR9/xGUYGWYVGhwpxUsoBHSvJmjTxI9YybGYV22oLEjbO+LlTCszfqETn0RDXX2qlyIMPBtTMZ+n5TKu9SaPYBpld1/Es/mNcDqlIrs6ZrqpY6VYiCqLHcS9SvcOoe0I12D860XubOEJOxs7iPfsTKDD7uiC/9CdCLVQ6gNO940cFtZm/NeoF5Ve6BSOugieKSL2yYTTy2tqD1yqoSlzatCj4J3jXI0sduOIkvPo0dMgH5OeBr3ty8PDMRrxe13BP0Uug1Nx63wj4pXedE6lCmU5eEkg50zhm+gwDl2JSEWA0Bm0gj+gGVXb7AuS3uST8lISW5R6BROhzGtvtfvnoewXXW4TqJWa1wt072JAVzAm+XVtB3u1H+5ujtA9kiwNLSNy65AO6jL3kO57LOiCwox2DKbmtBXE7/RmnpftBRfooE5GhYUrh8dIY4X4gVWbJGPOjWQBB92Tuoys3Gh+ZLkM8FAo44BkPdFv+EvjlNe6XC+CTEYq5aEITkWOeBzOONRLcWVt7LZBFp2gdx7wyv4zQpOSgMkGop5GwMuo7MDrzpESXKdpMgVVCrbXiN0RmOIU0heNTM8rn/OApzAv+Q3tPvJ/PjGSguHZys/vWPgAEJhVpw2k9z2yuARah6Pwtsoj418Y8UWSekndsSzOP/BOnTf0Z0FRf4OaS5DJQJN23q8Rqqaa9EHgM7JEm9JkJpzvWB8OJCzMoQb4SAZNpyiRIxxN/GYL+/2n+LBTk+zA2wZxTXEeUYXm52qGkbD+NtY/X6bgogsddiDX7yP2aTiaHzYvvRpfXoDnk1gKy5R0notmcCiPscdytSBNUAUl7GRjyeveD0E0ZLyUp+mW+Cj0Y+5tcdxnRdK7Zej6PMcW8b7VR1fSka+LkhOaPn2B/7dUYRDRIxm/7Xo0iYgd2/xUsR5M7l3KgJHocyj0YZ45htzb+VHB/jhBR7IT98fbqCMDwxTdNxuf9eaUFGa4Z2Ois/POoQluPbcx9IOU/YXzGZgDrYILlyxuFJyv2JQxMILwfVwBVDtF2gwlSndDEyh8ukFumOfb+Unq7QOrZ1Dar1MU5aA2+P0DBQNiKQ4W64br4sRCf6Nx3pB51IttaS11i6DPvkYa6/UEm4RzEBO5iA2JHoJTEeIpHw8qWcgUDHyXW7XqHA2uQvPlOsmkxPj+LyEW7LY+i0PYtgpfMeyNo8B+jRk8TBi/Wllt/2OmrGW2xlyU5faSCnUpN863alyVCLxbUZtlTOiBuwrpRwUxPaBXXPxT4ZuxVYwWbuoXCcdv4yfSfxDCrsHxnftKKkJlNtKGeP20xsxyfo4oJmBaLRh5I+Nb1OW1y7div5HBfT19bgdiwBiUrBYeuaaWQ9ishgQ1EQI7I/ojl8xGx5C/4RUT5W5S1C2fVBhhpp57Gp/8+9Wopv8fTRYx++rXfH4PNnxbees6kqDLUpdQeHK3az3WEDkmiLw50FbDfT7yoZJt2C5LR6bH62e7LUjqj43LIqzYInv9vhXalVb1mw6phRgerbX9Peb+rYu+QeUdg++Vq9eBSVki+qMuY+vuEgR/Wa2zfMf6YMWsaOKOfeiy2CFyh42VumF1Strih8aKwzqfweyDyTe0tPM2dYfVyyzu5YxswhcB9MEr7BWfq9+fkvuG+wIohWqUwseAW7P3dXwtT1ur/BU731Bvc5fK3lGldi9Cpk4i52MIDI0fKX+33WzMd48icaLQxzCOQHRJB6/PlYDYHlkKbME73zoCLF44bftnxt2nuBdEXJXit1SbFiN5Qowcbrd1q7n53Dk6/eSc2vQUTlzNatpuidnAGI4dED4PSJD+bfGDSCYaW1bYg+FRLAtozlT+3MCEabFuOJkMOiAYoC5KK/wFc83B+dzoF+KQInFU2CE/1vQ35HuNH1l8U9zYKvWOLiqe4bV6qUqM7jVp3iU4mCJo6kzc+8kiTooUH+1CiXGOUGzR0NNRcC8gRLqsujrdZHSageqV9tu97Wrx5JpE2UjopUj0n/xVgfcqbPbfu3rtf2gQXAXuYcHftawIhYK4WG7eRvUaJv8mTvwF1YZWanSqnTbBqrZ4qcfQJLtioMGQtFiHJnJpeHrPDqt3mPKksooPdXZvGW3dTZVizXYlGyhcI1SnwWcitc3oPFUb3gJ6ep+jkPIGU0fr5UWgliBhvRwRBb0Lbg3qJqPOu/rO7KzaotTmIcKopARmw6LhJkNFteRkPlf1m9Xfcpu/F8ynAECKzLLeWDl4/gp19OdfDcnaaJ9Ca89sEuwR3ARQNBkYxv2zGp6wMuI1GhpYwFR5Ry9wR+kSuK891zgUiZxohaDOn4gG4sac7iOTDZI4ctxdSLW9qfBtgGtqvJIaBHxsC1CdSmI0ZSr5gBVDk/0BgCJ7FTSY+X7AsgA5YFe/IuRkU4nHF38myCTwIEhLTptJ39ZV7pNwhNW1VpVy4pqg6sXSr7uYilys1OTLTvz2FGIu+U3bhX1nGytm1vQlHd0l1gpexbgs+mSyuJdSv7ij8sKBO0zAAD6C1ubPhnS1NPO73jG47ZeFz7GpDy+TC5ZUs/QXMuZAKQ+J9sGY5UMNtn9hO8S7xZEynigzJXveNFMl8dHU45tmYQ4Jy56w3MURM3XvbNQgpnHqpi0/m8dWdgzjGs/pLMCvgv1nL/CY9PzudP1Nwui1kYe7/1xLvBN7CAP1JcnEnMf7uhYMoZr8wS49t88a0Ed7rSsP8B6bB5+AYoyc/CUiQ4xDkDVAZ5z7kprCsAdHAFmpb8ri5boJnWf43xhsYO2cU44Z66ngQH9+ficaZmjAAMhqAZB3LzVUc/8rTiwlW/NqpbbsWQuiS13b6khg4Q35rTVgpg+Dr7TBjS8aUFSqiEZlxD0YDL0VoTEncpgcSJ7EybRwEhtV3cd7uj4Zt1fMJ39epFiqvnkE7E8aFlVgWMNjjBBiT4gXw1GNXuLQk0trzkpuNLrtHrq0qX1plhpaHGHhoDdciwqll5gxG0eA3vnTOV8fvR5aSif8Y9Gn72zwMmmrJhbQbYpjZTsn/uElFpf6a8qtrPpYi2kaUXLY+SIbbklFBT2gKq8sUhVGPy7RtNPNb96jUEY1dL8vGOg3JrMhM+5Qgcj5YGBORmzebbel3r8w8z0S6i8xuqYYIXCQZ5Yl8Vk42MxZ68zXvv0F26uXn4NL/3ga5ogQPPl1n5kNPh5y57Dq3WTPdV010Rh1QQcRwjShxjSg1FizZbVIK0r+dFdWBWneGMI/7ZKwwnDcxrm7Hzx+CN2I7uwDW4u6GpZGzQ0u9c7acxcExIjAiyJqP477UlF6xgSaOm64zScjFZcRrKpFgr+GBCt5iU12ql+mLDL5sRHntNxZMeib4EwzuGeVkLeEiShCfA4ttC+NfkT9C35HahQbEFWiGMMwKcYWetLVn3Ukzb5OfWbWfsJ47836M8E3DA1Zth1+SRE1QRrWfqWq/1TKSsu7YeT9Q8Eu1mbtJTHbaBG3F4qKLLfIlth80ExZNEDDSTsmjhA0TZYaz6KfgxLjAeljghcbG3MurIzNoqFospjeiLTQ8zK52IYIkojBScty4H5F/+9QMYYin8aTAiDUp3AxHUfHIv3a0CjOjL/0R/qzZtlcxmh6Y6WQC7QH6LcrtJ2sI7oFctkY09VeyQ7qzgfMKY4uj4nMSuJMQVdW9zptIqY2orTnhsQJqyhtf4VpuZXFFZnxqNEAlUipmS6uERKN4JPunU2WiQqpEO40m5rBDEvRsdu9w2oa+RszjL8ZOW65f/U8RzNJ93f1NZsDYJf+tI+AwUenf4LYX2yne1aoZwVfpjq+ZmhEzIZK1GbV7XZyQ29QNB2mN5pfoUijaCltlRxFcG7T/8X9XBppXfVXA32qGysjET+3ueKPIFVJCvayfN9catirnHFRlcZHzkQDdoVk3WdWPvhzGBdk/tlv6SzzYdE+mTsjw/atDStkADgdnN1khF2A2K6mxu8MH5kX2ozquc7r+0uJmhnE/FDuXikfFVPr4cOElooHQdH6oXbbG3Vr/nvhTqMdpQHoHxIsaA/0onSI6uWTxERj/CrQjCf5b04kphXqWn58Z6ozhrjA52zP7jhbH+7MKbeW4rjs2uELX4Mbu15S1tn3mYxH6Ue2+LFnSn41Ywcm/FprRgdgHEAcoQ2Q58ENZO/03vINx/yTXKzFaVSoPtSuvQ+lUsggjiZ7PaUyYJz0AaU41IvGT5/QwItHTwH9UjkgGOqLW882ydUTbWAO5oRvqRva901WXwzBD/AgK6ANK1V7ngqaOKgonxFStJbrYix6xfuvd8kUoT0myiYmLSfDROt65tu1dKoQwHFBCMlDHVZsw9fg0dGlFoAEmiNDRqOTVTbKp9GFK6sTzR4gjHbcBbWkaa5aQBgT2lswZsx2olP9QzjWnGIspgAWm0DAyh3XgHRyLu1qOVqYh5TQ4K1Ktq3g8HhQPyGUXUI9sK3Svivj4Q7k6M4I1ZSLs98sMVO1J6c8+QkYQ6TzUN6TwRe3sBJUJjpp6uaL2M5pmAlTfq/kZdxLTJt0HJbLBu8oUi2DjS6yvazavBHyQBhcSmqB8sF4OxKWTVCR9ngE09uGufCEMYN+uIit2ExoFMtMJrG6x11OgUXDA31b2NMm//v2+OU5ocl7H7GvMDyyqg5Xd7PHIsRX2n/RiKiGKWscx9cT7hopijpxLQBbNH5ZIy5ddhkdVd+OVFPn+YFhSjuHxcaQgl6pw8vidCFptbTXfsunc9XcytUAZq8UvxEumuxJNAmJhAJHYbdECnyvVPGbivF1jcYoy0CKvwT+l41mhFE5DWmp1/P6R2L9gXLbe2TwezZjAaDkCObCQ1D33e2KqsaK6nVPPk1bBfX2AIdu8Cf30wVm0oDD2ROK5m2U3zVobEagInmd3yL4xFFx5ddVp5CDzHbW1Y8+K3y/eQ96Jj0OmhF3PsNE5i/RrnMRurDbrOVdZ0K1/dB6dj8UUFPtUBu5kB+iBn5OQ38wQplJUT4o8A/0I0cQ1lM5ZJYXN8eJX+csElZpE84iMBUd50m0ts8GIh8Tc2vLbBNrWdDWhyaPLky+Wraj+paFyCSeubp6pFqbj6GvK2bc97eN73PjDdRJCme3RxkF/KfiedTiHLwKUjc5vYiiSep50nkPpjFSaV6VbuAZXkJXtFcodSE6OL9Up9jcEiBHSel6AmzjpqBEWauwbJlAKXgO8BxDbGfuETyqzDjVsgpi/rPT6eJyJ1szkId81OszuKv5kCDDoYJMUPDyrtX1iQgZegSpykWJigDVsHh46EFThotOE34G/++UCSVH3dfjYrdkin/6Z4mCQA+2/FqIUqyHveISfjXk6clf8SnaoSDe0kGP5DwgOYeHU4C/62LPxSZ58UpfPRNuz9kNjRDB4HYMnxbZZWqa9qT3o9+3j+RPPlozM/JlFtIvKpTzYhGFinb1UYPkFhNOl0bExa8AHz6DQfJhr4LfWj84RmdEAlEwqNWRb8oZBeu0wKs+kWRfbWZckl4m6WfxjHSJLQC+2T6JkykR3CLgHIzaXwkScSrnK+AV2flSpdZFBo8hWuc6Qpih5sOs9t1PhEHfSIq6InqC/XXhZ44rlbkXToJ3WSk1LlT/R0xmIoyQktkay7y1K08VdbAc3VRzJG3lC+d1VgVl5+zkmKE0ErtGlC/t31aHuZF89UFIxgTTXB9M6wAKBdFCBmSa8psWfsvYbq8u9cf4qh4zCxdWg9Ija2xS2IAAarhUR/N9PVzfl+FpYPR5V/bIyN5QHrp/Q3PpedaOOzhTOyB+/x39sRg93yxI38GvA3g+mp1lKBLcM8fZwfmNJUo4VqZ77R2/VONdRU6KR8K3dsjECPu+xMKWQhRoDMe3Wy0o7S2ZyQI/uHoBgaguwn/8qKecSoGz7Fn2fcq3/8SF3w7eYh9oc5j9GY7D1vshOigzpJ42xUa274siVVHCUDaRsbuHnd/gcEgQmW9dMO6NICt/q/1VnIP/WtUS6b6lILbgpsNz9FVUw8IgxYfAunnIkySP9n+acznHIKZUaLtcl+pqH7I3d3AAebU2Z5yuCIHDZoJZ1KLll34BhmdAaGph2SFDtgAc//7mQncKJC0OjCOmyhOroifWb4wHbcw3JmejCu99w3YYGzskgi0fJ17PO+9oLiB4nSSXPQl+xuretbwl4S7FGzqPdzrT3ZXR6z5QT1/sFgwbhNyLfp3y+bIoWZOjFtVSEBxCv0xif3nfRkajpnISEwfoqod7XukjmPl0jFZ88u0DS+spqRz9Gv6HEjeuaPtLHoxjPxmTBG4OH3UbKMJFJZepH/H05CLIN1wPPISnG4POscPirUgZIxn2zC97jTDhWd8BtqntKGUq/KOIpVNFCoazgRy260HWH9BtGCA1c360sVp1tI6h+4Rb31N8tZzFm9/1IIlA3fF7kXHyi/LXOadVcAp39MHYkza1O1IWrtXLxorMgLqugXvXLQP4zqX7BshpU7ciBgQJlssLLYu5GiqD3RILXaC2cdZLtd8glq6NIJdWOmid6xGdaeyJYai5PYlV5QgT67L6sPliViVwJTeqrJeEm2+mZRKHy+5LAqPjZXhYK5oBjnmbgOs0dwCQoCL/FRgff59voA1AkWMbNZcPVZvHWIMtASHgVNIY8/f+TkE5r6gYJHeb6bEisf4Rs4E+F4cvUPbPbK77F6hwaz838z52V3XWZfJgLG8ptBeZ4gtcMH/s9OIsmR6c1BsJiMRuoIuVECHYFFEF6dmQn+ylx28ijx07B4P8D19V9XOYsIZul1zcDoc5mMd5535kCLodonnnVzb5TdUyhl6eXciGf/0eddaRO7cQ03i3ZAKzqnu7bZ2oj+5sdJhUaVWtPrXIzWloz7Ht8uHxGRMlrEXu7eiiLl85tNqEiCNgXrUWMX3XNi4b2XoNha8RIAFn8bEkGc/87AX3PBsJIGvlHciRsA4j3ljhI1nZrPWzjJww+T6k0C+cHgtzaW33Zl2gLtXn2kt/GBFpIRSzVA4+z1cCQnKzatRFXhdEZ/EjW6QhFeDo3s9mgAxQN2iOg5SlnqPZdXzRRxUlfunmsDlt2dFebmOpVIo6bJMBUyNjvbhCE18Xv2HUcUyScQFRsXsg1BRB8PxjWJovvyO8XFcAVxMrG1Vj7ADR26J2VSOOE/Y8pP2TTP5ICoUlpiLJLSZ5xaeP+Z6PNKxXJY6WEDuIpIPoveYn/0itEbVpG3WQkW0WB9i3P9PCsf38mUlkNMVMlZNy6aTmiu53htsEE0Fz1xfU8sYSRgwGY+V7hWC9+ZsDzKNoqshbMt1Tf7poTDZFZuDaUFCnpsSQ6ZurJKcA9itHFYKUkd9pKJG8CQHLNUyZNz+E0s1pYdIwYli7a4gOnXFT7y42EbZKXvPUHIRm1i/sE6fGcVfdSfXZejALWSq3MPLQn6GGUPy0Lyo49SVuu8ZySj4+Um4nJVR1YjTWUhmcnIFLSYdAOwsqsSoBIpIr13x8Z8wK59AWKeaaTuN/8zM9FJvOfIjJfAiu54CfnKRIw/bAySNzlO/kXxRtO4F8r+9LNEEjKFEgket0XJ4GidY9k1gt5Jiv1mBeUrRP7HVKEPr1JC5HdHBicwAnC/D1dgwGE96LdlJ90APNQpXMLc/QMyANzcRU2ecMpeUmYmIwnmKOcirEWXiwl4/jL0SA0s5AQzs3rG/F+/imQSQnyYaD3ohQjXLZQ6+A5S2R9sjiJob3q6byylKNyD1tJaTqpL6S4ezCeuvilEH0btXN6nTATv7Mx796xkVBJFF5uM7Z+i0pR0Z9mWM2TZX33WOdeoC+baP/YdOq7747uY0QRmT2PgX28PjcCgQBNIXVTsDwZCB+IiQ4sOMntN5x6/Zk9jQXqP3RFns2/1/DUWjzvyxrzAEQsY1wLb6P33rVFZEFBjrgMo0ek4b47G1ByFPanAkmkbYCL1ME19xP9/+gcNdXIVwMDnm5cjf/Tkf21fDvn8ExmlhtPCg5PNBsj/2HqKKLbyUO2RRprS5QgaqG8E00lRT+s0ijB1JwQryoskWaloathTjjUYWL7zt3ef/vXwaxD+cZvSuCrZXIrDooWdwaB5AOgNKX5qbwnsdVyOlyLHheorru1rwrCdTkxLwnKB4f1nTzw+uHfl/VGGUWoN6x3dsmUmAgy9Flp3+hxc5iSBnuwh6kShXOVEqL0aUA9c9wODTxJ+yjwd40NNKlks5wZwTTS/xVfSInyLsLo4fcI9GM8+B2wtP3gjKnmic3KR3BH1BSD5yDOvfMCJdBf6NrAfLIG1V/X6e/MOmcz7Hh9FgCgIZxDEYLf7NeCv8q2vfbCEYrtFEpYaLd83x+QRU8qsA/NfXG/zmNDrgynxHtbmBSetkLRdObpuNcgPwENv/qbu7Cm+veDZE0qYh0n01//Y7eWEggHxj7WZ7SU3BhEeJpCFYrFj4ruQioag03URyV0xINMylBihu/JaWWxFAh0VI1OKlOFMBucIMe9Z8UsJVTSb4WLDFtDNP3lCOtSWGBudU6QRzLRLvT6jE00h2TBj9JV35XOzShvLUslAvlkW5xs1pE9yCVFF8OhiVY+XukULWO4aWMcaX2SGvzDhUx877SY1wi+PPusYD/e/C3bZPP5h1InwjsBu72p6aziM+jequxDkcdhyXFNjyBvPtUPmBx20zEB6bfgrQcLHRajAPWbKqb/GqZTPt1YeS1jzUgTcmT+Yvk7cuhr2Te4Lg+wW0Hn6WLW/KdMyIMBPQTLLqDLorJuOa4x2JVKKnrM4IeTYOrerM4sk71IO7BW86N53gSQp8F2NZ0tCS9SSxXMeCB+EXQ05Y1gP7hTu5SeAXtsTsDU8Pa+xP7TpX/vdoIzFX5K7zYOr8AjLx+f+Zm42Vc27LBQw88nsmfM+53nKQFjN8ApFil5ZpPcKnRceTNiRMeimxpCQkBK1F9xmRNQytu2/udR7YTlY5eacM7fIe0nD0/RPF7y+2KBbt8Jlj58XONVMB6JgglF/M5DmLsBz2QoRhJWVGNsm5xUW0UZiFqxPVIMqJYrY72na0iTz+UfmU6wUbbAWAsjBayuvOhqHWigzGYr6vwPU5HGRComhd9h/Lfxtg/WB9rzEuptMGFiDXGrRP/Lxo2aNyWp4b2HK2GWn4k4J6p2XiCILTATlj7BDKwT2H7SagrOYGQlRYlxixY1HT/ZpHcSh5zuB/rfUdfrKS4XCTkD3QPpi7+32r8flxpuDewcIZOAaSPvQnPExXIQnSoNw3esrbvbYXpL/fu40KVp89vP8yKGRVge+VZ1uNudx//Ag1N9EqPffcCR9bSU2VDHhv0hFQ6yDTFkpRX29LS0GzwtFjZ1c9C9/yFBOfkkhePuMIx610lG39xP0RwPrjlFpR007d7W3fjJORb0GsXPBa8qHAY5LoFu3PztktiFHqZ4WLaDLu+mbBesdZtV0a6SF6NqvqzqMXLMUWp4AOfs3VNs0TI4+tJn5GrK+NgiMIajsGx5Ics7uf8gAP+S6gXUX5Qw2goZy9mkWr38Sov/cPzPWbPAdxU3+GW/q9BabNMReCbWAXFDDDuMUn+sLo89HmJbrbLSNFPVsTNT6MXhlrZLi29cy2P3VAMW92Oz07/YAP7ol8LnE8osmNMTTnOHJyPMWLkLKsxBR31ad4kmphqaRaQ3PDD7x7PHq7AurH8Iirfj/sJ/b5j4DxXm+K/053plPpYh1boRFCyTl+ncRDJT/Ro9spvrqqtWdhu0CL+l1WDesNzPVRO2r6gSqzjcj/c7K51e+h/3veYQZNF05to3hgA3EVNCP2ko0nsMKOYsSqVegA3YdYeBlXqDCV2ihncQmBwII3kQsltjgtPuvB7vKu0ctzql0wSoS6H8GbKegPsrlpLEW2r6f4pEf3on1si0PrAY1+XnLZ129TO4m9rjKcecTtQ4+3bIrIcoILCpkFv2Q8njorWgL9DW+Gg5dY4g5emhnQ2E9bpBuc0ALAQtZnVmRq92bkiKCuwdqgO/sK9KUAkACLbN79HJNRcngy0CfQoQjStc4ptYMvwdZ9SovbXh608rkuTXWMQDFleFtPF96N6k5wwyuj4iV2MZvNv0Suo13tgRlEW5KnkR+LwM6yTdXTjdwO6BEnh9mFCnK7624KP/rV1rrs3rrO7IRbIavairTRDY4g4KpDWwYMUvEIvKdCZkvfZOQcAwdXlstb7FUbULqkRVDI8W5R35x9eT9DJRjphYWqjRMkQZjuAHFReaDLCk9g13rXoikCwNpKm7/a8zt9t2/oXaYt4sgQUc+Wj4ltUCTDXvLu1yaI51HaArHI42Pf2TsWVZXrea/JcBjLLersP6bqhbXaVwLj2Dc7UuuRv4tx/R+NvKwFL+ktRRZl6imHBy8cD3QM6IqvGZ0wZKRc+PyickrXCf5AmFH6W2pRbIGmUGVNAHYr5+DNErmbdgyvoM3TcoozZuIUz7uvAqdpwzM8dtRwVcZ8JyoN2Qv72QxzcZwmYLhEutWgsqWDra9cAX14EG9xOo1ojGHc5Z2aUgGE306B5IUAUp9e+f4jdPTgF/MS1x4U6WLeHH5gND0QVT1+f05o+fARmEe5iJ1++ECdRz2Rso7ntCNHn4yYTtKxbu0I1zc1JSKoHJFZxWwj33Pymo31S48MpGGVQz+wF88qMIIQp6zhOJ8p3NjJmDOwhPfI8pq9XfO3d4WiB9qxrA6mVxgWwI6NSvnDNld+LiSSI2NkCv/jYmKnzxWqkTIa/Ae1BUek/wCMgPks76qUQiImIc37D8IEj2UXcz3zM77N0VCTdy+6qM7XsN92NabTXrRT02fZ753cy7P7QZ56M2IwXxxZhwJeMPLanrAOi5YZL6RtrvzMLC4wnf6KYXERUBjEFOSf5ylVeOkRGkIgYtcXFnkFQ9/h3/YEIeaxkW41cn5Z0PBWET2R9BdFlZTHwDLfv2W71LDJddSPMA3DYMMUyICiw/eeAnroaG+xJp8uNamFrP0cNI1WJgDjDgUsucdsbspBm1oye9a2JilIhCxJGb+lGFF8uGvHqCjo5AZqgWlg1k4o7YnlwIDFUKCJhOGElT8sRSIElo2LLnhLNOhCtzkCskyrv8k3cpxYUGUBBl9UUzolrSkgJDsDU25X/o9y03zB0v5mmzlRDT0AQFWlWKEaQgC3ks02a9M6wovVjTVm0HAwvakyyARXYRI3nWCFLTP/wmaNZrL4tVA17mnmwXobWRq6ahfCo/v/wx77UCow4uPoXjo+bvkFXd6CmhLeoeYZpIMR08zjytoDizpKOb/17L5qqbRMvlV9Htf++4t2QBzId7RhgsiaEs9YsgQIfZXIQk1Fsn/4msMegNDaIn2iIBVq0YQ5fO/yqlM6F1XnOUU1wX1hf38kkkvrMXcwzM2W5aTV3vC862zh6s6/OfB+ZqnPFFRfJtWT4C/C19AT1Ksr8xxGpr17HH/q+/sJ1rkjJATwmVBMW3mnTrKW/puf/Os358rF940+3PlsnXVSxiIQ9vWRgmKfHw4dMDhvmNK14EmBC/ZIUGLccGULsgBnBIRgD3cMyFV71llcn+esBai2DhrMGEJPoqcumA/CR8SOLfhOnN7aE5oDr0gFLEk1a0twuOgIQJ5Tvtf6obMRW2wN+Ge2hDTR6/RSEpg1GNz8KDx6CGht1b9qB8NS4g/yFKdktF+wlKPjM6TiI9C08QOIhD8DFMrUzaIibR4FWNx4l0n0Qzv4gNFQiUIz7cdmCUE+QZSOugkyusX8dvSDc6M89+TwuZ74wF1J2cjVOp4HTCIK41SlsRiKfHa6MnP78CSYcssCjgXJr2rFgGpcTx9qJaLVlWTxY7mjCDdFiB+7Xu/5oZCD2wkSFaOvLWhy4Dk2Q2/AufFlaBwbA9YS7AAEdeFSvEmk1f9KcrF6zjym2M4IFDGs5RcSLRndcCThqToH+kJddydxKnQ7jX4B4qfI9q0di/N+MiBXo1WWpgun5S/snVXnJcoQUS/qDKER5+mYFT9Ig/+I9zYtV5ZtgmccDhcBdPyZ+73FtpCcT3e3/Fltzh5OFTeNuExFVzzhRiZy4MDcuT/kTiAwYoAAwSFQ3Wrp/pSZBJIOSOKUKq1RyrSU8rVZq2qBbD5UZG4xphanBSITq6EG49kspdC/YL+5xNhjr6Sge3+sIdNF9NTjjE7wDgdf7VYooH+kUxIyHSQLGILKEQKDQNN1JqJVoSNist2Q9XIAv7b4PHxNvWZh4lvXWxhNOyms5N7/UwM+QarC4ghGJ6+eFpvZbUCmarfmdeeWi4dmJ9CvkL49/oxalBUTi0uC7fwJBxPgbSNZZ7ge0vvZDLue08XNPg1GKjefCnvXpQFu/KSqxsOQ9FMTZ2XoEOB5w1S74i0HWUUe9SME5cyBU31z7/nbAhpqDQF0yeqDi10QwpyrW1S1cKgyZpMHifhZNNo4hNBe+7IGBmouUtRNKnBBgF2yXSdWN7mVNDxueMtHnGWVGSoi2UfPprRA9kMKr4kc5MdiwhsLMG77uL/AKlcQhMab2GCFHqVMK0zMiUevcgWfiNAvdcpg1Np041f9OiofxIKN5U49+iSHndK790EQIcQcAZaRDRyHJc9Ek3ehIMxV6S64gFHo6r2WQNPQIlpsmRfOpOlBzY8e03jedyfezAv71t/8bDX+WmhSttELiScBN7JZbttXGKJ/Afn4xcq/jW7wOco7+2FP8xIBrG5ooCUihKJdcvgk1DJ0Xuq6O7oH/PeyduD+AFSrpXhJYlQ41183S6TVAB+zSs7O4pNfFQwAMWXZzJAMZpzF6qRJF3R79SIGd70ytmFHoQGLM8YIMnwu7uETpgxJD32VSRIzBYO5vQaEw5K8fd0T7qG8Acmmc+Kk7gRB4i+r7HmUyRubTyR4wQKzFoYqSc2U1G53sTTg1Q2K3wnhtJXypaDIBmVSbZfxIefmpXbyH3l9CXQx+fy9cpQSOG6KSBqJp0QmKmBiwzipTjSZ6BWnbPotI0irEkVDhhR70G3g4Z3yI4UfJWTap7/Wwi7erMUWUcuAO2uKolJ/izHBv8EnZ/BSqNlBjQS6srP4W7U1rTXnkfg0r8UvWiizrv4/AOU6SzSSBEW2QZ3Vz0jNyHXBr8MzPKJc3igaHyx1re509kImgftF5Hnkn4Tg/F3ZZK+72vBPMEENCzmGtXvwFVJ0z9tkCIiF2D4Lh/qqBIMLwphvQh3v/vCfZy4V0FE4fdB2aGsLIfx3kGN/x+tzXJwxSGDWU0nad5UVKHB8iG0T5+fZlAEBVYL4CghhJB7UMDlDLGp+TXPK3/JCS1tjNhtE7OxfHFd1cL4pr2RwVvt2EBv3OCtxvEFK64v0dWWcE2lwCQ3HWNvVAcYQ7KIPXXTU4VEg68B3E9k9WsA7RXTcpagBR9iNhlAwc+kDa6HREJYyYhNtCGfai2W5ZsJ2BbWYcybVttV4uUaQh0thgMUyE/3wuselNTy8jibGRI3q9ovAZfM4WG49CbJAtcrG9dvKjiTW+SlGO3ZKM+gtx82bPg5616g0u7KgXDT4vM0iNTac8l3WbOTQXSFnk7prKsOQImFipdUz2cHNLo8bjweZjXHw5MhKY4Z7P16tNWcUdOdwz1yAqt8aDZ6X/lSiL0GfEion6E3L9NuAbWVohv/n/fE0ImAPTxnC09U+GmbJJ1T/G3T6h74zy6yF3n55cAmYZxWg3WbSyMOT6G1AeNLiVL5VHipRkz7EOctVglb8gPe+Jo5Wk/ddE75HAAGo5rzfr8hxKWOg0gbFBQ1erynZ7GZiT5SQJMNBg5y37IBdO7MTsJ/0eWcDTzmbwpaBWx0TED3ptflLt0aeL+b0dX8sRHzS4PoHGPfj2irO0//GS9Xj/qbPCzwTLKYuRngI/gsr1tRo95RqTKaF+SWH9SQWsB9cwsh5wemQubISVVQRj0EaR2rCrJd8JObYbLiiyZqf/xsBMy9EDw6zODP7XOv24IbaX4J4uBbWwDP+rh6I3t18GO7K3vN0KKNLBuoqRy4z31CXdwqhOO5BR0VMxwctQJHQIs
`pragma protect end_data_block
`pragma protect digest_block
7666c95bbe3cd690c0fcdcc9e3f89ce7a27a518ea5be20e25612ee7ecae864d6
`pragma protect end_digest_block
`pragma protect end_protected
