`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
bptz7bZ1keOh6rBAt3zKzR/JZ4Zw8sEECp8vYDlLe8zjR/KtUR07cvSQwVk+L/0UesF1ivfhXOgrKaeXbSA95tDWJlrxcV59DXGMjAfStUrEnyIwildyPvdxEhF9ybqoG6WW844j0U441rJrD2TkTTSvNUgosNT/rChMXId+cA9Edbwq5g8NSSXHUW0lOFXfzmUCQbdNV4EVOF8IcpTPAWp/0n48FLiLbedJQXbfOookisLjqG3Qx7jHGV/UjTNeorXM9tWFmEDaKMByKso38zSWFWhDLAtg+eLYrUJa8TWXSQ5WwzBxsR9SrtDTsmKb16iXDhnYaOcxYUtM7Sazpf21kw0ii1uimO0MQjseBzaJI9h7ikZb5P1M+2YNOcYHdtD6AoXNH9+kik0ToGj4kDERCUkzgplKehT2rL9JmGbBhUd8npBRSvdLWmHAbLo/rZUu/RZqIvAu0A4fIhKvccAjxd5OrxVZqK6GI3SfO4wuyvKvm4QozBWB8/6z8u4iFIPLaySVwvA6wTQShQ5TpQCg4oUcAXZ7RbDPIh/Rc+/W+9lttS6zSE+tcBHjc/97n5VRc2KUba4OSwaxyaslpMI964M7zC+GwGD+fqkrOaObarkTXdADgl1lqsghAUgkiz1jatyAi6eApxjgFefDFsm0PnGz6ea33MA2xtmAHQ9G1aDynVRd1t0QJDYu9UeOA1Toxtm/yhprz/NzFZha7qUXFxqOLUnX1QFggJhI/QjuNsd1zVpiH88WVaZ8w6YTl3yijJE5l7yyGRsB6kye7OCfvvpsCTRBZqOAzVXwwP58f5I3hqTretDeZSFOSKOCB1SFLkipyIilX+Crp44+b/OhmhPNuA4/MFzYsztJSHGGiG4oGJ2dgwMpOsTcGzAVOmucoDWYDvEcxmiyj8ViZCLgG36P2FIujrQ/ntB3bDJ/WIDrUVEL7COMyaX/1WPdFH72cVfyZ/hlyROvhxX8Sc/T69/tKraKxbNxhhpdmtxXEbyKKTF1WKYtawwGGU36OkTF8YY967dYhK+hK0pZ3fsaVnqWqWqW1g/QVitaaXhNwlodMXH78KnCRF0Ge3CD/jykuCin8aCLI1o5d+1mQL8UsHYyHxKIWHZ1YDBkecTBWr2gLVuTZcE+YE06PcJtx31LY9LFx3hG8/shYZHtt9rtv5k8I/EGSBX5tfuvY2cZDDdbM8WiUqQigyNQY8nWOlVmjfnxMWLWM72xjGFS1EuxIXdYIfHrrG0DAFd1lMXI5xJ560xoptMGNMzt4i+dEGfebao5SAEcAxZtN5KJxNLYTf3WAZX+AdEaknrnSpL7xnwQe1Rw6vGUddpYnLvTEzewdz+NuwMTNZx3EOb4t8WTyVVZCCYHXufgC10Zs4WI7L15V6Um22sFEeoqN4LJwquYxHYldgjwUAXBivjZ3PsVafh1JfbsnSBDkjecG28RgFCLnfaUuuz1j2cyGhlmKoQ6mRpS/DXQaqwLl4ESKKzQjNQMAZLhy1SpAfrTsoy6Cn+TYS8A5mCjYCz+aWv9QKgm3KAeJICjYhePvMSRCAz9Yvn7ttoAAd41qJblBB8t3IfrQ+mf66wo6mbsqNWfQbEbeoU+Y49XtskA8VkfrfnPfCnMJ4pHCTj+3Rdfl+1XWDdWAG1vy5XnsJTL+jrvasRW2zyePiv/D9S689SN9vwvfNg+dAIbjtVikTImJxZ4ZNIlQq2Yxsy6U8lT9Yf4XePi5IwzdU7lnLrlbp/IzHDJraZqGmlB18vwCaWmcOYfJtpqqHieVrv+TMZrhK51fOJo9VsvQvn4KITY9q30RQ==
`pragma protect end_data_block
`pragma protect digest_block
3484feeaadd6a2fc35dec22b15e2211af152d9144e881733bb3e7dee89f8e183
`pragma protect end_digest_block
`pragma protect end_protected
