`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
MFKWUdUiuEhM5gZpge4mouxzTZTFtRmc7k8WtecM7+cLI3o1UJn092OFgydL5HqsmSqGeADkpHYQKQs+KZfq3qg3ywcf59F3U0Q02kBGZ+5uSQUF2qy9a5fm69WlTC48E8rQTuI7E8hAgPDQlcd+7Yo7IwDT4lTB+rLLuUDjoAYyBJMebILKtGcIGGXiNJHs8eoJR73LWXMuTocyZ6xVcr638ja+Z4NF+53jMVXFP0jhRxJusAv64mXqnVJI+5VmomAO3AHyEzU1rvQy4d4BsXSWtZHCbac4GhPZS8BprhVswQg+lbUedB/gasFL+wJtaOVyk5mUdCzzVYMmZX7sKjHPMx2gngUU5ZS3bm/1IK/StTpGjfO01FtBVylZ04AznFILbyqubiBhs6+PG+6j+2MZG/rH4CHSv3+lg70jRXCAHvltzhTW6LRfXsoZVhLpjTAYtgLXtI7NBkmpxA4IXLK4PUnfv1YKYSrW8pT9MXNgolDlHOTbbP8HGrSkONDykjULiY0obl+cuAm8Y8k62be6HcKJXjWzUF+sOlV+1dxpsDw6ppN1pcersRWQWgvOYN+uF2W8lUw1pMstQW/PGtyIlcCWAviofhzetxOf4ymREYT8TQrEluaseY4KNapHLKtCqPiv9y4McRiFK2hxWZ8Hu9sQbvS+JZ3QaqxgUEGhXNuprGrvniQOaPQzLsqWFaeNq2MFnf4pD0qHyljxEeQk6y03e+Z5ybK3MphTpi5KYtFX1h6a14cJkqprv1lQbILIlu25L3zS3Io1vUGoMkbas2RRIIT53Et9JM+RCyrt+n9oxfay7QJl9kedEI4861kMEOTT6NUo/lDx7O6dk05n4aTM/YB0sk1kPco9soqLufxoUR6zfsSSje1xWnyRkLM+ZPTomNW2ResxaNx6vQdPCt/b0rXXRlHqqirqAmDrT42fCWVGEEhipARkWPa+AQJI16KrYgyNdV/pkOhK59NQuc+NeAgIEvDtNnccYDaMH0Yrvwbzq4dNppMu8A6mqKNLo6qSIesvvMW2/eGj9ectlCc1ZEvJ26aqC9p9NFMZ5okT/n/By064UI61sdMSocgFJBpKhuoLZ2zu7ZOeWFotm/D7d2zCuS4JTnWA8QUQggHocLskIb/nvnRzvyM1mFcEWIjAHL7AGzCKbKwI9kqbbLKUg8W72BIBGh2NVSJ/I7nsA3CRyft4lsAqzJc2mIXCr0wbpbRdmwF+ZLbJL79fUAp/Xk4KVvznYreWxja0f8PXFp2LptaSQV0ji2nM9dFeaDZGs3RWESoBh0qH8UvUyAWfraU5SdYDgjrwaD7hQ4C9NZiuYdoMY5C0XKvoJodz/BOUPNovhfQPUR4AiuVkVecoS8ASGuf/PuXRgsrfhGZGQq5+bO33sTtcAAqzEb2tkQBCQ5VWWlof1gRn/xKg/NWZLySuaLw7TK/4odI8VWyZ61YLYpjav6RoSNjH+NHdOkJxH/0y6MPROtP73X0OHI92hSONASbU55zBTmbZOzenOhl5oLD8lRa3ykuIPoriTmCrz/h0sVK1JAUyhnhYrGqktsLxWD5Afp72M2yliNMJRCDrWqLGtEIb6wyiUrNRYC4U9LJvFzGSMrzHbzYU7ydmyBCttFMZJvBf+13Kk+BbGD1JG2lY5X3j6MR7gG2URfgwYD1SXURGzdgugubqWseDNvEqe/gNiqhUrcHWX4/owf3sRCcsuOhGGPyVQyqKkyhTcXbZEPNCnHQbpRo8V0d8o3JRd4P7IwZ/KurvjMaDusKpYyLuLjA0ka4FR8sLAbv+ylSQ8IZNHH0dflWt7K/TFMcVU/ijLmAQkA/6QG7R7gTtpqGP0uNA3LIa/bexn5u7+AZTjgvPYJF+hXsU/blQCK+7FRRz2fju3mTUYBmr1qoUjJrF/qhjxbPgO+LK8YF0NSKhv3N7mQI/K0IUSsDE9I9fMAsDU0jCnij1ba9uD0JgNVSdb5ISupKYZWSps65uF+yh7tMT2rt3WakffVRvGxxEUZque2ZLyV2s4frSlBLjtpEVtVUPO7yfp953d2QTMjFrsrAmjBjTuBJpYkg1K+qh5wz73o/fBQuOauXDetm4NZAT9iSPFO2/eHPpN+vr9obhp2t6149rE5AtY1FzXqaqb7MJvzNvrjECBV9Xpf7vm3Uxom0XiInaoCaeG7pLuED1Lm4gZJZI2xT4OUW6Q/cVyK0jxeCI4rdlcxh88rTkoB2wT7vlMdxToOBJ0QnxeUelAVIe1APD5rdnnNaSqOg9k0G0Jsz1nmsRf6bWracfscXidnerTsJOVq3MJNvI1K7l9G8UtOAGLSiK47QoaTuhoXx4SdSPZW+amz9Pa8Vl1p2CE3SmQHCUHfSoVSOx27aIIZztBkp2gOamdGvhOccY4vIFonpF6hYzSXiwtqPIgUCvgvvroXMUMf5KN6WAK4+iCqBLCi73GAhNnDoSuXHDC2Yft0VFXyj+D8sb1LjWIvQFsriRqByQdopYImkWRUI2uZU6cltgOO2WXuzILEXtcsW53hVV47WvcE05JtOukgfLl47cDzccVmKBJEm5nK00M+bVVCxbY3ExeHasg5JWqbrde1KwhsFyG01+4sfxFrxWXWmaP2GZAhvIF1emfG1R6IvekQz3sS1GtcMlGJfYbc4JsRwc52pnhVlH2AbUm4SpPi6s3s5L+vuAR8UI7ogNF1irh0F193x2frdOm13k9GcooU2FAMfG7vpnG0wxdwhATwL/uuLrFNAGP6OI09JPtgTzA0cafwxcFk8BV3OrOH2gIuv1enmUh7FsYtd1SvZr/kTzxAE/DqR4X6GrIW9784BXbmR6R8ZdjkL84ih1ZmeuFYbgrkX162zeARfJXkCB5+wImsZLYduYah1TAk9dTtJ/osV6W/zrnuivKh789g2N+ER6j7BaqDBFgQvqPIVuBoKdG7KqArxXgD78roUDY/3vr1mImSm+XQ+6a8kW95WbNJTPdxmvU95a5qSNmUeOtuo2RfFQkCeVlPdLDJTHtvOetE2g8cTuDIQH0HDP6A8p/ksWkqKppkOZzyyftRzaeF0zLJ+DFe6l+IPx3i6iPyQ8kvXnlEUNk+lUItTUuBeeBuFAAdhfafZYImkFafxJKvMrWNelVeKHPRtHg4X2fh74IE7iJzgmGzccDQuvQA2ZgZ1Flb8WJqpT6rHkgZbvnfceGLur5r7ix0KCs28M6qq7gIuiAfDD/1C+9HYpR8bRnIZid0tzqsiJrbd+B+9ZPcyrri/5kxumWAOpu8vqSWeSl1czk9M4ERQawhzjsl79+TeiI/28Z0GzuGVF3HBcg82rr2ijBk5KDEoFV53CFq13JW5Oq65rE9ZlojZ3z9QtQEwY/pLBpj/GJCh9aMkbdAjI4hsJyB08gBs72GvMt63d0OYFCfEgv6yPXjf9fKRxG+Xg+TAs4ZfiD1hb7MCKkuvUsO4VfuZOzSJK6rRYRdIjln+tSdaUXAHPFkn19JWHdZCnHr+FosoczZyaxVhaHoLJwHPopoDtZ2bjJGtNC+lgYWBVLqtAVHxx3IOuQyEHmG+fgqJN7l8SF6ZXvb5t4TVvEXQEkKV0gWn2vP1EJnBlshLBJVXwjdFrXP7Ap2SE0qoDI/NNuVfYcyQn6Mxe1YWSbzzX2dcjQH0NwA8K5lRRm4jLnt8SAE5JmHqX/SBMR6t4S+WWuIIrSV7y7CxkxE3ZF6gKaSlw7pnfqOHY2jnx5ctqMT0aPC4Oy69Yd9ah9Pwiv7qN5G+HdeQVpN5TrzV/W6Z06WJ6ItIM95A4mWQMKvLFwY2jqNDuD8nmLRq4vM/q/GAEq+lfCDjYkdQbygvCOU33d/dKZDvObkTVEHONUYRuSzD6Qa7lk0OMfy9AjZ1y+irDoj8V8X0bK1M/pXlJwyLQV2VT+NaqpCZwTvSXvqRUiq1HDej3wAKm7oRrA+Ope7XOCupYnd22p7YtG/bS0HvHeeVmUe4BtKnpdnD/1YteTPxMnbBHE7/f5oa3Ber2UhDVyk6zoQ/6f89+BarGkFnJgLJcscrFdMNcJFYHhGMn1Cxb7HZu73nhzRvrARo3cK8P8treRINlTZPlbmAH8vVBwt9kJU3hBmavyw69YJWgPZCrsujFyp0/9A53E0RHZA2JVPebw2kDkfrD7//DrETX/7siu+QI3ksmigGJhSCxIrXB1DFfI7ZLmHbBGMRtiJTHlieKmyW/+nusgXZ5L7TAcIh6+V85Q9f0QqTDP3F9og2On8PVjpYZvR4HcDrMeImDgQJqALqfeHuKEyCZr8N6ArqZ0LZ4kAYt8JDt4XshE427FPQsVlByKfXNDhKcTrGIbPgcuJo9ThNxVWkgE8C1yRVa9ybo8bwUEcQagcPD695zLt/EdzfU28BAFe7SXEJRcY7M+cHHUHGdxtNnsw3nxDUUKXSPrdjXGgstM4AIoZzdsxDUylxGEfX3EtRYdC17VsnGjAcRo2SOvqfvLcWgHBog3HcheKFbfcvkQ+DbokcXzXNE1Ae3ja4UWQJKaPY7Oz4b2L6QMm1RkEZacBFSCBbzGBx4CvIIuMDeWEplMFZWvVJ6IKGGZ+C3Oo1vTnG6kLABYlgmPu1RYCY2qpbb2b2Z9FVA/TBrF8+9Gf6T37vDrVrmL/vOn6pDLR3JJ0n/iyMe84BqMMyM00dwobKyxPnsOhp1dVJbx7lV+fsthVtGSgS5SiHVYwIRQT3LaftZxvioeJ9mA15X8B+4A+FyVXCy/W7bkITI/fx5nVtUv9ENmF19IpYJcpESvHMkA9XBUhfE+3zCewfNrL1sEAPUReffzbBpGR8rOvj0sYcJkYpzJhN5WoRvh+QflIg8BCOZ0DqyuS0YUmxKyaP30ZeOA78WbfMqxBd7pp59DXkulGGeYpGLbymb3KaIvigU8CW1JHARkB5FiuliY8uHsmMnAZ4phVsoi89aDmJGCSE2h8ec18/cRpPvx2lSE/MLA8E1l8i1uyk+C/npkWfevIcdG54G1qGH/lYjJu+f29EL2/Un/qxPHt59atpJ+NP68Hl8QY9pSEGoE/IipZ7qTYfA9f0e0AZE8UxQjP8HJQtBgnLxXHlq7tgkvl8b5lnREAQoK+9Pz48dUaPay8sb6dVM90Uo1FGsZADdG9raZMzs/sRdfBROwX2lXe6VpMTJ6XwvGOv+3JG90OtZHZfn4HOUfRd1vkTc94PDbb2/kZV4GIDyksVqgwaj8GJj+YuI34HW5Ic6n6PNHGT9fBr8DKpzSlz5sNVohlgtCTMqB3AfGAV+6B3kcYK+3tuFl0+YY6B5khdGSPPAVWA80pPtudw1gZ2EZb/FgrXL3MbwWwA3vDN+D1h+Is8yuYZT/n8fgoiVoFDv0tIVHu5JoLClojYds3ielf6Samyq5e99+GX/NWtieopvJDWAQMIpqBMuGFPG/thU9ooQgs5j8tvZNeD7szsmjvPCLHBMBfIqqzTsjlWEbLjr6y9+q78i/vqFI8YqPiPKhyKX42np9A9+n06fAQGZIfrubREET1blRiJ0XEliSXm2kzVVsSMwYi1RP5TL4b1Hx3VoJlxfsRFHu3tHITNavbFzUp5amyHf7c/urSi0vdCjnQ+wHaYlP23T1+pwxeTj3ARrD1nxmE4gvdmuAPclcX38VkRPh3iuxIQVChAwTORKUhscluvYg/M1sMqSj1rG9Ks9ZmBHjcSUbznX1d3DtWxPqWt7DxIPlSLIkZtKerrQlJ6mP4QrbVSyhXCBpBFkuzLUA47qTltBbcbDsIRAxmVEe2nlNAT88YlhAw7KY6DoxWP2AyG+D8jBZWCyiZhgdXTObiLjY2zTYRzZ/t+D1i+yg8+0lgUxkS8HRudS5WCplh5y3jOQiNffHBmnlzbsoy8+6cxpfOYy3L6p/2MYGE6JG2esIs7VTL9tX5sP9vs5h2BKUdk2IExweWW+IZNPWrD1FrUM4mBkP5cg19EXNnpmi5RdA9m1rGp9BL+pSQ3NbqaWMFu0q+wbegdJESWmFDwfQtP/jQxo7VTmeykwuN5JGLhshrjQ8oWnrwG5qHQZzqGHsRqzrnGGxl0XsyRghBdVT+jl8a0ow7E0YYIlMCv1AqfSxWhLDAXvo8ODJQzyA9OBt3tctUDZbXB/SexJYpidWSIVmrXfl0VFYxJtBF3opthvCZ1ghYQrf3ntCrJ6C/y26oqKe/pcQHWsbdCcz8uDjKM7NhnDGCJHeIq4aur5fIEifbwi5Os06sTs25Q1Y8Iar2PcusvDZXdjHkFy+G+QeK5uHo64k1FMU2eU5rhdEs++LLcaNWOEXtfe7ep1bUKWXmRA77yqfvOJTB5zhxyBQpwCyvW7mmNH4vScwTM4qlCDgKuZduvhR04qXVrQUhVwLtFHG8enD8rkCjTIw0eJNclC2eIgUOeswkUeGzA4pVX3pDWuyzGkrT8AyS+NaenaDuYG75rS7No9+6DqPpNGPPVIqJAblmYXWZETyQJV+Ta81KnpKMirNnf4mNSQqQS/VOQO+B1VRzp6thN7Mf+p7f8U8Xr60OmOiWlRJh2+tIw67L5Cg9jnAamklfYHuZfAaPW6SgQF5gDR3LSLpi5JYjhVWNNBCPbiI80ToC37aKyVUiCSImFwqfOiy3uQua8H9wi88GUBUgYVoNsQz0wPQ3ZgEmZHVrvpeIlPFV5EK7LYsOAFzWHdHl5ue0+S/Eu/JYzDrsBu0tQQlj5PNHfI0qae2t2L05zkJXMwmzSzFOdaiUFVXrMCqTWUD0CYAE/l/iD14Oj5mOExZTUi4IqvzeJPx4EmHP0QUZNP9cdelPBcTxHso7pFpkuqT9NeD557wkpZeVWaX0CavLoqN792rNpv3MzzujJo0sX7rjLOgjYWmzyA6T9Ksar6v8QEx3EwFvUDJWNL/E4IkGhhO7tj195WbdfC97YClmqNbTocVv0Pg9vv/e+Q5TLHJPW4/OTruxgq/OjiiT7A8J5TVCdM+7fsj1o1OXsIF4ZYHdwQObEWpAC9a6hmORrG4kqwNzFTo4A42vqmrVcoBa7AIkhShGtMetEn5TYuA1ibXuMAWw+JW4/Va1fTgsiXSG3RAC6q6CuaCIK8SiZgYJb37e7kJZkE/MW1t+g4rSLQNC0m9tchYTcL7V04/fC07gOjGLYQimGL3PfbYoPGvyT+6jgXaynF43wAoPfcbTMm7Nz2+pxzIMbOlVQMP/42iJPHvmX/6jO1IieshnI36dDJ8pXxtWltxQTegsePBRqTSFzpPUy/xws2rmQMIsf5Ra5Lsz+SoDwJqk1ttCwoOavKNyg7m3Zr03OKShIOJaRbAhmhElJTioDOmaPW1MmOSF7tWe0LBdMxrYB2DafkqrlPk4EuyUmdIQ6M03jLOKhXlNKBFH7yGQPHLICrPEaPukLGsToDh0GywyQ3bnGjhSC5mU3aaWIbAW9vJKHPNn57m1w048RRoj/L2te5OsJXn/dhE1xo/Id2gPeq2bnhtZo12/2kGf6vuezkqw7tktKfudTNqcrZcH4DrBrwIMZSzBNTJCqoxNAHDSUX34f3PTXH9fPMjHP2s87c59en84ZDtL2guxxT/hWciGzhTVRNACPaR9x7wo7LjtUrX8egTQIQ7j8Opy3LZN11Uqfu3XsDW3Eju+q7r60PB8ghmTqQrn1Nic0yd+L6zMNYrq+dtGRLZ6IItSPpbPFlHlrbGy7QS9peBYhU4Y6Z255fjKhdS2Fgf1QS+Uib4ViR8P+opIkVuIGiFI/kiHGTiDGRxXQ2XifDyM5mcdfGXncJBJrf2duof65X2MzuVWRJQw8YYWrtSFJED9Hq/jSVyXHKxWhGwwWFSg7pUnxQciddPLGmSqy9I/TD8W6WzoHo/oxDn0+E3JnsJr2d8GhbGPK17bLbX6aNGOLtE6RrguCnrENUSZX1meurLU9hCJ16QFm5cKMF62V3xG4pW/uHYbb9Y7VKL/xn0OWldCjGDRlD7WWAf0ZKJHjteFEdgsNYK108XVE5AcVocxb61RPHFHtsPf/Cc5enJjzJp0rKz2WOQ4DUqkVpYfxMqamqXCE+ccD/YJSmpPg3CKeFWFFm+Qvl6Ro+G9d/K6LcIQTqvITNrw5twKNiL/5zMWXSdz23YYiw/J93ISYDMAnZqXzHFz/nkkQmNnzvUPeGR6mOhpF9Nc18a92Bloru5Oopw3CyiDyAfPoVp6iVWIpUzNo/XEbOI+IgequkByhuLCygnvzupcjYdQweHZr52zl7UyDs578A2zEyRh1rvicvyfZ/fTPtxf/+eGdoefEuR2V+6WSMETQCSgpW7UpVqAszJw/m0dBaD+jJwpqeLllkqQ5ybe4ZunNWAkADnS8Rrm/jYz+ZbGGofHOIl8oe/bGPmXI21QH6CFolXb7W+5u54r/fi1R7d39MRsSpwWu+x80gq63OE2XcdoBhxJOr1lFFK+TxaEIHcVtY7HBZDSiLeE9tZisAUQawQAvIELxxeNycXotvw5Way7+mzi0mQzN9JP60ZthPPk3LU3mChJQLpeMaGbdk49wp0WB4PS446j+V4gkrM/wx2j0fMv/zPtgcdWs9VzccfxUSlT5jTd5fVWIrhKA5Z8FhzuEa7iDO241TAC6kMegFeD4Oox8LZ1Vcp3QeoStKa60W/UyxKQa+k134ww6/JVupmatmC2jMjKyPd136d43DwF5uJuw6u/lPgmeVBGDcpaWkq1XOqbviU591QPuweruPmx75Ly5QSWtwAAbYjuJsbog7iFUQB6k15bH4NZtbXrvNYXCVILh4hIowG0/0KSgAgLI/mUViz8r0EMr5bXLi6dFs+OiEwh8JEfACe7abDjIxtnkZovQsmVxEeP1JO/h7SinW3IFnIkec1lAzdMq/CbTFKRxZgLRxCE+uFahnuljpz2c9Bz/bSVPTq7TOvwP+rnkOn/OME93nOzFvqGyDEl2JpY76693gLEt+Q8ybxYlB680Yv38hL+j5mC8o9wWDXIy+Tj6rhu9PR9QK7TPHwVn+VAefKd9RP2mcxhdtoXGS9UMc6JpVi5n4B0B0I2zlw7bnM1sTUp0WczS9DW1qykkaBdvMrpZD2D/TsblmL9w06aHQi+SXgPcFHdh+Ko2XdGcWxEbmcj7A8dpogj/CBZabSMj7AUfVNYFfa/oJPLTZSpcu38QGy3pIZkDt5SyDbZLacRCqYnoaiuY/RChKITw71R9xm6VJeOTWjVN6W1wzDFl+mgwsm9ivRxAT3nCItYMq5/gb8Umgp8JvT5JFpNEktoPayWhtSN4RQIZ+pFWWfm2+fHo8RWap5FkqUMzzhfaBXDnS/YyIgzHtYzGMvNojzYFzE0SCH7wPRFMQ4Qz2+hIZqSXIZHZHCJZ/ZgBcM/HQ9hbJKxOhEVJhPH6+IEfdPu2eraP04RsrSLZpSaJWwOCl7turoVbxl8r4urD/7v07oG0C8OyjUokHnr3jLEGnGLDUbehirNMJjcbZ/pmgwzg/1zKcK3x9S29XNq/01OGaQKpE2Yqm72WJbNRJx0/167SkemGJV3s1EoHAUbkOKmvUjdE36ofAlKxePWpufV8SwFAMLPPxe6+RF8koMtvqrTNECpOXhLSx7wrrtW+ALHOqrdv/AIAKjVfW5q1ss4WOEi/X4zfwX6cXJnyJz+M3/UKSxvOmqfMW2SJuvLBm3Q+cumlIAtHG6EXKUpKzU0f03GNKNUbi4SdWc4A87n7snlklUjJddEeC10j7eniRKDFeufF7nHWbgPDOhlM6jlCds5RzaDSDTrBV/AToAfdriE0OB40j+j7s1if4UUIMJrgF3lsHmydJDbqyTF/VNAFPsPe6AnOKuqlgCg8Bmeej6NkXdQVNMYIcXtJpyEWWLMYz+Z9nUJu+vueTx5YmDTrb2GxTPQHHBvobGHe42eNcC+mvMaLn7fUDpweeENM82cp8x3T4/bCGIDsu2GatlhHaojxOJntrKMfbyOQ0vhsvrmpC1v67olji9aJta2CMYzCz2AH0d2dFxPJRFRILLuOuVcJ7UgxQ1BnxoxqFYPL5bHgrKuK1EzXnIWjC+2eT4PH6+UGDnhLb1GNBH6awttuDmlATQk89r6M4cjFyBglNfpODPuklG2cpePvkIXB9TekwTxuyR1a3t+9XM8UAm2aesU3bxJQQZoP3ARwGmsmjBfOQu6k+AY8h2kJHea3fqXZsZtewkQ4TUb6eMZm1t3Si9oBW1i6uIFvaEHvzhFXAY5WamKQf1VY5FL54jRUJ6j1W5xzbo/yOnq+F3SaXVC663iPQYKtz3DVNHtQCCxiBiaCLKbmVX7z+RH3/ksg6o4FZMIdUwPccv/5F+kKsKbCQ37Wa5I7PScKRylvVQK4Qx9e2hohTFSU/jZSx15rWmhoqe7IuNeX0idMXwMPGPbw5Ip8LLA0R/aFhkw6dgd/yG8YZkyQgB3gz0OAvom4ZNjkoizuTiyYtz/jCqiErQ2J1fdcde+lh6OkEEPflnYG9tJzOZvqFe2wLsidN44nJPyWohYYX4nSDnf+2HdgCNoRsStUjxXQ5kIFCB6MiohVaqSNEOaAFxddY/MNhivWtcEL+grpAyK83tMR+PjdNBQzfc+o/d16czjeUF4rXjL6GTzpNTHYoPmxWwI6Ygu7jgQYjqFGfNyBmy9K2k30k3HHlNAVQEkmZBi2QCPjHD9w+0eI7n9CwBuGQTE3MXOnhM3tczk2Lm6xu3FJGz92PYwkcqlS4ZcJYPXTrZHsbgmPGgFAZ1T9IXrO1fVpp5GRu9rID7WXQgpLZhr0PvVBV+E25jrovMT9KNRhzqMPBuOil5xkDIE5WFUv6cWvRsTZWnITPj+ylGwpGOyTGIzuXUu7j1AQz5w7zAxW1GUEjaoNG+B508fPn9gySDuq/DU3Y66pMLTcJ+9vUr0lQpKSF5p2g/2AzbHhbcIaqYHdVpP8Mm0vbut2QeymkmjP4QaExZMno/Dzcy/RgpQmLXMWYk5ukN/TxfqdTQ3kZdZPs+zARH3g1xOa6mETWc4seQIycwmXXyTtdBQmH7c/OVkGB+En8wUcaXxpQKSFUJAhp2SRMLnewxEBpTkTjhCP6KgggqFSaD5u1mseFxNxKnQ9Iu82w/1hd7rNTsgLoqYbPxVeBzNj6iAR350dJcGCrZmq2FYMp90cXVtzQNxEJE6XU/HjF2pesJxzVi1xQA8TqSUnZJ42J2JxI5uTFvWjowg30jZTGxq9fFZZAXEds/uYen4D4zaVhAu/NVg1L3C4hUccszkf+CclXflUCZmRB51MCYTswFPE9PxIGuLcxMJ3lsILhhHE/XbGu5cmwRPvY3SBdm1TX2U9UnED1ITyd6szBNUzJPx6ZMTI8RbkpTrBSb8ePVeDJ7K9wv13mbjoz5QBiN//AKZI2b5Sl0NsXNHLBIYSGD1udnC1lEIALpbiofzubJb2Cx/gfuSfqA72954dzHKtPcGZFz6TxJO1ucaE/b1Z9Hjif/acjoPTgaDsMT/xIw4ZhXoi0h+NSJg5ZGNnugk+nmspq0vJK/wqbks/xirpamoqzwzln5KqmWnFOXllN68MiGiFqSilPmDIhoBigzHChgq6jmI4KkmXW/dncWe45c8TPkZAPbAe1czkMQyD8wxkEUum9ntYfv5lP6+/eeczuGfDN4vXCUEP6Unq9zEf1K1LFYuW7eOP+UdVqZwtXT1M+aBIt5fc6tTslvdsqtLQ9Qqdt8zktxAY3mQGt+UpWP6tE0dZB62tintJSzSDD1n6Owr6jlhpFOcswjo9MetwkOWesCGMF6zy0c/rh7PgU+alNyBt7t8X8jaMezP738K3A9Zdo4liLjspaxg3JOkthGVy1WpLcRPvoNWsPjG3PZPJJnLhy7VO0lm0HKni+L/Nsj8OU6KnJx27oUO5F9Jpk6tQ2MZpLXDwbH4ZYz1nvBaAVky/eRFvYZAaX3dqQ8ijQFUtmDppBx5HKG09jcL2nW3r/CJluW7S4BzH6J6mwo13UevN/BR10AMsXCjXEep4PrvFOA/B0HvkLixu802XDEt2uWqCE+yPh97wk1ZUAHGLIVSoChaY+o9+yN/qOOfixASnBhJYjQLPTLA9JIzE0bTBPzSHGBCxuD1XTy+Gw5MIiJ+NUd/q6hBzqoDZFpoNojp9J9KI1o1cjfdv1mawABjGHpbIx4oYMzffEmL8rEUuclFxioAPG7LWxw5jrVewFn1+IVAqpB4fyJ1Wg+yabNo2rU+gAtZfHiP+KK+tYYfkBTxYQuJBPDZEpZ6TnwCO0C3GPq4hiCVAcIeYt5vhoLonn4tjf7P8+myUhVLy8TtIgSIzVLrptYp8dHF3I+e6+g8ewCWNGmL8p0tEZeJzZ++P6sz27XJiSv94x+/NkxsL72cn5N+iq+bdu6XYR7el8rI3BM9ZO2L9DAvft9yLmKG3bVrSizOWcwjkPuV9o98upOfay1SlrIo+Xv+SOCwpChrN7PyK7PwPQXakabrdwgu4TAaWPjU6c1Sa2AqB+Sal7XEEPLLAYAit8NrNbNOAOY6FE26t8mZprFsyMiRs1XZJMIa/8p9oglXYe0dYnhdzVPWkWNYsgKCkSg/S/EImjXhmAT4NPpbniuWC8GES3nL5vDOd5O9LEA3S3gf6oVrg+RRJlKRr+mt6amSWqbRFkKChfaVjzcYZDjxuwjGeflneCrp4v7622qt11fA5L3rXMsAEsGJl1ufgn3gnApSdlLKsMn4N98xD3zmOAGyV9d69Ur3VGx8m47Gy4Gr8WlXju7zrWh2Y+eQ8s/FDrQs0Wc8pN1qxneFhFZJwAPT9KwIV3soiXrahtpGs8ZUdaQ7ILyBrwcFpGWzvqIlg5L1Pk5m5TTAKtaI5BOTI8CsAz0gU9IHQdgqMY41E1yxRa6i5CzUxMzSgtcuW12G/ZR4thyl1RJcsZu9choVVIjD55OWtyIfpXzHQSpzITVDyhY/UVP8E3HrQarsZpOiCHhBxMriV6ZrN8b1kl8ua/fFHd14bJ3ckExN6qxcFs+2FGN1YcYpDSD8rJcKwXgZS0TIwFho8oKqopq4Lo8LzOdcikd6YjM5BjpRDFP6NS1l2vM2B9j7vWunYRP2fWR+18OPniDPTBO5uBVzVe7kEh0qZWYcliekSoJfSaZ1tyuVv3NNN3V4kqoIyDGye3kAf3pC++a9TohwgaGpaFYgjD8pO6xM0el4X0J6zxYOfS8T8OGSwzCcfph5t+p7XpLfxOgbfHceAnwVHYrpJFQg1WWwUq5WYech2w0gzFQrEpGaA1qbRo2Fy55GwM//B3cOdSggepNoOZxJo5FsH0Va2XhOc50eYR6O7IILfClpb6SpxqV1hKzhW6mYrSCFVtvRybld1RF2MY73XBMy0JHUhA41Hl8UpImHDXwS8IVEYZjvTvSz9mUQqSeoynIwdW9FziI42hA2UPpGz3JAQt12pKlHRSVLlDd3rfcOV2iJv6IOUPVO6CP8VhQsg3aTG64nUXWlJ/cflRDjVR+uiZugj4deID2XGsjBPDc0cVU04wo4owcrPGYvq3vSVG+1yajQyS3VwaDP6XCQ6f1BeJ9Uo8NlGkeChqQ906zwir3X+oB2ICuY5YGu9a7HDir8ODi6eGSHuA3CkYlD3p24YLlz/FW+BC1AWqcNKQmMdyaXH9tyPO8ynvZWRMuJHloSxXCeatlUwbGPn0hYCq+0AOdVAs62HwTfItV0esB4xjUqFyTdfUSxWMKPlDhLt91HriPv7mqxpoItCvmHuU9DDx4xCwCHTjlIE6exe0x2hPIfhaD4DDbV587fBGgu8OGbLtmR+KmvEMFEaTUp3or4Vk9WEZJIFBYU8uqlx8sgBM2+R175RxBlW4QaYRPIjbtLDXxY28ansmZZWelfGFENq6V3/wM6dLNkOxy7nJ26i3vQ0WJmozbYKJhiunH+tisjkk76JdWXwyGLbomNNSJ76x1tPoyev1Sp7YREgSJQvSyKODgJ7BgmI55rO9tMyk8gTAEeaD+ca3wJxsT5fcsUIXW5jJD0FtIwp9YmPivI29eJXaM1Oku8YPR0+PkmN+1pOEvCUgjyU5napapDJ7UmHw9n2iQ2ilvqHgyvZcHJ2fm0LRNNE2BjmkuptrAnhJcED0pkeJPbCcQIK4mx4q8lTpp4Nw72LnSzUs664obOcYunbrmh61xoay4ahLg+b4hW2aAgbZKf1ilZ+L9tgJT9xbLcYjr2Vd+96fA8gk5wJoGGYKp1IfmApBVrWc4YdKw58GNFxVo94Pzr1h0LuK1ap8xVl8b3NV83kpaWJY9QOe2VuVK5wZY+3PTx6S69I5wh7JupUlCltpBBr2YlYTJYyN0imffjJMGT/L65PqJkPxZ5psmci1IKZM04BiX5voXTlnwcXyo/6XIsCRDhmCa4sr21ukm3sMfScOEkP+RGT1dO1HHGpqwgS2HT8HirX7IqtnybIeiyum47Xgj/5C/xBY7XjeGzPwTn951+/TpVBxV3dbKCmjeD0KOpPOrU0LdcTcs3IuLIuGwXLw72zleGIkvcbPwoLL5m1W7WnSYgJt7BQ8nFJJLS/acxJjbDtA2c5yVaaqdHTFr+Nc1xd5sCev5fK28AZV01rNbGAbGP9hVausp5Jf0CEQaBB711gZLRkIM+zWO8bK4ob0ACqpNkj3UqR0U/LYSQFOroaQS9y+1DEvEjd+BTEv4e5nWUATaDiWIrqQEoGUcHCODILK5xw93xWJwN88bwKsVLvspSPejAke2P6Eui9u7VVbTEWuqmGJYh61JNrJIvwd4Wpp+F9ic2RY2GUN0V8mNkVXLI0FbvWn3dIv8C7L8FOIUE1IOsVBfCtUK/WkysL8EIAHlKY+HZK9wdUw8IlaRwQGaAasWZhcv3YOB3TMF9se+ZuGS34GUcypfzIGNxuLaWuftT4qluvHoLZFyj/4viorVWmqv26eysml4qeECZ3ec57MsCFsWpTrdbuBZGC956BGsTVl7lXIyeDinYdcmfOVwJnfz5XjHTQp9m9+gNqbVbfxtVsf+S8FZdvOMP987A8HZyP+wfb2NFQfPZWmASxR18IwmKzm6fNh4pjgeXf5VOT48bPaKW5+7Z/fZVdNv12PuPIxKELWpuPFYMGZ7UTK2e82RQ2EfqPIMIuHZ6ciKqFmKbJ3xC9TDjBSAVim6ggSzA==
`pragma protect end_data_block
`pragma protect digest_block
4a33f84371a585d147cda1902c7bce18d396efd28d0432189a3807a3d761ff82
`pragma protect end_digest_block
`pragma protect end_protected
