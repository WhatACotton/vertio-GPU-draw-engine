`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
slu6f7B50TUfQwXyvG6B3GnKGJmtTu0lBRkoal6VNxjxoVnq/9lHHCl/Yv7ePIV/3WcM1IwNxp/XMWQnST0NU41KZ3eM8RX+1i0w0UOeu6upNgeB6hjAs9ZoaNYB7NVihmtShRqI79b0N5fCSkcYi/hPKslGTTZbgnR7/396CDfIpu9vZ+0osinld+CdI9eRA9rqwKEsQdX8Dv0bMOOyfs4alGZjB+vMru33MG6LQBnr6FKj/KNRJ19FveqCZ5a0Q590SFZoqvot2L0wkMlkaCv6KGUMzEl2p9HUOFHtZjC5SqLdBWNWVFvR+umVVZ9FqI5zNizpKYl9m+H0LsXThjWAT6ay8FPFoPsCIuIK5t0Ozz/FzEjfO7jB342D8bKjot5JBueFDPn+fcPkyDQVfBIyef+oB4eF3ut85hqhfQuI0c+AVeCwrshB7yIez1fNx7ePLNOx39rPxJjWP1LBu/uMnzZlVL+pkQawB+i4MI1m7BTSNiLl82fiLhEOzaHtMW6C7Z12Og/1JXa/DxZ+xcA5G6TAmexTsy1TliHhAAtTpME3/ODD7K20rlxET8cgIh+YR5dv6EtnG+wmfIJhpXTGQFG32el8Z9UHbkCJlX7HHfIVsszKudqicnWAVuJt9ACWOnWOGFxC0Pp2uoCKJItyp/GO0UDtgXaodGb5esnL/q0TCxq3mBDWannndOYI51YgkDB3Lnj1k6zVnsIGmvOLS+2BWRxZZibmvD3RdbwPVuqbRBWF1uKODzA2/69BrjPMBr9QF6DZ9K5MeuTGwxnICXcS5/7CJ+rsvo8F+6ONL8kxhE52PWnzZ6p6xQ8TZ85p6LlnjaaVWg1r9haHAFjBrVxdpX2GU8lm5zbPWp5z5wFmWN/e+VShgORbBkJmlLxr8HwV5P2K39d/a18qFlwjkgY/gmNQPvkrFR4pgZj80EcomD26oyCwqNq3vr/Q1JM3j4Bcz00lbQr9ZzAuLT8DF//6hxPbIWFWVemyg01ETri+MZ9+QWzAswh11IZPCWgUoyDYj/X2EJfTYOO0f7EJOPVx/wNp5rWEXS8aY2JQxfWYEXo+OkjPThtGJXILlFGJ19cHW6Te757O+ZD1qdJggyEYCck+/V3K/+hUJzycZj2rePbLuBH9tV63pgWmycRguIBfHgLWRheyED5qw6GqWaMlTW+rw2oVkSkR54SaD3f/T/PtqXK8PQlPmUJettQoK0X8Tr96lvYbzZlS2em8nrYY/ka8fZr0IVcE2lVbKdG7Dx5xIX5UBQN+dW9ra6egvVpD591PmLsdovF4ChQhOH9/Wp+MPcz0xG46mIq0mqyTTaMRDj+W+fnVhRtFA/wGIDq/owk+66NGBy/HKIAJfZlLBGwREVwtHo60UtQB1iU6KQA4z3fJUEya9XN+Uwd5F17eKB4xQvLMVP2sJ8UsDpNztA8nd3HCe59OzMYUxBLrmrQAYi0f7VoUI7qV3mLRYcsOlL6rANyQofa/lywlGaJzitauXoAfJt9nxLZ6IdGilaPzzK/Na00pVrqrM67byAv3XTq9ZEql0RMgScOF+WhOMgYeQR7WrsGem/Z9Asjab2cYxnp73gvLtHHWRZjd9Sg2zTERN+m/fC4dT25AWpDzUaK27DSXZuf0KCKpj2CjDTHaISKzmYHA+/RxUdWKGQ4YvDRF64D+iIhYuB38QWd23ABFPaPsk+9t+ah5dg+Y0dXXsFFknLSTr1IrOAZQ5uv+uVdKEYhpqyEOQdzNo197uZhrUNkT8NUO1DguzM2bva4tdxv93riKzo9FQ4BOOy1/PdNbbeMS9X78l3COF42/iuLMBPZwdT2CuWDQxwAPWCvQ8goT9Yv/Rpzb7YErPdeAuGv7pXJiLmHH4CWC3K2V0G+OWQsYaYP4jzKkCWZ87XPsjkN8ZuuhPiIK4zEAGfL/GOs1XITSAojwZuxmvb9J7pbprYMvh+pQcaJRyOJeFGGaRo78AqtkL0adaVoI/c78ol72UivAIS1SGPCHDej5COBYdKliiQjHO0LJMFPZry5CUDx7mBlWiWulK6jLsUm8eS3ZH4qIGSxKiPy5I8i8OR+mk26ddPbDpfAMr6udOLe6QDoKhIxXdgMfQ41PmDt7fQq97vIK73jPOX46isSoC0C3hEdAKW2sSybbR9aXYEQEjQ5lhbOur+2c0Mh6GXDbfS5y5TYawnkZlCyTWXz9jBu+y4UxLPlbOMeBkt60UBcZ6Wm2f5exFuC0C/1x60zX0dqtNo8H40aHoa9ZDvW2WB/CIN+iQ7wofst1Ya+jlRBrPxyxafK10OdxOgYqZWY4Kyc4ruwT/oTBhksBOj6VVKRPPhLJuk/4ICB7+blIVRadrEXITegrVPzmfRAqxCKpEPHHx4fP2RDpXedaPv9GZuGYmOaCuGbeL13pF/IZjvNQC20uL9D8TNDJErwF6JRq5K387+YADmAAwqEbqLgD9PPojPyG9y4kBKltyTjsS8rOsU397h/BTtuV1f+x0mLfKRzrOF0rduNitQyEw/pTGMYVQAZBwdy93HFB4A44xsGqVWn5rl0BGR8QPmndeUvHfhgg11zvCU87BKVXCnyXgygp7C/X3ewxFm+Fiyy9T7XiyFDGajagWZZ498XJ7obcdKWUUvGNO93Ey+dyVRPlS5L0WiFcBiYE1T8+yY5S/P3BkmpO53EsyiQiyZt789BzILQYXwii95bvJH36NV1VcYK2LltsPSz2vTTcMC+8fnaJCC9mqQUXxWs6VMQWUn4z2XFcV9///qjQIYzFC/WCratQqJV6O5RTprxSujo50TeH5eb9ZQP6lBHjcbuNvFm9cQdDfg1uspe2aY+KQtE1C5u1AIP9kvmLALn9ulaZCD9J3y71BolYITZEyx5Lv0E3BzDWaD7N1/h63vOxh3Os6VvWKgETnATX3ImePSM9z+93ApQtQuCG4ZmsWr4Hxkc4ticAQXXKGUMUYDDFgR5w10g6b4aDRP4ko3eXBTYAI08GgnsnIFQQig3h54OOUz8KJRY7AYlabMxmcFy1CXIQMUCmvlg1P8ZSTHo8hjkFyIMZJBXnmeJjS1hrqZR/FX+fVCaBeDSLVknGTtxyc9kB3+KqZ9BQXTupa2sNTefqiH4OoI2O5JDXc4kAT2f+qEvtyQlks1iWSQD625qsXiKu2ejCd/Va7gfiafJ5KM0Lmix0/qXiqV/iLGLz4JenPIKviopqqd9fX1YZxzORk88BK94MO1fcJGjZC1TKOOLyy9luQ2lPr1CAA7qlVmATUn964OElLXoHFe30boz6r3YVJQ23PG9m6lDUgTRh1PmWLCZfT1qAHkjJdd3H47l3MUfpW1I9N2vsnCmOxjlu0H2OMV3j5HLs3WQUKMOpDWVgns02tFOVVLlhCPxRBm29ICGOFDe3z4CEeea6ztyj85eNRHIRRtIszJ4S5FQSQRGwwJhsS2ROQKCII2DvJvQ+s2DkxIKuDBZamOrDUVSxZi4z1fSgxW5V6eZCg+IaO7FR47pqR2PQZ4J+5YWBfVMC4w9LoZdncAf36F5/3ioTgLd+KgEstMgvr1ZMpmB/79g3EnKKd9Lc/3tzf4D97TB5FOMjOSinWnUuomBJ7ZutEcr9opw/fj6EHTUo7cSJXlDz0gZo4K+bRP+rOYcPoh/clXN9El4F1IylMAKBkcuhrhaxMJtDP+z91VRMOLlJTXzMvIbUEB4P+vjZ1kQymlAwAzsSfGMz+ZhbDWWDxor3U2pabhDE99iV9adHVeyiNS0GDjnkuIowkWfVREURhn57bB5wOEVrpGKmx1vUOD9Ckabgx/YqGkNowxiRBBm474dmnqxdQIIOjfX8+wpeSuzQYnV636VlRNtRJYTmUIa32tS7WkVTcFRLy4xYFuWfWvMc2JcRNerbMYGkMfdQImXTjamNpPmPag13xBz69QNVbC8sHU7cWnW6ToMQUF8o/JIkViZVDYWj++Q5pOius7L9Jlvm//i0LLU+XrZiX7NPFisFcym99bXRFiz0cZKb9dIPPSfQOraycNd5fr4PXwExDPQFVtHMmJwyXkL5EShDMJnbvPDq3S5PdyDsxwMlw7IleKpYsBsxC8g37kwHZ/aE/0CfcuypTE+huT5Z5hORjMQa39rqPR+ab9Q49EuNtji0zx705CbQs0zmKR5wTnO4kR1Kxkx4tmloFn/9TZegPJuvSSNiNiEWWIcTEpSfY0f8o2WP17BGcHqJRV8vm+mzIWEnY3dAe+sN72aeoh/j6yn8A8n6+Hsdq2kJLE0NsgrRloguHuSoHr9h1M/HfQRf5d6Y9C9EF4VSOOkZ8wCxIq/DTKFQPCmPdIJ5m/tQHUTmM7DZO3UYJrVfBqwupEgqPr95QpjXTVSXI+YLur7gVwn4igpmgYHu12YRMQY97V2W+pWksoDZ1V7UXNsfaQ2MPOdPO7SlZMr9OEMn0JHpShzjBtCCP70wdmx0t/qhPsIX5TW4hFeZwdvreiNhkTfrla+eUtcc9PfGW/Zyx2nvq4oOmSHbulxgpZTeC+kCKxsu5NR5EMjBSniRXycZeBdbun4LNRI+eHm7iO4cVC4rBU1PT7zurZoUQlD3MY8tr0wr6w9esdi305nA3zqhYXsn8/fkM7pIRVR4Zgwjj3GbX3XeSf7oXy6XuIFyuASRGMDEhJoKsY9PC+56uTJC0luEqE2NsI0b6/bhB+BdgzzoZ5VZkGQyuEsYe+Lb36gsV5VddYOPc3T3enaUv8Q0FNPdJnje6TnzzqSCylDkfIkH4Vy5OOR6UJX4BK9q5p7I2puLaS5XhDJ/YEAxq+Tf911zb/GWJBu8ewRtqiervg496aZOSIHxH0kzRzdSYEc6/mW5prXtc4eS9EgxY1RedrSy4HrMHnrYQLIKgkPbvG75Koa/0zzWZKo2slQXB1BUooixdEqXvMZ0stFBMJUYNdrcOmCejhz1GvZoOmVba4+DZIaymm9aOr6VvWgx4XGzCu7/tHX8F0Mw0mJn0Zo4KVfs4q5TSyaQ96fa49mLdYT7+/zuhNcbuiY1OoulPGjmhtb0TtL04rUp5gFxpq1eHglWRAdBy+TU8LcSiKxO1VM+1mkSfRoE48Oja+xUGqUHby4eKX35BGQr44T8Kwj1QCyYhlNZx0CaHAfiP2oliwgmD83DfoS98klRD/4WW0PUusdWdbJumbOUlpuwW0OhxM7SgaUJL8v51XNTJ43LQw3Rk3VICJeKy94spkbGOmRHbfAWw2lBLO/dMvlI1Z9yHvcNIYl10V+RBrWZU3O46yT63Rv8dxMpWiKV8Kyyziz7dhurs82hr62k7NPRf85bJICO+TKKcwAeHf6+7voIPaLdNSLmVoo5And1kRZaX1yIaacdhRoyZRbftexsodyjhLGSBS5HJEJ+F7Knr0rpIm5PahiZVBNQEjyX/8Npg8euhHchexRFFVVatT7aOKzoW2fTjkeRPpkKbCRF6QLLoFmoRjI8R6pl8gr5UALbjyjTEnHU838a8Dafqf//UFrdpH9sPybpLyw2i//38PftvQCPkK++Y7TlWdz8xPlydbUaQoox4ItRIG0R9wwp5jDwK+jXl7/jNqgaKZjw9MhbrKq66Cbv/a4an4iawXSTHjVC4i0v0vmz9W/zBMmZaw+3yfvYnYrjspdG4XyYwgTNAMyirNRb6ySrLB/0UuuwTE4FlEl1uhEnUF6kYTcHI2MID1yjpUj89Tybd/EVvUT28jl/bKSju99Vb4irYMuVP5Ybyz4vvuvYy0YDc8/gUQA4rxPfLzZAe8MlNx6icuVY+u6O29dSSjG0p+IeWIYN1CiZjGUNu7D7kBHjqNduev6bPMwETFnyceR4U+QU+D9oO1gpXCnh4VfPnixVgKpy9lG1EFFcwv33f+TUgxaaK6pBQ2W7ogE+lt7FfLUEfGKmXWbZA4BKtgEwjnjhUEWK3jJ1bMq7NX4JPO+WOuehH15y5wsBqywDdhN+3YHxqz97WNkYhYd/kvRJwZ0I86r2QiEa+dktL7Q7cna02J176RIgSgChGYi+fz2/2nw+uDmTqjhlg4FEh4JltOSfh3NAQ159LmnjAFpjhL8BemAL7k4khwLYRPPIkX4snegOTIIn7Uu4PjcR9JJN7gug4nf8J7yv9y8a9SCeBJC9RHOPms1hLxR0QDAsumSPToep2/nee5vq4wJxOshiQcQyc2eTRJDeBaiOXxZFV+vVAz5b4XNUa6KukJu+z+w9ow/zlXHK8U4D9ZhfpMnXerCEKyDPNMcW+K9kXoDdXDKFoTxRHz0Fsp0plyjLLChut/3LIk37DfECJgpxykglBEoH3J6hJruPCy4sIQ3tsvZhy2RaFJbVHfLfX37H7x1Bf9D7Q6xRy5bLmCeDrncp2WCfbsl3e6Y0S7kYM20e70e4EhqFY4Taamuyg6UgVf7irQ5jRydh6FtMczx1FSkY4Tov4IT/FendJXugfQArqCJQDhAy9fnIkk75PYfQRKNoGZCsCjuXnMgpFOoYfQskXW52JDVD8UkIPRIcuOh1CXlkmHH/5X8xZLLWoXqpHh6G7z3ghtGENO3fiM9vtCAbVHpo0x/8XVrvMsIeysWxqmo420ac3zl8POzaJn33js4HF9hG4PdG8qMrlDl4FnY9suGdtXgFGtPyhpBgKDsxnQAVA4Vay09mgfhmyE2XFFTWPO3oFhP8VgB1YT3qt7kHWU4WUkT+jQ2C6dmWwuDEScKFoq0QKTsw+W3Bu8IkXf87EFFcU/AMkC9BTQ5zX7g+vHwWJ0Q9JiAfY+Cc46CZxXcDrwfmXwUv8kWToipaHqZFGvzyRF8tcGaMCo6oEnPe+MzvN8/72reLzhLgXFnbry/a/K2RUubMFNfeUFFomdhk2q0Ip0zRo3bB0Ji+bHuQD2ikUV5XNuddzTELC+k3Bpxc8xS/aVYcJlFGy+8z3wnlJfQ/a5XvewYkZgS0V8sLGxmrLEKxUCq/ak6dHL5+FwJkdNPGmrwHMo2+CGEOKUc3OqaqZ2VFcUVx9azmw38LZkOsboiFxcm4NPfD0TIhXKGyKsFxl1XmVSGQmjIBGofzztXsL/zQn1amP85UjslgAnK2+Yk4lWMtcikghVy/ymsmURQZqGWsPKccmxzuKC2Vcqdhy0FSycqL3EcKRvaUWALXTKStC98mi4FnjLOH6L8mHTZxZCbK7rUBK1Vc/fNfxvvf9YbMchmuC16Z5xqMKEfNJVo8yUrbojZipR++rU4KTJquqygZATWCkdwvG0YJNxIcjN1SWay/xx3dPUiUnwcdriK0mRSlar2FsjjZT+bLEDJ1ccDD8K78TXnaXM3v6fqZh0QFkVNJKJH5PqTCzng+CB8GrgErw2eC6+EVeM+El7JAnvNXNie7BrE7wh65VO33TRsJS1r4Y4dCBjIYWXoH4/JcI9cKVRBiTIi25mQdDt7m2iM6LCUGhtpH0bXhNkM2609OLsNGqdmg5MsymdCz5SS475WgE4yLESaxfKcQKa1oBzI5BE0mjEEyInHzChlodvR3bvD3WN5sYPC34q4QKVVeyx8op04nylyCJP8CEBUNCXzzibZ6shikQ42KqgZ5vcdVKNL5vHTJCaVauUR+MTOMTRfY01UANhfugtJ+wZ2EmFsB5rmRndczZ2xxo2E1t7suvNk+QNbAEbUhyU/YuPmlyqD7hae8EBV4KDp5qZ4iYnKk8MCoh9AdapzxihfKCsJXVr5a2ysXBZdwsK3PubSN0WhmhteNCb9aQ0QJWvOgSUjuARgSAX8bp7s2OjRNblDpZnnBaTAB43x/Gx5S4QMX3dNFZHHA/SXg04pWtD0em1Qg5jWqoFCc/bJm4zCGfUH0vwSu8ME+fmaieWG7pRlWnAJYWIVSyvobuPlMoCH3KKgN90hZNF6/O2Yi3NobWyydz98WYnUPxES5m6FNOl9J3d89JsdBXJ1G2fPuegEeuGHy3mR8hj9jNVyQAlqn7P6a9uTQIhgvHjWsGC7Q7Ynt7rJK7Mk1bAZbFcXgATdpRp1djimTF8nYp0e874IOmfhcIlqayU2Td80oLv0BiekgPuHWULt6MVeVBTJmAbpJLafZ8BIa/qF4uEN2GZqKLTwM+CJEGhNJVulF9UWnxm2m6iXCwOiVaL82hcEqn0X0To0qgJbvh8+hS9hvVmRIJcVsNRf23CIU3LYVzapvAySMKHD+P2T66BJ7sFwgN13Oi7oE4zUYBjh0NC71RsgXhoANA01aCQV+I6Bik7BeMSUA6xPXLJHac+G8pkKn+n9iklawktN48BZli5HTkpQ4vTM2WlKMDHgB7cnvhewl7XFTlZFH90/5JT+CERu40E430u+eKBD0EBOhjhSoAEVC1iXKFoAGNBAUwwftaBIouP4YL3XgnOcY4vfemJcs6GIPSkb0vKCsI4FSyQV40iy6WZosVdoYGbgDUyrXN6jDVsK/EiW7Pv3SB9nlwLUEBzTNoeNyetZ/vcXbONslnPsNwb2ku5y8LRiIwwf2DutIXYOIalgToxHa+pua/SN9haRO5Wo+Cj9Isci2q22XEooktQyUaDaJsHA65xuH8NmvdlYleiiBcg1eXHG8zu4bgvzFgXKFxNiBLxoTB/kL1t1oDpXDm7v90+CgxDMVftLz6B++0keADl9vEgCBLJ9f2m5gs5wZs/XNjrGCH8y9+XaZvnRclOi5djxy9j4voXmMi5/TPnQjU0RUkRgMgkPXtUuEnu01Ztdk+d4EfatjN7qWi8H55tBDC/F96NQFKImFoZzcCOsCZZCec5bRWvKonYzIhHRH7uoJjGImtP2xj7vsHuDjjX36xxYefCr2exbjMhUQ6WRBo+va+orN5IiSKfFyQozfw+VXzPTgiLkZWMCBUs7PTE6vQzhGJPu/gVM9lzUDLFsLoA4ya2UWxT0X/mV8+U4oUTiirusuizVtjfJJAi7+P8qykASelj0IROjwUC4fEWXYbpT4HSt0BZjaHe4SMWNWC7SUZrF3mpAGq+JNOwlXUBgBGnk3mno1utqQRjJOvn6HSytubkNxNcqa2sO/mfCUKiqFttpsSEvAUucWuHMcjrXO1q+p9x6vSY2MyxLXAtV/1/q1RYiq41YdK3pD6jM9QTYqRvXy5CRHTNgL1VUIji2BVyl75aBqgYhtbVfIsZVv9rHRqaFFNKf4Y9lbIdvRGiwefe5REdHG8lfUHiSBpJ6IFNYpkyHY9VPSVwWfokyKZQpFvr8gAtYS7viUcRUE8z1vAGbrgQM3U0w3PwzNXNP91h91cJHMCPhrJHGJ5cDVX8irEqZuUXrq2LN7QSKAiNSsMXg1YG5otCM4ShT+DopHcaC2ZhUIP0vMw6roQNgbU2QoLe5gsu9I/I7/bQGGPxHUXqQSbO1sw6U7MXhbQMTPMiDk8+aK7IVBthZ/BBuNyKkaM/YP75uCXGjwHV428ljG8LPpamMmT/s0PRK+GkPgWwDG494Y3ZkCiPp3IVxcIeQVjuYnOAXhyj8SG6dz/PbHv7FGIFjzfP2LQfKIO5Pqny/cKSWXG9Dw1ZetzAWFEcNRglCslhDC4t1Sf8NLQ06yWeglVlQSUNhhPgN4AvEPwBOySLNdHvli4xZI/s3++Z7ySedrgQ9CuyIvtaL8Lzg9uAzhXGlE7UH4ssaFmv/HRl+OWExva9/QXg95sRohw8PxSpTyEEEXzPGRRHNTphAoxKOZbpa5M/x8pj3YYmKgkTP+gI5J4w0qZfT+O6TXr6X027FfJmzj5ZIfZgA5YTCuupKek1cotu3WErBVXuhiO1w1iN3skA96FVCWvofiIA+5BpyK1xzbntByu4CRtRnpDCxB0i2ZoM5XMkdQuguLL+DgGRY4wAAUr7+Fzgn2WfA4lDCdALyii5UerMJCKUo/mQ3DqEff38UMQP2G/gqcUQ+7mVquEUuJn6W2Gn6fs2SMYg4PM4DrioZ38FvEENLpkOxEE5ZnvDgbC9UcUSsrf3IPMI0PoBsUloppYNrLdpCIw77f2om5tDYNgBJY1gzUCHIqDnWqD7pvrxGgPz+bjWtS6zuc5G6vhxQLMGuU+z0wQSLkw+WwqMle2ydDaJyuHrDxW0+8jhYpq/WhqLNNP8/uOrE+SibR9oS4Uxy57hhxH6+cXhUkYhz4oRcT7Yrv82Mfz2IvtOuavl7Ed50KsSi3ak2KTEZo+XBdYeNqgGin7R4WAucL15eATopuIuKq7nY57fXq19Dvi56k2eMu+F8FZmWB2gsU7BPyd9ThVKiFlcAggLxTtc8CEz8Ug3q0mtMHf3A0o6PJPK6U2gqBsSfj5ye1bHW7POu2Annp8wGRn7X9sMqry1Z9sWZXxR8W6mHVjpPt8mIjNu/JjKh3inUPdqaNi4W4OIMD67EY4B82BgZm2TqMV2t+ICCVreGQI2zxbWn+NVKjWupLAI1t/vubqpoWR6GSMIf8RuZxYZ/jIym0KGexeRtqKAGd1BReUpC5lcLKexzCwSybtFiqUmY9X4HFky7s7mLJhfi2I8qQsi9RraKDMr+JHCm0G2YyPU83zDo3FpOjdLJVI/8f/rjEiUDQJAxJCdemWakMKSyCm5ub0OJC1cdbSIOe4lfplnMh21jZcF87o7/FhTkWzZyl7B1UuRuNW7NonQ5dL14W+TYGm3lnPG3F83113ns8UCgCKhpyZcbhuxxOrKik+BjDt+NLuu/+0hhi9Plq2JNRlzzChyf2O+LwusdWF5KdEoWS7ZuJS7CLPJjr9NkOCQK8YtBEFaBlImoRFV1Lxf8223746E5pXT97E6leUkH77DaeRNHhEtCEqksRS2YcReDO/OhUsZnT7vtSZGbadUlkdwbAao408P3TVAYHo1IBBHYkrkNXJ31K4E3Mxe2zi9KkeboLTsu+QIQoAKxXLRJfySg1rW/tTFN9Fh6D24KQHYLrglbkanXW7CLO1BSjFWNcu9TSPMbBQQtMnIsQgOoArBssdf4e87WEDSm/FPj9GEttBpVo0ZIzHcyTx0Esv6YJjXzkLYDhaXnUcICB9AXamXV3c1/LnbqVCNW+yD1+T9euLZQSQSGa5Bup2YV/8ugILWXNKrLa0wfjxr8bzrcsKxJs8fAkaVUuDG0Qm5T44v99p+GQhBOWg2Pqzlmyo+wNZrOhwaie5+V9J4OXXsWexlW0R6v9cOFK8i62Wyu16Td0jm5KuHeUIxbywgn0VODLrB7K/F3DU70y/KB8mKNuktd4p4Rf8uvxK655UEl0HozAl+5vGIGdwjCEc4trokZSgH6rxrAL8gIfgDS4j3ndgC0tYIcAJmO3ezNY+5/G2WexaKIXTdqxzbtYe7VXsT9qkDhq9gq7pnqzd0423r5N9X3bcAZhx+MMN8RjgUGjxn22pVOomO3lLf3GHeFv4Mp1RdU0B/DVenOM9g0Dk7UBvrnrIxAbbMccQFTN1BZWR+kGdjsesySdkiMXooF18C+p6P7jYziegw+Fo7TyGKCubEjQWSzK9XzezL8VVnzacGd/XGYue4sPQ6gCAzTbLXU6PRJvj7dM2bhizYeVNj5HoecrLHnYvwI94DCt/Wy7nWWLZQCoHekbpJsykF2OapIbO22RWZQYPfcSge0p7LFKCEY3wPDPqtquO76nYzi2ECVnrkpBhjFd6BC7+YNlFJgmeXhfupHFc89M819S4pW6m05ma6PsutMFgID+CquaDzTBQVfrUYbfr32lDolM3pTE0ela3zMaDt/QnAskindfbAFH2/zOv3mxN+GxzItE3LzznqrZ/hCso/PlL5eWROA7gQV5pApY2jJ9iOQv6aRMm2+qePKhMto6whFFUDK9pzXG+uUOXsiCazrUlf7MEaUVvV1lbWVxziO7OF/7dsN0j19zZ/r91238O+n59TKzAd/MI4xESndOmRmuUkelscduu84J5+GKHd25MlKyyXSBP1n2tYluTaJYQl+36nOkg1V48/mEIp47GbSqTIYLg4yRzjRZtZWusef12JvkU2MQzg8yN4ntaz+QSb+GZcLb9Rs/W6vazYyjkZF4dtB8u3s0yb1b9B8YXJh52loml3GQ3gWfLoObghOUY70tDRF2ytZq1XTc2/dYvK0KxFhQ2Dh6irQ8SbjMUZYR0c6rba5+kq91HLYMTZmO3REucgxDDUm4oBZiRUq4/omkwLijfiU70xazAll4RyTxQMBn6zEc+tj5StUD/ER7xXMkKYCBT5LnKuyfctw9S4L/9tbnbqpPc+2VxOcS2GPGMcN9oGYqzGkFA/fdBkUALSRY9FR12zTUfmG2Lt5NmFHuNlTS1VheNkeiXgmbdW9rIIp4kVpMGWYDQ9JlUvg3rRQJ/s/G9cIdnzDt/neHI1MwbP68a/R1EsMGGQ68e+lmfI3M70SXxrvH+cQS/wTYBs0MJbqhAGYDYZwqnhJCV3lfyEW9DHUrrNHWJA5d7WgUNNMRYpdJLgi8S0C7U3IOvVwIQWkixeyLqklzmRCx+u0olHhn+dYV1BRQN8FiEoPd64/9yTGeOJ2ydYfW829IKibrOzxsLoPt/DRqP8YhrnrB3XxmUIJJ8ak8KDh1hcARJxwRCwy+QM0w7V3hXMvKr2LUw12wUb+hVlHxa7k1//AZeEHUGf9N5/LGXbv9DZ2OCf/Uua/pa0HLbqbRVg1kVuNtbgF5QpXBfl6xBCpoAO40NWp1OsOiv61lmrFBOfVc127B4SVJPpbq9aweI8cIZmjysgiOZwLYD4XrYWCm7gZirqaB0B6L8Xm42h+p7qekvkrw4suAAHd6PFV/BM6m2WjZ8V/7idMlugOJi+StIdk30Uwx5Lv+TkHbdd4jasOFT44E9zYvvbVGrxuSjMjCnsYU5OL9fDmZ/jWa0u4W5E5+6YWI0kpZDysSRwXp3GFRhQ4PybRcSAd75QLK6MTZawnBL7fZhqow8cJM5E0QcQO4YkVeuyq+QORG56DTL4cNm/hw7K39c2VK2WLZVY1nRjLupteL5f51sNbiM7X1i/mM+9455VptJ18KUlpIewNo5iqkV5xtJE1s72q0cOl33MEAXXfGvqLvZIuqkYEifYeBzraUVjVrhNGl7TtYGA+tTMGmt2MQysd/tYYd3ZYw964ceFT64iowBQRU85K77kn2oP6cf+TQEUBoVgzAdOT0lh+wKZKEQqbWLUlvpIz2x34Nvw0cdFzmbAjB8+mU1CtHkVj4xlmv1hXVH9ydCGBWKmAFn/1mdTeTXuXeaqHykLZ6HQRjBLeNM6XUWukfX5FfBtpLtfCJVdAHNwSuyAwplN5MufYTr6XkdTrNBmeZN5EzFaBRbHILpEh9u++KEcvRfyeDMWpRMx1mGuRlQuFTntVRtipAgitfnBCdJ+vewqGFLAXMtDkknrDlo2vvUJaHo5lDJuxY9dUxA2XsiaL3W94Ge3aJbBp8xu43TWb/yc8bpykcpHo8Z5lroHlpG9fIunybbf0Yt8bY2TAxScELZBP4Qu5jDb9MdsO05FGLbjXpaK+TrxWMVOD+5H0WDBSklV80xeXTPOF4QG1lTFVmH6kSgIC/8uHRJ26CeiBJ0HgGVvq6p7lviVsdwHtp4W9QouyhdNKagZvdlJpsczxKrqGnKJQojvhaXbUDZypl80Y9yxTvLw9kLVLTlX6GnG4HWBgQ/VZpH/602jBpCu6rYto3y3iJeAKsFhc55rP1t5RrSMGrU6/pxoXxIm2TmYdkpeeDgEwWuID1+5AHUKMofs+Zd4SbhtPZronWVVeOjc+JOTnJs+qPeulDOOsfFAdrIpbajMj3SzPgmOVgZtQpk4FlQ+WjZdr9DVsMolVX45IKJ1c//QmGoWlRZhIoMD3dGOl388FgqiqwqM7by19iGF4LFVojG+EFCz6hu9T+EWuJSTcVRMCNiEW+laKkB2Kt1EDis7R2gPcK95ctaQjr5bH9j01sYXedctzpG3hxIqAR8YpG62YWP9RRDz2oWTjCZoDBtpydYURHaeaahgeh0v5KYnWJf7rG+humYz8t0+Zr6rIRZoUjXs03S0q6aNrtJLhXpiLp0syCdyasfbBo8j0Xfcq8vOxIRLwAI5UwKfk73hmv97ZvFepYG3yFACDP+LkquguHVSdeQpRCH4Cqd56Lr5F2NKXSCjICTVTpjkagr4SEaSZbEzqPy4SpEvGvfVIAsfKFlDlM5lGCrFx4SVrJ9AvY7YMhT7GBghm9sLJAQkf37siJY4ZITHpHimCNR1bsKLeYzRYNaHpC15BvWItQ6LefcQNeSOiPU2ZplXIUoCCDayTZf0VotHVhXorCc+YtjF2St5NTb1hjRVd3pbTtVglf0Cl1Jpim9JzZiHydokGGhy6jDNbZeqOh5MBTyEotiRVN5IUlbDC/yW5/6wz4+qMikRAUvVdMGq2f8Gf5osrClrR9iO5XnbctpEaEMrynk/QwN3FRuBEq7S04B/MAcfS+UUEBA5gGgnzPbzFX0KDG4Uj/t1gP4Re/Oe2t2p556Yyzti362votji4LMMtM1K6Exox0NHDpMT4Mkca+27WOqfmvMP/P3qExhWQxYt8iX1kXPQsm+qtj5HfU/+LuZ/lr9fdyNbsD9jAd/AHaVnkfhGdvDReyqna5vpaUThHX9Zywfx05IuGoU3EYtp7GlZOdWScZfED0ENf/fEynRX5t/NOQMG81sFJe1Z0na0LQ5HVTmGUSUoOG2XQ/Vsynr4OEvO9SDiOiiUgpivqzrGJQQClgp5cSb9QffA/7jXxXuOQktVaIAoQRVbgf6tEUJ3SmQtVMRxqleuPKpMxIMUTWSW5cCNmhUKS1woeAiFIcmIKlgZo08gPExisGpsbyVjVEiBuBS9mE12tIIxQb30SXW/k5yIaMOf/VpuQvf7/BTNnOHK1vtI44gH7yDk7/h9tML7Ur2CnzP/DtXaCeygKSWiRWXq7eV5wwhMBVFgYrD30VeQtk3K2Qiiapf2Hef0DD5MrPHa2Qf2mbY3pdPhuxPu95/dzHxTFDNIOExqEz2e7IXeDjVwrhIfMSMqXIzd7Br3gqUcOHwrq+es9i6lULzfLjsro9HhLyKV/tRkUa0Ke3lg5x1l1pmzNwwfEOyeefvULDVjQ0LMsHtJnpdNYm4vkq2wwOhFKHEhyXdidb5VevOV3bbOZLWmlYVYT2IODGi2MLsQxUsCkPUvfNMAv2YLaTya3opvezlGLT/t5ucZ4IqMTc9jvl7fVi1yZcOs3Alkxdujk+EFh17hentuyaZ2rZ/SeGlNuffR7ju6bK+MJkUM6EgzTrzC4nqGMXhfGI6JGwiGszeEhrl/Zc7NGt+efsf4Z4A/GvS8bDicqMqwDOQTldPHgR88KNKnqmQv2RjZNr6xS9CCTwI6ZiIL2AYHSWLrLlCqHaojFP2+ubTjkRvzbP4J50QEHNWZJJDi+GSC7yS7tQwtAg3nBjtglprzSOl6WM0W4V5EvJNiINjAZsZ++AtO+GSeyq+/lAw+gMjNuzjyEhOtMPgFM1t0VQu6Ou+oBCbMxlkQmhPwCvmrG2Or+FnPO19recUMZghkdxtFgZYRCn4zonSMI3ijL1tO95C/ABt2BJsa183+WUKAb0iTxihUUhEKqFARiQfs5rV0LQziCKLie93Ydf1zgYoaHdwfiouEoWs1dFjLVyB9DlbA12IJRlmeZaFra1out8sSjGRfM2YGOL/CqkyDQZN7uKx82hwXe0nZLOYeZoXgk4vTUSsIQ2Np8WMGGiZLkz6t3IhF9eimCP2vqKpnvPxbPwH+EJ1g46HVojIW+yuDqI2Ulvo2dXX43I8GtLM6ND8w2BjWvpFcrgLKHn1Js+s0n1/pjpU/n2tzJtVoBL0qDdaoK5+fsuyrlaqgpfMbwvLGwrhFSQYKsELgOVUKRreyytMGk2le4N7Acibdk6i9ycAs9BIjb0JzgQnslSyv8KEpdDga7BW6K2u9P3g0e2suE7SdYPYXgHXcxSrGGMgNkFhngjncu0pDNCSlh+UcS39FkNUKZ1xHGIuPGWyKBNRt4aH6V740mW3xNN3lzvtganoaJBEpdbvF0LA2WkNP9Z7EYmsk1If36vgVUbp4eukjfq2fED622PaqTF3c/F4uLNYUJUkpoTxKPAKNZ9lpcqIgBdyIzlx3GMdzkYK0/IF7V+oIen4d2W2OnIO5EIraegRGfHQTQWPevOs+EIrmQ1cAXlo29L8ZP/+oCr5nRwpH9/FUBgTFCE4BMKrxi0ebJ6o2ZbjHHPD4OyujftrpBZYoRXsNRZcBeB+9jfdzijnnvHm34qAhB04gh3p3gxGTprELVnFaPrWgr/gSi4Cbkpe4w46AWH6Yzu2kZjZNkx3TFdwDPc2rQAjU3R+yKjoJcWUpUzVnd2jazFYV+2lfC7/5MRP9Pf5VVLsw/4Qw74Bsyb1pKAdeyh6K2QfN0+zQP0FEzT092sA8lfwE7MN98SwsCwne+0JIi9+9t3MRSPJpSH2si5iRlqmGpMqvoieeFcNKWdb8pzTKI+MtCxczSUPPquTR9Jbjnng2l+psaEHJ91I8YHWXLR5kTqBF8A5yf+N01sK1+wl4IcoRBgN+CQWgNP+chbgydNWy/GUTRDsLIeACjAI0jBE71YVactozsCs8CR3BeK5OngKZ4W8cStj7kuAMWkHaBDIiHmzQSsbIXpTPgJGu7olsrUC+cZnEweAOUWJ76xtbuoZUm+P7xMRa8TQVD3oASqViZxN+HpXF/Njo4UxV8/D2Hc3IlaQCogUSRlvcvw2xrdrHl5Y9Vdm52PK8kciWE95667oftwVRuaNXRcQ5WlaXfOld5GUOcdtqAhzcIuCE4uBhM+uWpBP0O8K///jgA04NCv+6f9TwFhOX/KC5BaIisSmVzx+8tNQnMa9tqgoe8gYna7iRehDjXrnGsuAu4D53+VIYIQjlroqbbke6Iu99vdVK6L3kOTOeI3PJZr7bZW3KdPMMQssGDEERIEYl3KKStFExAv7fShpHq2UfxIsHxdHcp6AV0VP462ENBW8/+JFhQkSBw72XpPulC2oaJWO2RuxqCmd3Q5mpiZaFri7Et2n6gp9T6pMt5YLwc9s6Su0/19uf2CT8C4bZrXRsAcuz/0l8oXlK6lmUyPXTe0pdAEJ+S+UXhuCAjLTq0dzcrn7/DeiztMz1/NSjPm1ZG0cYrrlFOcdlTKeSQfAaDlDNb2c9eZRYdFhaJsU1l7gc23K2kg/0hVAQN1342hREpaGG1yJM4SgKs0HM+05UNgyprLMzQfHQpyWq8YHCZUPeONOuoJWx7MXRBy1KA/EHVyc7gTZoigFX6mpriZf3D8jw9JeBS2faNBeLStJhnKeum33e9NUnOfOMzAkGriRQGuzXWzG2Yy55ScCTHd+IIXtomA1h9/3aVapSJB4v6YTFvf0hQA7nvANlHlWRdTqfgNMkC5COyyXLn5G7diqaR6rJgnqO/dNuQC7d4WajjRB/xrbaVa2FgpPo3zZ32E6bjXuwws8klOxUpAGHb+iKYVj9D1XwM/PQ/fZXbpOCe6ENaz8Jc2RbpK6Vi4Kgqwhotr7JVRVy4bJl+k8kCdJ/U1k0oUtRX5SbyuKfs0eI2MMkQ8/i27W4H2VSrM3VmlBOMqTHjarAa7fRC1NLdtQJagfZI/C5tuJDu6E9ChFRFksU88NqJd6nV0qEGKrGvvh4QI/n5zZvRDrSxs/hdto7OejjkN5xtjnLHBcoLaAf7FI+CgEn/BWiG/dfHnbkvQF3rYjFVWHgq44rCiblfoRa7ZXfRGyInkIKPfzQpJA+3qha/OY1NtSV3btbz+JDqAfUEjrF8hEZOpo9wpG2aZVPSzNlWna+9KhX9KAbAqxydmAU6yqhYDYHQFvplvUwkzZXAoLq2ro7kb+Em07GtrhjOYAj6E7Un9OhkYcrej8Owr2JJFXdxfv2p0YQZGFaW06Bpjej7FcOe/ThMSms2dJFIXWoe2UrxrSxmasa39D06L0k1yq7/E6Cm8Tp5+KaLnh5oOXt4y7tALBf6H1JQMF4NarZvvjImqHrreEN8kyihK+DMErL60qv8F+/OR9KGCCh49856tHlQrcP0OAz67LwijdBEnCtucrqMlx3LccTYVhlcZ2/1SUHVhw2iEoZMlHumcUH9tpNh3NKK5PKK9gflTIlSIbh2B6dR92+gJaSyl7rhOmIWwi2Bn1uqi9hcMWJUfkkL49fGVoLe19DaiYOqXbL146kV+gZGzyt2Nn0krfIu/nibDqjhnzi3wFMBNsCAtTpAdFEgcT2AtD2iFlKyKanm76NgozpnpxsNcaEYaxs3RnbStb7QOREtAJ4+uTi8K2yUDv/Dz/P9jUAIll8c5xXyn5k0XvgBh/uSqyqdnu+5PU6OY8JJwbWKhdx9/hBISLwwiQV6F2bgKr6dsZ66QW9akx5mskHmdVtbnb1yw+iX7MlHrd0JbiitAH8d+s3QSFQ1RxMa32Q11MpNu/VDzhsMprW/9ScZCbKUKQbjNjuooiDevkpx3zSV4gYuFJ6TPpo1rcB7Wv/nMNIIVZ2bHwrAjmVSXxaQ5CCKZJZ2sZLvtoyAkMhmA/CvDxDUeLK+FCVbPoXTPd1fPZYAufn4/E44L4q/47f3NEM8bcfQLlMP6GFAEKClY7KN8m93W7rr/4NhAFDTfZ30aVQYXWkrjJ0dYFp4sTlqOuoxQtPm9MReYwtGgOBvoCkh/In6GyOQG2A2ySC5Ltic4pSklPDc64eb52lIxGL1prNA2gR0aFnoriUghJ1xzHvH8o3yfpTmdg2Uapp7KeMA5rDJCLcI3irsN8J6P4r9XBw8f6Xvxyp9CsLxA6ywKX0RTY1p27mAtsRQt4sjaiTM8pjMAAibBZD7BRi9O1qb2fU5IQqh+kOZvpllyYxcHI3mEsviFxYe8+zpJrZeryjUxIbkxnWDnm2KDfmEvXQ47kHgqFW3R4ZydjbdEkyL/PRzEX0Dp6HScXOUHlAHZXpxDWna3j8onOhbkhyslxSC3BTBLPnkjcaX0sDIhZVwX5Ijyji/uvJV2ZRWrsHzu1z6ajrcmGMXIW6VxhORLUtLP83sF/S81B80BftYQvvYTdJI4h/RyubCmdSY6t7IFfjiF6hD2eLB1U+Nlva3rOmTPlFPBNp7ndRb7VkkkaEi0S3ZUEemxHQwjGG9y8P+niFoEnO2UQNPN/BxonFRVceg4/T643pzw2+8Wo3HNuaOzctEY2qHv9P6WwBaXAUxwBIbVAH0vMw1FyJ8X8Zvu1/1diWP1+gUlkm3Fa0ynaT6XG4aB6JNZlB6U7yVU5U9vvRxQ6bkuIJHbKyXtbse5c0IqVMOQhpD2K5SJfnN+57S/nqMPmvF/zQjB1zkRLkaffGDDZ93W5M27BPNl0vdWPZeq1Z5EzTEwJ041cDEXp3mN8H5WfUpY2J3NgErIQV3vsfkTZXvjhwWvS+EjmVfKiDRKwg/u7FIY1BrNmgX7TiCeG0An4c/EYx6n+YL6TNYFfOjOtqTIPRyAANCyUE8EisWokHCo60eBaaGRKXUrXUNXfVG34yJ+NMEKjH11qxQ9Z45P5oLrVm8NXMhD70vUtP1dEe7J1fvoWFp/rlNJUAr7hi7jLtz9P2IIUq+8MDgvBnooyLkp1H2/pOKamfafhqzzXKLSv+L80oUua68SRBlmpw/RSJ82f6s80p+H5f/PkWo1Q421wOiWfLCJJduAyl89snYNcM3ruxic8qnyYyROp5IbL+gWJ4SaIwCb1WH0afYsu+lafkNtoAEYX6mDQCX3nJ8yThMRxfBs998fnbWDDgzu0gnjeZX99neZd1645b/P5W6xAmhOmzFsdMS5guIluilsK5qWR/98+bYIhb9INeHdlnp45YpQRE8W9Hx/JiLDlZlZA2fUKiU6/aNYjv9Jz6/NCIOnf/9Gt6E8N9c2bMbY1gP9hmc+VGOwS0/FugcCaahOXGCceBdRyQ6cyUBw4VxFOpdDxQFCHL5z15nOr71OZ3mSUOUj7WPVAikRzLi262XeKt85S7FxQXuF06/jRkmFSMzbhhdkqcmPCblrp4SFEsNU60AVVajZTedMHhBgsNVnoZTAK2h22noYaK6DIUiDBudEBx15XOrMHFLW5M0ieQ27UqK2UZwOYgFk1RK5zoDkbuX1aVe0N6YluPf5l7QDPpwGi9BcCwXqoTatIL6brDgieGzwBt+E/swtxo/bCxpreUAGiJ59HTw8rhCpzPDdFskyH1jxogt3Go3TsTpIS+yE1gDPxWjrEP3uk6FAWGIMSlZNrpKfV40KVcRuvYsB4idfZeaCasa6ERMGsRtRDWWI2Q5sPxP4tz+WjZqJ6IIZeF3HQN/V4vm4M9jqurysmRXar7ChpVNtRJBct0AUe2oxKPuxm/B+sPWrfhkUrm3jawtKfNkVOnKkAPx25BT8Y8wbf6BWRA5qeVF9siJ631mZ+ZHxf9ThnnwzRWIB3c48E+HCjq/Zuelp0384l3+btReQjHyDhGl5N3ea2fCNxPePcYi6IaXeXEhnCt1Zl3rh/of9iFwAnWNJm24vZUmN8PoKsqXauxb0xr+SUV24yMphoweV+wOo+A07V8jKs8yYL3+0Nj8rGXV2CUl/9ez9XyoZYewMm0OoP8UrTkkgUD4sBBppswsBpXFlFM0pYMaG0pVZQR+Y3H11nfzWo4OvdCQu5B+s8PQ5YQiJ1Py+VhgCahVTvpngLsus8UVAsyqBVOMHLN5C9TOcFCASwPyC/wXj+FogAANrZdVBClazgbvaPbQWEfZ8aQhd1FvqNMjLWJHRzTCtI9iagSMJM+Jl98TfmlGa1b1vSN+wOJfrSKRKJowCyxxbhRW0Wl5mpt0T7kB2/5MzV8KuCye/lbfCfPz4AlFj8oanhhl6Z7YFfC8jJjD726CzMGNcxhjE9e+IMTewLMYqJBYVX6Tug3ntCxzZrS+Q+nzsxCK8jAmZA33qPq2JWn4ch7Kea0fntq+xjwI71wGakNyy9pZ169AfJ2SGeFB0iQwpMc8PBfr+Vbwv4QovptFBm3ZkeBqXFnJTbhawUd674zKWCzUhbkUi5zI1lnHXf0ZNY0zFk0zHAkkbVAZegqCgvXUoxGnCzUOve3YwaJUuoWP7nMZJpS/UTldIxs6C9OQXhVuhYqhbuYO94uSOecfgPiwDuPci//now1s++2ODl/8BC2GpCZ8BQIS5T+GBApbSDl1zBXj5e6tFMP2KIWTdIfCb5tAuKhKPsBr8mnD+gU9ZN0QwoExLy0MC7C8y2pWFNkQX+UV3TwQPvIOAENi/He3juZIvzVSUHTlS/+XTRm0jXsLl9OtB9cDKh7n6NUBkQNX9vJ+HO5sBQOOr+Ml9RM0JNaWon2WLSIcfZoRygmd9Ty2hK8cdkHdR+01jMipcHb/lCNhljFzcwwwNA9vsOMXmimrqkRCDjNrOwDGcwsFkdemKEN2+DEUqgb5AHK1/JJmrjggD4HvZCV7+85pHDnJfCWU7p+cwuk50+ITKWDfPEV3kwESisbO2RssSoaGhumtCqpKGEZQkuX55e07RebKpmHhTv4GQL54Wh1hUZld8Gtvs3T3j0OzJV/XRfBJ1volqydXSCxNcBkbXZKayXxdQzE20GHDJQT4fsPgd9gea/rlWbjKSdftBdl06sltrh/Ek1UZqVoNYfLjYeoZQkGdKO81DoFgajTQmjh078ZIo1/DvHteuMzLuSOlFZtIwK1Z4pnnQGHHIJp0LQSrsAaXHQES1Hbx3mGTvCTG/gUx+91iJHmWZGs8IXm3c1IFsr1HD0XVsLmzyU60Ytj6fK7EiRQYEEVnac28o6O4ooutZ/5C2c+4ofxIV+HkaqmPzEbHzqf2MFTjwwuevbjxqss2nYH/GGmA2A3vsgGkM8uP6aaA8nI0b5KY/SAWQmKFoWrhrCmx7WAq1ZVOiNM0Y7jvfOIvGiN6yYl7e/il7qDFTk9pR6ghJSiqEbRF2lyMGg9XVCxyTnT3wlPJWEAg94bb0C4Vpg6N06KZXh4RA6dPIGsd3f/8cfLa2eaFjOZceNGpUBdR42Ql8cJnpA/fWHrF45sM9G26Bkv/Fehgix8SYI37wIHcSaV+bk0g3DjuYhOEeR1AYqiyNXE5cDjoIQ1yX18/hSy2hdTi5ZPQbtfEGWD6PHZnti6Dve2MzyR2TE3cBCkuanJmLC89i1fwEPL3qFJOA9fMuPF1MTIRdOEr3cG/8Q5yUCINxw1M5Q8D5nkdQ8d4KLRvsT0GeiN91od8SKeOxWtJOIkSf1T+5d4IT0LSBsvfepUgU/9F9cLrhmN9EYOXUbWD2B4FProMd2tVdIP0gBZpSvrHXrMaXXK3/AvE75GVUNTiMEoBVSMfB6Bwn7jDCRZP2UKHJoxCcsgqiC5J1XkXrqGxFnxsWmbY/FHzj1hh6u8xa3b4WcjGBOcVNlznUkOMMXUFq5CkYSmyhLHsrylHfvtLIBj068u7s5hvzSDsfmdaMr6qSN75lX++vgQuqkTCLJXdiKGUbYgLKRaQTTbYQ5y1NjdR5+hrLAXFhuxLbrdlL7NP12SMb2hWWRKISg6HFF9YCwtOOBwC+X5XC8TmGqmDDUEusY8RE6Hspps1PqpbSv9vtRWSDiTqpTQirfBsx0kZc+9IbwxgPXbk0dC248MsP6I7ImWTJqZchf5Ngy+sFHnXnOJoJaKe9cj35q8XNxQOESTSnaRsjHK2EO9HmLpSDeooDg8beYLmLBxZnQRBzsDE+gnqmJ65ki1WSNGK+yGKcSh5GAFpMvlOxM4qpOBvjDR3uB/3xN8ZapxRKWZKpkBHsWb7wEXLZG9S6IbmHHi0DmO7huXqF9dAJaZXzkYepDBdi0iSmS3EUWrTr+XyWsTvF1gwnhp/sCxmJ8CKYLbersVvg7zfNNOxvLqlmgmrdxyti/7Wea7KeWIRMbvnoyujQHbUypcgsBnk87PppJkDrLJeLADnjotJyREnZRZZm49qJqgU8kIQImElh6X/e3Ave/lPnwJf3B1OUiNY/ReCqrf3tsGJxHpACcpqp38murDg46Uz3aMe6v6vLVZuISQhNeM0iwPZodUTvKlVRtU8TeAoIliD31sRJK7ADoADfPv5Xu1GP4YXyYUwoPn+NKAhBHSJuSALvu1mNaxhCbh250l1A7DUH1gf8SZyRJqBD1YMPsgom2qfl8yevZvQYbicOvB+NJOgDHUomTxoyzEbFo/Y59REWADKu6iIvgTctcRqrG1sUQ8mtPZTvSUQkdcV6PgeeziI6YT+u5/Waid5LL4u7EY5slY9B8fQtpNPnB7iVtBKkqMsscjaY1LRFfSvcXtx//muRfCx+HsiEyX+XEJlU89DVStNdnBbPk924pCVQWybKXTxq0xxuP+gyRTkyfzf86Mhetr1mWJp2s9c9sVFOLC5MigNU0lJok/qOZ+F60WfLva25ONW5zBV8UtkDj1fAq9DzGLMkyBHoUoK0j64RMdPTDNdxGEgH5JoqXkbWIpRjYLv6AS34d3RqYgWKZemjYg+RwchcjCrJBEr+iLJjfa+gC/ghyoiuOcLyBCI18OkaMs+utEWnPtOiS3+BDgF3WgX9qeZJ1RVx1ULZbrzAtfx8zEJRQG2sHItNTofGxVd/8lg/OFmbJjy3uFbxT5chXuE2xpthT1Jc15MEs9m6bh0nyTpMhNFof0lreBQoXWdmbOLMyZ0ru4MCJ7zuUfEEsbKP4sKdrL7dILa/5G8e3IEb3LAcDPCH11ZWyqmFiDAc8CiEOxQo4dFQYnWLjPcWwt1mQ/sxx2nDk9KX5jOMgp5kxK52I7YMnR8cs/TpN/RRgBmzViIQaQi49kIh13Y=
`pragma protect end_data_block
`pragma protect digest_block
83bad2704b4c3a39f7ed7e08674bb4b9b205b8ba8d437a7d1d9fa185a5f6187e
`pragma protect end_digest_block
`pragma protect end_protected
