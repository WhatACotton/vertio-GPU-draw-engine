`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
x23nbHVT0b1sFV+CTjF4h5qO7OWiCQWLVfsACdXDu6WWeQQhb5vB59DBdNeYRjJIPpN6RQiHj71X3PpLlhaN+aMoQY4FEplXFR7q8lWgmIkHHm4nZQIjbEkwB+Gf2SkOEIjHo/VxutZX1l9QH6epThWheDfWgKhcR0vgN616E4cvAgb8oORS1FL8FcSwnvulN/3QJZi29zKZTsQiDMqjslQSyJojYqSobcR8qYzUIvac/teeJW/+up125mlhfeHpRQMGY1GeFbwBTv6HGWjh24TQH4wuJJ3jmxf3lPpViexQGVwSuej0PcKzLpNS+5moPc5Hd7tXaW5NCXe6Uh5eZVgNHMTmT1vPV7v5Wutakq1ij++19ex7rAwP2t2r+FyPzJGaZNpy+xd+Luu3q1vqsPQa3Cbl96Y7FMhG4gmmqwjKH8qXg55mUlJMdExWjzTwSQ1f0gBCznpariMRfKbvv7YXJ9IOcj+m3G7wcVHo39jwm6JGt33aN+bueMSkuskglMdTulXJVzhPtQjYXt0/5lIObCQMHQ1YDuho3JRyQHdY9FKOdkPsPzp+Bvp1KgsNlTWnNS1Tv+92dYVI1LJ2uTKsw3fqSRUG+B/WR6YHz8pQUhEAfCvR6M5WFPmvzZc8Cm6q/l8U9to4R0aeY3nXUkCN3omETX0VRSwQeZ5BdHDLQ67e8c3l1J2D66JmKl0940IkVAYCbxVDfczQtMwAGKjGJCSvJb/qvHikVCeWdU8LExcie/4+vSGrEX4h75d1CzFh3I8xiZB8kwzixAc9GO58NbrNoA9w4pdVquvOGZ0Luee2NluCD5PM3PzzSd5cwfeHjT+zhYvUQaP/mwX5xOs+KYSks53qfXnlN8dW5eRgLDxB6SqB9c818+aXk1bdg9t/jQNkqxwh1TPpnMTdcRDq/6x0pr+v61hoYonCRtlc2QnHrnFG1LEkHGaMSToYm3m2LirBTYbJ/biIdVxylslDuhqdeUFDM/cUg7v+J6Frw9cT8vBd8JBzQ5eH+jJNXSp+HFdpF7o7ZFe69hyapQvj8z2oke2N1BCC+Ea+cBS4Tp3ZxjJ7q4pk+tMZPfUEoZ5bUNBmp5+rPBwZRzBSTDbN7uyrx5s7Y/PZG8Sgv5tP/25RVVTQ5bPuaXbY/uQKtD6GqBwBbGjIWUoB3yEE4yEi3HYusNvbtpduG+y3vBMewHG1ONW7hF3DFxXfB9Tu/WzXD/IKdAOSasuzn+1QIsYTmpExpYPEbWY36kFjQRIrV4GpB3CeXrz84i9d4irB8320+hgii7qECXjQW8Dug8ifMDQajUJf1egwUdHHoOY/iPDALlupjKu/4oeoTFijmVUkodMRKv85J5DcJU111wGvQvo9MGzSkcVv18sayw4In5rx70yv3JtOP5VbBfkhLmSD1IcViSF4e8EVFk5zXMYNMquge07s8Y7OcZxv0N22U3ajFfLsQJZF/S2L9M0pJ0RqtdwOcycedBwmninNK7MKDIxfPKt4+NR2cM/KuTszcHvW/V9Owfp5lZs08UMwXu3hp8ld9V6+ELHcC8IZzR3qAJYCKpI9e9R+KHK5dUrVNhuFSxngZdg+/VLDHDx3c7z2o1gyszkrA5TwMmVUO4juRLM14XpJ0aReCTXomXIe3Dl9YY+37h0u3zRg4Wds/adHiskFzGebX6m5K1mFGh5jariIrDcXpTLa4qZsVPtTXCkbJkbbmi2Z+dV238Ns7AL4DI7lHqX074Mm5KwKXIzO+vDQ1n9tGla0SGL0GlKZd3JA8ST2U1q4pASYuJKdHVED4DhLoMMqkMkYzkYTwL3YWdxVdl6fxUGSGCTJUKg2NnHEme/zPO3O03/ynSUwVHNXciJxHyEpb6ViCTnSb3KsCli4KtIZ5eo4awzNLPcGbJpqfxgHYDc9/7fROFg5kvNg1mvKmlb97cINpGvlLp4T6WJM4CdZcLNh8f+O51xUnCkwqTc+mhF/5JAckMk100LaxCtb7NK46Q1kUuXjKdDv4Q/QJsdxo95E1DmgTf9WdDMklCXqrHqPYf/YU8iTNQhrIxmbAWhjuoCBLE+VE51i0jJBPe+vbrFy7JbYvMDwxRhjaFjZKG+G4LfJ0JZtnkevTDywai7jVXwum+S6R5izq0d+geeSjFDhTWC9X3KMQK1s1XjZyAJhI6DetkIm02giR5ToqLLugUfIdEfYzy75K1Ivpqk2wSpz4SnFFjf5ifvtBDcMoeMy/Bz/HOerJQTYljoNi+Z+2+mcQJwn5IrdmsQLssPOfg3QyC52Uyhdt/8bnWWvUGEejCY/UIO63OEUWJx/AEZils8X3jEsrP4wObqe57c8Mn8PMECdC0R01SiB5seJzPXwfNLmJR8OV0v7wtRbwiQEMT0CF/n5eBy3WmpOo1GdGiy92JKBe67BF4FZHtxdvBeUxlEG3ZBGx2Tfi+3/OwS30NJbfu4xFls2zN+z3AIWbYYvQXpBxpOk8NdcJF8QE0HhU/zaj++IqJlcMRvAdjY6COeGm//aRCl4Byp4K+UF+QFJMboipdeFtOIIe+gBArqNR/A0ozh9dlOtpBtli5ihogRkpKeyRwFajLGF8xqS9JFJ2lQV/9TG4uWALsReCIffTjcupBzsn0Fi8KQFW4UzIWeLPWs4tBx2qCdh8omuP1SxqPnpS+xhiozB5wbFrfS1OrFUz72QeGBMTs3u4aubaZKPlU8p9gxZ6wBMp5RaWfFrO/ZbdD69fzvwoiHMiJNBkdm2ntnWfA8hUmq3oSaTslxSxUH2ac1ymQBXfVKqkN0N5Sfc3yLnCR9scPl3ItisM7ubnp/iGBGux3y5gTXrWm9Ze4GoYRo/OmPtxRFxmw3q03RY0jQr/ofRdqomDEtQTLfBv8qpNWK5rgGOROlqj6+3DScgt/LEQYVhsRcXUbBJiRdhCHKzmP7byfuqS/1oJfX5iq+0XJzPgPtlfGw8So2V74Ry50OMf/iz8Rs++Hlr3pTytjYWpibKcyM0wFO0smaI/XKyxsacxRi9xaGOrpg7F3L1mnSbmaFsYkDUeTUFh8pr34ajFCPubRw6VDGEEpaoxAzaIYwvgfv7+gx3DP8qtx/p9HC6xIAVeV5ecIutY1QkpnlDgjARq5cEmU4CtW2zGdFm108L3QZfXpn8gMWB265CWsIZJrT2xyYbo0ypNFyQtUm6fBJwq8ZOgsGSHUa7Tb7uNj6RZ6P4hJwP98YuQDWKIuBRHjuATPvzD2ujbCmX2XDGStURlnrwSzliw2HQ4RqcsrZTq/DWYs2qcmWXpM4kEPhYiDAMnsmEf4s1ykslcSNrnw76M7+Pbn7XCibzQYcwUkaYPDWxa1SEgAHWVWbSD55b5X4xNY2J2HQpeAUkeQp45j/kywO+v5uR0svnZ7l8uD3nb3AQzWAfb58YiC+m8BE8x2nKN05sql7Q4K34gZdYeSLQChJXQmdVBFUaOXqFyguOrL4hdqfA1BcK9uSxfbmRK8my2y1ZYYsGiuWTSuySAmDCAns6faQh45mxm81pJJHpnD3zriEjTBZzxBk2ATlG4k/V5hwjFzJh4O+ud+e1pYaWmmYRKkcWNMo0vV8yzWU9Zw6Pcjk1ufZPYlPgmPURPuhKP/JmOXNxHAwCWoAWVMzkwr0FQv8xDvMuZwnX4TMq9jSjOCqsQF78lesmRFBB8bNmzeUvaxgXxrD9a/j2NeDLfeJ+c2sEHLmVzHN+kGT7upDZ9e4bFmu3pBw28RHWww8cxB+R9yZX2XIoiDjXjoK73B59IpDuxcrIR71/TIPQpg5rBd4Cu4XU6a6fZoWFZTsDaMw2dnzOZqVbiJqFfXm0gqQMKz9FUdPk6DEN7ZbOaQU3qLMOYMk0/V5teTmR4Wir3W3WU9xs4KAIOkx1Ee01z17ga53Wo6VneLKWbggQ+t8BaHG29ipP6IkLjfcklwDvhuw4I+AAfObSnvIIjz9V8hybljR3N+V9dXq6HdGbPQLJ997Niq4oWGh4Yj4TT35fCZJs7Z6w1qKdIyJXY4iE3tkhkSdD5WECefUmK6WYyyds1J66I3zTom04ha9X+Ou9AABLq5jhFA/WW8YlfwkOFCB0V8PMFp217ZfQhHgVpRqVlF7DHRhj3yARg6UkpL7qA0J+Aeuk8U1HMoW2Q1Nznl6B8YO3wHLxTaqOzXBB/xqxX7VsvPX0uiANsBROU8BjaO/UfAnqpuSTICRtDJ6V68UYesdo4SEHiuFNNu2h0kTbBviJWthYG7su372s7PRu2HhFFQ80qJH7kYJe4DMGzJHhLrtdEBK+7+lfI3ZM7Y2kUop88EOSc8NDQC41SbQ/AhSYC/3UV4r0eLL9ZUfmW1RwnIuZXaswombBg+VivhysUQmYhrLNkifs8z3tLegVn2DUw5u3IGCvl7o8gMHrZm5uVd9KAK4VEAw9s/hR8f1299rAgCxpANX8Vwg3MJg1HfDcmWlf4GVPkjphYJ6ftMeX0RFbhaL3tnEpsSFjo+juosLi2RnXxfgN1zrJrfL4Wfa2UKJmTSdulnF/2GtchvtnCs+9ddRZqn6oNxKU9oRTNf/Q0twjE69sIFK2eHXRozeYpuWFtnjV+FrJlnWWltAa3PmUs0K0GHqVP36gyCjgJPnUIuvqybWpsHd0auDFHJmsyWuUANDBSymqPD1lcVyc89RMHYTR4e7aXp2fMX9EGIDX1zOf/UJLsJD8Aw/iqWTicYqAYPRoZa8tLsk0q0U6aFD3BvXQ0KMNoYVyWwtl32IOBnchOZwgIoHdhlZNS4l0fW1cWBhHa9+G0Hy9kGbFZFMcv6Zk3ZVpMn2MacO0HA8AJkkmeRpGtOwHWvVT8T2rogTwwKz3iHfU1nY38qwGa19jBCfqPXUDp8nlzokS0W+XMAyS+FtCVw32UQkx8CmOBntQPUDWh0UYvfrXy1+zBjrGMZqeUt3DIhRCcqCSh0RqKwhCP0A0I+7Lj3mK+PuJyAQWdY0FggCia8klD1APXSml2967h8SLrXKFqqDLQOy67yMzQTiTtQ1KWFLnjbdQ/eg8VDgwRqAiVV0C+aGzaRi1Bu+EYAwG6+kHXn7Cqufl4WE9rFJXKUfY7lpyYjImjOp5ZMHmjudgwQ+2yIVGmNMQg97T3peL/T44dabIfTrQTWxYJqOydiXzOC4ArV4WptZtsfSPCyBS8M343xCSESPudHzIwIPHOj/CDx8riJPdrYeJZJ7aOleHXkjzdelKIAdKeaaPaxo8R3ljvW5hmIJaeMd+d44/RlPx0W57Do76N8k4OxwT4EDUiRPN5qlzo2QyZCKeeT5mzr4Xuc+C3Imb8LeRAJBBDIlr0V14B1OOLfrqTR595F7mQAwJbKIIhGjoVIx3HfCqwCjbotBowK2iM1oHY1DpqpdfLvUyuqSh5X1Ve35kVI0v+1zDoLAxKGsK0xnWDW4WO4dtBAxURjOUO4FZZoVKH02JFINV9/VpWDSSqKdaEhsRcB2HaHpdCev4rOtyP5UCJvvjjwJhacaJOR4pvHy8ujydRbKtLqYc4T6+HV7hgO5pMgNhTpHECfAxR2o5grH/3iDZhh76EBqFt0cok2vOO0pUBFpRRwOuX+yv3FwSyrMhVIEER6aeH7hQA52KJFjUxrtcxcs0mgKzq6hTbh5wxBbNfYbesJTlKWYcmwHlMyB8vObY8J3AHpaOC7vSj8tY+D4rSDX5vTPY1Ncw+YC3AppnSVmL/S2GO1RP1+yDg+fmTzD0w3js2yP30yYEwiOyuCepwBtvZ+mwmLd8wdpRLxw2Ck8vlW73H2//UXsqG9XWtm+GQ2KveTI1xEx2QEzViYbD2yXA9BjobBlic8vqmW0cu7VpDGpy0NAYwD09Dz+JpYsl2tK7USMB0J4tsx1OAwdoAS52n4VxAisdwPRADVFmiO9JubsNCPtJw5odUch8DzDFYxoPvykrMEhyJ8hkBOL7TOjHhsOjupLVnKVYU4GvpBt3cpMkQPpZZ61VlmV+6eoaCCiUOWLZ+6nunkPQaXIUpg+uaGduWM8JZEAqpYgtkZBMjf1MvEOIFtNkDquSBN9nrMroGOFqtcUVVuUcYkyfaDvSJUb6qpY8ArxSbI2GlENbLME1W2Vp+Qyj9RkN1ztuGI68UCDMTDnwUstxVX4UF/NS1Wsd8zg4DOGSekawAA/zdZZzp/A1qUNERmV838BuK8Jk/rGGPNI3LkqfeRsplUk2VGFGISgHCpQFYdzgvNr9MS5RRzv+iYSl3LA04o20wPdXYMASrBkDE50U+wzGm1C6oVpLDDzwAy7BvIfCcVd2st9tkPAnyVa6ckhktGxY8IkrqCtCuYKifUkQ+t2bs1JCSgcADGUwBa2hl3CosdGXRfIfY5jTSGfUpCX7jGhaa4sZy4ejpOVpZ2LXcdnnclKfUKrZSMsGBEoWQo9EPA3kqcsyq0W94eCY2H8AQnWyED3Q1Cpx3GuDlmhBnTV3kt2ZUHtlvblZme6ArvMPe/p16f3ntL2hW/mgKvXhdSeew5qWgVfUqof+YWcRu5B696/8Vxd0p07aUlRxWfwiFcI55q/nJVLXMLnisww8CKYdiRoaSNyZS+0wkyY08vmUUu38PsnMhUUTbrBrRZDIAB5ogdshrKuHNfDfYsB0iFckZt4VKVTcaX1izgsAf1+F1naRknFbHHNw1FZpiB92zJ/LqeaXpuEWxs+bIS4V6jbihpLVA7oKJAkE1eY9ac9IdIRHC304pXYvgqqVDb3l5wbf70vP8Iy+N2vSc0DWd03sUz83dgbGZ85xcjnDtLoP9EffGutOJoGgpudo4liG+9yr5IIbpLOkrbGPuvJE7pLsfEz8DEnsj/oBHR+OuQkhAX21F7CgyZ6l/5HoCLM6QG8zcNWsr5yuAqQ/G880b34IAIU3m2lNxBJd1dld7JNgYCuyPsHZJP7WvaeOkTSmVYdpQe+JdW9qDv69Q0Ink9hCydQm8wh9pQSEBPd3Bdxc3+WsmuezJ7EXTdoRyUoPTgyJVt95n31GH7LesuQYtCzDCcel7Jt+ZXMWacIXvzNLrrx+aPtwZkpZRbEVkMCuMJsRnwg4W0ictSLNCh/aN4SKaicUXEUmTRjOzTnNjDJJKzsAaYRTU7FXO5zUNeo3Z5AiTeFqgyRmtNS7Y4drZgEqDMgBEalR5N0FUpZqp44ViX6znkT4dxUuAfiYLygy1fN+hg/1ypKiVooYVqQYj9/dJ/Ae9e8baZqHrthLVe1hfSARKc2lnMNd+9wLBJ5ZpFrW+N4QlnxEDlUjNO1AjvpeVs4PgvcP7tUUfEpSfv3rPcvO42F0KsQncvkaPAKSXtm5aL8o1fl4BZURlAdOdIRcHdojgJW1LdpyhKbgp7vX+rxsY6BSBLbtAV95vwD0NbGsxBys7aTULK6VW/PJM5FnnWgKGlPMhZvkgeF8VnH7tbabTwo7splYbWb0UTkMIV6cDuu7vz/AwMwoee7uePY+MoNI6Ekh5xba4+eeYkfsGAOQfAjYfcUmOMjVdfRWbdmD6N11cj4XH0KZ6T//l2zXQpuYxHasvW+UxAU00LE9OYuwsqETW8JC0ZK3ifys6cI4zKRVyndygd1f/t6VAnZDvtBbiTSVn5rn43CYu8+j1tDjYx261ySIjSRZ72kq7BPoo4ZgmdOWit3F6MxnAxq7asWcrlaYXocf+cF/GViCHU3+DdXoj3x8LGPwBck4rDgceND+cZXhUsFgWElXtwPScSKgkt42sNwkEFqIqvTImiILR+zocMHEouhMjfHokbOi4vz8iGgP+2d80LoOM+wXUbOAp3bvtxaZObeVJ3X5+3oCTLYbmlphBz8uXkSJI76OOK31wYKV4iPhXb9j0kG0TCzNAfmNviEfiPWnfMYA7GIIuCVgxEUbCTVebX1FkfMTE1je6Fo0ben7F6WbZpAnZRgKN8p8aC97zFuRppoJnu7f2AeVBpUhzzN0YEJRxojGQNEE4c6gbR2Uj1E3aDZqIRb7tcXugjczEOGnHxsYQpgO3Y1ksl5NODcNBTW/DClrx/7I3etFXfqfr6M+p4G/6z4dcIfDc+6vDoT0SGboAb+4X5ORoOBrRC5kf14gRSByLci1+LkQVyGpK4MDJAHX2F2jpZjwARz645FPe3N7He30l79gnKCbT9Fpi3fBetGOhI5V8iWb/l/r0O2L+o8JlS6I+kvskL1nK3i31GnpCeRsu+d9339++fxCK1sdyA+M4WpWu/VzTdnzMBtL+y3l4EGiIEPGuFLN5+xvCwPmoYkz81Xtndx/raIOpyMZhKvY3sd3ZOx8Q8hnjMAnyPkQp5Bjtvnma+nWiwiX84dLOc+OsTGO8vs7qxpvLK7BJ1KV+bFpUIj3azgoUsbGGuZDcSL+eamGqZkf3/x0C86NNsNVcgcQKy0wFAYDT6cbvWT3GjcgtxeX2LlR+ehM62d/j0cY+2qH5TVPu7HbPM3mtdR9i3kQIm99U24wNrSGVLh5BHnw4eOqvIEoMhN1PwZJpFC4UEdhERp4aqiNbfmtrXrKqukM+lmPR+jJzSDGFZ2S6yo/wrDuMa0lNkeTTarIZXRyMWjUm1Gr5WPMsxhDWhqWaQzCQDgVgkkWVY+5sGf6tNAk50vizM4AMnei5Md060KMlKUFUb+mmSHHXdYsr6UuVjQmUa35LHmc3kdFN2Ui4qkvHEY8nhmHGsxa+3g3B7EOcUK7lu4h50X5i8txJ5C9wNcgO9NcrUe31MEUmZiQQ3ryaQt45n35tiKu/XypBheIOdYeky29/a332W+CBLrtiSs+9Xwu3T8Snu/fYZSjkEEdft/gvM/PKAkXu24zI3Ok5JLG56nr71zJ5SAS/ULcM7yZ7YqccFJDe2rkVG0bST6tMXeQSjCrZW0IxdNy8OMVXljV6L6G41OgUig7lo+FpUu6MxAFvMwisSXwPZYcjYTZl17wPFb1rKKq2vgctgKOsvnxZBneRzv18yObSBkQHdTZ8w+j9UNkwXAv1ZAo867tKisS3E3L5bnGgplBAZzjMG9TOJSgOInsLS4aInuR6wrt36187SoLEBl/kGIoeH0FGZ66myqW1pPTVBhALcjJyQRKFuxEflGG+J1HiCPuFL9iYBU5TNZdyvmrgBT+7XDhJ8lOG5DgVP31wW7q6VYzP5E806xHUS6miLIhL59qmG6/0Ko7S1yH8rYQOX5i5ZYjNBJnMDUC8edE3r49u3r2m4N/QmK+mqxM/V9xdHSLmbMclZ7hECsVQZqfIoARUvj5saq2o3gzKc693+PXaVeb39Rhb7u2aExNAAq1wqmb+JxHuJ5KlMs/pVhoyRvUGdn5eiqtO5IZ/DX8qJSQw0IlrVaZ5mZuypE6/cjUkfE2Z3MBg9vy0B3K9x4k15iLKBNygFCAILOPC/HmTgNBOLc6dOJO9bu4L9OmJmO493Sji8zh951NC0yRpx3TZw025Z1NxG2rvSBj2cZe2HG1/RJ0diew0Go/PHPzIhm87qNoF++Uhb3Cg79qnO+GQxzIwB+cmtqiQPGveCXPt5E5NAf3Xdyswb391nyzvi2dmiP8fTHpP/qeBycoONVOFZQd0q9UTP+TDaVRHGkMBFoHiStgmfq2ziMoS8G08QfefmG4jxaEC1EygzDPtO6Cv5p5vA2eyWwM/Uo5bU69W9MfjIyEA5vFCaqluif6Jm0wZkucvcMUC4TsHfMPCuwQnHlyLcVyy77VkUS3Ls1nnmsDTL6smvAvFn7qqHn7p2/GG2sxj9qhAVmdoJmmxBfJETm3UZ4IA5FhojUMpHVNxmpj3C6KYdCKYFxmw6gLV9aLg3UXmjew1BLTx+Jy+xkAkJ6qAwEF2/JyndlfMG1yozQFMNQWzqvmASHD7xOiQek6PlzKn1cYxBEkq3uen2vIGR5giflZrZ3qYmwBpAvsrvHM5O55iAd3XR1b6crDCoVI7OKcwy7z5EV/NApfeR2jkNRNfD7DPU9eSHos9jKZ7qFQIiV4XtiNUs2Q8CeAB8GGbaJnKQTi0Z7fAtwUO4MTp/qABTR3Ts/KWSHN2NYoqC0HLKJ90lhOu7wx3TXMtcF1as2RapMisBcIFKL66b/7q0ovuEEjTpLn0VZhdhYPofRopTXfZSF2pOTCywKgbkRkyVZ41bC3Dn7Vc81Mlhtm4xdwTCyMC3Fw+B6m6zqeD0Xrppc8FXnQSVPm5TKpU1/4OnHxLntD+D5kFfPu9gGnSBY4ohveJsoKOEAlR5l7dfM7ER2D6clFYCKB1KlFTil29OfYnhLBcUfFINAHD2AjWyfMMoWkWQ5lpNr9fYGZoIuXn4LWTLDAeoC5OUn107UN1hbdvkrH7ujvu05W1PUF4v00svKSwKehq82r1QKsKbBA/4d3XRv5m18gDyK8oYmxkjwfZRu9q6ErHuiKLjZYTxVc1a/pIN8y4Qrj3OgZaDcskrPBr0KDwRFyMQh7mCqgzYtS4T8PfXrQ6RPMxbPTFZxGt50CDAjH3AE0naAx2mR9prtAh4zsxjdjkiP+r5NXOaQmjINmugwR8HAVbYnaKsJhq7CsfinaNKTCYEhspU9hQyi6aAtZKF7NMoK27QZf7A5AhQgBdn6Ma3bI3bUYeQ4555ZkBJjBLpWmye+g79KKnk/ceH1JTX++C8EfAp9UIRU9/YdBwMeBtKQopKPdCZIrQTYF2jubJHcnrmHKIef8KZgL6nfDXmX1Trf/twU1elUVk+KK2hro04OiC/cy4hAQbRbt2OoLWwmscXp+Tj5Eril/Y+EIM0zcSKYuQD8hNDShYt/rn8EjMTrKFxC9ZvzEaYz6LwM9rZUDJHeVrdB8gwtnSKyb95YajuO8icB2xXyYLmdQBRvKSujKR8R/9bO0d2TwbgHTO6idS1/Cy6lwkwE2sXjlIl1q6Mm6je+AnwC40qWc/0cjJqb2eJBPlADlB2qW68iZ1QQgJiwSoCyeOTd/0uVD9BElJblmszpNMa+xQXc2XNNPiKTY1sqwo5WCQCe6Tj6a+y92e+vIk0YrmS2lqONm+GG274/Q8C6/RCqnClsOO+cEEKzcZ6iJJAML5U+x3tOOuiIIZ/6UgRwEhrD5h4NSdG2z2pA3l+sfgI50Vk7waMs7G5VeW4gspKLJMPVGhQ0e9KxBzl7cqmE2SugT/6J8tLCcE4bVe1ddEwevT8zfdxzNhL44rVRPi1vl1zPHzleFIUaQa57lvB4luU2DVeVnTM+gm+B4VIQP2NH1EiasC+JaV73KTrSuCQ9Od6XMjL3Jkd18TiueOHute8DIPhcG6NUrTCT+zxOy70LU7wH0v04pCtq1RX46/I9Z40KRHZh9KDlFUZEKduRd8J/RCyGMYUbD/LX1No52Pln2ic/4fqyqxHlolem1CUAiW0bNnz5FU3a5ucW7Gw56/Yc/G8UpRdkRYd3oFunIDyh9jKKpk8onnX05O2rpB/xSLqsD7G0d1L595wcNXWJdtEclzXKy/7sfjeiyFzQ6NMqU7T7DWxDekvkuJF1S6Y1Rrcqbq0DZG7CSB+1T3zRXOm3zRN5KbvTN5TOS1kJdWpPK+PfIV7w+BNVM1DqImhRCKQDaVrO6DygCyvIR3xpkxkIVrbD07wWsnkeWa3N3wAiyZWAi2vqYhfgumUp8JZDwdwcXJZeqGT4GqlK6t46ummga/0DfEedPsR8PCYm4Oui0TgcabIHX1SN/4Sor1AF4JqWNnQJNT+R8HmNUDwFo1TqqUKHiSIoELHJL50rljvN0j45x6QZpjPbQk1qpiN3+B2zZ1sWH/ZTaEvM+YDQJvHgzKaO1oQ64/nj9TG3ZIyBrgIvssuY1iErucCOhNjwz9+TuAvGKx0Hj+zJ0J+/x9Zx4EAyQTp+k0sJwXap9oq6JsyuE7bIUwO3XYqCXg6ZilLvdYxjz7B4bp5uViMo9mvfv7mVk+5zhBLAatit/PSzXSvgD2JYhUU5bijM0PQmBRDAis2oaWaoWbRyjgkhknk31X9YGRd2SGPHaYs0/cBw2arviMZweSK+sHEk9ihCTcQectIIpvibIAW1WIeu8eNu776CKYXa9z5b3G37R4/dZ5/Y9h50yGN4N4tjYfK2KyxVZq/sdNwLajFMQHoa6ZMfqjmEvMI16/ir5gwmLMSpxWWTh0YL98XAhKgbprvx8CdwtGWQqZO57auP/ENzmE0bC9ndduGg+BFaSd0HpAEXB9xsU72iAAWplKCRFWQcxJmqmDzMa+txB3GP3deyG5kHYVBQDMamy/GWfi1gjFdFboZCsITbFoYQwpAiQsaqgzF2SWcnPdWigKP5L2uKLCErxaQxRdFw/gbxfJo3Nx7HQnUi1+H8HsqjeCnQgTFRzBh3e9nvlsXcnlSjf2QGt8ZdxwZiZoL7Crgky9O7trL+YJIgmtjz+mLj8Ty85rPaS9vAEl1Ct+woDcWLFB4EEBO9GsRircNSD1v4dmvrFKfzZ4yQbc4OMUGujiWymfWJYwkzkJT81iWlh3Ow7fAoh1unl5/CObcdtzjYQlLFqYzcpaMMiQflos6FsdjFtK+XJo8sqC//RLp44GxvGAYAj40x7iEwkZCMjz3ryZOQWh6pHLKDhaV8M0/mccvNCc1fMvyTGdFQPLTr5H2MUJSL+RvF5fzFF9HQaZbLYNmNBmKP6XWhQVzQiUCrY2EeUXKrDXXO8yzvel2ZhjBhAKsMv7UTeIyuGpI1PQw/nxbBrF4X9yegjwPi8xA/cyHY2Psv73gV0ktXNdNxg2vTUwkZvLWSqWFW1RPUAcAsZEhgocgeeJZBfUMFjvZInZpGn65Ptuchot1oG2ae+6WcfmoDRNhdB8P0iWMN4i19njdIty2yjzKFCOJh97EJiElGitLoPVCoZJ4nE2gL88NmTAG6kTUNFMXCLfTVoTxLiWdC4xJ5gDNbegtd8dROWsjzv3m2tJR0KBLxUEFapdNhBsl7GqN7JCNxfJMTKybS3p3G2agFkp5VvSJTkmsP4rFqVrA/cdbg25oEDs0ZIxVg0TFWJ6d73jhLDA9w2IrviJSHKmnzwxvdnJAlDs19BMOC21vW/lt7WpyOyrul0ebNTjIxhb0WNTmG/OLIV1SkXHdUZph2IcFl7YaL7T1EecC/Rd67WXeG1Dm313cX9A2n31e/PNWQafwI64SH2LC+qYkz9Pg6+T8a1EiZ2cGizOVNTNjWtxPxwq8bL9Dt+s/862UFWJrTEr2ng4XOw76LdZxhWpvE4Q8wKgGv5HxreUZr8LDWtYLhGtzIjOuH6SeqMd7jzVt+VnIyRi9FlBg4Xx7SlipNoF9n0KOOjP6SS88VdQJAU69ywWERCB1+mJJcy/EaFnFVewlOuTfWtzeTijnijTq8aiN3Bu/rPzxOt1V27qPhSt1pteKy4IWoBkVcx4g3HrfZBzZ3YW3/XDRhRYQ6nL4Sp8wV18HDJu6LWl0MNP6T9/cQZorCUrEkZbhFGz3Xi6ThexlkeFr4m1tRcHLNLAmiZJS6R9/ncO+t6JkU0EzaqH08k3Z5RCJyUW+EXWPTem5/Hu+QPbbYIWJyrDyLm2FCdVIjUnF5t9LKVHyerTg+v0SYYbJwPvj+q9vVirbwc38N26T9OBKGsVdYVwCeWb7BJDJw1Pvk3ddKf+tmIMhaKVldUAEOyU52ce5aUTZIdQ611Wtu/1THZiOIXUlvrcODlV68Bdi/HQSWoVVrF1bfsPtgCBM+HLwWOMzVR2NXy0BPPacJ71Xgb5I2maZKqGv85aALjUIIe58VAieJzWXUDOsdRroznKudJfT9JbmOq1F7MevrT61g9TydzwuSGraOz5W7dagBRHjLM4vGgoUt+mCJt1ZNNWjbCHH4wzr7E4PnpeuGzGPs2j1zb2cR9j/2KWHmwSilSHJEhKBUs0BUBi/omecBpwILzd9druynQq81dxUwISgVFPL7pCWJic1pJoltvTbe7gD9TGJQmxk3lGuzzaOn4ZxVtOJlE5x20J+pzeSycrMYYPkhCDst7S/XXjuXS6HCXsYmlOTClCxW3Ir4SKU+wVLFh0wn/g7Kkz5m5OM5efrF87WV7zOT9r7reiH7LRMNX2u5zMVUbWR8AAHHsmyZRFwtwLEDDs61dWSm8eZ8FB/YRfXjEFFI5qPYDSH9LzdfBb79w1O/KxhYfk3tBw8GFVvqj2R1ZK+ZaPlFLzo5q/rFc9NHnrTmNVDWxHem8mKMjO9YtZNliQhLUH8chyp61uJyAR/cX+afZho5jNhEJhG9dNA2qNOdID3SB7OGp9VoBjJ76ClRWb9ADgUifnfTJ4wZMFEqj88HBybIeHrgyUJonjMU2BXBTlgSJCKs+jQTxULxBt1LNM5vVxZnqIYtv6ilEaN2k8ip+VYbumgbSNA4huTI6OhPRQaQi+HTko77EfwPpCexFOhx8J450pCzS3dbEkaAaKIN+XlY1j5Bkcdv3o/9MXe3Ak4L/o+WcDQbPKmRrLxVMKrkgfdvGCH12gcoqsrb95sQ9pZSQZAmIvc9DnP6vLRV557Hslz5W7pqOocy2HAacWwqALOfO9FmGxQfj2wodN0a1UcoY6a7D3P9wZnxnt4CDdFzIrrB1H2QFHJzFbTSEFfmkxZhiEvz99dUASY4xSPR02vRCE1O6+Hz6PRpkGerFcebP9f3PO94BZj0Ql57YDktLcPRdwrpPGffM8npGQjXjBsK4tyLZPI0awmMwiWrnQD24puQ++ulEtADnOZqGmgMOFUw+NkP+crSmSX8Dfy5QFmxECSt4s4iNL/1FRwv6rwZQlhesKFzrZrJeT06/kwkqUkt6oU8YgTVRzl76EKMl40xvII+FhyvHI/xkZPgDHsZXGUkRiN4icEgoatoGRb4P4TCDK2XbCmK7/mu7MGnnPdS5ytnI8z0nwAFJEjtMSPhAo17uyuwgE/rGnq1PwwNuImh3dNU04zupT1GftaWAHr5FduLivKihC56NRvpfL9wHA34jE74oUq4uUwvk4c0uIV2p6IOKZWIiHtA0vSRDepdwOo+sPyRQkZ1PkvaHhJK0H+L4dQ+PnkhOvhmp5WF9nEj8oBPDSVHuxNTHpF5c5P0gt6vRrH2gU23uX9Swn4Xm8uICy6WqsGjGHCXOgrS95z5b/CVhXim/YYkHPfDJz6ow9P9X576GR4HhLmZcuGZOPDIKjJ08c1yvym8aH9olqwB0EOARIUCgtXDlwdPPVg40jt6dO0RQiGbWB5O75kaTAn2UxiyVI7iV48Y3UR9I4x9rsa8vXWAGVLsDNBBbMxCy2Zk3UK6ANwUFiU+hkQk5PttH1QS7soLbFVYBuhmBBrIQajPJ1lEhcVuhzICOIETXSzqPufyxfLniOqXG6ocXPHmih+IIaFYxmrwPdRT8uinE3v7d5m8aHaVdT/+dhkDccN+kTEVcETmVdvCWmdh2XCxeKNud4fhhmd5bM1nfMY4NsHulHcGa9JYYPsoTd0Pi6LNfl+BbROkO8hx+zQsMFh5WbU+pQMdpSUP68P6m3jLWMxHLsjoQ87oQyRkEDoRe+U2NeC3qZj1OnCzU8ELZdB9XTbNd0VCsX3Ugs2Aci754LmaIHibxZ/SDBORXnFQY0XzS7hjLggCVivfq5IVsbP2BgHnX6bECmOZVdPJpj/aME8FNieugn4TX+NgGmIY/QcbmRMnpYafScYAoiNwKwgDz/NPqos1p+rqPxKQ8L4/nXV6edkK3Aft+ULfI3VGnqV/00ngnlpTFCyXV211Z7v7ZJ/BnY+QzpH1VCH79Q5WUtLiFx7qsYhxrZS4VlWoHdSJlsfjY8z4Wvv27Hr8+0opCVvw5TllRisQNIsyVBxNXzGob3hjY2HRM40E5N7guaMQM/L7aa4TMU639IGCgwg3nF+SSeFVMVTgu+x4zZBy+QDn1/xkT+1sZxcZkXdXw7/+jnYCv48GqODSgfVD/cMWHm5i6gQxKZPPhiQRs+qwCiIoq34C9fcV7GV/qBCespXehJa64DMO9kTFYjoLPFCRCDI+Aq+xRByJCVqEDrQmxRihgur9mIIxKMTc2r30FBa7tZY6vOG37naQJfgI+oQ05IMp7WWT+Rm04aPrWudNS6r2oclNhwrjkbfxJ22ubCKMmcRHJ1Eu/+3jW/g4BnwZ5WtQYO64N0VwM5htvxVFMu6zFv6jeGi/0vaObAqZhBygVvnZWRYiYQ3Lpf9BSyLKwM6wRM2D3DV503oX0RcwT9j4kZUVictxoDtvEVj96nSmZQInHWn0rgG1Q0t5RIU0TVdfIJFeXODc4Tuym3vu2osUSIpcax1rzZhMwkAe3qZSPsLxB1Esv/UEmd68rhZPvda/0l8AVyKAu21/v7qHBC0IgdaQDTwXemnEJCEnFG7+a5NPNr3si6FN6BSUvLA1yj2AEKx/AUkqg87Jf7O76A/NZFJXS8svliN1gDgxVAjV1NMVW8JtX//KuXBLYirD4EhSgw1YfS544P25XIRJUJEVgVLH4e1WVmViQCuLC6Zx7QWY+CfZHwlIwCibRKDd/xJxu9OPP9LiGUrES1Y4sht496/5X6Fg/0NCC0x1DI8zvzFeAll6rOyU2//EmSBqLqdATnYbaB41VeVhCTvj7jPBnTCmHhBEyUvtOfZjpjW1cZbUZ/im1X6EyTxnnSUj7MvwGUA4NSVRzKQjTqqAh66nIxAO5QZ5tBWlULv6Uo84phcw1o2mbfVG3JByPywooOgULuBQac+g9nqyvV0Fwq4Wyuuo1wKG4GbYtNea4JANawYWKwjNPDw+DC9IZaL1T10XOGvOdAM+IysCqhMmZXgfL/3F0yl7eiOs9oxMf24mSMUhg6LP5t2dN2cvmNU5jiMN/o9yJMTlg5EKiFWbxk5ISNI1JOKNDBEPm8wsOsNYI51etOz2G7d/p9wrfkvJCnHibviNFcwvKf3KX8zgPkvAGVT1InRSKkaWa7DgNwAlSJ/bj/iVRW5ILBiVw0swT/ivnzlvrbhP4NREqol/IF+7bBudGCpZvNN8ERS8jXqNa0n60XlnlnsUfZKw1kEKRdNpAp4Y072Fs0/m9v/NrnJqqyu6DzhR6XE0EX4Th30JUJ0NPrGIpcamiP6lxGMmbOEQVzfPRtqkYXt+rxfZvhRvTYwFfghDnkmM8cS+FKJf9nXvzzJQrfAHD3y4mADUGjpexq95EkE/o1ylINfkL2YX3VYmgy4s1moKeNwqLLQTzF+UPhaUg2HHd600GTj5SJR7Fkvq84D2B+g7Ptu8kuIbVgMvQtpgEbdEJa3TyxAjWqnd3MU8LsMUtNNjL5KhHunxoVluiuoyBiPuM74ZHO+AZX55nOcISJ2xDWoYOlXbjv5nQ7wKm90MdgbqahitIkGLQNYT2RsQiHbwqgtT+4lma476QNBDFFL7huTLCFOX+yuEjBXO5fx4W7hxfi7yQ75xjcuvdw7l8ekTv1PyMvY+mnQRCSRe1gSrADztP9XOXm1UnkW0IOKs5XSKDMRKlzB9oE3mZdKNeK/Eau/v6eWsTzZNdXsryIn5pYhKqNv8wEbIUVd1KaBQrYJdWujx4XmqUbX0wmVMgphiLmTGIfe1wAZRocyrnizBqiXTYi3BO607Mvrn60ITTaQci3h0RBHAT3hZdL+pb7L3CCKuhh6qALMmPL1KDUKWumsOsU/I7JhBh8dewhWFBcKUHT2uSIo0kJMnxXYkmYZZjlO+ERgF5C4hopBhDjWG60zFqsM10xoENxjOhm/8PB5kYy3dU9Tpb3zc8wMjuSxy0qdRhUkD2m31sKz1pQMdss03Ks3G6hvcy6KT3lM0p5eQ5ROJXOwazG+xZjYFxNUmNkEB4pASXobxmYkbiM3H3MCMcCV5HF/2Peg4wgBt6HDY5jDYMzEbF36QN9BEJS9/d9kT6kFbF3QhmaJoOiJPPShEdArxP27em00LK8fdGs8/p5vfG7y4TY7cOMxLdkOwkoDnBxepPwnrrbpLJ4fMSt86Wu/BD7W2p+JVkcaeJq3thMIIA+yEK/SJ0xP69rgMWSQVKVaw9eB7I9dVIJJ7sLeFfP2OQDa0Pzd/kJeHsGQljwh5W8NJXuYOcQxXB38wT9m37zBSgXSqBugPvFIgRIgJp697DAocxRrYrkdj1SaazbsyUHSZpuyOpk50FNxfY3eCUcptE6xZ1VQLgme57GuSTlHdgOOTO4aYdUHqUztZLks/0HwqdDkO5xlxjcQqGHCBHb8lREDH08FAOm9ouK03mLzWYGTxgEybnCzhjz86fD5WqZNeadTlAvhRkZIdOhwSpjLvZf+ZcDAnby2YgpwKkY5tu5+WX0mrdq23GlXsXmNgM6TGe4Avi78bx2BMIRoUjSam6kXRzLmPvY2CFWb0tfDmJVRmOTMWLUJZ/JHy2xZFEMdEUZmpna3IkGGwFX58baZvPAWIja9lzXvuEo+QK5B2BZzg8Y4/Fypu7QHaVJTRCVzSek0wcixRN0SoX3H1czIxbr13e6+hxO5/S60G3r9LjZiH2f3Zykty9EnD14P30V73q5MfwtDh+Mo7TSPIjqbUNk1YGWgiiWmkYzx2G+C/mRyUb12sIkdYDgZFPF+zF96B1cwYJhrMx+zcmHJRCCVtNCK49KGvffZcQIZ9vJZ7zwQ/Ai5cGX6lpnoJiyW9EQGdPIiwxW/xEQCtVfH9pOvKyODXAnnYX6CadZMIovx9TTs29dDexvC+p/N3P0hR0gL8WrcxDd3uld5usFobqgsW3tSstVkXRDcXnFzxHxRcKp9YjhUg49sS9B57yNezXaHQwPCmA2K6bCGCDBXiCegVw963ARbexLvv8DEXJt+6Oy7Sep6HM5KEZF4YZO2olgIrOfoAZX3IIuUethA7JMPb7MoRWqZSFHuENQH0SD22djgwJkWBYIvJfGEHGsgr/fxi4TdBS9qu9MS7TJHuUZnBQg3u6HX9J50JTVAE4LRNr07/JKFVUS8JvL1vsNqLlmTmG1e7eYBk1h1J64ABHBQf3/WYdb6ktXChLW1A0Ur90TZjgzmUKyKE4X25TmbqvPz2ezY5PeGFRnYbd3WwddHveasNHSq0lX9AF/p6MJhX7BpmKdM/wev2rlTKKUajleMPaK46Q2uvFndAu5mHq3s17AOfaW4pEsHSA9cEFZIy/Q0dd3+0HBJApbAr1jpTq1B0PYq9hCxCAgYoRr954vd0xtutrFrSDUpO2oZp2ZYZo3OlbXpe+OwQnsSOxD5Hs0PB6ktC9RwO1Okqb1eirdp098hzzGaPST3vJUmAyercu1JZnAHLdeR0ppDCadam+My+wNCZlZyhGR4bWtQrJedlSwxUGs9nL+ji9mvYZbzNcGqAeNQ+b3m7ihu1ZBgC/hJs5ragwcPC6tTL/c0ia/8eG8Hafe19a2ldO8/QrRTEIo0aHNOAG+Jxs1RVn+weOnN54TfqNBqJ6HgiSY1QYQmQfai1kz51Nx5Zqt4178fKMiTRm0NufR61W/Zphz7UwOVQy7eCywAkO4Y9Dv7HPx6x7BjU/wL6G2IEoHLUaSDLIyypFabixKerDHv0tnOoE9WY5fGqADSsSt4QJaADSNgLoeFKx2eyeLx3d1xkS5S5aZvJdBRfRMbClRbzDrn/UhDvPflIGcSxYumjaBA5+clgSU8FZQV5myvqVn3BQoyNWQSGCqSpRFMzsTEidOK+Qey4vBYGci2ACkQAKp5CnhoCldexr9q/h9EyrI5qkkxzQ4stGgHhRHI1VNxhf5NfhiCj+kx3qBt6b2q+HNFUurikaV76LeAwLkMP6Wa73Nm3j8fIR8UQzHlw+SIBRQsGAjbNmWfk375ku0kt3CWzLfZZFeFrFafup0D5P0VKgd/KeLLIbo+T31zkFucmSnPqdHokHUPKue6KcskA3R6kGIEISipQ/kp/+bsu7IGU/+Riol9fkWn6nIJa1liHBpQLCL1GRau2m0Vr3jJL+jrQ589EibcFCEsGtGnullJG5l/iue0Y5EtXZf2Q+TB8cmM+XC3KiqlXdd8g9rZws7QhvRQ093UQXTRrhY8NvWhT44RxGOmW4C4tMikmwVEsr/yvXxuft/n2hhlWLUE7Hqa2r8K1cmkT4Ad1FEFtoMHs2BfTjIn1u4PmQPSdrW9EaawrGS6Sc6FIIVKfnQHfT8W9NjkmUbQTrGHM9Jjn3LUF162IYbg6DmZWYm7U8UC5ZJtxwUaqYx2HCsMH3RSVtaoq7gSN4+HTmwYVIQKj/Q/tN06SvvlMORaVDrDeAYDC73aGtGUTm4LOGga3GhQcQ2TnoFdV2G1cemw2dqAJu/ZyYyK5dm0uH7hqRwGYPQOjMly23vTEE+YZPjyHK4U9j/hLDjUewW0jtqvL1oaoZ7PAWP1KHFKkRUwwLqhUy5y2o9e8/svzeKRiOKXUPT4LHAXGTwSOefD8OdVqmAfV1ydjB6zicMVzJal1S+YjTxoASNOoEF+QbH5GrOAtVjm4AND1+9gSc9XGvSGMPYPt192hjPGwG6TAY/IX5H+T7Y8yvLyBR7aRx6YnWXGoKAqfQV3WgFU2BS6FkOkScJ0LWUQbSapyzAGHjRK1BgtmlBGqSFR/1hzjP+PdKs9S+LBxtDPUjRi1O41JS7u8jOlvrZ9dWUL9rUe+3H1GHvIWl/7KmI7d2cKG0UVisvhy/bHsQf71sbQazaq4kYY/d3El2m+YAX6cIXOmB0xVKm4LGC2ZKVKTGqcTRlZIEawf8zT9OvMpf0AmrucBlnNWNTcaBkY6YrcGTVfMt90raUJfG/teIWI8dsz+HPahxHnszyz2pxADDkmXaSXcmAhrnirOYK4d2m0Gt2I+rNt1+SliHSVNgXeJ5R+l/V9FXQbnLYQWU0+ALcNrlpZSqoDvYO6x7BUQghXVM0WOBmBeLoz61SxmYk76MMT4RtSoZykVcqI+utvbBU3zGaQtS78nOF29yIIRdo8W3xqtA+U2chpOamuj+0jstgXRD7XVCE7Yxr/fo/3Y0fQQB+vgMw8N/qqmiPWPx83jnNx4sEscPc0ITPsGp8R2JuxXHKxJarRfO91jieopjHxMMtRzcb6hsITlZ/l8Ur+io1ffqUCOaGHpIdItkZBkKaqsvWk4jGRM0JzM04zf97JxgYtCTQMGPz75IGe/bCHuStPTBa4li1YLME/lsZeO60i4pyiZoeYK66yR3lMsgUD9UjQPKGt3KabiMPo3CJUGhuLu8UuoRHsrqK6+4BJJpimQG16B+PTWq7T66ZbfBMTiCAPFtOUozPKiEzjC6twtuvxK+sDPXER8WD/fIdzL+fItlDVItWV69K3G+i9qOuJHQSNjXRYUrY1quYO8jItijvk+9w8+wQZ3Yq8hh1scHmD4TLMnHmDVopcNNQ1zCMs31SwkXLagp/AYgbgdkkB55wudYiwORflRgOh7naNTmueKwlc2VR+PSpXvT1tx1snAtvF4KXsPM93ZCbUx6E7O+7fplp4Vua7Hm61AklGOq4AED5pCHmDvFfJF/jX8pDLxkGoDIoA7bGt9ILmZoR4n+A9PUsBLAlit0mKgFtIcUJcZPkvc589M6TvV4jhyx/wnW7ObpBZRVM9hg9uF7e0oJQIopM2PjaKq5jqoIsZuMFPNaBhW2xYf5VnnY2JOBC2ZKnYBy9MwlzmL+Wv9WYT/YTuY0tFT2EcTQDIZDCnWEsh1t/akQ+ujKz4RlMmyheYbN1JqUY/SHsug6Tqr4WjwRsOjMH6P8aOo6ciPtT8t1KO/sQ9dgJP64fkRpv74hv/6kK8lCXecIIvohaaRPZ7B8lOADdCC1uxrVLksu/y6cjcPeUtJKQhBVjX8YnLVpvK0KUdhKDXI3XVKuVq3aO+6TzJCz39jo1xYTfjcaX04Kaoh70JygoE2haBDoHt8SKZ11VqEUZ+cYRrM/zp93pUiCWSeb9QwisFQhgo5TNzT2JaLLTP2uo3D/VqMhf+TjWQVSKcbjDZgyhdaFSlu5ksA2zXky5O9v87Xvl1Q1wAJAejx7qK0P/Xb+v9aIB+IrlDatCt3HCj9QJjUvxY5pldJI74qyVBQHD5gFo8LOhIw5nzALd2vtHPGbWiolWlI5ckBzAQsTd8GNydb83CEaeKQ0YnRo9O1DdIBhyb12z2f3NDkBSBta20fLRy/WAkd9xiDOYSn9RwmlVPJu01aosebcSw8fvmZsIwNRXN7TIR9bmlFWeUVqyRWphzW3GcvheKdizsY9d3TsRjRKxSiLs3wKY+LgQHYg54n5HX7T2ozFGVE/pGtUFOD5fygywYQWs4bvIaLrrx9Yn7DHkzE97vX0a7lQK0TczHVL3V4Tky4XCRSZpyBZ7Nrq7ifU/v3MUfgNgBVWV744hhl3s3GlLqedWCQyIrlH12he6YeuMp3aNJwUBlj3RZhMoGawTJLs1QtiSJ7PfmFMhsBnt9b9QLLaw6EZSt2NktNBoDX5UAmtY79rVtEtTRWwj7AtQMZ47MzIFnk2CAk049JEyRqZ0p7z8wo1VlYMLLdqcUi+CEpCxld8ZWNtoOaEfafMA3SSYRdNIBk2E85lRJviJrys08jYiKalG8kpxOuZP1YsWeCZT/0IXreHXSk7BFv1nO3Pkx+xoMAULRve1CuqLS2TmuDrRt9Am+OXiOB9raul6odr9s9Jfw4EwNW1B5BxJpHVokKm+J15CSclHmnAf2/Iq6hjQlgavKrArZGRltUZ6Z84ssV3xqC3nVeINWn2KOz2za+H6ckXL+JooAY2PNXXZSp6uio6t65Tpf18R7jV8Jtbv+LJg2KFxNnSzAnilRnU/2ekH3N0KMEVjbheqC+jh7Xu31zDP1psJ4BCKIVKZLW1TQeReqNHhYKSWLn5Vmgeds57UBl0k/+988w914tMBw4yz0qKK1QeR111GFyrpEytJppr498xYfdU9+wuxGX8hGwf/HaN0O8eKTLI5ei9wpsUVwQFS04NjET9374QAuAhDYJTMT+VqxSBq7SmAVuXSVb+R8L4BVpLzzbnjnFcSzO4U/mzanqNJP9JYC56iNEh3K1LT2lsS14hIVUOBeAGaMfVJgGTkiP9p4a1gFEfTKgbGun2JH3QyQAZPZu0EL8WzDpCuBUmN8AGtrfmpUpnwSfb2fBt2Rc/lTz4o+GB5rf0jQ9m1lMF+if/U+k4YE3/XMymb8kxTGkRsArie75QL+ogqJ5cpgaGbMbjASEefMyght1ghj7SLct4vupq4OEfK8uehlicirpAad++i//q1eUxeacSn1gWfY7ye15FBUIU1hNV5j/HNU7sMvyoeb+R6apBdFKbq7I4tUfIjmtWkdHC/p0WYUyM20SjaDHORSxRGLh8KBcVRyCh86INFMLNL1HXkyVdWyf2NLQ54+kA7MCuxsBUAp6l2kwr3IES/XEhazOY0OzCNvnvEcBy7OPXAg2kxevqrZgEx4Qig6ipOd0kOzHMlHyZVsVAxqVtOVq+lAM1Fxh3NMjNEOLAmzCBvsYWUaAr3gROpCPLcs7H8ouf8W2DJFuwWjaSDj0HQiO8bRH/daNIrNALj4DJtX0EbubqzTQNIAT7bPBaX7+ujy0e94WodCjJGNWVVGx0c/4nnKYxhDFhWFZcaZ1yWo8q6XZ/yPj399cNv3BpkgCRyfz3IDGQ5+1qT80DKZFKk2ED4RxvHNVXZvjmsJ8J2eQHPHEeScUujZ3drU5l5yHuakNzS9SpR2riguQgRapEwfkEqU8d/QcqVBcTG7TPnSmpwHerviGkT2byf0PqbBHWf3dSjsB9NnvMgHKcy2EyG0pe3hrW+1fexO6oZtKYdpJ1Ecf7kutkVYcYOV4xYbFzYx5z5xu8bC5U31ySRBeCdwKJH51a4TeMrnuvtQON5C8T3k7VCmVyf7sIjYKlB357TwpeY2OO61/ieCFuHNwUmvD/vz0XG5WpFsc5sspj23Wf/e24deMzm3BFavtQDnnykTBXez0SbHBhEIoFC3b6V6cXGnRJSWCjvhRzEPPAssuQgIwb594k7Zcc73sKcswH68I9051HSOiodnbyTQklDu5Fo1RouybJQlbMKWqOlrxz580gXtI3TP03JnC9jAm4BNpaUn2lBO6fTASN8grcZlvl9dklz5fshr2gaqduNoj5RZ7tnKHfB8qkUIoa6QLAomOno7V6xh1WA9vCbx+fTcuEzPx+/U3pCzuWdkDaY8EwvAa6vEKWOY5UF2695q77qHVCHRHVFFq/Yj9BU95VDyL44olHeCj129CAXLyFNQTxUZ4f6X3NlxrYgc2EZinFS4pE42DB7be5Nvi8YNJ/PVz/dNG52EwPovH18wPk3/wBhg1y1CANAfriFjis4nM361P9AeigO/ho/YCzX3urL6a1FrPCgaDB8SuY/NLQ+AX6j8jt9QZt7/0k51H2SODIcprETEiq8SG6ELZFTc68QGM8xANjcrusPKOy4Gid6KB1RlzsSeg3nmj8jex2nKfOf49olJGxY61lTVS6V48aoiyJ9jOP83hwwZg3vitLPBlNfqTYwaO6CRIM8aofgu48iTn+c4gQnPIj6NmrWbK5sJncHtUMIBoZ0PFyIQS5bJwOo6dw4f825aNGF1KA9p0zkl4GFoLUsvPwvRUDJiIKgJEYDMLsTcqTPxeUzWRJo3Fz5v6wf+9woy18pTFn4BXvTFhlpjeJBtvYofJbju4gjDPe1j4jhPR76sJQRNb9WEotqQ71QSCNGi4ELbxKttKd29y2BxaNU2B8sJfwScKigOK5IiikvrV/tbFw8Ge+PGUCd9+vxyYRf+M7rmFeHXrpbbL3X8bWGYJNz95ovsfHERFkzY4dHof9dWu7708jl23xwiJOKnAYOO16IBfg3T/gzIuFpDvD4A4bnvsFyQXiUupK2pZ1iDfr/hv2vl/dAC12z/XWrmAL15s+ffdp7VHM9W26QQj/epkZQVzbEsTM+qNemb+YMll9ojVGNeAK8hRpjvCJpuwLHlvv3lPzx46LaQBU/SYF4eTn+cOYvKMHE86kiuf4QjEaJutjx06bmvFBjbDti0w5fMmH9W55U8iTj79pwJohFv8IevJGlT2ma+lYk5j1KH7bbK/pAbs5DMmizWu2H8+zpYRc4Amz9ugQ9lS985CP8mAPeUEE4dsXC0Jh8iq5ytD6Pc775BxGrkKR7Pm4dpi76++kcpQ5Lkn7knzMfMiDfKBqARkD4Ozxa6svBEIzZKVkrnwX+deaASPU+ysg5sJnWUh28EDnmUCs8VbQQ3ei/DlE3MWNTQgjQqtfgoX1f+P/TCgrhZa8zk2QMiH/f3JE/bxCLI1VD9pKE74C5gUg+/P57nLYHas13nhlonZB75MjfrqKOtMWpb1UEv9OvhmtnOxNCFXXEdogznOBzeedZrnMdzX5C1GoEfE5UaGdDAJsLmICgOhg/IkF+yKtN2kyHujDXwI9UWEV/3ddiekjlx1oyl1dtbdc6O2GMvsIUpPd1iobVujf7W+mJa4GrnH5Gd/kmrboVfzAC2FvyQ8BKdVOMK8piyDgkfCdsZu3rPp0Hd5VPpDwS8oG/ELnuLq2vDwarPEr0iVpbzY28wDpFOtED35S3IQ92E5AWy1isvmpO8zNRRYOuMmsPI2spk0inh8dMMSb8fGfIOy8iX1Be8isSUPPTT3GvLg13sB7a7hUl2CZ9wZFVPqeQe24BVOgHMlSBaz7S+V0Snzt9x+GlBto6LsRQ3bEsyVnegWpAq9GkgeSzFlH4UPtI36x+R0AbUGs4Toj0HTxlE5rLIGHqV5KSa1DpARbXtvbqPLxKw3P3v3HRKmoN390LT+7QUcQYGW+TTj7QjjvahKGlaBf9ryTNFx7jDzO/NqjXNewsqaTuJe0FtWUMIwBvQNoemvV1lzXD3Yq0yNRLkPkUapS4Z+pU1MlHxkzhaoLGNW3TCuyOq7KJXg0XF/bUrMqn7NxQlhFVnymPRKJUChxsxTQTslOwJJCeew5r+tbKaKohr5eLriPCteYap8TO3mz1Ut+8BK4VqSciMuDSmirnI14ADsYlUbCdQ/0Mx51tval7qKr8J1vMUq34YheoJpRHBheKDPekB2neD6RQ0d6FmFmvEo3Lc0bvhURwEqsVFjwowaYIzDueGHJLCC2LDVQH057fELrHCEIIlXukUzYXpUaUcedmtqhijRrSCgwTLWD9MIdr0F+tSpd4UOxK12cd9Jm7tfChdZL8dbRBCXVnqCjWlxK3o2I2ckVVsEWaz9UjS24LLJs3axFrB97ay4QpMNzjR4HisemtfOKJ27MQrhJmARNt9GdfwSgZBeIcGx2QCkHevkCElYyyhf3X/M3HYa88+UwX8ww37xoq41R0LbT2MSJ604h8Mq+T3Zy13/tkyGpfv/Vfz6sw5f/uESneE3Wevr1joCqPaIDWhk/qIAgktl1zOIMrzxaeuZM4MwI0d3Wg55R26cL5N3dvOgymM//dnZGzuuwj2eySz0ABmyyu/M+fH6r+aHot/r46+L1oneZ1+DJb4SG4yy4DxW/97gT86OO56Qfs08puqK5riyTyVmXNUl8cQlqi2Oq0KK34kbcFq2QRdKVAi6LB7kfjFt3jBJ75JIt7saHtr8DMHBjfisHKxhksIi77YOmdVtc+M0AaUHmg4U5LA8Yuwy3En0cgcjjv+eH7mSGkMRG1KzAG9e8tOeKrUQGsxpzthBuni2iEStRCYv4rIQColfQ873pcnb6josrjA7kKK90FkgE4g3tZZY9A/CvuPKFQ9rbxqaYHiYBJrcuuABRjG9lco02GDMToWiIZ018/ReeSKDXcw4fVAijZi5LTbL/kOJNi1ecFhOtpkb++E2/4a2RLEENVEBekWHJJH77SVbHARceRJ+ASL8inPd0y66pvlnwoY8jR+gXg2aEfdEdZ2FGO7uKBRV3vZoa6NLiNvflTiiMM4TQYqApBX06cv0Px9vlNd3lEYYw0hS1/4xD6r8eI0VV8oL3H+JXm9OMYf0jiDgIjIBZ/FreDpwZFcuGi101g+iLS3WDJQMcwfPP3hEH1Msa7J7GHxVrgr9XkwPAlSTjlJnpap4243WMA2eZv3edXK+H6e29Ez8d4P6RTwnKcoCVBGAo7OkWITitzfnINXaahBgjLkJ8s23BmwreeE+KsU1PkCnvZteJz1rm9UA0/ORIIZy+2ovYqHUGupU5Rjrnyv3QF846X3GjoH9XfdZrY79qNFuc0MP2xBxX++SOgZdC3tMzCUsMNv4BQx29Y4IweO82pzZRV56UWVWd8piyPKhbknBuRoOFS8fPNG7NQVrCPPbsQNrXJqqFGnDF8VZjleOikzx0jcR0zKwBDmR+d/3St/dbO3THsKk2qKA5QXpXKJi7+j9sa2Ib300Jc7NKA625/NfQU3Q9R55sy/NW4stEnR+XtYpXabJBCGuH9d87Ciq44HvVeA6xFRxzdeIkUGKDBbaM0zz2EvA7o9JMiHuQu/9e6v0k9JjNndQyXsI+sNlucUmv3eA/WuKHsg0KVuaJ/9rZlAD6FeVnmvtePOj96civDmEeut3sT5RxKMqQztYzZ7YbPxIosgNntRLN5qf64PyE9tkA60sU8Y/HgNMNlYmauq1wif+p+2ea2lJLJYWAUqZ9St+nTNdpc1leqy9XYu36gqdaYgr9EnIzyacGaAp5vw4VNWT1pGu8jHwu592URro4RwQVgiF2HjwvxhI36W+Im8fWJ4A6K1bYFydQmtpWzuPx0sJcZm6UuhLIyICeSMKZOVsXrL9PLuEE5F1r990Q4a3vS9HyaBOk/EFT0++Im5CiGwjv5DrdDJozD39C3Tv6sgDCdc8iJURwaozFsIyw6aqIoSKxwatEOcj2so1Kr09Wrbj5xbgBxPgM2fpxFk786TlhN/7RR+Mba58NXjrBXN/ITap3gsknseFgBKx5zeyexCKReCqlempqCtVTy8pqX3Pifd1Ok3B+3ecW6Em0GGxfajALXW3Ikj4kcfczgVTMT/17lwAIQEDioYaJiwzX5JoJfm5Bb0pOaPC9F9vrcPF7Fh6XXU1INtZircpvczLIn/TNAtrpbHJ8ljccEow6KEmI8R2+vq+aMsGwTy0IfLP6+z6Sr4OT6ZZoXOUwXhlx5k7rpmcLqa+yMMFPoo3oLaKq9GLRrxfJTTVpn6wsdG0ReLA3jb/nzjJlvJOZVAh7eIIb6UWJJS7vYzd1l1sbXVz//8ZKvZL3ZEtQ/KTa4ERnvJwfLYmcRo9uZAiYeVs1pC/zWYXueC9GfwrqoIMsQjy/6MYcKahRKbGHRU3I4B4lomeJf51ZiR7GEn2WzGEas1bCDidiq9wxPBC5zIQTQnDpuwvPKg0g+N6BWytWFgwLEAxI1HLd4Bk46ikNwOYcM/lKdh7CVWSZHwhyuYSqnMsMpb0cs0YsrOu6kY4ri9Y02Q0gyl3B3xoDnaqC604r2xQpWqaRKRtLWOZSti5kOgmOFjmO1SIQJsi5MfgvVSnzYtLXetXCXu79Pr9qzTYRBrvoOPeTCgVDKV+NXnVg6UwD4uRICEL9q4zIiBCrpncibzMBO7jAulZk7Ke9n3m9eKnoNoz2puSnl63ujEdpoABlf+iFBvsi4XeUUUe60TszQ9v2BB3YIirPF/91nCe1iQ7tXH3kar22GvCQ799xW/EkE4rkW0E5WgBTw6Ehy0lpVHWcy6OvaDQUJEKYqP+okNhMYBV4cA+npoxEG8YkE9HjzXLg9I4H9aB3XLLiVh5lpGj9HwJ2ofYQHMZynzKPuQFkBwaxkQxCWucDUM2e11Ae4CmgBx6ntPI6NY15lHEOztsevTLp1S7eJFENhv5nzVcnjIV/TAia5UOFdvsuSwOOoc2tCTKetwX1CxHz5Tvrn7CCZDWIZzRw4TJS/0qrnGiLFyjGmJDm3TCw2WJRFoI/nr5MhKu0OEpc/p6dIWIkf4Q6BA1qpCYuXYlkp9J4CAONSUqpSmaQNe9vbGS3FI2qD41vTZs4ohU0dGd6MfEe+uY/Oz5fKlfuLF2CtpRAR4gKMXxC/YuDHBFs4mi501bWE24Anvt5MhW0X1VIG1h3y+sSe2ordZ7IMs7O6Csh9WEjEGUZZp9Th2WR2GGvsN5lg9y7jpwAFqwH12p1CmVUG4Ha/AeJ+6Yr6GumQZ2mT+apmsAIY27KboFZatwQD5kJWv/+M1IrcjyGVw3v7bTVBO/OWqQiQpHLItmZIT2IlZ3zQqQ8FznUJ7M6CMIIYhqyJaGAnArqiyq0MHPwuuyEZnXSu6MlahuQTijjJPFWwmphBY+L0Blz3R1Nl16THBqtoUNprkILS6CRe3kOf8pDgAcxKcfGPsWa5xbW+2dLjG5SBeB9TVriQhzgQ8a90dkhRjo1EdYsKiz316xl4T7TUR4PQehf/6KsJSuwDUJMkpk2ZSzb/+GutIjZMnXVeYRnAMUgPmaB6b5DLuGFLurKf+o/9SOraEaOWS8M6wfRN5vg09OM7YsSPH3Std25Y/QVEbKcsr/kzEFuvHxWCQ97g9DNGUgtUXXyREves1rG4VDremE517BVJXIlJKu5wn5HhJdVjdIcIZYt6liVhvl3WwFWd0/2B6/gPYFaeURDfrYSI63bpkiSOJw/P8DwdwW9Mt/lDcMbbpsdqYNMXf5DeUOyVP5GTu2C2HNCCi/UeS435cer0WwX5dhEVjgVFMyyBM0Ur/A+Wvu6P8neMv50Y+Wv7y2xmog9nEEWWNFjj+LHr5fMWB0TsJllsU6zo8cNqcGViSa2k3okbjas427eA7RbatNEP8J8aQosN95qxznSf5PlvS00bWPScs6FwdnqMrliU8DUcdtvqgR9oDtPA9L5HajAw6vHtrpLYQY5N1joGcu6Ez+XvJJ5dNj7p8/FoaXfxsT4Cn6FDkLz5iEyKTzjAZR355A4ockOf+AAmoyJmSzibpghdlbpflEB44w9WAGfnCTkzG5aFrAwXwlOSnvcuP0H/7PQh0FFKsSLMPN0kym+4+HMeBKGUxKX9QM9d6sdUz3vRD8iGH97a0Yr7uVNiHyZezbbVlEm21F2sJ8BJD5FszR71r+intC8MDhVGgqvYaYZfDmNwL0NjQPHsZ9nzahfchLKQNE7GQX+91F7p95mOgP2do1VKXKaFqD9zqUPR2aGyyIJGZHUG9Nbclmfv24Q7iKFJANwsK18Hr95/D/sX9NkuAucJOCMAhNzDzfrkZRo+MoaZCJs5Ol+c8733AzDThxRcxhvISj3NJBs8pKMS1Fb8PwwkWG/kar1rw5Qk7gYbsHIAwPXvA5HhLkPWHUV9CXkJoA4n9GT5AZto7GDpLH8qe7uwmdxf1jAahKK70ryWjjIj/K+nFTTVbRvtyNZuTX/j/ht6GP+wXP/tYB3ehToj8j8PCS2P2Aj8TFeSJiRpftjkPcTevposGS6k67NOB9KfVIG5kZrUPpm8SoqSofPxPnedxLJY1TytBR7dgwIJFOlJQEFzdE5RLrTCFCDAV9AoLGRI/aOs2FUh3wfJbsNTsRFQ7vwAtb+fVfdwwAlOEOgskC2tbmgarvoLcSWqvG36qJum/QjXGRp/Xc6BBfic6zLZXcIyWFCxklTSRlgXEq4wDtxLczgr5R7LiheRVtHCtxrO+2V0pF3H2YkrxWv89jiqCjX/VM/Pfz+Jw9PjUh6LI5pWGktTMabzMTfgDNP8qSASlBv4b7TqkYQjGd9aUHmw3wVm5fOf8WRCzrwReiPvIq/STDoPo9xEWKkrYiMoTHd5cp4SYNrhq3fdoZkwspt5b1buFlYzFs6kHCwfPg6IwBVk8xkjcYtMdy4vgfRUQPMJ0wP7BH2Fsras/emRLmwCNXRLHRQs70cZ/BXnyOLw6NE3zn6ZZju+NljeCQ9Ws8TaM6xhQLnasMb9y92OlbnPGO2GbDwLLLNFT/RTdm1koX/1sog1/1i3zll4QAMQpLjQDJbj5rO192YdhAoeKTapaxKL7Ly+ZvueKCy8iulvYZFoH0J6sovYRhd3SSbP+g/8hD406upnNxhxhocucO+0nxKtDDEP6v82/MV9eeBMuF86h3vNe3luQ8P6Sg0Uh9AjosXKMg2/WNPNndBfyWh1rJ0wYlQWWWAeziFTYdk8/CMAAqn8+kZk6vn2txr3QIblTXxTK02E57VwvkUdkk8+tT5ROOgVyE5+MvK9gL9WSzaiZJmk3sCTzuOS+MgT814B8VrDA75T9lTeQxcgnLz7npzSWO694NlK3FXNFQmumzG9Otj784pQIsSDQKe51ef/vqiXVsYVSUXQuj/Ximg3xZnPxDLbB36Z926L6DvuSfU9JMfrO3pcdabCVbkyvUppX51TNqB3OilnaFPtJES3B7H3pwrbS7gOPie819J3nw7rZAeMzUElFHcqnJGOhycyTqYDO5u8t1fRikmO3+MlAdgAbHeKMuhigCwdlSJWJG3meM4SJYDn4SagZaQI8xp5HOqCaxSbcdlNN2lKRWdhJISdfZmIbCic/zzyEOLnmujr5DtFCaTaS9qS6VFw6UO1n4PbKR/8MmeNvNNxZBGv3yvpaRjGGu+mmvpNDKtUkXLfzx2FWGPbf3qoFpxyMFf1q1OHlgXm5YJH6OfTt1Gd6nFmLDstjhsXQSoJnGUm6bLyU7ssFFCFajyjUpLvtInX5KIKPNpIjLlpCwKxBPftIjIPW4r/USATPAGIri8grMTddKPyWjsZmnaW1bXEFXR7/Vih7lw00ff9OwgGryt69L334kw1MqbtXGZCPnDlVifVm9xz79MBbLznErGMQ7fTZnp/OrqCTDkVAerNWFBVsEvRbvGhEy7ry5o3niy3PE9GCLG/WZj1DdwB3oSiDTq8nvTXQa/DKqEq2yprlO4zqSwOS3KpaZa45a1V7cua70Ls6qOS6emFm2fI0wprosoUSG4B7uZq4RHXoI17KBxliQ/+Bu86O6bdhPfQgRIPw9dAS+IRsfcHgsTXKu8JR4piMM903f08YbUYckZYwNi55bDGVn5HNjfsWVJ1wPIPPdXlPjLHY0Sv82rRWujI/m96pKb1NJZZWNwqe3MSbBr3u6HxSEXE9GZQAnAvqXES69GgpmNYdxvPviCYHgDphT73lMqETLCVMccLekXwyLBgBsqPX2yK6RJFWW0JUtMbP2p2wCgcROWTnfjS0/A+4bY3yUuYkMyOLdLPYwMMI/WfWupYzyYkCqMppugSpKsoSyEHhWIt9s3+ZJj2kJC08Zz4O7j6/KOTYCVMfEJO/tyhVo9Ojj/nifZlZKj7brwytzSaJ+djvq6WkfMZ6JiBY8P6xyMZwc4wpRXvyiyk/LZMVqOgZpzUjCxdePNY7Cag1USOP/Gj+JwVjhuhJoLGnjG1eZsDCFiCX4InqXvc72wp5oOL5XxEcFkkn0416KdF/4KvRasTRi+oSzc3lm+ucQtOqenPKQc7cnOaspsao8ryUfIOSc8Dv9+B4y5cWqy2lcxZr/Hn9AGfbB1Akpm5l3wcuFCG656NofDljulTT8PbPqBu55RyZPEQao3HH3xlEIzj09RgGGc8IwFkS+Ft9v3yHMGzfD7YlDQiNni9s6dfwr6W/Oe1H4skB05bNcoocDfWOUqMwqdmoSIkd0/ZJcaqTq/d/aFlZug1ZQxvNNmPj9LwtvwvSXUcb1a9uw/nCCO2Xxt7MMTQ0bcmSqIiepRJNfpeKYTJv/54WV5m0K3MFepZOFM3yuo8k5tiCsfnmZQCEdOTCMRqqaISZp1HWYEQMlH7Q0QhvUWHyhtj6n3LZAK5qNtXLaRwvoSIMmZtamJbn+bZoelgtSl92PYretUc5HEDgMAn9Ukp0pofiPLH0A+BNli/Brz7r15FIODqW7NEdpgg2H3zzDvrXj7ulMv3ICmuwAWvALtOS2y5lF7NUUh3Ab+VSg0YNPE5gDQvAMHB/QQ4MvtXb27ZMJa6O8Ai7KfGC1P0ooXttZVaMYHWXaYf95yt+f23qtAglnp0QNmY5Zo679vKIBP/IESW9nmNWk0EGwskvybTrx5pioCfgC3xw5EP2GfGSVrpZZvP6ygHH4GYkqCZVX8HWbdl+5tkcpnEgDnlOjMw7yWBkn0nEceGjQGkVwnSipTYu0XoRgD9RbNlnMy8tGRyfP+4m6IoyyRB6xPHl1I9kV7JTt6sPordtqm8MHBBc2vmjH+KHlyDHedeyxJ1ZfYqTpBKnzH08i67bWxPvue2L1pXWQTGU9lHifNbbvsYtbpX1XOfPNgdroiX/um78wVLIgS362VSp6LBIRipHnAwhqahjm1NQ2hi+bEfkJWwHV/t9ISjvS9P/lW2r2wapCWv8cjJ6W/964QVCy28A+CmFoYDqVX1iFcmZPHwbT55D7DrNxnv7fAnILCrU/aRScEalZKljhT6ARMbMf6Kj8n62IRYebP2I5H1uSfZrI1uB4l3S/Z38RyzjdI88W9hcoBRfzgBj+lhbZ+TXvtnqpV2ZX3kwdIhtJmpAXlzKOGrHZlMJI0NjGclKpvlmQnLdKnZFIF5FWoM/CpkXvPVKDCdTaPtUUHgOMpjwRqpWh7caCE4XXsWeKgZj2lofvgiVEncDk9zD/6xFkFp1wUW8GDou1YnxG46G7ZfPDf8u/cSib0+o55zF0pT2/GVKdmtYqAeZr3QHVKtdvBSzQz0wcMz/FCekOdEIAQvJIp4NMG4QAhVO1D+9VUhq3eEjwgUBKvrhFCOSLYnSbcIPpvd8mIGNOY30WlEoWLfKoSq96JZE7SQheWc3w4lUZrvjJX6LbhZso/NooiptPpctHoAxvtDlNVfClMLjsClgPvQvCbAijUCF86jox4/mBryT8XLje3HYhjknCs7oDljBiKuZP7/qBi7fuYcw4BzPxCcHPE5QmhOF/ryKO97g1FHEbRoWGQgFXwVlWPNWIxdsmAj82zx0CGQ7dMNAXAA5N0QveawGyi7HAvgqx7kpzcEjyBHbTYE5PHscF/4kgAPhOrG0rdw1m3Eut1BxvVly/SxinfTiUYrzH2JZS/LDHHVz5ysXdF0ZO6PVAFwF6eSV4uS6AMIQDOaBBMYFlPIBNyLJxUd6SbOEw3GRkNJLfun0NeEWSEYfi1craYwLuWOSepGjKqTw1opV/5W01djGGwXHEsNeW1ghlqqWT9+8YEFaBkmrNxrXhmj4L22Uc2oYrnAloVilRktXR0MqH8qYfLKgFDJctP9e/zysAOg53fdqVhBYPGIYN0Sk6t5/ykL7v+Ldp8ZmncZzr3y4k0giEa4RApjz6Uh48phMhMoKMbOp3updgjPCgw7KLOZvE9Xg6ibNCk3CforllEhIRsrx1WBxs9jypI+1RWcv6nfrTldL317KH1pJ+pd0HkEgUZUDRgIC0z1TXXmd1NKOuyWDvrcRHwrBBaHshIVqx3SgZhq8o8O87JF/dQZEJPZXykjeR90/wKycNXhRlk8CzIs369SKWF928zJAkl2Tdk59+2/FdY0t/r75AKRGa+Y0A3MInDp+xexZnIs+wN6RaItZkzkzqSuX3q2XzdXtDp/nwFCC1jeoYFqPNQ1bl0Db3w5kBsQttHhBa99fhoZK6OTrV2Pg/4jc1iy2Fq9pVbsLcZpciKDsJwv4PcwAaWl7HpMS4K6JURvM3ePZo4dZqSIbDbC9Zoyl9Uo/AImUXunEGrF2R1wgpSkzqt6rrhMB4xnoGe5C5bAwfgbwMOx5twlC85FlGg+uvdTfvvuYQ8KNhV+J6Edp9GuIh5sjg3GmaIRTPdTO5jDn/XsrtYmNGKNANjrDcLi6bfG9ZCw1YdXjLWMdlU/XGx/dDVQN/RL+my1Dpk0VUNLjx3Wbv79h20Xe4kS4o9LWJJgzEfHAYocHecRqeeT9FF+E2SF3iEy4pN2R0WLXn8a7DE3taaPgFrGVIJF+jn2/spPX6SpNzB+igXvBekJtKbC8TterDe3W0cRowBpcsPxmZ3cyv1FccmtrLt16Q+EXxvpfH9bXkO5TjaF3knQ3VzrCdgtF8Lh6e6coH4FyfiQAVD3fTe1z7lbIM7YKrTi9RqRNLuMGhJ63kIdL9yKPbcK+VWUV5i7e4Meg8QO9UPAmHSSzr/9sL2aJGRY1bZ3OOtTMT6Wj9gOK/JAC/PEzKROCBTqfZxLd423hpZx/wSv8NupgE1uhxyHfjaId/jbvVQid1jndvl+ftLXlriGFPYGpB5CuOyP3eroALx0gmvYKRmr0v6KcF9sForfrUboY6MxAkQuq++w40DkPojYWicCN5u3tCz6h4rh9USoT0CqLhxdZvgGFemeBQ3le/9ZzFVqsMJxAwH40vxnP2tZ1MEqXfdtnzyrz76HKR/KJ/dFQOdlZFtWFKcjF7vpl4937n7poX561MW2vQZMAOq5GNLL0CJclnukIjtlkvRrE2miuTPXSMivzYJSl244CkMJFXv99IVGuY0DvxqkRp0hysYpmHhTJw+G19fa5XA8JJZ5Hxp2i4UXI850udgCM2LLOxXxuCWgAfhsIDkXP4nSjAJANiyCCrd6yNB8lMuaVyGbAZoK30L6qTMHSDcLuubqh09kzYi0gogILuZ9+bKYohMz1Zr9UdwF14yb6yrMQ1dTua7BYCbCB0HYMs1XV/tsvjt4Zk83A4ez28ug/JJy+6Gv6L1cOpUwvlq/oxB6zaZJ0vyR8PVKnl/izcUmGBkxNRCHHah2Ep9BjMgzFlPb1q/4MsiRhOs5yNK2TWPLWAWwVVE4BuT4GN1vWiEMoIyBsoCYzXjSrYvbEANMXlCkeYHbWKNqs93Howulvkt3ygesuw3AaPFzoPTxicrIjQWNHZcgHPLdHVP9KcFyp2KgiHGL+n6Tfy7caM+COAq9YswFTglJxinIflu4u4voyWqxHVTJXBnQcgz7IHseI4yTi8QFJG0kyZU80zAlFOvDuqW7VFioF/kTh8RjIQsHIgLfTUajXN9XxD2CXSsjKnq4TSubIiVFFjmFU249FsYUcdH0dWBsW7Nt/3dQM4ffpsvGl2q0DDPKRk2fTWrBS+Z1iYOQDq8NaUC5hBlp2Cl8txuYQLf7dkUPIY4v2JQ3He2uyk4QEAcwxlz7ILCS0Uqq/qSZQol2odV0HoFc2kVYkNOVVu3T2BKmNJZODB9q0YuZiB/Ck2yJU74n1oFqgLrulXyUHGfLanfavz6V9wirtKUtUf5rgUCIqxyIrz4e2IfKIqOxTrHuCjifkqkkGDb3YwjrmJ0fl5tcAsSH0DvzrREeKvdKHgEDKiwYCsMVIzmK/Focu4rbx0qZDT+PfndANeCNXEdhpIfVKXGE4E3sSKH8NMquRY+O6YwG8zgKZLj+SJj6b+zFFLI0yYnGYRQIdEArXRVcs8Qe7uVy5H4Egt7O+ltCDXoHLT4EwlwbuKuK3qkymyiyHejiWMBjN2UOL0cJpeJykfKD9bDxPirgmwTgD2VuyJtd0UWLo5ZDs2+8SWVuNm6F2sJNEaYO9iuuwdEIe5ZA9Xw827DEMR3MMaLuF4MAjvlxlqcHJ6G67bHH1CIZkwxhPbVg9TgkZI0GPhcNrv6ssz3q/xLFBeee54rPAbdT2pGtBiG9EQVFvK2Id7nVQLrNdHY1T0I81CTTrxwAUq3DF35fJ5XTo31QKbUR9bt3oNHDb91ciif3zeT1EryLIzuUu8w37GfNgDDtVY+jo5JWgWZmtX7bRHusUa3PmMsFydCdffxOaVReY7fuqurKfsswmHbiTj7go7S5q3wt5AZpyM1lE1V0lN0QgsKGi5Q1AOsRGDLielk/1cBOb+4mT4wAe61+dNsOCAWUcm44wlAWFAk6RuxeLT2btuYmP0lmrIIJIzBw0IPog/YSTeK0+9KSW7F0Axxk9Q584/JmOXv0kPY7AUo0dbFKOyg12HrJCqkP6/WfcdjIFSxtTAr+5AhBD2k6GFvexg79syUidOXG7uKMbRchhs+ZjSBoWWLmclz3YRIrvD/nD/JKUSsfeUgZWCZ1vcI7ygFgDcyG8wUb6AO5is0PKkcDm+04/yjnhlJDeHiKuF4wNXaTC5CFKUlSLpPizzWT8ljK5419JpuADvIHLisOQ+dGh8MnyFm7EUuZrdEKpnYveipnVA3MpTM//8GtIktQ3lNWtFlvEIqFOcytSgDwQeMayZd9wJHH/CusxQqCJetPD5I6C+IPletozrba8uzHUV3U4DHA8n2Q5/cn7eFvYUrcnaFEf1Vm+YagM7caDrrBpdMF5eJP217sIWmJhNEB4yH7uYZ4ynPSNqfEyAxAEpc6z6ucW3OvAP/KzFoL38ryyeE/SrID4psfCK37V1OLN4hBjOg8hlmHob9mr5N0zHoYSvnynB8LaQ7du5rb5VBRodBEDbDTN1tOPQxxzkteLQCcd3tXkM9jJIJQeX/fW7fFT8VNlxMTnZrlEAJ6eKAseqZ5UwxFzo7MUhFRmUqlaGKMMI7WsYx7fqktljeH4v4Dy6T0KXcnoHzN0IK8vKXl0/UG5/i0Ho4n5WB1IGbJE8O3OZ4/CkHzZzcy4A0DDiUBS7ntZToQopbZ5TEdUqXma/jyGsMG+Dx6lKRcs3rL2aIontJl23C6ZCxGGY1vxNpwpmrb6aASTunmULxKqgyfoC/smV7spYfQ0pXhyVvb8S8KH2mVT9Dde20l9ZFmzQ23q3tDEJ+MMVAFbsKriYGuiozv0LOEek+ces8UmOV/4/qvQenUtTpXxTa0XW9w0sF0LNgS28aZceoqjFNz5GbLvWwOeX8gwC8jpUvL4/lUxnRuoQDmdMhNnnz3ZWmSQ4QP6vDK0xW20CrQ7hf/09MxN+mDFgvMBoyESq2XfUZjKbg0i8x/CPQeLpuXt2YpcqREuYlsNAyZWp4Kx/JnQQon/8KB1qQG8cHRVetf13alTG9D9tIibn3rFR3uYjc3sDUwo5kAMATeLNoSfAZPU4+S69yjCeRQfxNkeRw+94iw2y2RkZgNZnUKcjMC/KXbf3EIPltFwNc+41RwWm1hflV0j0Y1tncBirqrIerrjv8loHSOMpEkmaadnFfLPxfLBJDol0P+yQ0bsz57NLSvraBqL1LP4vgdldOCzT1s1ud3b/9vkx2MyasXcdr1Swf7nTyVH5JfDo5t/AdN2dK4H08JnpO+Zspuqk8LP6az0CtBGxUAm3TbqNQqPO9+U5KUv9DNj7V5gGNZe8qhkeRcY9//c9TQ07z8+6JNQ9XpOndzu7K1ThANy5u7kXogw1Bur6cpykU3FcmtDUcQH5MdisQooyVmCUf/HT5qj+PCag/itJd8otQ8AlgHKyaGeYy8jKQnLef4EooK51XygM8K8Vi0dYK/Z7Y/vBBzHx+2+nPtL6zpHMYEeB2/yMXcYPCSUPJxke2T7Eln965WZsyGwnqB1c+gjsJz7i5HhK+l0DDgPaezpi0YRmPNXobbTnEL81RjMrgWQaFLx0u2JAMnfdn89cIVT/bypTpX2EVzHSbbV09QHPze+A+bmZW8Gi2HyiYxJQiB0vEiqeFq8JchvpXazKwYEGUGFmJIvWsvg/aCGZca3Ac98b6CLvewFiNr1RBCXkddNdRhxG3pGkiDGlMKopMDOcg6S7LGpVliuwGrgPquaoo8ijOAN2i7IEKCQWemi7iJXvbexGwkbBQgmakc6GWwDXsNvH0nGnlOJ8A8QCYizgorMFwg8XjcoBwELH4O03Tv+P9bquRWxj/rLwGE4paMT6WwiiXHzwA8Gtw3Mnq9Ro8YSMsxAeOp76CMiEWZPpu3a++ASQ3eRh0Z+ZNqcRmPDSqQYkVufflxr51JRhre/sUaTDyJWVpzD+EzX2HH/tPPXuxu0dL42Qz3xpLJs5lflLWmwLaw/dOAklrwA0Khf5xHjxFekoVCfyNmnSKyS41CGT5xVhEPbhF65TI2PCw9hdGxzz2i2ervm5fQbK1sBhQRxd5FKz6LXxl+chhaawfVCsCAh9GMnMVbQEohS3Pd/TbVfq3wVgrryQJQSx+vaG6nc/ODWmw+8rmvQIVO9RrC6eGFgOYqJ4+ovFiaBVOmmyscEopBtALFyEpYbcAM9qWvg5xlHv3uK3qVrXgNYY/07FFEs1kt506BBSMTLTVWgIhsw/iNT8ERXT+SSIgyUgfgVIpkHn0COulbDjztXEV4XZq0SmyR6IJkq9gDVfxuxlhoya7BnOZJ6pe/dwNTjcYqHGYx8LyDtEoAScPyvH7u8Du/n14YYmOLTCGnJXRMeEuLP2hCjvVGLkdD+TcQLlFwNvX6/iJ8FGKvckdK7GG/f3RLQOdiS9Jpf6hotOtDdClP/msrxO8QWAQeyMoTpBjYH6TfjDqZsMBkrK1cJKkWDgjXo45jEssc1TTMfCAJfp9mKoJ3JE04S3spEpOwUI2yAjR7kcvGAJp0gyKTJ9B+hZq2cdhpfQSIFNi+/OJBAdNdoIZR7Y4el+ER8DlRUUdcSTh/bR1GrsYkU2LUAIuJpQWHoCwPua3jHjf9bz9R8/8GkTWXcbVEP6l4UnRBTu8WXjRVxGxHW1YhRJPO0nwlWF/IJIbbfoHcoahTxlHycCvLQzTXg0mAVQGiq6NkLwpcULnQK8HvlCDaT0iJIfwNkgFL9ddFbzIadV+SG+VzCiOCIthSSiXD1cm5Q7lSj51+1HGQJq3ujyp7xE4mK64BdyMV+m4tdNlI1XdL/P5CyCC0igPBfUG9YcFNkjYLjHQeTE+P1S2HB+mhfWsBEJDUpcxfwN3uWc5mRCGpRvw6zKutnE2yA27dJkwCDrejeRZt4ewAKAOf1NBF7uXEugyc0b+PY8XZqxW6KbaYgdDB8C+9jwmVTJNnBqpiU/4E+tIWqWbmC/Je6OivZKcYkyeSZqRVXfYgB8q8Bz0555rzBaJfNPpM5H3ZgPUWtTAOfzTIe8V67trG7RYH5FKYthbB6xyJkIKXohIc7QHOW8OOIthSghw50Tp4N7xGmuipsrSP1LUt7WAjUw7b2tEnQhvmQs0/1Siu7AH4bIdjmtzJ6/dqx9vAUKoxGD/XWQGdIA2tJNRhoGiruZKCjizcej7UnQrQ9dHa5rVsUu/5WPEJ0Awgb3U96IsRx6PzSfDIA6yr/L1iqEdlXoKWzNn/HuTYdJ3/96TZKEia3nTnvNbhDvjgo5/nLtDL9AkMTu9Yqw4mtzaoF3MJU3lU0JCHkl/anA+WqscuDLTNqpe1zIG1+INnGxaCXPsov2oCDdkeYt5LC3i48IaM8oHcrKnoaIlN/BhfiMAOMCy+MBP3E1htMZtwkLxiTl65o6rxELf2mMV4s8d8EJKcxvYvD5IrhBoraTrIALGMVqEVZpc3i9LoyGusIjI7NmKxcnzmvsVLhfVUjUc4L250iQlthwlqXEb9BMSeGmh3sgZuuJo7o/HeNr9ZJxhYQLmPWpx3r3qD/q2lx8KVKPvO8G/AqYSTmjG6j8FvCNoE4yIztpSr3i+s3OX4Dxw53IjUvbKF6evAb694dIYZ9gVu51AM/hsYaGQ8dgADurqptiA3lXzs5JjkqZKxniNBJ+AeoEyQQ9qAcyzxvzyrZC26FcaLjoqJr4t5zcyYLo5hl72Z0k1yF86ciqecLqZ4odEkVBx4UKQuo3zbaWdz7JM38ijxtImcVe6UisChfLImZEUdwGQHmyohYws0x4Q22eZzanhBkQsBEzGTy+XsZ8tmA51rRIEBxPbEvdp8+BRihQFHqHC2yipbbZ224FeQj/oo1YE90xChMdEr+WERwMlVoDFqdtAfS+Hlmi88lQXKRwczOiPtnpteRBU3IP7u94bRf4XNFRSFkX5eJuu9qAtFmE/N7lqQPR5WSVKGlz0V8p1lSBvcui1lU94Jgb+cTO8fMYEgcpzv9ZX4sWbZ7BSuowoMhmr+LLzO/jPysRD8tiF8lPof9HXfiiSzzb1XDnIiYniupWuZr/KJGoHAtS6JumuoP2uz/AeMBZ6uwXPWpUy0Ow10mFffK+JuqMYAlRGVCD9L0ndbksZfNAPWxz2WOnn8cNbB+PzT0lRuBUxVIta8tnGRmrltD5Anjqi7UrBMnxEDj/donVkFS2madHt71hLcHLtpdXPCPOqAYTR463UPvQXuY2Ewg3Lehkbhl7ksVI7Dur00plpEMOxg+FwvlcB5JPXWWgvZbCRLiMAnV5T44TaCMCkvVR5Ez5LPGhrwVVRlWIapizx9PEZibvMOovfTIS1jqcpgiQIe0RCQgShIHzS7ECVTqqq/xDSMs5ENpgNVq0O9t8nN2IEr4ui/ueM+Z3tDZO3Iam55jqsA86DAcu8Tqx6ocjCwxCx8zRBvzaqn4h8O/MpwYxvSYrYz8He/sdVsltzlTcmnJfFqng4+uXPBLKhdSbWjir49kr5Z3SPz+LaI7zZseXL+UB15bfl4XUsEMG9sIW8TFweiyTmF5Md6J2pOAGn3sOwTWTtsJVcggd0in9/JGNNlVROsRffYo5iOs1JtGyVO/wHd5tlhW9Jr4fk8naULAk2dCIUfO/itR9DOFDG4R14q44X+wmkzjjd90P5x7IZdhdM75bXNPYSRu29Wf+iOPVYgXG2GZQ7pkbz44ppmd11Vq0U7Gv5gg+zlGXsVLVaO6/OnTaFg9f/Tc7B7huLW7yEPR8mlcYb5DhOpheqXdoa2jKgrCQ41OY3se3FaZ1s/DfS2AXKZFrupqlL1RwciLMOxQlLikfjp96s3sdQmiZg+n7J+1JI6x8mheRT3Ltwl0dxwGSUereoznIV/WzPhRrM3MBczjmcEz2Adl0Gw9ky2rdmyu2WWlPXSGHT6di7AUzE/l1ktpMQcL49Hr9OqEtnW8ukwERL8ulNm9WquWYKNev0tLpQSqKpZf4H7K+qbahwyoh/Kl1B9VwJKJxvNqLcoOUHU1TBYrDMXAXmMRhoQDeu7GR7+VMZMgLn0uY5o9FbZ1oECkz7nb1d+6nhu9vCj730/ea0xvykey7QBkiM2XlPdS8sUUUHS5jXwVLJill6GC1HeX70Fg2F6PFr35Wr/LSMgTDrgjYnKdhPdczmVsvieiG2bXm9n81/hUnZNwIm1fCaaWKF07FfCe3eT32ZIKK5dwCELGmf0yKSyaWy20ErhdpoDCpoQU1gCuXv4542TpGWN9uZIIlyiV/NFWksy7lh2Pl2EAlrFPuY8wMzx7QwVrIFEUdeAqjqU+O0hDKM/mAML298IR7wjXfFkQWpPH2BC5+nNJrE6+I3KI7Aufzn+Cv7bWF2POp0BZQorDjD1n6reWY/V+DAnuvuDlogFA74npwMA7HMSZUI3k1CgplC3Re8z2Go+F9y3e56Hf2NNouf/9M6FcSo3S0Z27GlzIIG060rmDGZgi3mJbTPdxg8uXVknd5m0+NgFxBubrqg4oAWp69pYtuG8MEIK5yKNFXIE+h4gdpTaUSzSMnDDLe2wBP4+WkknfWGJYFM1dEfvXQf601aov8WTVazbw9+iWS3alyzN7J+3olsWJkbcLNYRpVvvSSzEoegYHxEysq8VhHylaZDo07gtgOBeX6ASP8/aZjsgRLCNTpUh0pGeOZQgQg8/E+s4qKjQG7U4oNKfrDIOnT1bpHAy7uqGe9IgUOadoM37LmdEr7RhsB2NT6au8mjqwuBog0nNyMzuTIsqLIE/Ut2otdO7pjZwNHpE8EVK2lkC5A9nparA7tDg8W7v0Rs4VHLXdXzDshCkiSI7HlOxPmBqbe1vK2aLSDy/U4nHy/x8I2qdlURSEXMyZvO3hSotKFvxYpXOsTg3nYlwqnhEp/cnzV+7AwhQpIAQbxCy2YK+/h5RSd7i/0mEFax+vWbbzH3sv/XuY8Mj7cOKLfA21r2/2ehHv2XUNQ3O+N0amrQg3hGaPV7OXN6tTEGAt7rvrskuNuc2tdU9WFPuJ7Dz2/lZ4o66nAOdtlMf9R5EuRP6hlB88EAp8Fx8l/tgNLcbKwWaRazu+k7hmAvmqhGNHegAIhDabRY2cjpSS3Ih8geAa0tfJ9JyHE46vmIBhj8Iqm/Z+nKQHG+JiWNS8GRJu5ysUuTDsAq2g1uHeIGjs8/A1fbU752Ie/7+iYP5mtlfNm7Wz8WBTJz77HLa3U/BxMsFN7+XpIg+8MIlNErQ0EOANz95Nyb0TcUxw7KdTrqbiTBnKYolomOQhxslT4eQuo7iWKmk21wsM/pLf+9X2OXfJZaWu3KEe7XSno5wPZjy+puKeMxB4ItlmBLzwegsxWu71s3++GWGG3sscKhr36rzZ6RnGjFZq68FBsWY2mdxX/DrIuzI36/dNearmGGVJBJ5/D7Jd8xm/uYOvP38PYpkrMWjppT7NRpFIIdl06fnlb3x8JBrK5s7PVN2Vnx25ov2umF5ys6pry3AV2Z1eoL2qOR5Jys2vSeGpCcLJdJSB/fndeBDKlsh8g0S0uXwvd0L0jWgE/Pynx658PV0MvRK4qHmphi4AwNAFawSFPklQlroFi/Puvet21+1edBxKUS6CE5BUonj7ioO2Z3M9gsbArSzjRAtH3G2j8GwyTHytOffMux6rmQqotjIhZu63LwW2cZC6R23RYt+fmuaWpRfObacMeocv7SSGTQqoOVBRuexXl8gs9GZ/SvrWiEGN9QNcwCm+QzFBJpGW+EnhT6+8oDkGNg9x3xXb5KXrd63s5JYDxes6ef74dwSrF8VEFWBd19Q+Loqttz/3iyZyax/+R8w4DIp64SD847WJ9XVrIAMWO81iJVTV6npZBjhHn1iiel45Q2Rq8cVgcU5Wm5iOxGPL8yECjui2yaSutoxz3aftADdWuDOp4VIaE7bwjVVOgzbDUjHtr5X29b5KsThbAxuJ4k0CpDQU3py4gFmpEx7U8yCSqTDS7DkJaqWNjbTO9uwfxx3p1/ojWUnsq1bTVOHelTGOId3iO5r3OduWe7PV5FCt8N/hA7e9jiXpbV31A+4mcvZSOMZ2RonQPv87SGG93+ghQgsIkv5wtNv1f5PUG9XJqr9epxCJ5bMJVIZ1Anb7V73hzEa42aKqY1SO2uFQ5LI2ruswDApROyr7wRzQ5EdwB0Uin130YQHQBS6H7oqIGGCQBYFUFHHdo5S6OJJ/F+22miDFFTticP/B2eNaIQ7NoE81r9yAb6VezrT2Ldm8RLciEVwMCutzxcfEZGGim8eEkmXHbzynV1dzTsYt/NeVqgX5mA4PEFwgjET59gOrtQgK9u0eS9/mKQshpcly+Z65HvgKiWs3HbMmEOqHfcmDeWv6mTEwohU79ye4M204wNdz9h14BQeVqfDuMixu1zcuFNiyV8FGZMvJbrQIwAVfiFKyrcD3hUPtMcxM9uzGp8yHYOyTSpkfmX0BmO+grGYNgIayo5kUxePiPy+HySlwEDlLE0UjYsbp4NRycwBxr9AuM9bsxGLPnCVl1dYLfAiTHXJpIanxl5OUoPYYLPw8emxeInMbUzGqy8BjeIeUHNlFhl7SItpPrG3+u7SIw6VBts7F+o3iXQcWJLmRwYrenewioB4DKZBe4QE61ozchFsSA7RD5CHBgwnz2dslEV7pK55ye1yDyM8nvZMgMLlnsGzoRlakgGjfLMIR3NDbRJhCFolAb0RQ0/cRVvwOJ+gFVe9e38X6N1MVZZ5s068nrFxFGm1LXsLW1YWKNLtp7Ds0JdJEMkr3eRwU9GshQRsRyGXJjjBOzzHvTjRpG3cOmtJ1NOMN/wxdoUpYCqduA4f7YBgMuk+A3CD9jjSNNnhCBRshg7Exwz1JkDq2PFpzXcHd3W33p4EeDglvTuT7y3Vo+42k4GltF3jRquN04nvSeBpdf77tJOqqSKqFarv6GF3hLmPKToECY2XjE2FwyQaHmKUTYgl0V1y7IeGTDqDDltkBqtIcQzEnmyQbkDLjbrC3EDOVWV+sHZlbFj9C1R1pYHJyl7lllq5ge47uk4XKPBjAcjtjSH2whur1oAHZ9jWEKZEKDD/j4YXjSdRuhi9B5UNPCXnDDqnnr7a5Xgk0mhvfy18XgNuPWQBKFUk/XtNO+Zcj4WTLVuJvZH+jLwtNgwWF/t8uLrpIz9AZVWezdwdmABTovwNXC/tDt0s6h6Dx7GWSV/sEMwOcVEztM1W0qmEW3fO9uoALOYUgmq8e5yvroIWSjTFUE0VEa/sOLO5I8fxra5dPDlyB4gG/tPO+Xxn9fnTXddbPxsGDgVgH8HysD5CJhjuXofqa5ql+OjLJTCFerhLPmo9JKSFjZU1/qZysyCTyi8cQVui/FEiV9kimGzxEOQ99g/tuClOC9crbQS0qELT7HjksgaVfHKs0Og98/ZQfPx8oRVFmMudEpKBtK1iIAqCyLb3ey+Htfn+eJfb9JR0Tof8Rgk3hIjU8VD/E6zNfhN7w5qiE5DfnTs7WTDHMezyWsv/yjkSFqaXdG3zKiaE3xf76U3R0Uh9Y5wHIpPBj5rjSJtWtxn2puSUfeiG0tCswHcS1jFNvekBB7JwkVWHrJf2R+At5RaGOugrytNPPssWQ65wUSkjjrd0aw17461fcxHBOeiKfue0L1ICzPIOIHD/SJvtOMI5NGCR7vFyZloXGmmP3j/doDD69aP2/NRApD2KDVNHW4cqD881Hmp9Zwz/3wwFYRTrtdp/dT7PeaGL4/pJRsKC+o4pjdBTSxMNDE4q04+9K8eIyQLKfpkbCRxF9T6Unztcby7dpHIGoDY4D6uxQjwOZfAGsIM+fsBvRrFMqdR0hr44fXqB9OdepFThzvi76pdtQIApfsKH3S91KtyxP+bG7/sOTTLIxUF6IygT+bGWRiP5fAdi9lOwO7yM2FkbTbu0J+vZJp3gRKZ1MRvOAi63qnuva7PcZ8G7Ea60vcvcKQvaEGwhWssa02fTb+d0d+pH5yiiCBfJkuPXjl+4yRTxT8GYBvG0Y+tJuqMUrkB0UdYChC5XW2eb5eknxmYb7cDpcfvYb8KBFpFnIFG7HuWRJyiiy50+2vp69RjYcqkqRdREomXPWtZ2CkANwNCoBBpE9y7JvB6Fudl8i2IClSKFpjBIg8e03sVbcTlzcGiYko8SM/qCYm5gB8FUOzVkpthMnC4t4dds+wQ8C0dyri6sirXYurAm03Hl2o0UFoI1TGds3wKYqLzNpP5b4S4CKi6mpdm3k2xk4dwAO5gJmiFRKMRfnXQTPy/iTuuSeeRUyYTGCk3MrJp/Lj2ZAxGeFgV00Up38nF1V30aWPridNZpSnQsOv4MAm4JrsnCy4/Dh7wlFvn6suVRMFpHFuPp/KZY7jdz2FYo2aRINnLZ24CQJ6bnbB7DLeN1YRwxhJjoLw79lEWkGex+HVBXXi0Pxon413fIaRDfXM+DnDYUcQyvqNEkQBbXM4z9ohuFByKte4yA1Mv4vSQ5b+wv+eeoT7m50Edcyji/hWcw92E6nWwUKhPCGBY0SS0tYryas1pRaUx7x+ZFTip+KQVgobV4WBUbo8RmjJP+b/6z7tZjH32tk6w7Pzgj237ZU0MwM/N/7HmlZq3rVetWY0esYA5raS6OhOZcLxSuylcUBY+SSImhWBFQjPBrlM8Z5zB0ewzGkrq6Ruh66S7nRQ497SBOLBSj2y/jrgotpuESVxmJ/XqsUk8uAGL+ezyRY4rVaRrugu10zyW25cZsZsmFYCxtoBZq+zlyKVFm9oWpAPLmJyG1FrgKlmWDMWB2AuDow3hEoZP+RzNml9xSvHCXFyVyvjHnX2tfdOWKKv5hjN2N5gz4z2+00PNks728F8MGFGXDbIw8ebUcAac1FHGGMhzNmRqOzTEM8Lqym8EtRUUQD9l1wjHJUzmYgFXJJMRrIhIEYZRsNKmTJVzPsjo+fIsiHvf76glE8Dj9bL1oJ7X4MCY+88VELdr4FUyegYzjpmP36AFnmJMbiRIrYCOi1ar4X8689r/lfjdMUH5ETQBNTqL7kFUNZovRmuS3zIa+QuhOb1S5BZO7BJfUTtgW/3eHrkNQK9kgG+KlfKwMDQdh1WfcIVsB67bJjKtkppZTofjhKojklo6sSvw9ph86EJGE80t22gHUqJ4eriPx3bDni7ZpKwJO+1bXAdtoKNg0D/RP6QrmFe/EajN0b/8FJoBuJyxfSC+hFZjT3f+DsgCqQil6xQ9tyfigTOhgM5bMf0PL5HmWTVj4nMk8opMntUSJAI9k8hf+QwLzRj8Xv5rBVwPJM+khDYh/ZCCBaDAgSk0jxgimhDzX4S8RZLUxtTyi/0ysbxFs9lVCh8ZRCtcls6ztQ3HK+EUzizXjHeCWL048ex+eh889xvQan2T4hW/0nJ+IlpcJF8H4BtXiPBwO0nh3ESBhZfCGEUHnHulfgfKzDBH8ReYrm5DzoV/yCZdEI695664+xTEfxGdZ7FmOklEQ4jT5nvXQ5e9JEzBNmQyPBr6WD3MSoJb7I58EvGgetVo6svriyem81e3fNXDcbHyMOOO8+513zzNnE+Ep3h3kQzWLtHE3PFKupApHwmxMurpNCfVMt42mXahJ/llH6VznUeOSqsJbUSIVeinEuufbu+3bCSX7qGfZElXX+2Q59ESmPR32tzNPGpKf3+D010dWlWQI0PsiC4zFk20e8uQT8AAK6a9p1Vfqp6VPynngI3rK3oor8+zo64bD1hEdswHA/gG5WiaaXxR+BDxYEw2DHb4FHhgvWuED1g0gg0TeCBleSumjUPKcvFV3idicbLqKkmtrfCVB/hskX1+Jkx01qQaFLFAGmRLrFDuSYsUwSJTZ7/SPNf5RI/5W80bSDLBNpQp/2OblJSk+5Zi3bSoAZMtGCUUSCInYtGwkh7OqXdG0EGyRt7mmOuB/64td36oE3ziKf3Yv1geIJfYnToSqhSwfC6GflS2aMFnkPPqOSB5B5wJsjdC2zFvzOoktrXa7Zigun4nMn6mLbQXa7/kNSXBDxnkBHYeLX8s3P/NtfBNIiOMhvCvRv+neB/q8m9lhbBye5Y31HDUJAlFLPaujCGw3ZA7c9h4OuaekXn9KgoMEGFSasE1r2ojFn5tU+tCG5ISd9NWOI/mvwyR0BEkM1aUaaulipndGiKrnCob3EU0MH6+mcXnLcZz/0iAhNh8SHvUQl4dnKzRBFNMR7xltRKV+PG2TeeK75agjJmfe4FmzhdcnjptQIco2VFrgh8c6wqBCJ/nRwQVpRHVMwS++yoUnI2P7pqw4tPFAcSnmV5EVyJS2BKwJ1mXxHQ0cunpO6TR5Aq+6eUZgD0iL35Jvl3NIdNBj6XPqasPN9oLvDjBaQ713voTYso/cvUKpo0T1WenWB71GnY0Vue2modWz7fTCtMSvZ+yT7yp33lszUQSRoX8PQOZz1HFhRDQFJB04PYPmdRQQ5QuIPD7COKSIRaQeLYlikXUyUbhpbSQc1KQ3jw76g0CNeoqEnnHIXrY5EPVoWHzgMiIItrxGnGRCLnZp4Rx6v/RMLaloZt3qsZDHtboDRQfuS0K5KCh/Jh/aCaQEycv5//a6bOVzy9o213kAlEOdbRUdkw2e21VYUx0v4CEtgqj1ZfQ0ztXmT9GAkvpv/IkJEs+shjN+Bef8Drtiz6gIuCv2yrmuZq4EFgTBzCYtof5fTlCKubHjlJ3ndSVNp/Le5YofIy8Uv3Cspp8TOFESf4cWjz/qa2CxUrr3owp9bqzaHqpb9qo6x3ChstokrgBE1/Ln08RYYflRbCZK5jJGDkjiEthA8AR2uTRFskAv583lmYvSRolwwNSGnf33KShTtfzUrw5zv3d8T7LXPAf8WsAmD3jqa2Cgkh0V2pxfiteZsYDUv6DpFa/yR4jF9mCCHYoe+yT7Yt7Q0mHGP/Z8yTvHlft3aWA0+VXNRW00CzwAPGQyszm66qRGeLdUjFZ5FFPjvttsJcwJiWbhkDygXUBROTzRZvaUltxKaqm9WTah0H63qGhON7lxNJ4O/EfgWmYX1GvtyV3GRBauolO87cgjsvucj/oG95LlVtgXGgZrMt8uMhzyGDadIHnbeS8r5RCwTXfu2Qp2eJ2Ml51Vr3kKtgl5iA+zzs1JioXUfHWaryXdxtHGAsZUR/rO6Rfj/Ogd0ENr09r6NmT1bTZ9pQtekWxUfSeJ4luVrM/YQLAMEG5ErGHlqxWklk4PgHScsMdjNBcLBnfB4aRL5ROi2MFsz5n66cjhYWO+kQnnUiGjupg5aDYOUPjOx8DB5x+Qsn4kbAySRMa6Hvjg5NJHjn8GQS3Il68AZHxfISEFrZmE8zspvxBXiL5YJJIOjXNgA7vuIPjWHC5/9/6nAevFdXErBeThhXKw+CBhQs4ywM6xiffyIoUJ5jSYB40J06jmOebtR0PQ/CMruSM1aD2TKtmcJ5rC/m6qFMteAW0hDx/ztxxUGHpMjCqf4Lb4MjczP25gBdRGVwH5mZxCgcbg6FzqIfWlPYgA8quhhOlE8k+8WnaW8DxYGE2FfPtyH2iZLXXO6wQVV7REAv4LNjQ1SeKmopAD3DNYXuwD3hp4enWMtzoKHJSYxG/tpHwAj7WIfkNe22bpJxZ79VQsszWzOtoRQeUqLSlySQijxztE/KIMr7G8YpV/HhpvtUgvAgT8ie/QkNs/twnw4ciM40f7fa/JmQhRRsi7XRFV0jA2HJrSFLF5a+pWl7UcrM5saKJwEaQJTVaEdhq8ni4YmRU0wLmVeclSJqRipwxSyPCJXRCP+NKnK8J/wV9Wjx1MIp0022mShg3TDt+JSawj4QgrceVOACXkvBXNHE0opB7hSeGHqdQWU+IgAwpVnbjcwPwZTqrASRGH5cF1xpvqU4U+cEndMK54f2sEePAR1V4u6Ls9yAYhInyd65EOnTC1TAI+oYDisNO6FqxD9H0ZZZlFPB8DyS6JAujCyCPRrK9qtp/9tPd+bVVZmUaegBGly4+QcUPzp0rkWQ9e/dEOXntweUalZAB/1hWa6chapp9hxIZaik6EN+0+QS+OOwcSAC/2oPZYXRGpgBeAxPXmLYKA/De0eBupIMQmu4ZRVcuxMGxQM8lCwRwV/3DtDH9zl0ZnV0xkmnYRyxCzvmzkWtpALNPqxAqgUQo5PW1CsUq6buAWEkjE1ZWDD8NWnuSd12GXeZWdncD70Xa+LvLWGwLeAxIzavhaf+eYI1ltbLyzwiA646M0gOcJYfYCBLtSj7Vuo/0o8IZ+DWhDGLiYpTMFJGvfpxe/x6sUUOnP87W4otagKxe/sqYL1AESVGnTaXiXWZ/egTJNaAN4Kb1mjr3Bmxn/Yio2/S5dVq8ocHPxiwrTVkH+NIjVG75Ew7g9GQh/Enp58kSEkZbCTs0eGOII1ysDAEPdQX5EfdXQDbACCB7NdV2/FbwNl9tXWi+MFfqssmeRiBadeev3kHEd7Y3fmyzfFK3VegyGCea7umXFSxM3txMUgfANRwTlABb3JErPFKRXLa/+T9WGoH9pCVLmbQrG/q0BXtcbrgb85SX5Ir49BZ+tAVCj6dZhrvzDl5E5DR7PIkmioo4rPNSNSIiIaj4KHDKMptbzVMyHPFssrA+PiaO2ai2m241Tk7MejNSstJAPdInDnewSQEZi9kdCkzFXi7P8enUxEMdR3OihT/3SdjklaiDjV4L0/nPD7h8Xtz6a5VOnmizlTsxOCbAO6Bzo1NIMUjPzpWDb9mTaqQp1gcwdN79i7hXfmR4uaKsO+gGq9elLkMx5vHwrf+3nfcUNXNUfgcLIkC4kdosSwPT0SVqvIVyG9oCQnqQp6hAU1LHZhimunRedF5Rl4DPA+OXbZPJU0OXPA7TEDBfOLaIbu0VF9OVe86L2ScWABZz3aBZJwGOp1CzfD9Mxyf+beJITMmrYN0h5YV1tOm0ZULHtYHyPZEfWrfWKxsuw5K0z7erkuW7vIlTuqB1kjOa7lr9X3l0HwFdVTtZBly1CmW7Jf5ACRhrJ8r/POFk4UqdqyahH0C7Wtta1NaMskbGGGa3lnZdGO3ELgsexb1pzeepBz7X6zIZlIEHQul19694ry16ZQMK1Mhy/dk88EQW6sVgJ56FjBWeSW2CT3QQPulxpfihxTKfDInpv1aukXhgqnCllMR/7cxKsEKE2YVLukqyntobjov++Hfh8M7U2+m0im1tmDDD0yFdzPUoqxkYMgi66UrBPjBeLcAiYL/zk5fypMk8K8WihS13Eg+qcDd6Q+z12/yy/SiTMOCQIhCExj19vlMpNRx1HEK7tzt2PJgTEMvWacujhup1CLYRURaTIgUo3lkrwPG+HgQ/3ouzpSR5aRklhY4AT1M5r2/7YoOPhxPHiPULADGqsodZYGyk5KQlU+q9AumprbTTH+Vyg7KMZJUYruZqvOEvtIXd87PsiFdP1DVxfdhfvW2SPCVkBofJY1TyiSTR4of/+PmOyn9SYq2HCpTMO9fT/OjJX4wO05oeD8lAjc7kn0hpIhGdV8wbG7k6is5D5ntcixJEP4D2Yzlu3wnJHYsI42ZxIJCMSjVgYLQZFcgScclPtakZoJQZrX4ln1BYuUiA5du2VF1CIy/14IqltiwXttpG3NTYDLT6HRrOhkAZ8vQigUyS3NB58bQJwfmZKDLYqDVRqq8maVH8ZND5FwU2O157j9rJKx+7xAdaMNsgHDvSq8wel3HyLW08yD87R5aJwmQfiU+HKok6CiCDgZPZ099XMPk3KWdYmxlC2v09RKyy63u+vwvcIsGpmyZi44z1PiUxqIA5tjmGRib70T+JO6HyuEYeM3np1gpIwZigFfJ7eAe/cAjsgwpZdUXadBNS9WMJkKiE8bbc5vmPhiECbnE3Cf5mM+uesPOM+TDBD6mIWGe1+kUfDeOJPGHdFfSEpsFDQ3EB1o6h9/Sx8vBOzWWtKApUIq4nqwzLrLCAMtprbHzy1d1gOftR5TTZvo4Q4EqtDIWyfJsJRXtle2Kzv0XjI86sLRmAQwU6s1AbOZpoGOLqZElSUn7lvRy3SfVTEHT+LndWFbQW/VATL4HRmDnl+enhDXal8AvRHVuCFMp6D5d0hIQ51RKq1JdcPvdqfd3tDBGHXTD1PzVlNz59AAu0/nebnGHiONDZr0M9Q7ADO4E8+6KZTpwjmJyjh+Ji0KGLCYAYS91fLABA5HwDI4tr5FvyBpickhDmKlo8D0rDETWPEhMGOb0BYKioBj6N/FJY9HhTW9TAnTgTFfTbYtHhQBwPbbEMSMbL+FkjVfiXozK5N8fUbmNvqW8GLjGZShCMeOsygOm6dOEdzYpBJJoKiv+ZgjelZfMAsWa40fTzUOIs2K93KxULKk2BaBThy2IhaDLTIeQDSXQkpBkDuhXyFPvYL0uSxRsYlO9t0kjj3xBL/d/yE45NX2G2YAzf7HtVo63XIxG/DXYNEK0tijC3babXkMhcbqcILLTc9hcIjF+Fm6ndJBL5cj54FBQK4M0OfXW0d6AXrMq8eEHF66aKcvbBw7dW1h00JKYq3wdgS/KUjVmYIS0CeZrS5wUikAFVf2QIajNl4kgUkzkftxIjuPLyxEZOsXoo71OD3cTLRAcvOl3vEB8oAMBp7iUcxA4Y09Rqj5ariM8raNLqbDsl0sZ4Ryim6qsH0Tek7iLzKhuwWmVxEuHmOkiGig5aqwRyMM2Ix6J44VvhixsaK3l+dYPy3SDipi0uarAfQjtIcYUXLlan9flmLUADB/SHB+a2Sk2Tn+8ZVUPMMXzU1+qj0KNgNm71gdMPerp03XDqYE+qB7yrnK5bDAD8EBenh0El7D5ftgdx4RlZFuJJUxJIaDfZNLV207QPLWD/pqu3HNmeuGjZ4Xfog5ClF7XHHWALvKgNd8yIkEIlD5cVWk83XZzVx2O7QPhTg2FBbcHnU4Zcb2jFT8nVZQlcWygYkrtQHzDQM4A2R3QgQLEP59LUqwNKa2dj0xW+1HR+Qan6t66knHiNGgnDxUU+OeuaZ1uEzBZapCUSgzFx1uG+f+6tsCc5rzHjE8AWtVNU7BRYwUu6uFhVLD5/G+EZc9Gy2RS1BS3p+eM10Bhf2Df4d0re8RE4xtNtWQLrHo/IcaedOl/U8DoGhVpVX4tAcOGqz3xW9vyGiM4wLUmnA7k08JaIcf+8j5NJaqOdAYttsWErJdhIQGMGrYMfrJhYV0VN0AbnIfK/KIqgWmzfh0mBt9V60H+6mhyQmeMbqEJRG4DZhefCYLOruckgfKhb5gBhuGUwKcJ8BcVjBPSVqBRv+gXSqSRl14q61RjtJ3awdw3e1QphzRcj/bVbD3fqZp80AKuAs+fD5sNJz17BVYTKKytX4lC1+GKf8Wd22lCkIZtXWYBw7MAs8FG5059vTUMsvW9igFh+p7Dtd+GqMED/EYi5tNqZSut/1wHyCENWm61YPs1tR91GgDc//OLkbtgrFPpYWAf2xffHpx4JHoV40p2oQxgk4uJwhadto09hJ9rKz412ySSBl0SYpGD+UE9EO3NJcRTC/GaaA4DTOOu277GEZdHaZbn98sUQ8anhlLJjh8PdD82zZvhrpZoOKZdBDqrznlJERC/WDaB63IIw0lp+ixV9FRBT6t1nqFc3J/hxsKnohbpqWGdWpzGvhMxwqMTCFLEik74c1GfRfQSZC9tsy7OAP+szkx/vLNEl3z0uV3rPZCUHuRfQSVs/P53p9Ivw1JN9tgHOvMkIK4lHhJG7po4+VMJi5NkReATRt3Nm0cOVQ4GfwBe3dfX39Lwka9G+EWC7bD5vM4hEDWnuV7f4noXAl1AL1F7xwvzHqK9Pz94QZpEwuPJ/Iqr0YCyTEsJ3Ju1oRMBKSdI3nst4lNhzY4mx6VtQupjrpc/m4fNjE3s1ayAkRfypGxS8TXPEQHjz9O5zE5lFmeGb/+zIWk4t+BsYxjK0DKOUsJ6I9WqexptzVFdq4gd5YZ+NlexFN3IU7lcJNI8m8/7ibpgOmhKsXt2aYqYLOoVuewQW3AiOXWdUvbTWgsaOfW8EvKbXF5FyzOcf/Gd6vXNimFzfvL3qqReV0FKhenGd4KwHZP6WsT6triAKsdA280MBnMefaKzIwS7XvKA9K3TjPa1t0zM2gTeVzOXRu0MpE74qPM2+2REl/RadEauGBZHojfk4vGz5Vl1AioqWKFykOdMSW5g8TPgg7bVfcFChxcqCJ1VW99Fss2AufGASEGvM3+GQ2xtlo/2423r56+VBThxsYwSl41isseHvYyesrc1hEN1SNnUSQIJO4PO/3FRtzoan7cehUmLZOQmuErWMLE+BKU9HTszSBeErhNtlMhsm/5dL42ZTrgHi6TR3YOB7Jmbj4DYvqhcRrxfuv7IXk2HfwtZxX4M9QdWPUiYMuxmx7zI0nSYREKOeI5ejF/FRiCaIJuO4BAsNzRnxoDXFDxJp1/Z0fC3OsbbY5Zl+wctA4RwbdV0qQulx64LMK/ULTMOM/iPyltnhUqdUHTVi5qDAtft9pURg3sks+1t/V44zuRImp/Z6awku7hhLiuh5uAotUKOLGOacM7z0eTC+J2aAVeloxgADP/LV4bzDc2xX8RUuEH51uXpn3r3zSVal58xCSBOuFsJN8Vg81ENlQk4CDt/+XEfkHYGhMuqSjCqRcA02UMUBki8Q9lLcCBsVkaY=
`pragma protect end_data_block
`pragma protect digest_block
20459b596f5cab90b54a7e75ebf51706888564787979f28af06d03e9671a5f0e
`pragma protect end_digest_block
`pragma protect end_protected
