`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
qz2hcTKrEXxmrHfNMQ7qYgJGG/9c6yM3jwJuTQWagWRqRurkyq3TCFnvCh85gBd9W5iM5x2ufqAJsG7n/ElYkvZNFlHILNpIXkNHnd7Sn5Y4RyWQByHA5VlEWjucnvQDbw+PH28vk3VvGqYsn0noZE/rBmippzF9yMVNOEnq/v1vsNFDTQeD8b1RAHDSOxeHeAUW4Do6HANTtJOGdXgIRrxooQXfpwutmMsbGnp6fFrq945iZ8f/2kyT2oV5pfqIcnQ+SKl0EqLXSkeigYZwF7d9n6qWn9tOAMN+wSB6gkUwfsCP8sHcLhFgToSaK9ANo3bjHTD4x3Kahik7P9mYv8zkRvLpjAcpAe9PvLq+1N6+DbgoDuZcDVJQrTH/3lIJn+fp0bLncpZKBMnDzEQ+uU4r4aZWJ14O4eK3FbjJZOYbecVAeeWPNkY+V0dA84rD0s5MU2yeSyZhLkeC+VXkAyy2trquGoEE5WHh+a15qJQnu2JCy6DkVlg8wM2b8auo6AphxCFhPE2InjP9zn8s31ihD3YgIuJ70UCVMX71KrVhKwHsHqOCwak3Pf6dh2tFo9OWijX12JaeIW6BGw6uSqd6O2kwIHZqUzFuK9D9wMIaA/TQmIDf7uybbfxrLO5OPCcRTxWVh7fJKp9V2ZG4aUuCX/GetvrD60bMFWcV4RGbfN2RGtqEkO6IsXVGLib18e/c65EvNEhj7tAUnUxb2qTVFkVMGfMM96vuYhOiGQu1BofF50XrifYeMcZbghrzq1Il9JAxS0Y3uo+x2vTRl0+3CI1lT39xRyJ7zL10R9hf/61kautBScOrU/LIE/NWRbMBZ2X16S25BGhUsPREFoGmfY+8UnYQ9YrUNASu85Z2oQaftgjwOnpc1jz+A4X/R8HVB7TeT+hLg2iiN2IMkHyCxvH2HNLky+umBHAgLQZBoDM/M6bM0aaleyGGdcTMe75xIUX9yxzn2neUE4D6tmS/sAIdpRFjoYDzX1d2niHBuUOyHQwM3arGvH2Apwtg8qnq5T6wjDvMMVM4UYZdFU2mpGWOu+m/XuGKY59VVoLHa/xyFA/+OEa/3eKuEWSrlgpRhkrxaBXq+4lRrBZ33vhN1MMpXwnuOTWVv8gDIeRTpnSYPnpt4xMWKFnNBQearfO8n2Qn1TtIb4RQlbDkkLnl8PAywzpiT4mR26veKf6EdZ4jZ4688/TrDLjobt0CJ6ZtYxX1cgGRlwZcV7ZQKtV1lvsbnmU4YIHYoA6iiEpeSE+TwFjvFu/fkpuLISIT65fGAs5mp6ttZA1eKZ3t9qAfg/51rNyxe93EjQ34FWDZx6LAhfyxjhYNJQtadiS3AO2Gyhq1eErLumb5fMWATBnc0AeEgP6iSzH6K5rpu1/tzxifcqIUkwG9rNmZv9bizmtf0wZk38xyom/Dth67FJnoLA8YHEF/3gHx/5cUiLdZsFSdYyT53w86Z5gwYxGa/HL3dYKifvX0CHNiPygEnuGyDyiG08+Li88o1IcZQpj3IQ5Z2sojyggsHgTUOSp3kpnbCGvLXkEkqY/CxzrsF2ytSqgdZdV+Oj0leWjR4dLYQMbcZR48Wf4Q0slXPaUhz9LuXnLPrU7Z9oL1ni3enlqqplwt6ZgaRhMriVcBNEfWtPEBPhwaQ9ZoDgnV56aGNmxjtcLidDicgpRI1rhJ+izxRhvUy4vvnMxxzwRfZeWjcUebjs2dZXGhjhMyaPVxJF6aiaNU/7vFzpPv7fy8+BEt4fd5obqZpWXRF4V4bQsi9osj35ceUZ7BNz54uaKB7Kbc/pmovsVw13IA0/+W3yl8KzKEdtTiVwMPVgcjVKGPjprGq/zvAdRfudaZV+x6bLNvx3t0I8v6Xaqq3zAaZRLZ+7fyPLUvtygjRC2Z1ALZxSJ+vFI8txYf1OnyUMDmtm2lKJwWx6LXQsJhL1ddM4kE3Ssd6ZpReNnppFVx4kggBQrAHnEUToWWEJMZA+RufejNq2WKxIcGWVeeANq2nOMd0qQdubkGASW0aRt8Q/dsIAWip5KNoF6tphubFt9NVUqWMLTt+3MJykk9ce4BEWfU8wwQkNUm6fnzI1rhrnI/EVQvQNBe+6zVtPNfHGO89enNKZa+p2KQjK0xC5luxQiqlXQ5gAQGys48xKa6xybtmFwYiv3cfLtxdxaFtLzbW9KoIW8j1L/6fMckLi1AXmoIbTUVIIOcElQ6J5DP2FsTwiV9vShoyvqL7C01mQuoa/uI/lOKXHPK5dOs0fxIMVPFpgzswwl7PjEBPfn9aPO4pK1SnfQW58xRUMJHNuYiYmvlTy+ABsZR4cNP1P8DRayk6IXYYBpYQmwu5ZcivQLbL6ZaXYDYx2VsDTJidaxu3bACehtgUDwQz5u8KkedaYcThz9PRq3SJ5xoMF+/r+f5c+cBSMO2q2u9hMd7wNDigxZ0FVhDhFO+cAnkQsnCbK8iBqnzUCpzQHy2Ewf6/UDQ4coVp3q2jGfNBudutMxjgDLAAv4ctUe8InQakLpBpYobGt1tSXYu32E5FRDK8ENQ/a8/WEdMOzLMrXou0JylyPijU3iINzERipL3IRmWPDg0aKO4oC4VuOm+QTGfGLOVkBxppd4qbv3Tz9u1zXonGaqKFwFl21Y5Zyv4tvGmIF7Iw6g0op8gEE+v+8Y2YO54o3OAukHw1SkBnYxV/x92Xbp2t+5hBjDOnBAFdi7FMUFBgNFnMJe57F/tAdhyEKelIiE8WLFC65t/DMr/RIPq/edEYQ4JocneKuPKGqOxVwdYuZlxYdnkOM1/0rf70BOyUNFvibDVK8/jmOmRFGx3fO/oc5RKAXufh15E6YlwmBhSpLBfJy4DL+bfawl6dKslnNhreFVUounj9w60bVxJNwso9D13how/B4WUnREuZjJtBsYJf9vBGjgelNtsLuM4dtJ+h2Nmk5ajIpz4RfuIBJ0+arcEKyaden5futawChv9BLA1ZTiAuhU4xjRBbG/GTbK5UOiXbPW77lROwXEe+Z3PuqFaSCefXQ976+gyeHWKivXkoQRsTwnAT9ER58nuTsHbQ+xC4vX6mO9RRCe2ODAIa8wZzaL1nOwcjROzQwhenvM361ImIQrzNmW+XbEWys1o74KPPm+6eVx/JEBfqu+8+zgBBCcZWABy3jJueo6S1RSZXVAiL9+konJW9DfAGDXI/qE/Zf3mBNdRUjUMWZ/eIK6y6QqpQWRfuyfuiPlr42VbP4CxR8zZACCNcr8zFUKb20I5C37qHThWKTYpWdCAs6AoJGazjVUThZEsPf1Uu5nmAtkZ4ZV8gil70e8k+6mO3K4tNBFWBqDXSSzZe0bdEN15mFWFbQc6Z/lr2lXu8lx+cc3oqZo7wwXgJVw2aeoaMNuT/GsVzgiSlA6VMkXmlAG/kxLclOF2P8nserEAxBAGcmNT2p/uZUtCnJCxh7WezP7oBLPXFBvYMDp/VSYJnYtx8mu6Quf/BUV+ScOzeGK3uHniB9FG5B6PmUjXjq8kU+8UtVg142aGtkiIYgAmt13uQ6VGJngaOfLU7ze+BKgG0yaxHhJ4GYvaniUWUWir1UC5QE1h4RUUecIQGVrcyeGyYbq+rBiIszce5VLE0rQ5v8aMoEZEQFj1NCxvq60ivw9Y7fy0SDax7YuuuwJbcj3C+zWUawoWvDMQ9xfYOgGqsDmu7vFCRBTiM6Tm8SXilg+sOqif1jEmCLZ0DSkl8hysC4msGRLOIencCTrV6gDXW1rlK3/MEc21nhy02kkasXoeIYyMrHTPPRxsv77Fma45r05hraR7yl7/vskioskk2wXDafkTGviMHjm10PrV4fMSF54lI/z2wznxXaLe1i/YEome0+/gUiXuwpjdGq9ILzS+6GEUCNQHTruZH7EHV9AO8lggwOvA2puNQPiktG6BYc8w3to0QfNT9VTTgo67mwsL8oVeU2bk/UW/Q+hVux9FsWgaoWrIJxU+gjO43ya7SdF2PDzWSXf0WY0jThODOYO+jKOs5qE7xejHIxylCR1dCcaSJSygId90Dalz92uGwxHUo2Nc/gHYvm0VXFCjFsaYCjKm0+t3fBaUZBWAm5iNwfjB3U2niD1AVZc7kFZMYkfKNhSidxyDMaMdAplaViE9ChZgmBilDuSOQGmfSwDcZKb+3zfQRVqLtNEh0LQ+CnNNZgP52lEeU9vta5LEKBpTbFna4LbCOD5UxNqWAe0m0+k2W7WDSNzUGI4c+UiT3hfWHdZN6BVe88RAQb6TAXJkanw7v8fcHMBDSf8ffVzRP5xAtkK5xIRBxvA8JmC7YuWYdXCVqcrRgbYFF1U8CS64rcgpGgwTHCtD2O8TE7mD3pN2HEPlMdwH+GNedKc1ZOrzBDInV2InwHS+7ksytHkA+Lv1KJQODghTnH89U5UKWU3oM+j1nDgxTKtvVJxjLcQc0QeAp8QhzUP1bul+2wuNJSlDO2WvgdQJnVtFQKEs2XmchdENg4yXGjeYLUzghNBCPhf14812zKAtplRB/jgS/jCveRUpHQ1X51WGYUQoc8Adqtk+jaJNaGZadJQR0IQ5ww3hp3yJA0ORhZW/rhO0/jcpfh7x8nxpr/uAxmT/MY+J+mmNM0gjpmwOi732uv1TlJiWydxHoHJohqoPOLiqM7NslkFXdJ468R/DtxBTVhwkoTvFHVBJOU2Ey8myQGAEiGYCp3gyDLaWKZyM57hH+f3JJG+ulW+RP++H2TWbmyGG09VAcVtWNk9EE8Y0wW5gmZhS12il3idr/rlPuVkz7u6CtJdiM3w6bIDe5a4h1OzyFhFRd3wd15HeYzMCLoTsAgqU4Kc+9QtBw//lEElWakCZgoVO2ZP0V5gwbMW6jfrnvwh2NETZSSzRs+15/HdM6MlVYGqW75+9NGEoB61KcC8gAprds+R3HwlRs5QHWpZY9V2pPYaNrX7Zmve1/6ca82/VtcNxqKJLDFfGpIJvN6Sx/jT4euspvFmoZhm+xMaT2ohzZYNFFrl5+LyUSC3wrCIuuq+53qJwZ29svlF4Ao3sJEeQNLgpfG22SBMuSUNVEUHH/reetJH49Pjnj+KC3A0SGw/0hCOzprc4HWMdxxb/64UbyydvERxEiIfifFmUzobhfSoGAqHJy/nf4q3vbhKSOYzwhesvVcrxTrPTtSa6DctP709HZK9FkxNshrzahVd2dADtLcI0pk9QBqaCQOVd/wdC6guradxHJECAXKTwhCW8Jg3c8hOAlnu68thmUN/f7OblLsbEWWDD+8HhKLRa25VEHpOASK2tmPdlW0tj6H/Qh3GRsIz5FQMoBTHyv3XDEzHgrWS0LvDlq57WX1SMK0zBCn5CucsBRZNXNk1JwaZ35JfREos+ZDLT79t4zRBi5lqwCTZ2elDyCo3VWjioxSia8U9AC92BzQ60kVXrhzzx8N/v7+LVgl64ptZThCYJlaSfC/R/+1mBJVe6zXCPAutLm8N8jBRhqyuRB9jxGLtjMwlxa4T1MfEbkFOKfVNaT07cWWutiye4QwoFo2Z+Sr7U27pf+Ox9I53X7Yn//WKFN5ITljJVhCl/Ey3tUsIUYoRSfrqY7ERrTUCkW4tnGrj8LxYW9bJDTKD+pBEeXR+Rnss5XMSk5DQeZsSvEpWU82ZkKLPnBJFI7HD0kn3h3D4YNbOR0N2zdj7/cTjIB26oZ+NVxmvAW9XQwogqTBBbn6UfWs8lvR7LLT6nCdIvOzVIoecQVe9Eb2mgQb7OnD7+p8prtJlA5la/mGsDWNHBTH0WVbuAg/nQAq7W9i6uIFehMB8a9jC8buJ+ctdGVYwMADA+BRD6EC5GyvhQGwD7o/MGeSBVoJKFkTTO1dC7s1Q4an6zvrRKIXo3E0U11fJaAZa+5lKM+mn4SIwaryW5KhMmF+PpRcL4rcgjCf9fitHd66bNuyk3M6Ux13I9JqRXJReiwNiktyfgNl9wS7iOWTHYGfH8HkOc0qFhyJ26s5TsoU60yRBMf8qc4I5dYfhHcldT5FhpFavBjx2PLjoHk35NBaEj+RZlZs5PCKLb71OE5vZr0UU4Lr+JMX6qphi3bGqIsEjfElW15n9royvZo5i/MmQdbRqPK8k+3Q8qJ95J8RIR5eCbwL1qYpkirrlwDwqZzUMB+z84HaxWOe0YGGEp80n0EcJcPLG5bgkz9kp0wq/udbt2XKuqmodhaObHn6ozX42qNT6ifxEU0XLShI1lChz4hRIVmX13rrBAAK9WL5fpnIqhHKX/GdzKeSzpXyVvTdz2AauzNdJveibceMW/x0bHaC+q/FGC/SzwiXnkm1kaXBckQ1hL7/c3IC3pF1jSmUw/klbI4OEjhcZTtb/UspVJH7YEB/4ckTKNkbxucmWHJbeIv0QcZMppHic/gbzX0zaaXM/tgIguTXJqitLTUiDf5jFcy5EieA0ms/s0dZpjBJDk+BWhyZW032Aa4NQKZ4sedvktSeYqMxgtrYoAqYQdobM+5gTnv/IFyueHTAS+0A8J9lRNy8i6kPzg/v8xGjbAUhdBdsmjG8eS/p7CDZd6Hsbq/6mHlG3TZjtc+uOigwSCxRO95AGTWyOwgkQIqoBfPrY9UWbE4X06lGJKpJqxyBkY8SU+lgT+oDf8wVlx0jxscr7Cd1QvOCIhPaJB5g9wB2yG2eOlUe1DvLafygkXgrNxoRnY+Jc4f3RZt2dCiB6QI1ENDmT/akV7z/h0OvylB7uVcHc13LdGTadobWwtQx64m13TagAXqopbL0npU0dYNHLIrT4jQWTKmEWcSlmfAKe2wspO1/zpXWvQSli0kAg42i5y7Yj7O9LUDsio76E0E3/Xpr5W9B9sjpk1Et282lBldVz6sUcZtNNRcF3YznYPVEEwK2XDJ/Bw0WCaX1JLARZUJTq3DdEna4zit1x28SsBb7lcZBZReQsIp9XgXGa0pgDbX+Yxa7WvGs8yPKh7xt8Xr+A2XEo+pzXQp6hcsMe+vq+2QWhIjuZD2lHogt3702I5JpC9wqIDyEirNzhZm365JO3uYMk94qgF6LvNVGvr8E5k/GxJwXZvHKtgYDCWCj3nMrXxNt9o/2zBdaEWT82Nq4E+ny6ORUXbfMvH+saiW4AeXBMypPRUDAOMaAWIs96l8t6aAIF2gxGfKvM3qIGfJVloVSPrUKys/wrCd8eB6XLkMg/ATIhG0+oOwNaR1Ouq9IdNlqQa4cnD3Y3ICol7RTUZFSn2fK8FAJ0B3ABUS+PVr/FM9yg/QyX+bSXz7ZuG8pHJn0vzqMq6r3N+GVUkO7gsl0mawsLVALijdHNiPCVSNcnWG+Vu3s4Y7/C1kusEVz00uNObihJjiBj9kelSaBU42XXg41XbUED0dsxK5A5wXof912JfUcvBXTH/I7hKhGyfhY76XspTY4TbF6evu1Ns51u961JNdpFi9K4ja+bdQSjiCi07mqZVyGpZESom5GyBGzuTZCo6xJ3LHJLjcUiLEFKvgkDW82EG+jlRSIR8UjsVhU0/U2vcn6CTxRjyXcAfuwED8F+3CuwIUL9h8X+xPHOka3dPZ6xB4ZUk0lgrFZ10PrOBZXfAojp3etXOUyONr3ALa+7cy2S4mM2AHPh6x6oD+1JJ4Zza1i5ywMAisC3pGM6seD0ADqAbbCQA5mDBLpz5WxSxNcGXhRAnn2Y14Vfk0wM/szZW8OhTxA9ZVfTsZwmhdq4dYXRizmcdWqt0ebxMWNVqyx4HJea+W3AnTRM560Zga7a+LoLuG+x93vJQGoyfASPgFt6Q3WLKgNCDwE3taQPQQ9MnAYnGchnompHWQP8/bu25jjFWkXMe+fyB0Fg8Cv4AHj4JWVMyhNuNZdxYKOQUAgyMLbDy8KH3etTtFeF9xgno4bQkd45K+Cp+IW7zK/Ug5gAWsiofSyVxUtHe+AGwU3ljjdEWud2ATxKnT7SGRsi3uZS0BHaZrwuhIKhxCogNSmm6+ix6PAPt8/OqdypqBD9nKH/sk+YNwEjHcKBQ4Jskz4R4NZSL0UmTcsf/anytwwIdzP1ErQ16KwoMPaoodebvAUCZrqpHkaAai96JqMwxZVTy8nM9Pos7rOX32JyfllWUnfqoQxRNOu58sfKL4/5phk0rGwWzw3LKkThCGmYLr2NwGvFsMlRjdTlTLFnFYVfykxEnXB/WZlYtU/OVTzApdzBcv+Pl2bmln5oJ+ZhTXVSx0yz0UA7tw17jYGzrh2oWQ6Z2W8Cop4xZf6zxFqpBAUmrbD/vPaTPRqkMFhkb9UIbxXKzA53RM/Wh5BaxpS8ScBr2hzvcTSkma89bsLn9PtChw8b1aoGZmgV/IcUpSwMgwU9zcJs4HOqvgzZ40aIIsiudFeFc28xfEEI0bRd7GsPJV73jvI+/xX9JEapkIj/C0e9fKOiTKonmTGmv3m1a+hGI0gRfv2EN8WdNBx+IzLvbvKeXfiJM7zEOMu7F4kzH6OId6BUGJNEAOyR24WcvivpdXzEwu9sW9iaNNuv96YRwmYLZKXkI8Eov9VYUoHdh+d9VLxbfl92k9908jKxq/oTKzy3qfpyos0OyKxKJ0S4JLV+UtiEMYMVQl+xlmu9Ltdw+7ruxi81x0C0WtfdjrXb3B+b32JcEGRaQS5olTkbRZyMTkLc6Qkn04fc94qG5LYETrreDJdu0ErZiPAZGWe/AI3DbUw8g8zZY5LcoF2oMBWzGcxWO9+Q3X1zqA6Eqw1LXxzqRHc/jkjJ79EYEuDlprSCBHkpcNRDRGbuNYUKg/Otb6WQWUCaStcNu6HYb5pGtqyIPgbdGIgH1h5d3B+MNHJVStIDprAOu7CvKpGVSvBX+6wbGvDcjXYZC9dMs7hCT7gG73qQaWGYnNPnRd1qJ2FcAaJ4HNGixIgNLHWz2hzL9jaFarD8U85v3vlYqw+23g900j34FPSSHRFXPT5xZe3mRKNUBeO6NOkiPbFk6SEIqiyVE8odVEXDRYmc/NaRKeBaFyAi3EYy9L1PJxPU1f+XbmrUPvOc6dAolI+2aqWdiPYo3QW88K9udclJpqqqFVy4RWNsJC6nqDFXFJ+Zt8u/a4go73iCpdkzf46XUd4ogxBqSFoucLC/l5SGz8VfrKhq4Li212mHfgMyTKk93KzSDdD+kwJrH0B4pPaafo0MjZBfbRLVS84XEbq5ylRepXoLJH5wPs7i8KzwohsoElbIGHtQJ3lzspsqvPv83CS6PEjv85Dr5NDF6FVup25SiqZYtfzhSS9hYbFtZqiHeMcL0vlCz9z12dVdkawtOrALM46eamffARyCpW2jRJUmU1iulNCB0+nnv+7LozCqxvlIF31lZTwhasjT1M7BTEmKO15KNMik0jtXcpujJoQB2z8vG3LlUVUXGh4dni5TVtA+Ylr08EYq3KVg5xVEIkpHkBZ/bcwFg4LjAC3zZajRTS8lBPbXHywyTx3LGTq4fAWtJz+ZneOggF15xTfsV54tti07DqDRCqlKvaFh3DpJDXJFT237BpDhW7GP534d4rbq+e5jUNN3uPYFWqw3m/KWnvQfMe40TDZiSuwjQHKk9fZtGPGZO+0X+ITVpG1EVXA9hCNO5HX49wB2A0DZN7u9z2iIG5bF07WE77MBAMy0raoSpghCa122LW+2pibBqBBMjsNc0imECd87QDJguiqPJuIXm3O/wgWv3rafJUgrxtl6+lwhsbjAaR6LGqu+XJ2aNHS/cg8pU4DK/8cszE4pQ1aIegblgIL2EqrcbVHPwKnGWxfkoGCnVVqtnQV4m+Zgt6icRvGy4fZQTwzfqrf1qjKjHBxTShH5IKAfsGQJdD4hBxEYLt/SqljlqmdP4EdrZWMCWD53ku1vIjawKKogo/h22AaTupdRLSZdQ8fSY8n+lKZb7trjNYtWfU/aniCJgueRmQLbDbSajJXJDZGPS6cOaXjiM8MoP0lJZVjoJzrKhV+vtQzWtROFXZeYk2olgabLwxBDsC6YoIAyw/XhlpCtQta/311HVAKGRwBqzbeXkxhkuBWTGh6ErTTjay0etYEx826R57fqBIMk967qVooKaBKJ/mVatinHoYx/jPYRlRI7T55dCwJAoo6kqJrMiHJwi6TYhnkXS6qBYvXQySlvGGXR/huRUY7+uRkDOQy+1cyeoi7j3SaFAt0VVUhD14eKQF3yFqOKv25fm1UDYIE071Szwpz3h3pMyjyA8WR/UmATO79+JjlSavyUuep1VojjasfcV2wtpDdK7tNEN0b2sHI52n8hSPbQ/JOe/VudvsDf6n10A/l8s0Yi/Ph+cMt+fZl3t+pNCrZy7MGMkdJRRKIeFN2ixozW7U5hZ/pExuBcBu2hsrM5e/AvQzsnMkDkVNz+zehvdhSYNumbIF7ETH8DgybdjwUoqmPnQ6esW2uYdK55PS0cw/bN5Z5p6rwY8xQZjy781XaV4JvrVABV+xSmHlns0kE2KZ2l2SUoFsXxWOCfMGAYVV69ILYobqAfpa3VWfgsxOzidMumhmEqZuH/OospsDdpX4d7QiMYvT9oQvzTcFmu1u5U15FA96W3iLDJ3ApOCYhKd6xFOzdKR+KcE3cRBoVAIQ46guD7IQPn2u1d9NfjNZULMkwtvq+fU+7XyHPmy6ElfNe0bVDOlfZ9yj4tGZFY5dLrlPe+lq0/zYSFBogpDZ/UZORD0VWTXsdNiCepVo353epPardr4btBsz1IhWkHVDJZYVMbMNL8CIRO118O+hhgnfJOM3vXkarbM0SN2ymQLuWX6d4HZQXrNYXp5/UMmbwArrrtC2OQaYT+K4cptP6l1cNb7FTgAjFTRTsPsad5dDV9yteLFg/rCl2RPoDZnDgh6boMlI50qjXFtVl3niLu3Ky8o3DV/IwqKm0LPaJRdhStBPF+xfyFZBxkjJ50bsZM4/6oZicop9A5CU34qIFpxK+qX/txfS13XstD0jJJYwpyS+dZ+NQIg9GW7Ry0SCZBueU+XwMmgvGT6dHFrCFC7frBZ93q6vlGnyQaPn+BJZ3+qhDR4DeucL53k1PG4dzQxTMBEvr7ijjDUn7y7CQkTx1o3laG/LnKrDNexM4q4bYsJTeNNKoLv45bWhkT9BeDQCM4qyX1GEqi4Z+o7RP00aBZKONB5xQF4jAbU3iC2Bvf9enKabMr9KxJL8+ZFXiV593VBNw8XHNvXd1HwV8ZWyfBslE7bHZII3Z81u8ZHZZxe2uCKYwEP0YJJofvOz0GcJn1XupmT/+kS+5B+bj1XewcFyC+27XyPauKGFpyJkMFuAf9FGR69A0iEQ/nsMHhzB79RcR2a2CTu4smMgOpV0tckDg/HVKj5bYzR7EvUWWvVkjpxG6Ki3WELm8R7m7tqz2Quomy13/QfN53kgjFKftnslGfS82sp5/4xtJxEyh0vr6fbBDpWTkCIv7faFjjgjbCpQg3qh6knKNN0aiT9S8od327+U0s3ENPztiCG6AxS60mxGlhrq9K7ZJutbpL8UUm7ER+/QUlBpCDYRy9MQzD/ZmO6kKj35ZfshlnfO+A1dcit/5PvRxAXPnnaPvwzpLQXH18CGAWwfuPxJRoSlXhVUFiDCvhjPW2ceTDs7bMUOR5Mzq41ZlBbdVCAj57WcJOqlB9M0a6pB+08f4L2BBJ85jCRJpIjwxqzcdOrJGD/WYfWc7zkbHX9YqESZT4W2pKf8U6QXrBVaSuQAh+kWXMamsvtdsh1giq4aMbhhB+Tr27oBBDQInFVTVW3i/VWFQ/yYepGzMkVTCCAGfP4VeoytNM6cBkYc0d6AwUbWCyGDEtxjNT0A7xV4ReF6ut1dEHBXlS6KKjk6NkXGN00UV1Zuk62b0UMmWeUybXOXUTdqn2JDjGAH6mNg4qaYUxGmXV+kEEQCTtJNvTKdqlNI1QCfxfBj7CC5SpAIqSCDS/PmR0DYSkFf3AnnhzA6Y9w2gMwfrhEVkK6BuoJcnJ9Xp+nA1keK4szew8EmkBU9Muts7ri3E83/++2BG+HFyCpnep7s5negdLrEjOem0aJ7z/clS2qHZUZ8GMRU8qo85QroKJy2/bCWdzJfJHv2c1eOrbbbKUJcF0/4Nls27E/LRp+HZCHY2YS7VG5n66P2erQQSFX2+p39Dkt02EtCJidyW3uLHKlQL1/VygSZaUdhPc74469QI3yfjVXOeICFzzC5u5ypzjTHYu6z2ppe8QSkhCd1KZhZeGjQkzN+71yMW8oCCPUYRTSsMVGX2/oOJBaOpH4OoMvNO37Kh1+In+a6rs2hTQmzIASr+DLxTxg78KGHzOZrmVyQ1143NQA1Klt+ryailZSptQATdN6rmlmlIl7OvMqgU2v0WyLjHmz3esCTLt1+Ku4Gl/zRDngzUzJaAYjByc5sntUUkXWLKbNlIaPCAorJEwqGOpI1T+fQ1SpUfnE2XyaoEOJe1SQbJUy4ZFyFfCMNZazuc3fKokyi0L5oxJLeD+3PeHGgDIkIXlDu4oY6J0MuzP8kD4OG/Rcxiop8Pg90a1LVuFsV96znBqdG/nK47CpSbJMpxlJyGfhIV2ih7FmVP6OaAu7XNPzMbXmdb8UgqCEnjnQGZYuciTCOYoQBh1FPidah8kOFwVtrgaIGEg5MnXLMGruJxM5lvshgsC6v156K5mm6/8O7NyMt+alkksXufOclFlO/GYGXErPcihN9fGKKCzbytgsY7cFP2LBdsTku/Iiky6pYFNPvjGyDmOw42HsWpZANxv91fIQLuBxpFavQkhLFMkfcmd/UAyjg+0vgovN0DfSf6NFTitoCWtY40gsrnpUvQs9RSL9jygSMH4dIgAMOxwK9pWynd+PwQluU6bFYVfFVsXpNrIwq2GbDptdyKRnkXZq8jnf/FnaI+Ph3EZ3Cfzd+XOwPhYJaPs5ssMQRvEqV5uZearEu0HLrQCio/8W1TA6yWMa70mdKzyeYwNm3wI0Y6tWAlICMbsY/8cUw4nBy8g4O7oxwNZHFOadKsCS89IB/xQlOSwUw49pa5TJjk9zRJq7/a8iNz3duI8ekKvknOzbsMIG0OBzwin6eEWEnCLx1fU/Z2URXX/YKHfzTXDjRt7/2Rg8eqtp8bKRhMgkdj2/1CEZr8pFAIx3SPHLaM6tktnpY661+l0yaEk+jUYHUD+G7mPYQnW8RA6RI4H0t4D7S1ZD0BwBuUvIWcdgJV9YRbLlU6hMoH9+nebWhbm2vy2PVzCQNwVSILqsIj93d2a00j1ircdf9u6kibozAc4ro+baYbNZMx81PyCaNCdXIaymzUYs+QCmYYtT2sGz2NagPVJembUu9kgp1Z/sc6ITSWw23h8DMElpWSq+68t1sdu608zngJ3g9Q8uf8FrykERtTcw5lpCDl2TG5dCQCHERJJGXF6AGSMsbP4wS/WLET5Qrde7nzK+3NqPvAWHA7JqGgjpmKXfDilnMaC+lfTM1ZsQHcFHAhyGVkgQgPHgYJ0gkQLXRxzLZGor07yZCxS77myBJnSCNUQfPuHZ9XJ+AOaeBrBUtTqQdtkXGNNyta8BsKFn2K44VXZF1xT7CNXRT6wVY6qdTsLeYbBcYGY8rSWvA5Xaz04opiT5inv2+BzFAaw+ZOOSf05w4QUb47uMAinzgZAFiwvbV34dOGToyzCedSKPUlUiAM7rdJw3bl9BwsHyZVcqARPmGW9lOizCxqzLRuP/JJJa9T0nwjFkUi1hQHa+Bf7iXPSSu+2I4GMO+4V2eE53PlS8k8BCQDdfhicL7FGoq1mAWLP8wbKEMTnPiYgC5x/bipDAbdCIXUV6/h6vsTouXZD7K2JTGr9kGKbr2N4CjjpzykSDM50AufgZsKPm9hElTCoOuy1qIJSxMQN3/X45kKj+PmMOHX1twZPqT47l8cceNqZZa3SN6jZF4wr6Y52cB8e8FkHJFjgNXvWRx+OIEHuUMydRrRD1rLbZbW8cSOi0dn4jsehgzrsy5sPyebnUKnTT8Cg/vWlQGxUfn2W9vZ6iPZ/CpKeWC4dHM9VDtCL9D5iCfDasw7rWheFA/p1flrqi+5VjYz121a9d1RNjdnx4K9myN3lY1MTC/LVKknnhDIkY7t0K/7KNar6ii9duJusIPWsSFeiuFXwHoySfr3Aw6aZ6hyemnjSOQcBwYOmgs1sGEkkV4jSUVjbB2xdwIgiD3UxhVRUU74zUHZKXfe46N0Rxz1UWqegp4Xy5YzGiLGUdQbsXWXqtUH6lbxXQfPpP4z4NxOb6MMzvy+wMcVvp3FMhq3Nfy9D36mK3lUo7um0vPo2vhixKPKVtqFIRexGPyIZfqJRZNvexROaQOFdr02Ew7JWVFRMVScGkpMm4hUu2UJg+1ofjrRnHgrvVUkNGginjKfNORS752JDU7GHIkTJoK0aEBDq9oWEYJyh88whtHLoULQoy7d6yywJZqPWzkQ+s+buJYkhYHQw4QeL0YpBTZgZgUnEMRll0j1FGPD8nHi1k1jGChNfmrozQpf2p8Cs8bpQ3fB+OvG7/pC1WjPoK654PLaHWnLI2+u7uXwjak589SScZj+bKLFh/RCF7H7NmI1FqiY5sbxCBhYVGW/jdO/P0t5Yyd84J56osrm+KmbanOvUzCsZ6VU8CItnYf1GOgyx3vEnJZsNU/iXl6+6NswlERUnf5EFof5L/uj0UfNQcY0VwBhwD3rtGhjwWoth8A/V9oaYg8Jtu10Xczv5dB4LMe7LiX+CrTACRXn8zx8jPJkvUDSgkDDxsAoPGmVZ3fPVCQ+JWj1+L05rgcVaH7VwJ8zy6fnJVytrM8EFoWAmza++6yCG7sKcpmGMX2kRGhtROrrIftX5kQHR1flpGuWMtVcnsgvCzhy0yFOIl4xuUGJ2CHEKJmKNtJNLdCBDINAPVyxeeCzr9iRqaZf+mEYW9acYzmmSYd3iPgodDjMkw30zwjnv1Rs2EueWAhuzM4+ZKSpjcVsxbdUI/7R+Nz2IV0kQJDgMOSTH+/P23VJDOeWVL5ow9d8nnK+x8V6ThwZvSWPQWyinUsL2F/FeIFynSv65tcUdtMCvS0OReX5zJYbzduGrQtFwWU09CYStRNIrnUbKT+N8KBi9BrqQzxx77uXCte8y0JXawD+2gGpGQRKZwAoao42zcJQ3ok/fhDlRQTLIoJp0AKXvuS+ttjAjA3b9UfIxQwzQBTy3I1qa2yG68vNTVHezNv1ACfshCEe4ByfRHt6CveVYTLOXq6e9AZ5pld+RHjRcPcHORnWJ1+dlbUUvcgPvaoyVpYxx9zlgN8KgjNAFzwG/a0ZYRhL4GeRYS6l2vH7Pv58Xep75VYdflBYFIAQW2xC3NhoxJ1rRu7Ln+4W/mnegNTn0ONcsIqGqJqcA4rhymeN5Hk2Jqyn8ls/xShTcLe9REfRyE7O7etYntrQ1U78ZSJte3zTEj1WOv78Qf1MMAhCNKI7rxDARs5yLhQtotKLThpjFshkPxzrolsrxQd+ugle9wBrYN4bCexKOvDgi4/MKP9y+yTTllkafj9IOkl5EpryZITOCREnU9UnoWOxCzUH+YlBtH9SQogyZBLTM3TDX2AKIqu8qF5ymmmKI1XwHr/aXEPovk2zGlHfLqPDhzAEp6OjIqc9k86b9CTqSkRbIFsdVhFHfkkuQqfytTJfJo45vR+VT8NaNb3R2L1Fqalvt4KzLcvHR6B0e73DXpqQy6hNq6UXmoSgZIvqEfBrb5wvBqfelauYncSb4OaL8KKnD3QXvfriAprg8hBbBotytuLu0wbY7Seh1OoRlhrAI0iI6oI2wW9tLGvMqBPk+tBb7aFjgRCSTS07zK/6ZTkBV9G5I/IK2qBp9EbFbsGcdiM0NU1rbVz57bI0eaV6+cZja9nDsvEmPuDTdlgEDAUs24KQwIdb5jvGKeIPXMbHbFHVHHaMxtrMJ/A44gE+VqXSfQKlGh+ru3Rkm/Y61531VJZbVsIFamy/+st0963iFmJfaAEav8LcC3Aug1c6x0TeJMV+0GqVhTDQtYBWhq+6B0skhgkVIL57MzWnFziDMd8iXcmZswUpfhVhlm7Y/LE9KJ6VNqLLlMQn2jP44VwM+SvhPzSHY19iFernMbNzu0UB81JKtPTlc28onbdkijNY5yRuw1TmXmbF5j8FS7I7RY6uV1SFixg73mAdaeAZGceBboeJQGsDYFs/Cu/Imfo5GzGhiGc03GcoOV61elZY91OIVEzmbSBMx6pR1EisRng14jCgMzHG06UblgH4RR91KddVg6qscJlR+JoJouf64BzIHzzdTVoo7DnZd3nq+FuK+NH6P5M95zDpDfaCMHiRQWxs0X7cNKPWSEmNoOn6kIV9l565cAR/eopdjVZdYA10dsdVbrBUfexoHhc+lH+hPDacYyMvrZaMH2Abrn0lgkX0BAN98pEs+TT9j2oRnUfRFscExK6XVtHtfjlJC/+yDroWpgFrG0ztznHOiD9LlHVRy9Bc2ChGJY6O0JNn1pJDF5z0ZZhhil8vWTgjsa2CY/RrC+rza2djlatCfiD+7qSZ6qb94Jd0UZ19SLZ+qywz70lp/q/Ldhk76Zc0QV1isXLZsL4y4VQ7eH9lhxqTmgwfyM23VMggiXOp4GlEoorIYClkZ+VpgjPtUofxsXWukrucLt8sN3GbYNGMp3iBVi5Gs9i6gZaK4Fxsz+KrMn/wA+41ZE8LjNiM3bORywcMAP/V6/C6TaCf5BtfM5TdduJd2hOPNyKexeWqQfO0C1XShHHT7npoR96Q1JBoOJ1ZSYkvnfAg4RwJihFkIoZA9C3BvdPYEU+wIavHhEAd64ZUHeNZymY46TtbJHWn3D+Bn8F+Bf6R80sbSB6U5cGPrSYlzFtBvpau60qWkJQMCBVsKtbiqBEkGD7LvbkTE4DPWIDQS5XBl4S3tiwGTxanYaGDTyu/t2hvEheQiR3omgSEAHlYNA5/DLK6AUH4A2l/Arm8av4yTF/GuirBLsa6BEkaqETIfQR5ts6Iz96FzT6S58r+DcDPOIayNbb4IZmdFmasSmTmrtNB7F5lDm/oKOVHIwrOfBN3cohmlcGxOfm30xGBMjua7CD02WNj33wYPTDUkrS1SYtq6rw06NwhGSTdpGZ8rXRN+9gdhas45RIL2hPoe0dhsCzRRkFcA8HNTpb91HlcvAlX3IpyocY63Nb2GSIOMujSleahGlsA7O+d4dBJeIsGM6GBWhRAcz9irsZ7v6HsFoKY4NCg4ALUqJybho25r2ByefLXPI3C2PiiMxCLAAMlslOiT0XK48hleiuBM+qhEAlS5rf8Z8s94aMTLkxPUJo+BLMfkRK4jM3rb7+XtzBvPrBfmqrr2pR1LnzBWc000JJBcOpV9l360dH42HyxZmlRV/PC73UfmNF9nGj3ELk9BUHP8MXjmMCp4AP9M9RvC2ZP1EjtWZjfU5ELqhUpMdSPXDD7jkx1ckAmBJPZNtHExFhZkdUeDwCOsZQ01QXNz75zYQxgFzF0k5eP50/QVPadTFt+oyWfU6StJUeIlkS2s/tWri+UCR52U+9t3TjaBq3rJDrQ0FuNuod4jx2H6gtwxavhq3d6iC8Ay4TTvDP/fpjHa9TeIo5cG9OVTC96iz6xKXSJ7AFALpkVXeiLMdLsrj6IkePRoUDm85mHQO5W0PRgmoWgMjQa1OAjze55J+6jrj7MH3Mwfz7QYB3+XQ/y3Z8CF0b4JZ0CQi+Yzzm0UL9ELbekH2BpY0x+g6dNmj2sm+KWl7SRytqpCqEapsQcdPc8/xaz50/X7HDctjoznSrXzYWhKrU6E0oMnUbMG6ev/Qdo/NOxaOjJRHsujW0sbSxAZBPMemVfYAD4UVD9LK+wPGNC0V4q8S8NZY+6B5gSp56mffu3A5ziH/M4jmVPmOjU01oReil4H/DNkq1Yb2qTJqLrJggzrhtava1xTtEbcHQRWWxZc1LHD+WeLR5fc3ikGLRme9f8x4NEXRftpUOjF3Vh80J90qbau2Yp2caoOsGZCs45Lwg2tGgsL0XnMfxQ1kH0PuAYR4tvFOuWBSFi2TXvEAAIuCmmS/EyS7aSE7j5cxwe85YxWs95oJo76SLZ6hjTuhYrkZyd4D9cbCjqWLcLAZK7xHPSZJ+ZX88Ywj8shjb64AV9Xy9lCVbIgPzse9Z0XNMJNrmNXO9enmyWnd4JrWFuswNCwzmTtplW7B/PDSbQWcix5/4WjsesMyJNtYpBwuFdkTDwRkhyUQvDWrCg+Vk37mRfeFs9EYWBTd03p/GQunGtrLPGqLuZ7uvUI6z97iapHcoVcsLAwa1iiRnw67gFG9pw3MYi/DMRO6MOVjlTtcFmEH1Q129heB1/88DrEuzZPP4rVQ9ClpoPa90Ra7I0Ssh4ookPLkRT9wBopJaoRS78lAtOIy0IMg6ZhYELHyIK1jWRDUi+TggFK4VMzFN7z+xqAzphMwT4w60evIx2QFtYLIFd0b/KLwHTW07q6rtAnCbrmArM1cFiKfjWIaMvb0NQcm8tm8tOAfD7x+K5iuJsdZuWXcNGEsfA/suWa3OMy4PLQrqIkxbO4prhGXYaQa0jS55JhOWfzVjd5nK6JHaA5lPC4TA4NUUHCx3XR9HycZl9rnKLw+kwLjGVkgZetSYACSePTSg2isAkYZmxuOusvbn19anazTr354cM0VbrqOTYxkj4xOa2Btwu0y4iRR76b+fyt6V0IH73XDNxiIBaHYRX+6uP3jI4LRts6nbSmMGBuCnaaSts4eXXIQK80WgNIQrrH2hqf8YLtEjMe10PEgfoANqdhMwPLOuoPJn2lCstufvqR3X2RpGAEQgO0caUjJ9CmbWFVFoYglvw+R62s3JEJFOGr3vjdkTNOy7gJSMtxjjuKNJWxLOZStuRRToQD2DHbaDLCZ9oV0XUulZ84efmtK9wZ7LOMIo9T/ba64WfH86BfPd8oLyqmPQ2CvlJmnJLyAk3jV8evSau7x36YwX3TWPYYA4CHLW2v1//uRoqa1sF0xzykw02/ukcfFFLfbUMcVfVg6Db0mRhrYittFbaAFD3ZnfQZxKq+SuSwfSx7nHZkr1biJtB9/sRYgc1gEChiXmSEqrrytgiUD7fLUDhhN5bOvL0jlXBRoz+e2Tt/fI0LKllx43rrk0FeGTGi7rCNVy+nYn/qwPrapKD1z4ivlNbohF6AmP2IQFeZIlpgkLXf8zOjdiVr+0IqJruxhNUCnplyH3K41rouuAerIczl3pcouMhqdzYTIRlwT+bha/ZvRvGeV0aNkZ2PXtvMN+l0788GUd5dWCkwq9ZS09987fSP0UCFPIXo9j8epr7ZmWgp7/6ZzldvVs7SVC4WS176Mn1wkC85InrHY5vXzg78pUOrusIKsMR35GGKuQF3Q48Nfvpmi/eXK0IwPmA0I9RUhI2gMNwFz5rjdn/CgbUe8wm1tHIGE63lEtB9jCCsVtttQQ3JvravSrSOcfsFPXPs9lnzG5BMxFpj0PtZ7+RYkvr4/w1hlEregN1k0lQCImroFVtsEw5kBDB+eYnUG5lyM0uGBqzIzKlvJwPVtkL2xKInEOywINQwtNnUNKfeIUYv0NRdTcWUnoyEJN1kS9yxmbgc2o1n7K3CJpnqRqFpnQPpAdQP3+Ont36XFqJo2HiFgVatxk9HmRZ2Kt4CiLoPs5ZwJ/uNXRJq943rsZQyTqlb23aOHADpe7oqi+7D4q9Lik8r3cBatwIGSlNXMZx0XddkdrKd9GlzAXGmWl3F50j8jWKn/YIApRNJaLLZNEXkj1mN7FFJH/LU6X7Wi75XFsRzqGulxIhzSVY/EkkYBp3rtXe7aXXgNf/gCJ9aQNhp00bF/9edevhA5ALZ+BLBD0QC0j9a2VnKBizJPmWMttNeT72tPbuzM64dlGioaDPM6Xo5owPV87U5gNW7BRmPlCGO9XiLrNj+Stv+9ipX9FVCb5an3IIBw+K/FEGr6EpgXFjjWlzgQQTBUPSrs2XVtQVRc2wiVirtmjrqRfksZeTj3dCteAw3BMXhtEgc9Yo/N8KIWHNtuEiuwS+cBBYN1xbpUTmHCCpBMQ4X55neXIlLjADaoLZNVZWq0MArcj7TtKb+tZMINjY0aGAVEfcRdG9Tay/OPQabzX0uJ+gIo/cw4e/EbtOfZohQOirPT4lGfVwaQDqF11DcRq4ysjPHr2W+FnehP2Qa4sHh2pMKRixy7zIMOhF/7xU4J26/8SzDs0clvIsmWcNsNjZBU7ufak3epGTM45EsCx/Y/fqDICktysrz0XDAwf0aIsODq2jpvjCo0LuSWv0IJb/IvGJRy4NJ95JQ7EjfQXLMauroC/ONw0SOldpAsYVr2+zxxMZwax8ocDk34CZEcQymZaioCUSDDi1agmn4PPSv9G/PyQpWETlbBBrLqNjVQhUXIqzjdMZ04jKwhygXskiz3kAm7gInNdAuZCrlykFvJ0u7xOJ8KiFhZo3hUtF7htAeWP99SLWgeSKJYFtnFAjvVWhfdEpXpOG9nirUgLQKfpBQWpszyGKjFOPCnB7+V61/nNBNYU0ba7ESbA4JVe3SKJ8rPM8AObDwRsx3+jWv2+iyUEMTTTcOgiqANPmHQu5BCDBxltmYVa8b7uhZmNMLMuJsMMgeVm43x+ARbZuG6SimSuG6QG5XgXCHLl0E75cXk7o4=
`pragma protect end_data_block
`pragma protect digest_block
7790cf0c4692e08bc5c155c53407c4a37b2c0b8cd647d9412de2002917218892
`pragma protect end_digest_block
`pragma protect end_protected
