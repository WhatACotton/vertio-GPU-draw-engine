`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
Ig5CKps/HcNxhfb4URgpxHjrEO0UxMqA4tt7jPV2vEEVH75Mu1XCU5X4mBT8H5HCBdTT49eEjx1F90SIdJ6kKNBxco69PuTxGH42fXM+GOPpn2GVX0fGlUHPE30fh2nPPNRdKuxY9VIrvYAnRpSYwM+M1GwmA6HE/XFSuy2pDJyY8P6Td5xBwgd5dMVCUvF7dQqRuPqewT8VwrrLvHTdD67zJxv/oZ5cqy5is6hoRhj3PN6+r0AzC1djJMUPsz4J1rynTjDNqeScSiiLcJJOhaH8NrIP7wD4u/HBCXI/im2FVQTn73lNzEVtC7lTE1eJ/vKetdoiHGliG2dXEglb3RXWqvZ/jqECeDO/DitJZdWTKWGr+hVR/kyFJMR5JCe+0uaxVJSWXbKzCWnt8BNAwEYcUTbl39c+/8F4AZ3+0IxdwsIEuMPNHddoNNkTpDz03XkbYak3p/xlLsvBsHqZxsaDeVgDQ1vHPkhLGXCFMmSpyzZ+jdoy9RFbT+2B/cjPIVqnzjnVI77I+weFbm9uV7zCST/WhCYe1duc6oJ81M1MuNLVa06lMvo5kEQ4PXKp7zABIkPLZbvVJ7SN8aRIsKhtlEjPsUXilC9+s0K3IFEUXuHXyn7Oqsd1J2r4J8PL3FJyRXj6dVB7Y36Bk51ps91nuodynELJlpgTUZ86+p2XpXRIVKrhrDpr0L4F4+2zZtGD9c4ryKyks6T7ZZgBK91cZM+xn6g76tUCqJrTHX471oXxCTr6Wc5+T9Dil1M7XXnRaX7M3CTdC2XtAtdWEb4rfIL1vTV9Qmqk8ChArKLNoDM0m5wSKZv+ki1fL8dG8JkAGGdAXx2wtdOdeTeV0t3xWe6T6oAJtIMjYmBk/+O3xF2jHRxswaYmoczP/OIIUdvQAm6YkBqTOJkn+1iRXqxl6IwcZyPntzLLBSSlH+rJlaNtgPaKTtnyQMRLxtu4wNHI23Vs9wtW/QI6Q/QUL9YilLIJsMyZvFtlPwlBR7mxmj6Ub6Ob/Di9vNgcxz/wQHKMGzCgp88s9n/pO+YuP3xy/AKq9bqNHcqyMLtM59gEsaULkZLU9NA+EP7InAFCIAi1csDZWP4WsJZxxNol0fGRdwJBpmay1H3ZsCzo0gSh1Pn6z+glU5rzBSkt5jOAuABTL1PF9VrvEYvgG5IYoRxA6TuigL8oOHPalpWnOmKNu3BeWNRNbGkzK5IHI1B9MXh3RUP/TZRfa9USVsuVie9+526ksTufqAvzA1PRgiwXjgopYCz8S1PIKRHNg/9WhIuvYhM5NJUMo8UxUwxiwB8z6AzG/6+2ZrM3juwoD5zV+yFimnMNGb+JsswOZ5esFtnHfuNjPGrTd+x0VE8B6OQMui1TqlCky3CY+Hg9whNBcpzwTpv78P2V6pTTQ1h2DXOfJEGZ0paMiS4kACPfc/sBtNVZXdr8hqXIdnumGp3F5pJrQQGwdH/TD0wrENNgQ2S2yxtW99Uvc/rZ6l/XEIcgHNQzIinXi1UKZZLDIBfnnfOvTlKlY3YJH/CTVcWIiUIeAJ+MLRXRNzRo00+nMyYl/zy/FX3Wa4+2xKLrunsu9inDmZsNwPd8ME1pRmCMzLGRT2l10tP+caRvBVDAhMxWiGnn3GVZfwVgibdHOMfPuBROKcb1NWl3XRLwGuuv/dIC8XDvN6R1tD2GB6VaYk0PURm0Dg4PHD+VjBMjHwAy+QSGUZarLPyg6ShYJKhin+A6eT6zJcwFSjbgfBNMx9dJt83aB24YHVLJy4g3ZNZrdeDcTYpc7Cn5P7srhuUpnM9rIz6iPDKPMnsHGyErvUNGEX38W8j1eNe7fnptscNqdJueqLasF2XfPvZlJJ/+JYFHpgkaJHfO0N106EeWb0Ce6sXNIbYbZ3t/Y/u0f76Iw6j5U3e3j3rh5TdOqx2ukcBJydy8eZ/ImEK1+1WXWoZan5YSlNLSvD4MsnPT2ZI8s8P/HJbmkCgIvNAUQflmbvdoiy/NK7uhhp9FXRLwoYh5UqVZRX09GZxXrl3AzZ3MgNB8y4LYI522I9E3P3+xgHulFBWx2rnfjCfr94b3HI93EBOJ1uNonbWPl1hUUaszjQ5sjLJPX8LnkjmuszqBjdqBxOt6xwq2LM5qElbapapbZxnHySLIWhweeTkxmlUHvSHuqyJtizQlXwyzGsf3beJDioB2U1Vx9wk6txpS/EImNjfQYGalvAlqJGJReDqX4MR3uAy+zK+HwlGKuKyfaxRNMDxl4uG+i57YSL/sFsKwmEE2UqS2Gf5F1Qys1hu17ex7/bvijMhyGs4EB1PBcKSvaeEfUBSiOJHgcwltkcRESk42162XQYIQtI4/Py88vDh2zIdpEDlh3Ubsp6XMnl5Yzlio80yk2K9JlpTQ8pocH349UeHFfo6dufF4oz7deG1SjdrOEaP7gY0YARJrz0oKmFG012tPnKNi4DJSS3H2lEEWEw/ahEKfBlAe2AjnKZ8wM4KUyy5WYHqx3nfRd1jOlNpAqG6lNIojSzHFyRmTaj9Js4xdoVTH8gGMmdDO/U7i05aZuHyRDG/gi3O2NRHxts6BwNtC1XfgJJYx7nzhecGV1fzd6vDKvnRRShY1WenavhasTfoEwANBwgWq//RHjXqXT01Ajl669l3QgAB/hl14k4a8W+yZd99/d8W/rpu8gROUiLZyizPtkUZ9f2i8OsR+8TNMqgqcLCMtdiGucXnewvaFPaDMEOEBwAiTPLDi8IQp8IENPI3BQ3/7JqaR7VugLaCN7UoyJgyWavPLRwiQew2S/bSt4riM9E+MniOU4s52NNuPeKoJiJwfnCWOPC72mUIaJGbneH9A4leCP9cz0kTwW4Koca1WOnZ13Ti9hJwUoxfHLYnbeqtHdo6AgjVPxqeT2Qodbr8wh/1NDMIDAroJcjM0inO1S52ueYr8YrGNGjSMw4VIAK1eFNOz3PcTbkSabKRGukDVhvlRa9t3NfXam3thQnWib1NY4jMu/s9gG2ffjgA+y+7bpLolVTlxhlgh7aSBTUt6HplHn7jvtMJu+TtBtL3yb4+E7DvH2HoTQiM90Rs5sUvPxZfNrFei2z1QZn6+89W5ly1vbhag0y6HA3eY4GqzHlsjypdowuJCYcuhjByGmRj6X5F1yDXKzYAfkJYF4/hE60gfbjs530Sf4pEbJH+W6vKXNpb4wrXjRF4wON9aDdLM9FuX4ME9ycPRiNnUOo3M1askev8zIi5aL3VCkivQzmvSqzlUSrSA0iFnoPAoEM3kKiXkxdqQC/KUh4bszLK2aqXYROJYWAyvLpFjcvU8thA+yzkdTuxaH3z9Rzu2SMmMGtBPtSmWx2zJhxM6owLiPNUQR1mUqXU9Ujn+LXv94n+8AAZAlV17AFXqUX429e2infI1jvXdTShEPoqYVGDZ6hjdcqjBjAWV5sgH/xLSs8Ip8m/zTmysq8E75Rbd4jwN2QfkHY4FT/j6764fN6L4IR/hV4raWd+OTmTGzKB8YyTVI3TAhJKyE8gxWM3eL3AdJHXJ50tXT2Fxl6PNWuBo5yx7TRYZa9gjOHxMwUWSWT1M9MN/GIm0J9BiG0a3Dx8a7nnkBpBqGONY4XOo2NL36JMORMmT2r3HMRG1fM1wR52xcnXpiP6ZOvmEt+nBuIjcBuOvXFd+MGILmiydQiFTfZ/pYwYbayrOrQSDk3knD3OIl5b+fz6AfCPhIuViLWB8G99Y8+HBMqQ66cDxHOo/XeVKol91UW91Hk3yPdVroGytDzz6j0Vx24iwh5dFRE0jbYOm0iyIRveYrnBs0gj/p0TbFMe6/0QTDyUoTFeNodANtPdxVQiICVhp3Dy4NexxO3DrkxJLVKoxgqqGk2JV/ZMhJjDt/LbSRnuTFqEeyIpfWdzQ3Db05A6Yh3XNTIdFvUmEUXMM8Xoiwb11nuLeD+DFwljiWNXTF1n6ej9noVzIv4QOwhHPCULdyIKDwtesLpP18YgXrQ1U/El3JPqELSTNYLerAzrJ/J2nOYPL6f5Pe0TFgWvaQGiEOoDoCNci2Ntpx3mbbfwOe2Oyg7cE8TgbsWdbs5hEau6f16UQ/ABWufkAM7f1WgOjaD7dtjl+QO/+tavbwcwsvAHT4SgoHCw5W38sLnJfX9R0Pyk0BJhbpwhTg1TITwkcV1mvep+524UT4mazvj5ejvdXFHgSLagL8blI+a1bkwGvJKLaVwRKy72KkcngVaLh5oHUJsgskWxPUGGFPOchvCbfTwWPEpNjOygcJHp2O1wf4IU+x6UPIcJZEFyLcGhsi4uKOQAUHZemcvc+z9o5P5nQJ/mIs3JK06KD4/jzoIGiORRBlVCIiXrYnjnPFJtAPX8z/G+KPvO/53gSfzOthOY1s8rAqaZE5B3z0Gym/sC+EWqns/MFFrceYmBCnXG12HHvuBD3aQUg951bJw7xD9/GmG03+7hnDsSRuQtFt2y4axaaa4GlV26bhg5yJTGHbObIe0DVfkKStju0R4fZ84D4S1Rd9dy2dqUImzmoO1OwyNJnvaUfebW3hcPMHc3RQEXXR8O4P9iiK458K1T2GNpl5UoKUSczt7MMmKuEUh2iP20OwYJqTZxVuKDgGmFRwR2NBV+QijAzxCplrHk8N4ynneN90iC3+JXnoeN+5DrlTrfSO4FOVmDXI9sVuV0GqEKxsGxRMe5cJ2o6QYwc/L3iy8rmOJTXxqmIW+jmZVGQB4aaZdvUzMMTqz//JdnEMB/cGlJF6czzvtki5WNVIkJ5Cg+mGBOwZCGKlBCR0J7SJQVZPFuZQIhYH5jWzsydQZ1l8TmFNKag/ckcJ7FXIiTrMwyPIHtLz9xxBfB+2rfSpD7SXpnXCaLBa5EtCPZD6eOd3klKq+jSOlx9MvH45cM936Kt2/cpHdsQz9ZKt7v+447gHjvyPUKG+fMXNCAhV/ijehq4LA1rfMhhKd5gbdhbvsr+5YZ/S/qgh6AtNma9BK3FjFAIeq0lY6DvG2P6eOGyQ7bB5c6ELjcGFrbCY6F11It6nWJh1IvY/TN/rcCjIFsj63E4v5Y25fDZ4zs8TIqX9EWKf1aD14CWwoZK5NviQSw5lDMPcDyo3OyIaMCZZfI6yBtoEjxixwsv9N6Bv+KVUhb5MqZM/LumMm3b/AKwe5Q0IFdtD08TZ8cxnvZceznzKg4BQxGrE2zrS2JeQj2j2k9d2XzF89wYpOMsctifZiU0YhKBU9YVEMCbUiRaFGYhdoLk57xrF7NmbD/w2aCoLFtnlgiyGiGH4m5JNLClKgkvTVS/80x9SEVizYUOKJdoxAHO2+mdYYTgsvbGafZ2bne34DWwUCo/3u4ck0QS3Hw+hzit/axgwTIoy0N+kpzM4bF0GPMqQmALHDHCqkMpjQwMoSBZKMPWMI/uis6hkzs0htSEF72YCVl+5PZwbaCGjtpuaitJ0MgW07AJB+DhZmmf+iUM1Z9iKHPWrSNLTTeRf8MFLsP5ANZGMAgN+QnvOfuv8kxY8YYzUufEJ2zq9XI89zjfavr7INpvie6AWINp2hS/DsP9FCkJRCQ/6JI6aWlsvdxiWp9wsLjat1kanLQ8ZWc6GG93z8jQ3dnL/31ESQZ63VDiZvLuZZF9KCnf8EpnSP22shhK2J6r2fMPsQeqhegMfW7Vcx9kV9G80sSQLqU63v5cKFdVtwJfmZwiMCgok1tYhnzmYHDOif9b/Hqx34Qdi7H1VMDRcJqgX75+mvHJiLCxinTUV9MbMvH6hgdaxHW/rbR5Udq1AgUbvS3PvhEZVGmwjQcy5ddUa38QAcH3iqZWuWZnH+gMNOghJWhK5DKDYiBTmc2othBizPE59uM7JcORe4978+V0Ey24tWGBi0y1itOUZoe5BMNoMOh4Ow++l7qC4Jfar9JlKgpsts7RmEssMTlurrBuhcgWIjtilFqFmIJ6dta0xBsgC2T3+EaFgW9jadNfKQEs1d/8+2mIOclgJ1z8tCPDfdBWPUnSOLIXqU57Yx0+qQ25k1i44ibBerHJ/Ycez1ABFykCJP/56ltihSpgLo1MzD4IftkLHUfuEOijoy3I5l3E+C4fXVVAllt5hz8eEqMMYcpdKo3sLFPGShlFDgy2TTjlP55I74MCHuUKinux/f+hP9j6DIwU/1PdvYIq3io7KFr1Im79Qh+iLy/9M8CRHJzOQepudWYSWIO2pv+bHNGR5cFu6eApBcULrb9uu6cjZfghNj+B6BllI18Id63k/pxwYmKDGsyeYjd4ACXkt5O2A5aCjTRKXL9b7/3/Huw2/iH8I0y9PoutNKDm1CI/n2dJAkqsJU/0x6xiLIKIFSt6f/6lmVXQPC8EIWE1NN1CcilcFv/+h/CufMAAaILcAKsIBzigyS7hX67hq1C8Ueb6iNUs548QUiaQTCFDXyDWeCPw7UetRg8ebKtK6Wwo4995M9QyGpB7yKMFyGfGymHfCDsyBiON/1jv6p9MbPE9EZxxlSyhI2gyy9jF+ZaDoqkmL2NUQHmJIOxSbd37tBtDGgoq0Hb7aYLhZw3PDfuTv9HI+RvfxpMVbnmS/ZlFdCeMY7FMKSQh0Ja4O12xfsheEZluehqZDbGSXQ6DHWaP3JWUn++0DmGRjEr3WfjvhqdzpWncNdVNuqGtRsj2jgc8lJyaPuRUQiDv9czhhlCxBZwpiAzAKG6eNpesxmuzTRz/RAka9QII3GwY42K3PPES+eCsEEfTKwYhVIFi6ESUeOgsu2EXAYw71gSpfk6+Pqk0+Eq1luQfbTvjGYTKcg7R6a+2bggonb45jNYBw2At5dBoxorlqhq3k0T62zQ8aRgBhEI4A9IKldEI8XS1ob9nREEpwLVbgVoue+vW38EHdK2AcrJp5QMZ4gYyjlFYPE4lT8gx8pM4xD81zlPd+iq9dDHBqIs2KZ7U96IySzlQqVIFJdG7/x6k8dCwFTDlk97rKayp319dHY+R7bSWmBJ+KYC3v5dJ9tj3+0kTJhTnxk1R7gvVOq9iE7DNp3Pq4V1goBzB99wwqoenUvRwvqJjUEgBpVMGn7aoGdwQ3CIetJ3kQHoqlg1yQr3ngnuu8O2a3cot9WNmopNRKZZ6qPsrez2oRLWqIbJeJPoIO+WVOhgPfuM4EF1nb3NRSTfjp+4vkLDp76jGe6V6j2+PmLAgVDx3p0JMyeEtmfsaSTFyCfrkzpJoDpMHSJoYAgy+f9LuC8afE77zmIgY8uUh8k6AP31oszCp938fmxSO9y8THuBd0n9F4dGKR8BU9d8aUj50YlX5QuvLqbOV1JgUn5UajYcPE2ZUbMTw8B3QjEQWMnaeEThiHdzj4onZDaHvZn0yoS59bmMBhmM9gU6Z6i00TeOmOF3hLCQykW82zIX3KrGzGI73r0YMEC0I4Qqd1mD1RGN4y+ZtMF+np7nrjd88SlTNi38HKFRK9vFr3pLSrKBZJuwkZ9RGdzHtyBcpxiaKyg9cmqoWg1iZeH8DASjbWdT2hXCW3uSW/f5Yj8SOJiH+CAGUi96W2zG9BuNEVPpUe0owB8kzwXaYW/psVr/7LvM0L8HC7uBP+94grA8iwHxR+ieQM4VD/xPHnbewQeHZgo6woTV6OO60c5yQqpwvicdCdUwrXCFql2f9vKqwiuJZJ5WuM6nLhm/7150eN3O7uywy5edJTMhJmgmuU2lvsLNHkFdUEcZlaJSCccy6TztgqVNu+o0C7SdrkkRsDBQODXM4h8DJiVPQTPMBtnqTq4DR1GjovgS9KxKnd8GgzEo0Q4HbPuRpnwhVcU/EcFgqqGVGDp5lD5dXe0rdVyBEsoR/8vKrp608baSEjPrFKZohpZrA9J8aapgK0n3VQKoZhlw359tji7LnMFqK3y1L6ghR/sxk9dPJL5GrUJqA6qaAPyHYv19Jec1x7sVrZWZsKJpDC3CHX310jEDsjMIbu4kdh9ygFOuBQ+9YqywSmwHyovOBIjm3HrAWYNjDU+EF8VMGbnI9dnB8iQN/X353BEj5zQb96ydJFzPNk31ixRJQ+Yguy81+8DVMM6u3FlgY14vec4GUmCabIcauzZmLfNGrv66jyra3XluVJbnbuqmrZWfmnEDoi0rkKxyYUhl10/BI8FODaXu5EFJ4TCywHZXPxzIbexxF/AyJ5phdfTqeL89VIOIEpZPBAAdqcBindWmWYyGD89w2Kn8L8hIzyKIJ6aQ8f3i9x+Srx/RWx8YSkiwTw+EYbbF76rswkyvstgM0+IqJ2pxvBbAaT4SWHgX3ERolxtreV20s4/sc2SZrXe6VnbhG9nzHXxR+vcASYK3H9TfSa/c5g3fgk/WsdPnov5EknPAms8T65kRXcbKnKH3kI6OyhPFU8EW4cvPV6QoBnFkoJAF0XDEA7sKywGKCDGaqVYIHQe6buD+SQ1fXTsY4l1z588oykl3xtVNn9T7xw9fS9csaXqVqm1ID0s6RoZpFtb9lxTGgIUhPd0ZFeQ8L0LgWodDG/fsKwiKi0jOQJTbIGW4EVQiFSICBcBOUzL/UKlELbxaf4TbTuzyMm+ejZWyYUVV2WbmCZuHMeSpsOqOViY1kx4aFOUnE0ARP/G9aNt1rWIqc/8lxvks3K3YeTcNJc0xxmnCVN3rS1hRPTYtgqbGS+MoCGj7jie1L3nnQQBSmd47KX52kW91+rRy+lF8EcRUephOxaFVLE0y/0QtRfnNJCjwUH5ygvnAYqnshj8KOfS70VkHBzFvcmRThltijK/lPsWeu+nFxQB3PGvWUbSgxnDVfHcw27ndpEodYczeH1tLqD9tAuGguVpMTT/NV5cDl5PeItUCEcDLtLQk4ia99NESnfpVxkV6OCK++yrVlfVRWUww70GuHwGuJtqL9U7h38LHJ7CYnWyp/eXLCHcCjaCHdf+d4aAOOfNJPtFK9Oy4e9o932WnlTK1mTGg6nvZfwBisJRuGyzxIJwDYo3e9QCxCs3OEvd60DHnjBEXlOjxaFY3rmpwkPEGnILL3hckLcO7gAvTlkwJQtgxvbukYk+7PM6+pJQw6uxpxNiBvKf+KgnKjrQen4dJdaKxjLFervmnzeasqkCNdHDjU6J0qmIAGAoKvA/TZydZw4F+trplyksegmJI07UR/saZ+tvT1QGvqOttK/JlI1cv68niMpMJyC0jzlpHfhr+LxjM6f21KniiyUdicZg3v3yEyk2k0vxYAeZ6ql4zAtvdhxuFfpL3of8NbJFoaouLCE5eVMLm15k9g9plv7U4RTmRmAwMPlV3kvG9LNxn3UwqhjLrG51wtGIqIAStNe2cCh6XupVV6C/Eg7TAOc18mmqh2p0l65xLEFWsPStOJ3/Q8Z6ERg8pVvD5/Bb2j6FUX99zoffhXiwjz8b8GfWCZy4813S5PkZ257rG5QgbuGKPMN3hkpDsWl1J4TNAiSXEsdlGUZ/7ex94wLxBMzlH5QWWoRAt/V8pg+mnuRLYhuw6ZBof20eIQNRFWvQIMPL2hUYasvaP4Z/FSh1numcQ2aKx/uI/XWU74DMd30U62ztIBCTp1ekZSuGMr/1XGR0eHfRxiClcBcLZKVrMEk4Z603SVwAsKzM/prWha4KzDD1T8EEvqbkkDkjqdnEayqi+rjOtxZgbaG9ikdZCeiC4g0qRsooyyYRF7lOMRAOdLNY2eoqjllpiNGoqq39X821Lq6ka2XJFuATEstqCZ6Fswh3xqDv6YwTIs9t89UcfJHyB7Y8Pna7uCjuUomYZaNnfvNwn2vs9CABdoTrSK/mLoA3Q/4z4IdHWsbe22nn6AMjMX7gL1tdIqpq1/xTJIs3HSZ8BS8VzEsl+ajA7XpXsbaPZkb52K5w8Zb6Kz1XxNnwqNknv7Ota0nb/r1y3R7jD55GBfVPgQz5fK+bZzRA8aAHb/Ht1GXADGgM8U9a/NWXKZxryACMh14Zdq7+LpqJKYCM9a6uJ3JMBehQdZtS+c7+DtrTZBkntqAixgYvK3JRHRM54CZfbsgnAzx24mwRqo7FGEY9SesPsddD8RmPsjD2rTukO8AxqB+UKS8J3alBvW3Vu8ZT8gojlabnlAvzXmwb/Q/tbdGDn9cCusnN71vG83xZB6grYP9W37SFh2Yjp1R5ZEIq8Zi+TAHRlLqfRtBNLNxJOyW5WC2yf+akR3punfIXBkXOiugjyThpFNW4RDjWOlOWj3l5EIeXws1VIaW47u6+mvK4aS+qVME3BtRCFWPzaZBVbkYgcv2EH48M/7WoCb5PlebfXIynlY5/LQnVZIkuKqMdgOw9PlaecqgUyFTDGXBhC+dDby7e9yHQ/i/F3jdSyxdP/puZkN+D25Ll61ts19shUTNTKXvJuDAIiC1QVqC9915o6zOuUdm/1r1QH2XYJ4+YuaPofjFHrR03bju5Bf/eCsOvKg66pgXYsdH1r2NNoxDooPNQ2/o2yXqkA5/MVhvAb8NpgvyMgs50KuSFG3sgUjEd6V4pczjDYbWghm3jlXzeSo3M34DjtJT8C0WfCd7k/SoI58VRwPwGyQ4Zid1HnCTUuQ2MjROu49xH8EvRvmRaZlaeaD9dQ/XI1rcQX023lLvsWwpqlIUyZBabWUfkev47XJ54lGiOWMeAuepeRrzwc/7mRlbfHA3K0On5BeWo/vwYW+d4P2KNOJIONau5NYWJnR/xB7RUxiYLOoqmDIFR03lYtnJz5Zpp+epRJvUqSNdTbSSeORK+Hr/8QKJBKAp/RU6GEIh16zy4nhJ1t2DFDOfUuzqfijhtBoitGUIXb5igLHaIVZj3p2HxzLEAKR+DDqtrVVWUYez/gUj/Ff1jP8Xij/hEwL9X+L/i6ue62LsYTKLFWTmywI8x6l2QTSzwfPOpQW2F4RfYisdBTVbLw9OJiozGvNfF2ly37hcZIkiwW3n8HqBK5uC/5dFIJc5qRUWYYQsUc3lfaz00ppKswY30uYhYx+u4FT3yyuWSIm+JPm44nMAbb0oF0SNp1gj7TUZhPNY4Z+z8B8SIcBmnWQTT5RSnHFYiZ+9SCDFn4AWrDXLw5boYuZFgH2/w1wZSb9W0w3wEBCg5WiDKtFGJ+D9fYFpRSacz7j38+aGNZzQvy9lzyB/waLKYIXX5RYdlUmfrOUvafAulfCC9rW67Xinudbg7/zdtYmqHQlO0CWgrFw84pzFmLMGj+4B9RuowwUg1RZcKKyt+v4GPFfgvTivS8zy/Cc2Uv9lDixwwJQhnAsfy0jiuBKCJ1tnyiMqKED6t8MibNzQ+CNjW5+HwbxHmpfAW/q+7aJktm9JpHHomvBewU0PfYEncMPD4rU/3UZs34u3poKPN34NUNaWTaP/K3KUkGq8jsG5G9MfqVto0eQtm8C7zOJNQ8ZngGFwRFAYX1I3h3uGkWYqyPLE+jgbZkIGU5dKngg50CFpazPd1mCleJByn90dLUkE+CAw4OF+gVQKiqvzxNrgnLITSxACg5vKpz0x/3q/6alN82Xr/EIvJ7JFtEYf08RPJu9T3VbaEKjTj4SoFpR3lSxPSlCzfkTpOBD1Rg9PSjEHh7FyE/FY/ftPvygsCwouwfBrO9CV7zfrUMx5QsuZsS0xlOuDUkJffeSMw+0lS+cTkd8Yzwn9Oh/Fr7ptUSXOaO99Dq0vIQzaQ2s0oKSpwu6dS8915NyTlWqToPclqBxpELPX4qBo8qlF8BD7TYId/kqk7ZU4eB/xnr/bqVZNvqeAZc6nNp9l9LqUQrjbsTpPKqe1Ppw0rypbQlYOx2kqtZU9CjVtzALXXnehwZg5lbEM7XgCK14khBUDY7fghjr2OZnW6alhfz+Ge8V1YKcQ9nBKEXcUPUqJgOhmaF4FmKx8Ncu7WbFnAAqswGazTnELQhR6+/zoa10dQSYpVPH38sgL8HkZMhqvJn+PUDwSwiCLOldgx7Gpmf9F5iyvckIJU09IBPP4OlXa5jlzDM+CgZiv3Ow2mFMrUBTey3e9DHFBowGXfw4FMZ2VKESUwNHhYJYC2hmQZOq2sAFmkbA//pa8qQOfarMe3NOvENrSah39Tof9AKxheujwvgeNHBtFNbFXSKYGfYSw7dWawMd+tkXoS5TpQRBgdFF6R+ElomnMNcYRCgTHAYCqNmvdad5NS7wRC0HfubR8+L+cPHniSgI4TnZjEySh525JJCL9kc2a0xP+9CSlpSOrD1zU7D/rMKEsWm6rqUsluL+FWvxRbrcyp4kc9WIluDPwJS9gzphPbvLhyMed4CsAtsLMs9eXYDclzGQjfZks7d//wnO+uKL498W+PaP3LMGOXHji0M0z1dRadDaVQGPd5cLTmfDWOrfhInO26ycvIenUsgIV7vNb/StOKISnXIaulgWP78LWbdu2BWLVs5r/30UcLC+etgeZ/cbr3L7pxz+NROSLXM723IDWXRraaWOAo8nwOnV+gYxd5pNRmtrzXgnRQf/00p3I5L9MGmsXSSuLJtbrE7nVP9AEx1A3vhNvYMRsgJL4Iq9LFEWbTTVxVxmHHxbW9XxJVYK7Klrorw3+tqzqFO5+5MW2U7QNA33AYcoO0M6h13Do9VtD7YytMCxwpzncFQi8kR/rNVTuYr1P6boM4XjBCrM2+Gad3CIrIMgXwGEpxI8CkKhI/bRf4mzs9sd6YEABtkjDHH5umWhlI5riehRD+ngek+fLM+ScnT8tna0aB/6NEolw2+gb8Ragfb6I2RZxwFdQkfNW3sM2vsrmhnufyHg+lBuCPN2oEdmXzcyNSyQuNsI4XMN2CIf24FAtQudlE+1xeAV5gy3/RHr1ruZIXgk+NPcRPxxknLzofO2RxzGJ65ulCTp8RvYn7LtF8FiGajJY4diRk6SeCPgGTQfBcgtQpsXCwCB0mxY7ggosuqNOOV9erUzhcXrRDqNAJ6aYqhbR1QXnKm4iT7DDLZT6Y8gkeruWVGyBsPQNjzmC2TtHif7sJbsEzNFpo6CWeo9jwUIWpNOXW+NSdW20E7Bv7dIePggDoeMdeEbwZnOayr/1Vm7+NyHfwQ3GuZN8Vkyq9e3oo/1Ju3Qs+d4y5M7F8PShm64bC+kOyZFgMAMTrt3Zrwek8QYIOTLrI/vGoHRe6+UUOGKwm+abvbW3mc7Y48oSKBDI3Jly18lVE5CyWClR74650aP0NWiRxCHlzjEwvhciNVF8PzB99odnc56w51ue7IeQfZYgVNNqsLoJvqPPzcfsbgOf1cRME8yzr8X/u4XJmhjxvZdsgtLV5rijC2kgmEEbivpsB1R6ZDdSuQEgjbAKNSnlreEEMnSgRPFcZniosQT0qz3V+ShD5T689A/loKy9FdQ/MAz3gHG9wng16ffqDH7y7RWA2KhqPUkDZFJdLhjij7yumvC8O1OIWmO0/j5mBDg1q7SrIS3vMGstMhhbnLc6o/IpvVHhwvxGd2lLVbJf4ZITxf8QqxGRJ0Mhbt37nIDUF9evE7nXNyFkFSa+VoIeE9KNpl/zW2dpvwgpwPb264gPCDIVn3E2sjlUj2SKpMY3jGHMBulMAfuo04fVZ0ANiYRsFmunmNqivwUL5QpHvp2M1JD0k7J/r017kF6XGJTkHfFaQou1fhVkusrHZcJwti4pYhBUXtbXrNzhIXR66lRn2lNSzXJzo+vua3+ZEed1sNp/hL4ydZ13IQGYB13NzsFyapdCAkd42GvI8WtXTQNRvuO4btNl+7QqcOhaCGULKFA6eeRABWVFHLgIuh9l78rjINblfzQxyl+NLeVSmhhh3oRzG2IjDfXaImp7GOLq2mtQ6sjlM9SuQVJdwDyJY6uJVLuwLkLya+P4NZ8VZCjO/rg8juW6ZcDJv6xA0q3+zuwgv+CsuAP+kCYJxfzPApEJySknDnyl4p2LETO+4omcEeX3u1Ym3FwTDcUbUNMZaQPsQAxraMj6Tth6LIbZoEIxka9HfDZwZunTwmOvKvKiQ8yk2zx1RMJ18M10TA3q2QteX3bbhR0Mo3TTX0yoMBxlX5UCVgV4m0vKoNGp9RWXTc112REfNpIU4otH8fmos2EMa7bp1cde9lroGZWFNtnx9h+tiVrkc7IlK+T7ky1NiQfn2eR//zVxfXpVHpluiTQZgra6Ro+geb7ZOp2JIc0qVilGqWmH+K7wMHwUkIxThuhEzI0QSNxZPCTvT4ibjjU7cTlUEZ92hiaBXahVf42Z8RVGuIWf6qXoLhYTHO/Ijrj9eym17b1PGhuqBtL6v7+6qMjizvan1mvaNtTRq+QKxQW3zYfEwDCZ4Qtd1G9fiA+djeWX5IJRxYVJICHvz0fWZF3ZpXYNjYvQ9ynivjkwsfk0S44uTnkMqnzU9gqFqpSAJqZCgFvYQdyqDRYm77UQ3ra61kfLpja04iEmWpCToKBpHz1pFjLm4XGzt25V3eewtzH2S4FMEn/bcV2giPQOHpfAG8n0JkfDaFzSeA0sJKcDKtHkZ7Yj+pboL44TkfiCzCISCbY8nSfDNDHhB+o1xP9fqm6zUj9aHVp7D6pI/iZT9enwDfcGSPS+9UvBRMvGC3xTFi9vwga5EpDuHdL7vltelekQf9tPcEiBRF5WZftQ+b7e8y6LtqRDY6p8VPwB+XG66F8NANNNkxi4iRDOhvgGsrbm9Fui5eV+BuYW2BKpS8/434MVdL3Fqr62JscfFHjU1Xc70eJS6UQbEmrLPj0yhjGrQ1sLwxDuV3ScIhAyup7a8xuNBWg8H2Fy7v87XzFNdGqTTjMMWqzQg+exoJbUg07OQV2jrPyZeQdIs4XNEeDMvh93lALS8ZNCjLeZoTXg+oXjLHhl4rEciLDld1gcRIPaw1OUqPWLY657WqnWjkDf8prcSlRCOQ9mDt+LgQLuD19rC/uwv5ZgMiRxc59LawR2TnFww8ffjonI/d8Id2z8VCE6H9fyjFQgt73yoVeUwFyZ/8a6OeQ49t3uqM/e3MnCrxYfMZgQRYmGDzlOwh0CfEAp9Wfjz1znLrYz6pCHUR1l5XmcE9dY4k7Y9z+4zLB9UDu1bnLZ3zouyuq3eQ2NSPl0/BfoxKvur8CN/SoEKGRXS4uYdbWe1Z3QGWtOwKGzPITxzltWTbntzDGuIG28qVqoMSws7hOtCOJXE1b9wjB0XocDEzvD+jxsoTRJ3qYnxYtOfk1iVfisSLxQFQXIA+kN15f8vPywowJdeUorZQwtyNLzW2jQJLj2fUp5j7nlxKWqaL9e+M5nWAj2p6feLI+nXaOS7Jor0hwAgPJHo3If1plH8so5v83cSxbqOjWRrC+IGDixofBdXGBAMo8aJcwAqTOKnNwg/5yjfYgfpQPl1XrGot+lzMkN5PtjRS0q/AAHgET6gleF4dNSvd+zcHz+OK82tu2rvjbyTaiHcpYhwMykim4W4ypzr/g3yQxVlIqsIHLSnOwaLZcP3p+/Mr1s67luRy/EdkYyd7BKH/7QQdTnavmZzqR+z85DDa3EnKu8jDHXLMS/FUIG5X6M6OIuEYy2XbSK+meD94sqaXIKA2Tb9B63vqtFzDB7+OmmvP4P6xgQV0Kzhu0ONj9pGiNVzCo4VeKlvrlKqUoeYxnQ0u6SDgdkyFcvuFrhEZZrFPSRLWIUxdh5uVid4pw365orwYq7F1oW63aFHi8P6vP7nDK5Wz9Clw7j5WLlbw5T7Ujz53SwcXxAB6A6QpkzwL9xP2gZJT+bfrJKkqBsXF5m94QQm+nA4QK9HBX9p2lPsOi4unL4qvhI47e9JwC4GRXwmfDSsovqmI7nKddCpSwYl454l27+v9jOuDOSZwUawJi/vBuuGC0vKpXdv18PB+hohPRtYmuTM+mKOx9SBfahYdFDQeB8ERtDBCL+INIcetG6hkoPn73qTJjOYW3bXpHEhiSqdN5h+b+Bz0odYBNz33faByj9GIOxNDOipf+kDIxmlYWtIeDA1rWcr6NpmAoMfkvET7AsfvqcUTzeuhZntriS1HWpkFeZs/3yjN9gCAGaXl0EKtrVdtjKXZRARtSwPyOBC/8JOEK+aYRx2NTJmCO7w+81uhu54LPuZrAIQIw1s9kvlQ/CSO8H7ZvjDzRWvSxsjKPZyKRVHV+mPjmdbYeWIHjasHABnc07kMoXJoMIPrNBozRijJWvt6usgN8OQBBIB1TkYTsw4HTeP4MI3UG3/xpKmd5U0huzsOatd1n5NciwR5dTtof7cGmSW6jhXscW8GwFJe6KaP7wZBMQttlsf2Vu9W1ihnZjS5CB8yk2wqNtuoQj1qNnl0M3IkZ0J2I4OesJ+zOa6SyQz2CamSEDv+XgXphHL6bdoS53lEUEuJtqR08VVo7E71yAPAafe2UQYD94kMv3vi9eUcCGih+O9cV5OnPI0hCJygKTTFeJ2dseXSppvFYvpf2xJsnrwsVPPogUJD6Ysp/B9m0h04rGR0nD+IMKbk4lMHPZONTAHCZVUeyMIspRhzrhCMUeHlAm93N1zNOj7l+3BbxF1Th4Ww237OcQwmjH+7g7hKKf1YB6aFos+v0S849ION99jeReOgAYEsek2PIdXaPe8z1z7tPfBEcdXMvu/YgnJjk0Z6ohod0zJwHHPBebSV4VpOJEuvE778UH2iQkAFIXE1Gi3utzxI5v4K36OGtAWg6LoSy1meSS+B3TWr1aRWqSFqXg25991sxk7aafbglK/YUR5MxtkQePAnvuE7/aeTzqMtnOmL5H4pVjRBzD/x8VZ9eKHR5aLsoTOEotqdAD4aXHKeazEeW7bZ2nAkEFIL5ywp/GrusjlK30cmL5TwMgafKb//xTh1ES9S+LwQCfPReds1HNvGCmbZT8czTelzUXSuJZga6l7Gh0OAR5dT3TyIpBb+Z5jpP7CdbGx930O4klznkwD2vjOp/UgSlCO5043XT0477rmBqs75Cx13oeSYioTwYehiAJ6nK2cjPgRWJsCNcS+/ZNhNMZ5Sry+lR071kAZIC3HQYUgSfTf/zca0epdqgzHV79FNizmA1jwze/EKDNvDAHtkVwsb7gS2Xz8Rhdirqo1pzYNnAH/mDQqv2cdnd+6wz7a3wqq53OrgAhKw42AnU+STJglx5rr1I6Wq31JY2U/Ml1OcR8cAQzpr0Cvc5S0GqcCfnqznhJOuuVYNv8kAZx6++jKQe9QM29v2+LNIIxAfNCXfm1Vz+8J8QCKZuQfcrPbs6TEPh/iuPDwfXrcVy1/Y7HQ8xQHYOdXAuegT97+hGTY4GDgKmn49qI65HqwHvIykT1lzq9M9fM6En/3VkNMdScIB4bKr5aU5Td5f788O+Y4TaWE/1/UrqpzrKAgNNn6xlkcGRDDM1Ll7F5ryRPpH9KOXmzP75bIELF9hl+Kunbyr4vfBQfxsMGnqiU4zb95Wzwv6wemLxueh+sGYbFk83uEiHncq0mHK+oSG/xVA3CfOfnG9HNkzhOSrgjfbyDV6OexJFB04aKwQF6pKLZ2ONO5BgEknSUFZrdRksKPP6vFN0MdCAjwcT3HzShDKB5lFjociSPX/SxjsvfnoL4Tlh6dfdFtJwO06rXI8avXR7+uCLmMDeA29omBTGE6opkDK8lFm1RbMEz+xvxmr/FtJCC4E48qmefJEADxwsKviARM+LH/nOCOd7zJGiblansQHAd5UNZoYw1FBeBdfcyjG3Wy2FZqd+3yS/GSOwFOjjrjl7gZLph16cyFxvfBN0ofYgSsE9mPmuhSmAkVvRPpsn0ozEsaLVcpM31ET4D2n2jDXajGf6eygdVwoAIRVWpsUHOmwQpncMrQxPDyQp/CKI1y0PVASJYVnBk6uLRIFzXglfEOqDUIhY+mn9lTCaiblk8f8BfeB2TwHN/VATlOO9dk8FKynzEAcTK5AlLT/msclUkGEttBZg45Oz8cw2iUA83l0otcEZweGuF6njLpYeIBYdu2xkWoLI33IbdFVurQvjavxFCml6N5zm/3NzW/LFnb/js8wEr5/YkmbH6nSEpr7F3CL5C1dnPMAPa5GrYJLklpoNaRyzYsuc8meLG8wC2G4S56GTulve+NvdEjCWjLhZG0ihvyZctaQUbyax3z4h8q0T65RjD3Keaw7wq5Hpe7GWLwaPiyCc7BJItB7vCSi+B7QT8igY5WKMjx8XY/xyjI93yQoj9a51mgFBvlyT3Sqr2nV5+pM4bSNxIn/NMX6RC21JcVpP+SbH5u90QdYZ/Lq0VyD2VJ8FOR6NijY57rjlH0fvVgENMLZ1+zU1ki5gxKTPTLBqdOhcmTyO+5XGw/0znQYUYp+HKshDV1nSs9VB9m+2RIhAYT6hv25FGkSYMgszPqjK9TvlLroheQMeA/DH3GQ2Yir6ODp6mgo0LQHnodaxsRKobfinKafbyIY0N4PYmjgjgZ1mUAyiTvhS6nwjDfuOpd/SgxnS2vst847cH8x8rc7acEfth4+8/nFgxuPUebwSOuWnBAOICxjOZ85CkuXWoLiUtJLBxI5jJFnq84IXcOk/Nf8ugxj2/zW3SG8adOUcJC8vtA5+WiVQgQ2CXEh8aUTVESV7UCe1mxRk+D5PLOAqLs7tSoLlhUKxZvYj0aZYYigo4Eu1BDYuz5xhzmB3DIntzGOhz7a8Sh+eVRfiEK57E06BFClPEq9DhZp+ZoMwUOsgs1rGoQA4F/iP3ODM55M3PlUhxuWxc7EfSKD0zEr3Epmes1ZB2ST6pBsDxWeHCx35xwaElmCbRE6dkl0Q2fVIz3dJr5YrWKShKGDS90J47Y6+kM03C26W5RtTgYdoDHZSSCEvPFzeyS0gz7tsGInkQrF7pMx9Yv9plEP4FVMKziE3CagTKyMxAatbpakXNekH+ahIoAeeTJSYXYQYlcoVggitx42lBKLtjzmcgnnHyJRzSTilCzJ4h7+rRbleQgah9/0bp7KCH0N9YYZ2ZOqRFvPv3WbKlX7JqJ1fs+PdkrRSfQGcx/I9ryAZDUzHCbgfyBywUPkMpSc9FgW0yZKvJAIiojs41olTPJqsaMSUOKLt6fdsrBRsrBSZv0FhGE6fJfHrtaCSDyKBVdz5wm/iVwbZXWQIHLaT3q5NJbZ6HOBs1IK6RQbhXM6gMLCwfvlijptoY1K7yBXirlWswOtRz8uFEKWc4oNn00jGx3pE1RZnaN7RIvxMp54+LAP5YodGNHrHqjicZQ76QWNCerAor1trYjJCZCO/1yAsQsown61w7u/v6IRCzpNtsWgMLq+3vbIe2lJ28LN/PqAxqwBb6R4SpfjL+t9eOA59A5DzzwFJB/fau8ekw9QAG0zd3BLaIXZOApPk9sDvKgaj6NYBS11mIdKMimi7HliRNl3lMirasQtZ3ewgEMro6KFExlbbFW2iGPy36bzsBi16RrbbX7rDIm/HYI2LCU3GJuXV20oUsJjyJAW/txnksNXgPLdpe/4suDXdmdt8pibBX2MDxsWeDI06QjIBNdUSiv5pCO5FWwVQW+5YO8zWakKzVkYqZ6f4g3ahiN6Vxpm+59oL4M6GrcIG98maZ6NKrXlTj07dDlaZjtn5x5n0RTxguVBaJH1kKFiDu1Qlo7Q2tnvUSea8RbwzgbOUuBaO6o05T8lLnhRuY3kl68n9U+dqq5TeVPHwe56lQ2vY4/Wj8BExyywkIz4FA1UgjFFxAeW9iRdNzYfzn6UpnZuMkj4xpIZq3oPIRNgwu4un7vglo3t2G5J9OtTLr32y0y7ypVumTQB3/heCp7uUCyJDtU8XF3nUx4gX+6PEzFd3xpORxGyCow984hkwU8n1B96IHtTdf+JRK97qfj6yXABFTrErVHhb4kvKnpGzGKx8h7mfRIoGdKuRpbqJPr1ue2WiDvVpNkFldK6hW+Y0ZOa6NJsZcw1910mA1IAEEyBrTwCoxooMLyfJEP9xfJa1/m1bntk9Kvua1ojmaPjEEBIovEsUtqKn2dCaq3RieeXPw7pkfi5Psx5wTIPoERfPohqjXQ0xom0IBkbRbP0tjTWUTaWqkfHjCtdwM6JJfkosJELAK3oHVMjBwnWR9ISi43rULSCHMJ7w2hARzi0nvmxv2VOs0w+gSnQG8mLIeZLjoJ5TaFk23idiGTwrkSU8Z0uJ3/C38u5IaZyd581PbwfKGnFGoggJVqDn3cZ+CXw=
`pragma protect end_data_block
`pragma protect digest_block
bce73179d3112b72a3d1d3ff7c880649fcd1071ba3031574d1100bd354608db4
`pragma protect end_digest_block
`pragma protect end_protected
