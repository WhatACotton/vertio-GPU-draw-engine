`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
d3mThH1ApHQ20nvMI33hAC6ZdBADp9dykU++PGc+ZwwQEnHCCDAEohe2k6ZfNkNCgyvqn9XA4zQmQ9WQYeO6uyTggOXmwwJTgjukWAUm/313zolGrfGVznh8uYmu6ibD9dNCeX3M/sr1UyNqDnBvj6x5RCDfT2NJcLvmkUlYLX0OvoXW/TOXuSl8riUnTnuUysIaH3Tw7k8ZA1s+A96QChePMkrgT7oNYzCy3a38YmMl01rbcFuujNRrezSF2jnxNxBuJObf0YlR8GU4j/AShIkH28DZ8UVaqa2D/oNaPKr8FCJjFeu7nA0RWZpU1w5Wc01pdwFw1+R4mI/NvIVfCKT39iNj7LWW2pGlOunqBfS2iQ+VsVF3IhiT85siBoxc2tgX6WQSjF8QDLmVUKm0Ia69mE44ehKV2kmdFWbOUBj94apxPLjDSUEOiczMjdKsGP2HyceNw6RvUxSTJrn2xxkS4xgrR5E+nzhSmqrQmdwUElmUgqe/Ill7/567VJEMK55+4pKh57fAM3tvvAyhyrYeH/GlMFsUkpv4gTIlu7wSNrBwvsp4XfIIgo4Mwje8YPAu7/8G3ezW3/I5aIBoxihKB5IbwCAn63n1lqpnGCG2oTwYs/dUyLWSnD4Zx8zvN2HW6+Jjrb4tatDeGHsf8ZGKHJiyedDhPP3LyTXhT3gff+1qN4XHIs1It/VE7BiNcjBnYRHLDydW7wbdxMAK9ErasiaGsf8C1vPGzp+5+V2piAAGRWE/nbmQTb6VPbd1DpdBvxERfAfLERe38tiIfwnJ5ozfISKWYMJNpT7JuUCxKyQM3yJR7F1zOspbHxDNubCYTCsdnMaWIKEvPX6Vuheli1Q2l6qdEgX4eVyhavymEyrVj8HCwhAOeDYZt7/HIsD3vbaBDTR/bOxq1HHmJY8t8NqJPAvMd8cepXPysMgOMb1xoAfi53JTrdMZBCQ0g675xmdvcob6LNWkZoIKy+0syfEXldWgmmBz/lUOsvmsrJLY/dhRuzmW9w9NoPqzga6HWgc3hsMjknK1JzsYON4UuHXQ0OSS1T7q4sX+lRdMyN4y25Dgm5Jtv1wUdJHlfh7m4h23GcaC5FDV4pB+UgMtjt5tdgFfiikrUdRUvIXxxKmDvUhd2mpa/swx//WewHDnIKHkJC4tiRR3JkKRELg8CoURN5OdqUqadynA1lUYGXhlLfQUvztMF2OTIN2YYOIIiedGHPJi2NkCGc7meUTcX9dCyqY9nTpIBfco43n9v2S7T1BlpUQlK5nSRH5Gns6Cn7u6tDOnnDrHzDeSnrtmz5LUvbt+AR5v0HvI7RGwnjUIkF7c/LFneSuoFDPBEmSSTJf06IfGUcSqUv1/MZ7EmaN1oFtznhYZHYw1ERsTnw4rzr17woExf8OQzvU/zTWfbvmiepC9KiVsp33MdQmyGWtkTaeT3w+rFH25J+c=
`pragma protect end_data_block
`pragma protect digest_block
ab8f9c22960944862346481db0c6a8b83a94d436de09700223bfbd4736573d23
`pragma protect end_digest_block
`pragma protect end_protected
