`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
TvtN9DNxMGbmNlTEfbSma4JvBlSIGH+eBOz8h+jjiNmJSyWEAlW3yQTOgbDTUYv0GHOEZ8HK52musiCdJC74j48Ey9h2j2EXBkLwkJ3YBPsdQTsj59iFY4RwdXSLnikp8UH+ymfd1ywK6+Bn869FpzRbgNbSzewHaiELTCQiMod47XVzVpkqgNvxz7pQY9yS0prSsEMmtR6DtuRpBkOhVGCLqJFpbsUwT2i0H5Xm0Mh8xF2MSCC9TWdVfuqYNOcwaX+hzfGwNv7V7Z2CSIUkvhUDK1NObcWEZZsGU2y1ttYo5A4iPWXZJ7lrWmAS5nKi4rGT7iXIGAw/Y9h6nTlOe+ELteMs9lPfmSBV7iuMjHLPRy0BY+aPNNLYqATDtOrjeawgafUg86kUAz57faE5YaIda9k9Se80RBIkKg98dsyGb6wqxG9SuoEptnhrCY7MDxnbDci3eyo/5+RLedAGsGqh1vvXo0oZm28IYlTak7hTSUJkjvGkZN/XscnkeiWE/jgKhYqJH+3009KQ5yBKiL7l2/Rybs7MoWmfe5s6eazWYFSiyQ3nErTycdLIP+pivEpEgshf2jakx1IrBNfxXHzrIIh/ABkt76ttP5S3HFA7Bm4Ja8P4eVntEz5snPDus/kF2EzHH0JPn1wEQj3HKl1V0oLgbYIfsQ2SEqNmgqTvmbmcEJsQmzEWId8VmWdtsKG7inTNvr2zhVvp2TruWBXYopAMRunf8X/2wJiX9C4hs2HL6FDJaWWsq6G+vFbBIZmt0QNw//OBVBk+08nsCzhbcQ+lODgPoxFun4ZDmsJbcHnJPZlvL4I/m8/WehEpZM14WvaMTy1Rssi2j/iuu+zucaeAydtGF4B77xJka2Zo3ElPArNrYT0HgCj+WUiHiglpIG+4Wni6K34u+nQQGjTr/gxSCH75Qz4gt9QrXhmwkG6R8tej0h/HcUb/HiHVmkV//iGbyn4m64vGbkDaRY+KBiq0lkXNUbCRoglgHn8uAPwBoTENYHj3LDcycnGqX0JRMZZAO8Cuj9rDQkFtkF9PrpPlvUGhN5VF0a284MZGJFmp0xcZ+Ovwqi/47M5HtgJ0LiCzSsW1To/BvAw7H00kIhKYClWMCoDWo/Syl08n5qcy/a7MA5R+2oxdwN1VA8Hc1NDevJ8OLLIqFwRJt8m7+bKhumj+uvoWDjasU7c4E2YujvTZXkkOZf+SbH+yezp22Ihywsk7Zvqh2VqIx/ulFcd46O5tkCfmx85gUytJ/N5InGFwr5k0euw1Rv8q3trqNWY1SMjaoo5UHpDgp5KOj0o58sm/16B9nNBbAwbYsyxVM1xfvxs8feW55gF/X3e0OToEz9gD3lgVpSnHROcgJ84IeLJnzJowfLjV3hPUdIzOscc/J9fuQbDPaoOCo30XzzmzLVUb1vF2+EZH40U4OyvtJ8HElNpK3y39Hcz8pd6iqIn/EJLkoqPQ+5/XTSCSg95Gj2JW3oIxVYyFZnxUJpqI/VZDg186+lQiEwA09ZCZtl6k9cr0ARK5CqRUR3Za05u2yM2uwbygihowHnNhvNWp73tGd8m4Koo8srSJO4oT2xB+9N46aPOTh2VtmRG2kRq9i86y4IrN+KZ3cgoN67oc34Brm3nOSSrvs6LKfEygT5ijMfY9/3ZwXgN6dwKq1629aoNRUNBWWH80dvmxW0SSIo3bu+F2VTO+UG5YYMUpv3HVHUQ9zpO2B9bS8LfcP/NaxSNyPCz1Rg4FGxEwCWgoWfVUzXM6jY7G+oN8JmZQdRR8p4FIhw4+/Z3VAL3aLhjePGc4p2zpzPDfm5fCXEkbVba2ywk4o+MW9e7hW3DbA1P4auv6Hz4qGnU16U7eS7JG/P/7fYgaQItlvO6E7Rsq/LU7Op+87z1atgIWEDP4lXVgqBsLGag58FTcNwv1+j7qt8JOPXQ8mC+VBq/CmX8QGtfv4qadpYRN8zZtAcOjZhvN/pts6dv1XOniXirR9Z3LdBSVzprXF6ht7buohtjXC/2ac3bFt+rGayb41ZUzW/4k6tNIQgxQIN/E7z0eqHGZkY93QKdAJ+idyzwd77GxXnFSQcW+WtgOW8qre7c23CrqiLHvOCggFPVccZKKKfUeP9btJWsFpVzPZ+4YOtw3jPavTmQgKkvbabp/puMpFwPWGdjTWrp+wgK7GYOtl9tOjwo5bAAV/djQmA6LRRVWS/aawtUWeiV4QooUYLeyaMy9IayeHJHEzdTXVoLWq7aJuGMpR8Wvdraf7w/furjNpIk4e5uK6FND1zT8nXoNx3806jT3J0MenSeR+UA07ZdIxItA+pLvb5CFFvFP9Rg17K7u75YOZpX394f1uMs32wO1PG1XPh3iGpmGIwlc+umN1Fj+sjCS8K/A66c0xWByFwpmkfm/hqBX0WNkwPCkrbB+P5cE9A1c4yvtdAtweEpyK9DKC5IRZRaCIokESSQzfCl1gxgf2gkAAF+X9AXcdIuw5ZMNxVOWV7XQpL0Npr5XblI6UuzzFsM7dK+kfzy3ccdf4ErvCDyWaIRzSk8puC1L+EULtfmbT8PDf7oxgsxtMaN6zsf2DDbmPSTFQ6to2dPFit5Py+RI3MHkmevZm6HPgtbIFDcfiM5os+zw1NE0txOcT/Fvt9trLu3S2j7F45RjdPtuGQpW14e0mwpHmYT8t9jhFpr0cmpjHCKGyCOBoZlvnn6GUFCe9mPcmfdOWev/sKxntzfe71kU45SGG2uZ0EHI1kC764obIvnqAin3hqxg3b/fYfH9k+kWPsQivGBaELNTXHPoOfeLA6BFF84OJUvrG86369tkZiH6cAmJaO2PMgRBWqdKaWYvoJfdCIILzyjgMxFGiGFO4xpViIbe1BqTqlLriouZXZC9IGL/IOFdfM2B41ivHZ4wZREYWlQ+31WhCYXGhytDqhPEpfIQsdsGAYOxAL2NWxjnjmDmMiJeMjYaBmaLBt8RQ8vV7ppJ+v/+0PmOROZfwsx2nAeHjDTbYtpDNIx37Iz5Q+EvV67xIHFe8+tlyrm3E5RQdEbXrRBZCcr9B3oiO1icDi6YM6s/s6p95c90Sdp4I/9GXTkxbOF7Tkzk0+/4DFA4Yv2Y+jSg1IEeR4X93Je2Uk5SPBSddtyNzz+GqdYwUJ+8qNn3/1zCNXfw1VvTO19lF9P+E59X+mRPm/ou64McR/gZi0abkG5VXASJxZ+GgdebOGixU59SQ++KH+/H2homGB+Vo0mcoKiM7iOm+iOO+P6zy3MKBlCADYOVJSlcn8ppJJSHInswouS/hm9RMMmxPau+eqSGiG3sowPAiuNZbDWUnHPbyhDkSFNwVPW6ZKDOQnYsMCMThHXCaa66RRmgm7lsHM+yRbAp6JtMAUrKSwKhefOPQ9cZ3ouiTri3cN9lzHiA6sgaICHKbdlGYDT0qmoDzlASJ1VBXYoBka7uVljImdYbN8RbwMuB3R7wQo4/1foQm45aUzMEqOVTw3hRb2BSVu+ebr1O2pZqEgwrmqtfDpj/qf91X/s4MCFQWAyYyw49+8e1kV+cmnxEAP1dXOdfcHIzpH4af6CQ16fXexz2NlgUsdRhoHLWXo7X8OP8mbgiJ/uyGVir8YHwO4cTTcbpLMIqfV7kgExHE/3Nv5kMVPVftWcJekFySW7uE6tmhjRfQDeupzjgYcS5GnzOCyr37Vf02R4UjYCCQkLkbELCXiLnh+nBZ7K0RN9JJ2+EHAIu89A2ySQsczkkx/lS4e3ngGfCn3a5zqtLekQQ80iC47ENBcdxBVuJX+VhNEE9PBIrK1Nb9BjwBHDewcaXT19hhaz5pGYExH+L+XZTFHFmmHt+STWnL9jRZWTkLnaARP4WTSSGcv1vxPMvyf8hQ9PUczOYlxi1z3wjDMUn6TW6XRduA+gMAkltH32qKOjD2RrH1yUfqrUSJdwHxwsHLB5O44JM1qIp0pWSfru9LV85GfN9VujXHffX3mcFDu+db1tvId+gbK0QEbecwqQhOleLDJ8YvhyzmF2LBeu2A2RXf+2qfNVz9ny2WA9q52wCphkMdesamycXtxTqsoG0REjaE/ORYQSGTP0BT91wfWxWgHED6IBXWwTpZj97kvgDNrX04CtoCd8ZIkuMq3eXRh5qVO9d7IKHV0a1qftRXY/PWHol/QL3Vayb9qQqfxaHZtfGEjunHTchyeHS24iTVRw8eoDAd/npmU5djwCEDowU5Og2QckU7v6EtGAV4v8jrabGsQcBiOdZCZ4zLXa3z9OB9EqoXQ3olxRzXFoOb0uDPNYNsWqP28AKLgwAgWDIPrwd1rFemfTDfirEGLs7DcbGcRXJZpU877imqW62FCVN37HW7jKnzSBvyqTVDpK2w3xCKZgCHMPf4VOaJ1ZgAq9toeNIOCvXzBhmEz547sy/vEq8vxz7O/YJHbkuxO6RjQpHaSgZXmdHGSe5D0GjgHxGdgMK6jvgwXVjbJZavO4TiWayuObrMkeJLPgGgaPoigTUjrkzeol5jMfWZTMvzO0Q8ZyOB1+elCZ3eFYIBkAhZAVadO0tXoZST3ynj1AVp2K54JGAt2CrYWjGVcsmotjD4QgLDt/By/xRxWjzbbJWwILFcjacP1KWgePw55maqgzAcnT6eGroSrAvHYI126N2UVvzhbQT/zV6mVgyvzx7FTjertez8x/6CLT9rW3C0H6j0j5GwMZt9tEgO5eyie3x+HL2Voe9kMQeYKPhy1cVZdjcYwoQokb8eR8ClEzK0ildnlOlRfTpUhDc59Tnkn4HNwn3w7JJYFbaqcDXEU6vqGxSDEyCtnqct99YhXEyhZlFeH/gHYokcJVnWa11Oy6urP1+FnyLhoRnnRFr3blR01QrzcXoEgxuBGby9jMIQa+hL/9eNx4W9M2fpp5Zo3CGbA1Q7+GxJOooS398AqxbGLV6lGjPZEB41Mbe01jEILz5p57O56ASpAMe13l5l4rh3HPyaCRefTvWQhuvWp9ClnIBagtKnVXH55peaqXAfp4RADKg8uVAKU43OynZKvt3NhUL6LcZoHzY/5CCjKkClKAHmg0Ko7YIqmU4c0QkWUoVym9/8b4XlFW4bHemsYeHxPXWkOF+Mpl1zJ82Zfmehd0vDTK1WQRGo5ENaHWEU54a6lvaGX13Vas7RrhuWOrKDIPz0Q5W2ZES8/a22GnvPAgJGFHGAN6kOtKmoh1BRulZYHDpLhTwbrkxKC4Jit3R6gyZbD3fLuJnA7osI0hLLBgyfyPmEvURDni+NYW0cBUb3fVQWWhzjpn0bUudiefGo5d1HrCkl7XOxsxJiLQEM21x3amX534zzJpURlfJiRN2ejutqUh3KxbfOxV883TQTUGmesytAeE/623Ex8nJd0qovxumISnDObStjJev2I/2BBGFq+kCJC1NHVtTMdmS6yXqwQy3jP65kG3+F6idlTWJ8yb72Dom3GmsibZbaC5KUun9vtE7MGulEcGZwZFJhBwmeCdW6LWSDrj+qJW1O0yzCl1c9uabJ5aT0vqGNG2D224TCt0gH/GsJmzdKEo/rzIlgRL03YlvVs2sDp6s7nXxdMZfIeUj4ePMfJ5tVJUpbyzrOT2zq1zqhAYTkpUAr67lJBNoE9/K3xoj1Ae1e6ve0t0uFrwCWMG7DQe+lzcDIN4VhRKqn4DhR6hBlaWRtO9ZvdOvHkTTlx2iX9mXbwQfs5n1199Cdn194lPIXgOp4+JU0gBlxWcTLMdACMYk++pTw32pZTRd2BDaS4+H84Q9w3/0JxTMTHjmGVq6nmTK2nTrli62vB4KkB4ujNTtrPLjFyI/UsT2+YXdDpblB8pjQHKTcJBm2n6Y0XKUvXN96nr66Nz3m1HLPZ0sxaE2YZj9GaDOAPZgNOwTUsCTBOsjqLp3Kl46vv2maSy3rcSo7b3fnvF2EARKNbAtm1AouH4QkbI5JBsTQdflRmqXssYdkHHp1VJOi1idokLzPeCqPaTGFGZAaLsqGCp7veMMnt4z3Tu2UDzbsk2LCdjfp1OqDEah5p0N81ibSdU+XfJGBZCTqcBI6RmQ+3Mb+lKduy4TEdZ/ujmoV05uAULryYtHWqYazN5Q5QkYlp58IrQ9YxpmmzVXnRhkruSadz5D7Vo0uaq0yTqSbCiFThQ07yBiSOllXym57LKLbQKfuCQ/2f8i0CqL4rzgZ3oFYONZN1PEboG8Fns+UPdGD+ksqt9+qqQVV4Uw4EE3YwStQJFhtoLGCGlRiGLaYyTnafQpuC5zKFn4VH+N0x0tDqW24YkfT4bls15vg23/JXAywMCf3KPIjqEB5/IBqLGoYoManI1bcMl0W41tfs8gafXMBS9J8Zl84kuwSlvcNKvoryAGhmrO1CwBa6XiokXkDrfevXl4c4qmE0DMHuC1KyL/za7zWzJF2AOaCt/KRIbsqITWmN/INUpFq0VuZsN6zc5xvabhsOQekBrgAfbyq+5pbXuk2VZkuatkvkMnn8yrC7Ighm2wN2NH7DbYHCjiSB84a1F6dwpgNIQk6I3AmZ+GVSC4mxpa8NIafFwJu5mQhTiGpZKpKBcI6u3vJU0ASkAbHO+qE176g7deiwHUS5LOQY+F5/hgfyWEN8m+Ry2NWLE9jBMU5YI0XOh9vIgBf4uIaqNYGJ/laziDRroXiMXO77Hc0WNGT7Sd0WTVviMCwnnTp1hoK/M7+ltK4JPi0+1uG26fOYVAmswT4lIJbXhauHC9Ni3fd5SqnTNwAuQ/4wsn4Nfoi+K3W7q5/n9cRYKW/gc5+UlPjqGwx1+/b8Ct34fGxtxg6TBiMmxz4+D2Go27ZXeJvqZ1tHLgn6HeTNyvWB+1PM27/cRqAdnun4pzmwjg77pHBqZRgBv+SZYZI0rmCGeSLAvc4dvp+ETebGMJrJsoSDj67TpG4i9iR8syAcrXFotlZF32LlLBzbXLpJnR91fo0yHn9inZs8c49mEPAem6kIUcXExrQuStShnZAjGU95igQxvHMu0j+PEa3+Rm30/OYZko59ZKzSa8B/2u5rsQx8tER3SO3qYYaeBAUhvjikyMi11ntJaeJwttdP98Zn8zz5dr9WRBuYqFJdKkbA2LwRDskcCgYzm1P2ninax6dvORHqkUnJucd6D69eGHAnuO0+6zLsLaANDkbTGV0MSs3u6hbFEGhUANMZ4DxvCtnLYWVmGNDi/b1EskHFavSi+k4VF6lYgf3YNBxkkjyc/add4cri6owjYxjWekMO/j4A4dpyJ1PSl80KP9vtdEeUq9B9L+Umy/I17iY0AggP1c9aYb/OBdpUkJm7QnQuw1gfD9haFvb4huPf1kNUOYxqGsEvFbSjJcYuET7fXgZQDDFZGE3TpmZD2BuBRSl2/jMPJoQXHUbhzYhAqkmyIdlEu+S3vxJd14yfxqaOVXS1ZvkIe3ogD7GN6KjPN+I8XPsTppbgE7rbdkhrluM2NokO43yrLTa4yj5XtENCXEMcUM5QTreopOtLeWVoGm4KDIv3Y0m7oYShPZf1BdlEgf5NNjsOIBpXnshEaiHSrs2uEc664mV6dvKy0hCEr18jzYvYS4Ustq0Fv1/RtySBEjC8GYqiFAK0DlnbR52IHXSWo4l1NYVgOflrFiuFGe926zLxNBVlvej3Kv1+RnBFAUL3nmUAjm+rv/XURiecj0FFTvOnXL/FHDqClHCmHfGEeC7Wlrk2S+XNJVzjdrYhD3uHL4hSbj1pd6/w/tkvw+DNKt/XVqvDl6SqFHhdOYho8HuMxTyTPN+KqMNU2haTgoirl3tTf/3L8zmm85FikFKKcWhJVHpAj8R9I/6/yK1v+gklk0Fizl4b4z3CFLb50KicuR/q7R/MasQ4v/MIAD0flV5CTSYm/ZfH2BCEDEq/Vl7MyGFLgyV7e459rhSdcTeCE4oQO8a2J66Y9Cm2WJUhWF1UEpWhTY+cqWUAKfTNEDJ4qLa355hPG2PYreMAX0QDWHnj9iUTbTezsX+K8vpV2a5L+JUqlCgcbaAY23l3eZydRSbh8kUVgDAKHNqRyYMRcLlAJMexwrFPHa9fVkMfacGOEYq80ITngP3/4HNbrBgp56PRMcP5HOHyiC2jAM8J3QlWUuiWllbFIZytkYQr9aDUsnOG+duhrTVG2PTH6gnCX/G4GCC85RHEpi2Ct8UoDZ38LcitW98fqFn4AAsbheGoDPcUCBW943/nLHQnrZFqTUtH3jTXrJw2CDM8a0hZh7L3+68X2ZjlXTHOZPpMMMIkQObE4f/4FoQYWx16PdwivgWgafTlxao605x1DiAYycMNZah/PcRvJ0wxkxnHtfyNXYEDcb9E8E/G7Uar/GVL9UfwOoBfDoRbO1y9kJsh3VZmIkF0IhUBnrPJ8dOBZ2KVKu5jHrgK+scANIK8eG+8+ziGrHtsGtce+jSGyRmpa03rTrz5sW0bMgLn+Mhys/Mq1qSbSZoO8LAKIvtOvhpNIMUWay9RbcuE7H7ChjX2GRIT7AScv6m+uGzP3IJa2oBJY3NuSTd7ELwSw3hjW6K5c8Vm9IrbxOv1VN9ydFMIlBGdkzmrEtyHQYLc1dIPXXVQaTtFsYPruecnAg8JpFuffWAAN5wd8/98lQdtE0O88Asm8Tkl8JgCqjlG3azDtlZ3ucI3Fsy0Zl/AdirERJZ7z+PqFU/W91JpatwXoyTEv4VFfkP9MRjXKSapUHBB/3xSEc3P/G/294VIwVxgCYC/Beq1/Pf/Hb1Zyx+LS0v8OUWzZ7ATJ8V51f/3U452w4v/6Mau0a72yWY2GyeuVpwbtlrkMpS1fzOlnxS9acEj+x3dU0kppIEYX6KAfJzI+hMtYdj3hk9HpN7QS09CyRRPesRhzzi4LU8eIgVV9EUOTbCJcDd+IgGSAWXB7C4CL2jNNcSExAgm8xQHcgKvB9NlOAKeXALMkiuzV099s/3J/6BMRX+FLzEh/3TGru410oJL5vCrmUEKsa0Ozbi1uUPCF0ZpcAomBN/kxz6yFmPssNyxE5eSMp7uf852CFGzP1VPKbGRsM3t/Y1ysWngvB0Ro67cNhoSYOHzBn7XFhDvdeNPTFbd1eADuz4E98/0lbB9xivD3gdPCYizT/6BzcXMXXGJmduslhkDCrxPDstaWPzoNjFhiKRDbZvkZQ0izrp/MhwXQY4ZwthBn3F9mC/BijGNxR2fyUuJVlC008Te0UXJluDqV1ZnFOl+FTMLkB1t0uU29/QSGP3NAjiujKT/YOXzNJm7nFN6asc3CDeDFVqJXcOOI4YD9cAxelH75bDjnpk3Jaagn0CtpSEZGlwhVdKRu1Bh591qqTNRZOmqc9L3Z6EiUHWQEnZ5bCuY1fa3p1CLyF7XFgeEeWZEWtw0THCYGiwFb0DTYxW6eAUt3368dsmCbZj9KN44hxJlEIk6YlbqHTCJtERYkFEMq+yfXKP9SzJmSKxn3ysvUiZfS+0C2H1ZMj4vsNCOXW3oonfkMed15WaTaajI9fQenQ88jojW86V4AGAQ8yT3QM4lt4oWIKNGvGPVdpZkvBvS19RdLIXhfbR2MIFtEZ7AKycR4Hv8f4sya5vZVpjWa9KBN3btY04eombGtSst5hXOkQBlmc8RZwQM5xeffm7b5jCVLCGSlzbvRjqcgwfd8tAaF7YdjNl12hOMbol2o6mnon8I/0KPzaCobMAIjiwOC4sRgBWyQXqtoz1zSEo3tYaBjhkDMpr3ePjAha9LDfdFrhUiILcwwqNlRTvVEBTxCt+oS8pUDSKZ278WMn+KVxQsDL3mcKGc38fpP5Bpt7reLdZNMlPd/Ozo2BD0pHocd3/uVNU/WUnFKLTGg9eh/Mmq1btmIwKGEGqX2mpZOxi/ZA4dGJagAyQ4PvnO9jsuGN/5O1/2fG3AaIjuxVcocx5Hx6KsYdRRYFnofsgVsHdQOn69HBYHL1hx7V6JACETatuFXvKIcLXlCkHY7yRUYHUfFlUy8C4xDcz0Vu9VFVtzfrpoehkDZdbWnB+OzML1Bl1Wm3b/8p02fKY6JmqJ0YM40DopZFvQs3CPTVrGDFpGb3jRt8JrPTboBDQ7N/domnXNKF12cebuiNbPQfDeMrWMtOwEZ2BmIUOzfE0NqTzelVVwh1Z4uUOn5mBDw5vw0WTfURuukSkXslwycRYP3D3FuIw9oipq5DMEZDVYydhK/heooA6yebJtvQ0if0xRpZpwetGHc8uF46Law5x4ZARwLxrQKaMdi7fqHRh3aMUrQ7C8PkFRu2dvmZf11cuP2l5ECA5aZ9xFFlL1FTy5Ed1Sq9DSPf4bLo/tJqfkjW9pkAyJ6XQexEq1ZKbTiRVSIuaKEAXFt8b5y0ISXm1rOah08CVZvOxaMvC7ChsGZ0WAC6PpOH5KgJ12EqRQclupwwBwfRyx6F+XY+95m5DKw9H7me0EVmfjak9Ph8Uaz3d+YY1+eep8lQ4Ak84UqXsjRJ+f3E2p/iZV70WpCgkWxntdQQF/93PgekOZym9ZsSI9K1d5Cx/GE+bQJMFMiDFsCRq668mw3Z7lxQB7ilPSnLohqmUWnKhnAhLO7t0+FuwEnbk5i2G840CbdgpHmnWrBN/4t+lccTWQncdNTRuuZz3/9jvyGRr3rX3+690HvCYKT0ZKUswBDZNnept0S2g3/a8BMhIYjV0FNGu+B/PQD1t4QnYub37Melpfne7gA7b2kXPSySXVYzHPxSYA06rBwamG/hZllrQwNc6V61Sc1U9pI0GricCJtuX5Zbyy7ajuV7dW9nlavutYll5WFa/DXWF3tg8TPjMN3gi7DyrcRxEGmqsIe0KS/mCxizRyoHv/syOW4fQrL72ogysDc+ystFit+0g+C3ur35BMLqViRy7AWDhs/sZG5LK3QAl/zFGMhOJzoMXqnr9P6Q6syDDGLZLnVD6xQ1u4i1MJn74anA8wD8q18ukilQVkXsbsr4zGn3QffFf3pUK6deDfsfLfuCOth4PT3IWYTKOo4goPzJXWHK/QRLdzOk/MqbF1SgHzjnLzn6NOwLfxWI00Cx2zG93L4BG84LEWE6GkuSZqS+6FYqAZRJl4kQyIHWhL7wBJQr3ZkcmdqunpuO16So+2RC5r7ol3WEHml4itXNkpmsUn/AVlHblMOAOUEyyrt2EnAx92naFqqES5kzP3JNv6MpxfM8pb7ff2TdkVG0mfPqqKMU4/5yx8mQLodtdnMLwB/SO3BriOWWnSbspwvDkvXEA1w7YhyeDRMoN9n70H5CsnAoSFfg2Z/slE81/NGvuwr8kd/0/2V88rYpPlquaxSHMPDYlimwZHc1jRYeOc1Gw638sQqR/aI4xDmvHKCH93rM5vvdhp9D7lLhvRRGim7yHnvC+4o2WLnd46yJx4yeYbjAhgDQK3mnVVARxyP4Mvw/SzDqeFKNLeI9loQC/VYYRBwcsxar4fdBowH7OhvvFBt5mV1eQ6exKLuAVt+qgNhlspuOEL+hlMKtM4wIVm0zXGWMcosViv6pHxz4ONvLhvnqlFlLId4fLuaePWf4o7rhQaOVnMr8U3qK2SWgGhG9uQe2LjUvklDjr+gpWcozuE1om5Ec+s31y3AQuG1IAlwwjIbNLEgOZoISNVfJ9kGttWqKJPtckjkcbHqOe9bPyzwCYx33RcwrUF5r/UOcQ5Z+o7vCzn02VdEp2s2YeU2gy20Anim0yAp6Qsb6Rl31nc2/rMBqHu/qNWbcIc21/BrgbxV+5Qb/aI9k8Bz81+huxz3YIwSV2j+dQw1TyLK+Ua9pWGXWEPMcGQh1x7Py20oKgziNftXzUxEa7FFV9dOs/ClB7BSxJOTjoiU/uNBB4JcEH0msaj5gLseYLr29y55R0ore4tSGa6h6ty25gtlPaevGM8YYB22J3XToHyNPcsmXS5u9eJa61kEvVmSTayqMtBvut3/jAxo7HxlBBE6SKC09fIXuCf7jedpG15UpQLCKpM3L6asovGUG/SynlNESTh8wNtUWCJfQ8yoGwcL3j1cmhqx/PNX87ZXgO5PO5A66b/8hDD4bCC8whjXKbYTCCuPOSQxHyTrfc0REbJAkMydEruQA78wmarhaLUKjuJOWbuUN4ahyBgHBuSytr/Vtyo7BuKm04FuvDt3Ulcjqs8/1MzX86Z43hL40BY1EdgnTktutR80N++BHCog/NQqiB4kcI5s5w8VqVNqAMKDInYGjFjUtixYkv4YDtZcUlq+sARvpHfpI4nYs8whSwNP+/1BXXu8oZYev2Hba6ifhg7BInCOS3c0ZbNyK9yq+aYhjd4mXSRDxzRKN+TwdT8FJ8Qx2uYnyrycRw+0rT1Ln0ihOKYnHvvq0PxlYQ4EWzdr/qTdCeigD0HDM35b3s2MRRf8ZAuWln8mMjf1SW2y81PKgrbpiGcRv+ucum6ks3q7+eqf1JYlCV9NvlbL5YLi3O359bxBVfUjYowMToA5dusamFWX3zeZLqkrmjoY3Dgbla3U8uwPbf8DPhQ1gzJBdUN5OM5JPNYcHwQRDJrJLDMfc/62W4vn6WP62zBOTlOInxko3bRMpPZI8KLzTkO3jZnsCmseJTT9e18rWX4gwYjrTvE1nhp3zLwbNGNn0fTo0cG8Lx23eHpuwzvCA5VLyKUeMncP0y1auozwZXpKC5SkvftAyI92gi9V0LXSJVtRCS5y7sbnSbsu54ca1R3yQJy7J8lKyy9mFblwLTOY4dKGe26XNdRKiN9860quXxbwp+fD0fNMQ61c2GJ6lm7BdSE4oS1ukIFkftMA60I6hUGADb+YhAF42i379Vc7kYbj9PaBEQrXvTdAuLKWIRY8g97rzThnjZyc43rFalkrLbiRLI2ov0U/qf1OVHMp7I89Y4ygpafvSKRWouNPxMtmZulEkVz5TJKeoXT+6PHVrT7QakQ/02g1GBE55a84zNuMosrkIiK4d+lIJ+EnOdsuPVgCWxBD7j20Bf9RZqYhA44GVzBEbZL4H4rvV8oDIM7oe9pS7ij4MTN2ielq2fZLnQKj9/LQ+hpW/wGM2l/S5oNMhBQJw9d+y9YPWgTHOBQQ7oB2Kx4ShmqjHwJixA+RF0SePNB8Q9MsvGeA1byfxocqLrIE01vU5R27BCR6x86M5nL0zQl12WygthhGatusezs1zOmaDhMriCh8rz6i9gUQYaucVKlPc0GRod3TquNlOmOQbXj3BSwrMWMJTNjJ35gsNC3NvYlszK28S2BuWX2RUrHEUN8tMB3CHH8bfhGehH9hAGg5IS8xNoURYERLbHwXXSLWifIGb+GT4pukFVT0+9P+nh+xO01WtbEmP8Gdi7gdcASmqJN+bxR5NunxWFccX3DwlVOB/4bm7lt9v3QA1I6ndXMsXAz3s/PcOspHvWF1pcFM/Ht3k43cXESSFbKtOujtuBNitP6CDhxxQCM6kFVoQbZu6S1HzoKGk9tWgHYXuG8bD9LcFDQ/XtxTEwSYfOTsLZ1Ez910o5mV3azcLVMQe+lUPeQ0RXi1MOc1nqD1jeo2slBj0DPRB09xLfgTAxEcrcOx9NO6vBQ8U1n51HBL3j52G3+FM4m7Hh5DRDjgATub6aKVBlKVatZnsUSh5D4d9BzmPUQC2AlJF5SR1ht8u6iVp2m24ogoXYux68kFjYJnQPfoK+DXI1ho17GVzg8JjMiWQA+Dz4CTd2n8BPgmhT2dA9T8e8a99zgTAKyikk8ZCIXNUQH4v8p75/ba/UJLW29/VVpS6KTFYQRiUhVMpugpSyAmVWcbCdg2f4dESd/veSwNm03cLXqsrxyhBTHFPaYEduhUWcOY2AXemGDtiiLCR7dhfar/YfmXEWdpULLA8A6SxcsNQShGj37gixkQJD67axQylTb89Nrz89rupclA7/0ud2T+50VnXArqH/ABgcxIw10sFPK9yFPieSxuqOcfZdfa/aFiH29KJ/o+3wb1TPLQ+GpufSIcDs38NTLXmHHdiGyejOcTM0YaHbGlV4MsBUnxjaSG5TU3mLBfMtAm0fxWm+Lei6O0u8ZvRGIqa3CzEnhTjZvPZnWeR+oqAIIrGhJOdNxy+hFU1mz60uW2klIh83SBpD/FEG2jXhUmTC4IytflE2a4TtupLx2Wn7pj1AQgrJKxC15AGsaq7GKjF6fO8mJ94eYJOAFlITPLyb4sVmZaxL+jasOhU66lcMOAUvvwTQbEQEKe5QoJTBifwI0YaYV+CpVWbG59niSJO39Mo8cRMBUQYbQ2Wg+P7w07CwsmAhDz9TUfuP6yRzifziLzjxdMbmZT5iOxKY8m7KdGk4yfRE6SN7d5wlYccsPCp3QCKbQcibHfrqnDpa26qa6igTTd1FdxYkUSwhtcscOHJPlFBL+PlPlbAjiWdtsmeu+cDrKsbBuWUJYt+nLZuaX/WhOE9nLmflINThqul3ie4T4z8xr6uiY2zWZtju3lgRbIKQlOxCxcv4rSZPB1V2ZX0OBBr29yp5aylpJCRGuOkRmGIBTYzxXxF3ftVbDOks8qqKaHhreQRizJe9HTgM+Wk+4uBEIcSVvqOy0PbS3juxS2hNDor7WTyn1jLZUBdg4HxvF/VmkKZeAN6sxn5Ke+pABzIenS3oycybchhkVFF5yL6re5fK7YnNh+0JqOX1ho99ImYF9+AQCgr/iPVAthUt2l9ip2XBqGe5fqV6BV97OEt3iCud4p/w6XcsBNboA9Zv0PiUMcKfpOWlezeNYp3B6Sj+5bLwwJlQpcj6vxcs7EyZm6LBX/wB+F0bPTEXGbpVa4+CVajLH8oCgv68bNKvO5HiolWRxe7OX42yYEteJxOb993r2H6K8Y/gJELXKhyOLgendaM6nDPXHAjDnKz0W9VXwD/+Nefu/MQQtUu14jitnFMTxU00pstOc35EsQsrYVlL1b7hyfyF6Z3YZq1vbzpQrNZyJ0idsWCP7pYNRsa3qyg4c+v+LK+V+rXAlDwrTy1ptQlKelouVU2e0v9IDuFP+8Tf6HKpK4gCOmHst/jahd4+L6dKs0WpAOL33wgzUcU3Xf6dohmc9lObL1kA/7w8z0onUql+gK1wMtl35KmbP59Nd4yUKS2A4zYfxvvWC6B9I1r4jRT37Dh6lOqNz+zNd++5ZC5p/SDo7KheDn+x4fg3Wm1i7UDZ+OeehasWulu4vuFXt6SvCGBVtX+fjvyEAzxoExks3tU9RFODRze5d6X0Kmdk2k4k98pp+HYBhGuauTI9DHI2DrJmv+7D6Dojd/3J3KwwHzlyWSAObultwSFofpEBXRE+G3X0Zz8ADk7iQHNfDSRVQtOeONzuKvwGO/1gtVMfRzpBMsf6hgUHESBtTQUxUCWT3Xf6Hgx1ti95oIWwVJWIewNO//0U3nynaHF2K5eVA83UXshEX28AVzAbh7ZrM01XFucQdbSDFkq0UOCp7kSbJLo1o4HCy/EOaej0FsOdw8WVkahQqNS64iZbsY9uuGI8a5DgTpkSaKrZ0jzRb7Svq8mZxUNXuK6PJrCO0ijoBaW3aTjnQU2nKXS8W3UG+6ptBe10rO/iVjWDtNm1t6o9mIo4vS9JQiR9jbATrP8V2fn7W8+RbiCoJ6haO66gYUmjT/sMJbfZjwRlV830k7VHTX8D0zdQm9HDvWnUmQLbBv0BGm4k30iBlAqaezE3hiyKDpfq6ZxLIVdc3dQjFIwJjCDC8xHxDu3ERKdWKgfc5NBRro/0YDmLk3A26mVi+JlX4dLmMkyNQHQ0hTR1+eZSbApuigYoByZWbmt/JJ9TlAGUoIKzpL/TpM437DwwBqB+g7fpmkqVVCuFG5HZq/f6auE9SgwxJEl7YfmANfTo46+vgR6jPgj45W4d1Xr6tcu0eHbT8f/zn39e0bKnUuSGqDuLN3hj/c7ADp1nV7k9ceJgyDAA1O3/Q30xM28QQFLdaojj06bKvyHESuXGSnMtejhEA62vpFGtAYIm/aNmRCz26UK3tSFC3vOKfsflh+l0In7+JwXFThQyLR9bG0KLfmQjR8ame7CvZEJUodPx0/5GIE7h5guizJMpgpP5VHX0yfeBW5vYhrvdA6pbcDYq3Xnt/uVfjk+Phb0ASPkjAiQLLo4iHON3kz2tdQuwgoQhdYR6uzmTk/iQHOvKKR8Fms/LxEVoUq9DnpTwqgu5eHBwS58GaVauokxKjFfd7hc1HxrnNWX3iblbo4n4szNmuxQJlKuP80FX2rS2QabtRCWvOFrf137cj/DcfbVhn+4Ivn4LgRW5p0f/2WPcwhqqQy0jfW/txZuGajI/3MvkpTVsBun9UwjB2p3/5Ai8tcXumWyBVkyjFPVrgg8MSAfPhi8QND8s6QCau6lRJR6OgVkWosvqVTw5w/sqNPaLtIdB9oerKMW2Ozbt0PrsterHqDU8lTfuGApfOPUeZszdTOTlIIwJbWZh1tmdlya06+Xsam5dlokhv1f0YGZePaU+hrzJ3B1M7Xk8azOv/TJtTiuRCsoiaD9GlWabV1XbXE8t/6N9crtnalxFZtp/9JigQ9NYKanZ/hhmJLE7+MCnQlv26PgTilh+R30/TloGfxjhZOw4Qaf7e1Vc27IFqX2TqH1NWySqU56SQCXhaVvHoobf4xKsjWGFkljXFRaHu9QaHq/Z+w/PFeisfWXJrGHcvPmsgmxvj42cpRrE4cwQEYX8/7ALYJ1cHSMdUHwx7Ry68wtWmxwvOHLnv7K8ikDQOVNDmFwSSYWN/f0ehAOTP9d5S1BT1TBvRpc9XcuFM8/SLt575nr+2cklfXCJV15qDl6C7gaOCKvrH8AhH6bq7+oQKNJOKP/VJKzfqE7biw5+cVQx4oigY3vCuqc1lXn1apof18qBKKnjnwH+GTTNdGDMg1S9TWNlZl4U6Sr7OOXBlPY1X2my8okbDPtoxVtPkcoYDUX2NF6dgk/j8h96mLeo96y5qOOSX9Kz/82Nr6WRekdSjgr5LxY/GGzLvx6Nbt7Ogs8n+6nB+ZuGS8jtTlPpSNKOZ3UkykkzPoTK+uTmam8WrPdAlzMCxZD7ZMwsM0q2RtbKJ0Bgqj8/ZqPzcN9fSXVoovm3Gz7AgXlePuFgIru4IPcTCxvw1vP315YlkqM4gGg/VmhDEV5BK8hKCAWmHBm0aoj431U0Zd1O3L72kI9R4pRV+VMZpbQ8NHSBQmnt8jZlaUYn8xoVcWOrhqd7PYs6aiuqyCrciY3NODfrVrguEoHI+XV/hjeRlgku3TPrbPMgJTAzu3RJDA74KXSSuBsOuA5kOqSJC1J/uBgi7GsbxdCAM35kfI8siBXldLuVmTYZKz/ZqWZgcERVKhQboGI+FFj/RREqXYOsBglv5dP8DRgsJh0JhWeixcE8LR1vwHkgwY+xFn2RuFjhzgfbMYoe2ecXT2zSO1BRt1CbR30Qt7fUiidoBOj2mEHviuhHYwjtPt37yJxeCAbreO9IwrEhbe7d8Zbrt7f3Jv3pryxbrEei6frt+5iSCd17VES8wYgrIfj3ft5Poj6psYjcB+F8Jk0/GLencQa0LcCJezn4+poqGmqJPgJ3CM5bvGSmrTn2H7jBo8ev87pQIuOqoMKayY3GlLGOvAR4kqXIlzaKvt5Xew+HI3B1lSCvgBLj62geAkHnZD8lNZSleLFNjFR80t7KS6tj65nEfs1hVKgA0djii2uO8pSMJoueJejmhQhbPj6poQk6OiiorwjtJP/B076wlPOaJfrJC9GXpJPeaeNS+9uG2U0+BiBDv+rDRu7/1iHVpF3g40pfBNTuyG6ybIRxJ/pjfQLXOy5y7rnPeDFWkaYTinLgy8dbPaKZAqtntEVe5tZRU7STSmxzFP8TwRGxkwUawlxucSjdLGU3r/16jiaGbzpWE9IsPiPLoPGrwi47gmn4xgJ00SL11QXSLQxMCCyctfIM/8Ekp33H6K9PqCmyAQzhfOhu5qdqyR9smnM0x7bx7CFdDRImu+nPPUu32o87bpbRkX3b0vsJKtLYB0jwLliorSxGfUdcLQBSzauzfOm2hOEckQo/irPOUDPrf0Y/vDTxzqlLyMO02WwKXWJdkw+VDzVsp8ZHxDFtj2X5zpUnDSq77mhG9TsWzehYDv3IAXq0x/va2aGffJjQE0EZtecOjBg0QR7p8lKfK1giUQBIqVPvGGjmTR8K6MD7QYpPL7gP39BZ4p8vWj4Nre0or9YiQfJYWGoRSiGrnnuDwUXeg593Fov1O16H3fSFbyUFemiIZtnSyFWax5cpa2+xm0Dz6H6jJ6fggzM5EibUiCxSCs7TmV74+b5SZuQPs8MrNBkGvQqqjswtJGx7+W3xW+92/fmOrT4acVuH+MBffw49JghHyekefHI0oU7TVKz8HKBbLJRb0QWwj3z6JXrfgao8LyapF8P3FKMjd45WIqBsm21L2JHN74gjycOZROoVSDegzoMkpKGg5mnFASUdF0faEe7QOcTjPiOIsqZuitc1Je+RoEep22nW4lrlawKJuDpo4quxOQtngY5w0j5YyILOZBQjXmEubULbqofj83Ejhj3fNZ6QA/hchZTWBzulm3x2LzTdxIm77r+pGJ0mPi3hcf2A2Z4pbkLLZRKl/lDMjZrOshOL7itc19LZicj7EhKsHp3dR/mIg9EDkvKBZ17fHfLIt6Ey8P69AOVwe7q+e6KJtdOijUYcmv8eMyffS2hrEdQD0EmnMCu+5OHUTvVfyHM2l45sZ0cT2x8qFdKV8yiREhMc/b25/OroOiIlzHS/RbbUwXyB+aZvCtB0aHqQHMCTooovosD2bPJ49mRVHV7NYecBGkuGbuy4taBeObiXUDbMFIndePgPx3hYV8UBeXCnuU7YypnGL6j7HVJ0Bd784OxhBSmMp7cTwKvcMNxKlusVdnYQUj41ECDyVuhrShc3F3NySi25ahF8MsNcrbexk6NAMar0J+6Sl1fJA8yrOFBwtUOHCrm4baHdbK8+O97bu9CyKc4dYH82ny8OjqfkO1fUhAnX1qBod89GuBAP9UFvw9xyYuOe1g5881bmvxKq3XPIqjaa486g8AD08J7WBIMF4kT14fGBx6CJ2t0WHqw+7maYI7Gh1Hl+ObcYQiaYDc+mhm/QPagR22yA4hSN5PID+sYH+4Un0QLbOVopWyDDMxqEbCIVI21nJLsJzJYYIGioSOonceWSxnsBFcZYiVeBDZ+ArE+29/bYgdtkH+UdgUyR/PMPSaZfDSxVoFWohMzsBRQToEbcKewiuQpdWyviZyj6HQ29VBT3DUO3+nFceX2GNY7ENkGFp4N+fsFF8vRU5UmcD6HPeNlSpuB8Hzm/zQLKFbiY+cEacOXGlw0j0xkJ3WSXHHwQjXsMom9tXHk8OT9TqG/lgqH2rHd5NjT9eUT3XiI2M7wwGlgUqQFU8D3SPJjTi75X2WStH3G5KwwerTKkwc4pLMz8+VkdwbDiM+SLY5yDzJjU/11dBgUevam9g5GgXhmDgmBJ9qvxMP+KPMGtL0FAYrRGA80poenQJqLZY51JoE/LHNu3cS61KmVZ1ZJu7K9d0pM9zJSpl8uuesEMQWCxyNi7wRZWXZfVEp3tSQowxll9quD3PAxqohl9rJgt4cXcNrCC9EbeR3nN6eTWbIv2qmFk/NF5OQdAezl7Ti98ynjmQ8fG5KkSpxT8nrLzmXeLS+OzD0S1D+q18mcNHtMJ5rZaDc1wTgwa2j6rEtFqZokPuHMxDJc/TD/tRFfO8eA/sigfoCs6G/MhphvCWSyO1MJDoMuceLHMSpdQuhZc0uI3UnVZjIWTgy82rRI7LqjxoBzetrTt9FcpZTlwx5cuEgfvncsL9nAFtA0mMGIfEAec2+lYAPH87PndDcf2TRG5Kw98uKKNj/PtyeX+9zaYJmBnYla+a1tgvcBXs62LMCW0yS8+jV9eurv/g70zoH7hNQ65smSSjNHu1BqYSg+jIgUr0lyepzK7gTE/yubXGzCoDgPcpX0feZlLsjX19jPztvAKMRML7QMuos+QDKlmvQqVkZ6PMjPNNWFD8jO801MurryqcxY/LS4UevAQUDVxtfL/xCsabr5VS6yuNQJBKXzXu7eNlvGcTO9E9oDwJ27c7Lc98g=
`pragma protect end_data_block
`pragma protect digest_block
587c135c5600594a74777631c06cfaffe66b8cd4966e19918588fcb37aa51b36
`pragma protect end_digest_block
`pragma protect end_protected
