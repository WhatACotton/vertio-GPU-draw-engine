`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
nsyDgcYvEKmUVUSAqke9np3d+itWZwYBJAq9RiG/o+zBoBYCqx4ti9jP7xgOr0eEKfp4iZmPaAtKsvFFeyC9KIlqWTHVeMYthPRqqinXGoGN/0uF2kmgzwjV8IvieLRJ4H39o8jlhvyxwZAJzRzXej2f4qxoaKeru8QAU3ruA09zqrWGi49Jj9AMRFLFtmu8QV+03fwQtoAOCheAU8rVwAWS+TxxR70O0YygNQfuGu96fiJEAz3KsdkHtu9zCHAGVFJxDCLRLoRYEB9JzZMOIsUFosvZ+u9Xda/OpXLM/hl/f1d51b21pDS4A7lo1YU/4s/bxa3QYJSipUe44wQrntp/lewA/wq5ADEF8d8AN+yaLopNHk41UAr/sr08/uOnFE1W/FXylwImWB7ULpDie4GPmTVp5C6Z29rh8BlRykXAGb0iL47i0MQBqQsqlve2omKdaZQlXKOyDmjudyI7Jz1LHxsNommb9hzgJWVxFYZXNAZD5bojnhCyzuVzZGBR+o56lbywQHgEtPO05HMpvDboSSTuvHue3cxxIXRAaC2/OpwNNiaLpyxKX7qzrWE3FEopyqk6YL4z88INC7aQuzLbqybc3dZO5JTRbE258wbEkPkFensLsZbvWJWPOd6C+DuzNSLxBV9UU18mlyyiEc2CWQyQJvGyPM4/GDegDDvR+TYqfOvHMPS2KO9UY6yuVrpjqjsMEdP0HJfhqSI8v5GFxvKdLzWKmyHpRL7G+apisK6emjQ4oARTUhP0xeUGncGX9njMXMBKZT5soUOGDgyxg4IOCEgNml96KCN6KBf8ZAaqda0Eus4Lz/PawoYnDa1p+9hG3GN48EEJK47y8fcU2zx5zAyG4C647l0pxXB4UgFu1DT4WhSrFbCF7b9MmuNrHCV288XjVmoFmUdZRmTxbdQfaEXKZZpNgPWaT0jZwmJiOq9Bq/GHMC2Kt4ExtoT5nkqJoCU6ZDSJ6/jaIYvi04Vpow2ADbE1dRszEZ7L0talGfVrtdU3plzJKdEXyyztxd/RNblaE56uMNRVWQq+lm1CcLFuQyr3lJlv8FyVcRbbrywkg/dI4xWUU1bCxynsgtd6b6+5plOHpjtJETE2Z8bc6pIjLtY/lud6yvEgyyi6W87fkYNvInWlQ2hkIi/tBh8EIWHaIL0blyGamcN/Zolj8SmH+HxAG9U+zKAEcqwTaNV20WAXhw+U1ZH0ywI0bRTvXIdf6MCmI465rNxh06Y1+DelT9pHZNEwIgNOdsHX+YsQ1c2OJoeX2wIED4r+xxf/2EOlu/u3lD2XvENHXLqivNVgVhcFhdQz0rSbdR+qiw+1ayEIIC2GqUsnV6fUyWw8TAkNoFJmQt3LvHtG6ItKQWhUYC6EWNQu1Y4gKGKdiLi//SJQg5tKte2VBF26yti8XOQ3O3u5yWdVgAPM59FuaLLOsv2SLaxGhLbdsuYnUZyza1opjynVGH8PGhku50lXvczL21yFyNQLFMy1orW86inCIHBAo9qoeexIu/cwzTYYXPcJMgzzvIxTMokRMSMo9Xit1DBGj61MwnALssQ0xXATQgiFIiAgcZIYRS4JhSshxG39NhF0loN5bHhRODP9J/CbCrw/P7IPU6r6fEPvQl/PxmA06kW+qA2mXQ5+WUQ0qTZeQVBxiKI6InF4yqv4DtE7lYD9b12a/q9DudUZlLcH0gjie2NlSpxWjS0LEDonFMciS2j18J8QxelaHnvr8uPKAmXPDtKtJlNvjiH8WSis1MaNFkYfKR0zooStY0/YeXc085QSufsqAydD/hkZc+++0uznkucrMELIQudKXbDHTUEs9OtS2DKcgKef1zdhLNPB4Xup5kLpIq+GDUsCJ5h08fhjAuV7y5YOGg7VIlIGxlUjelcbvnnf4GiLt0od7yjFPwsF5UcRMqMrKj2syR1Ka4Zo5nBK6VNYiru2bYa6iWfVylbuyCRvOfg5R34E2YuYkKCxtAcT2KpBUgZm5m8KD6pSDXwWodpvx/I84Rs0tLRFbI6rdO3l5Bw07oB38g2fccoK6i4Ldq3UlNN7HZbCKmk5a5rfG9I//c9zWuM2PQA4uqMngPLdX84zb1eIycGWdgoelfVq1/qR3E43iPKUchidI2gJR1VRabO5aRJRJyE0Xfo40GmMX5gv2wzAOx4dTfOkf6BKB1DDlhxNdMwmnQ1wX/jc1mSdDdDQN0dn0C8yMeAIs1gtLMSC9vo8rG0uy+lpR1gJ00+PIfdR3Ll/+NhvbRKZOdeVFyfxMkZAMzNecmDh4D/3wcZA43rtz03wsdUo1bZ+XzJbbXF+Ow9no5goK806g18GXFbgDcHQDCYMCK0DGFQuNsarR3tmpzHZUXpgeVc9sN7EsEWMEFWZYhZs4LiTO7wNyggbZft+JyoBmikCyNT6GpleIsUH/trmp5LoedbYudaFCZSUo+1YVkfHXwu7bSU182FsdbEU5vzQh4OiiwAKRPO2BKlAcKtBJeHTLpAoEUkUC2V9AFkVNtiqQ9nsl+UG4EXbC5cCqbHTZJMx9uVmOVgOqohBwU7Gi6rlT/X9webZShUsqHb4IVn+GXM+ddmbeV3R+0LJagTdQh6+lZPHVZLpYvzvqFbH6PJdOse6EukgpiU78bqTL3cUgjE2fhQH8KphWbByV9duXgIF2laV/5YRDL/4CHkYCFZv1mWGiXfAauiJY6slwxI1x76ItsfUr+6YDVyyOopDiprYhEJo2Uh+Z9iRifaLgOpv2bi2PXzsuo6yPAiHfK/fOLwI+3aGKpiOC8xyltjsnmUDxkYIf6vyX7TTZnruzA9NUkxfwqZ/P49fQX07J/L3TuCyxF2byVlyaErOdPtaVcN51bSY7OBCs+RZRYQfgJZgquDVZ23nGsJmj/ioO09U/lg/gBA36FwTXAg6W3RilcbsJXzRftRCwR1b8xBwOC3EbESBfCSOm8ffP5kzLvO45MxOj7nkz6SHzZ+KghmVMSS3bu/A8GbwL5Kmwkr29vPuPbzo7QiiPuTADv4KmCecwgolAkbrOsAhsfixRN8CZUtR3qsW/WVqSRWzix61RRt+5B3Q2QhRYKwUv2vyTEHzsnkbykY7X1rYsXPvPZEQ3OteoTGFUBxo//wRrq5pOq9XtIxJVs7GHhUwF1HVBn/Hx8E/ljig7G5FjxOtL3UYmxtkYDfh0MfIEmCdw1FMycUJTnYG5xTE//+6hk0Gtp8aNVFusoYekRfvggtL7oimF9BMU+Nlhaq3zsoIr9psCzQPDO1HW2hqxf98j0q1PgGaJyVdu6KMZAybyeSki+D7VbWi5uvKLKy+T1AadhMKPnx+fQuBCMf3BN8ifFHgPxUlNlm5GBYE6AAYjlBRCYJ+/Wq6HungaUXgqBqr/mgjYJcxUJ0nwJhWoDZqYbu9qWia9t3LzWqyv52hjrM78q8IYnA8CZaL/2IZlB4yJSZiFs9Qu7AStoUWUwugcTQyqgsPQ1yZeceWfx8G8ShBx9Pr9N/AwZM=
`pragma protect end_data_block
`pragma protect digest_block
e1ca5f1d8327b298c4aadbbb45ca73920ae7ba3dc3ee40bbc3baf1eb1443397e
`pragma protect end_digest_block
`pragma protect end_protected
