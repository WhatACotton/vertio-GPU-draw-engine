`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
uI3JO4E6wY+TgWiCRvd+WgNyVKFR5VpbUERJeKirwaZ6C79jglBFnBpOQ4BPx1G3VXvYr0q6kSTTXkUAWL3adwPIyflpdQJgrRip9m89P3l86L7ZXBHzE71495qqCvoU7FNYatxKrnKh0OQue2O/rcdO+wJcOuVIb2VNjAeyQmud4dGfsYT8h8IHrZUVO9OWiZj3DDdY3wMrwUcSBXH9pZfxS8ihzZ75bAXn+SnKDt6OGTZNWuisGGXy29rcMZjjRVWdfBiCWkFQePxDHbniZrRnImvJz0YMipwHJbQTwJ8KSG4ngXd9EDaDXaVu6aRMvRyzeH5+OGN7AFxeQi7g/ESE3FoEWbA+zqWxsR6gm0faL2+V/hbea4+vT/WmUuXbGcZ/EnEWB1Cw8PYsqjMm7Wy4bfqKngVR3lup9Fu+vQH/go/cjZkZT5gHA6upA2oRkQ1EfuxvY3I6N1BVXSFQenp5Rrj6PP9AuK1oLOXXjevNNS45KvJVuIhoEpEMkdaoGWTmp7JH6/m80MUv4mwOkY81penK0otOintnf/CEHfmITUxXy9i/vjiKw5uuEbrlpk8tvaqd9l97W4yFl2IbXm0cE3zJni3i6wu+84yAH5/lQ3+dHYi7epn0taPc93gaBmh7F2my9SQwxMD6AIXS+dba2KQjwE1WEP71dYpyF9+VxvUcawHiBYM/Sl6e9CPsW0OwSOMJgKrkVwXiYq+yTljarGEufgaNmFXSoKDVxTItWYzSbRKIVmctkmpjkxXbd4v3MdEruVBx+xCrG9X35EXp2MTmeOIwBc/4iLaf8awnBohuZZUPb3bTztvm9jCPPIsQ7eEBZNwKP5yC8RR+4qq8d6OhTqgJd9YviMxzduFFO+5LsNfe4LncGZqgRAy54bQzbZ7JKVYjgI5cn3sXXx0rLYASPxYP/LknWgLk9mbvpYTe3KFC5HJBBbsL1PXwo+v65xTJfTHSuYabxkkqKOJP2+kkV1AaaGu86e7ASQeywzrdagh+wM4fBEqvEogcabdO16KLxJH4FvTBIDd0kCadxmQKjQQYT5/wV+CVfrkUdJ8TBUuHLGKbyNP9hvdVprQ+T6sDFZCL0t7/RfgLlG8k36/GUi32SacIagwtvpX0Kta6M59ba/2nZLbUuILa7Bg00F6DVxQfhoTtTXKPIUMoqRQu9LZzfdjBALEGoZ9nJDnTf6KxtjsJMQoeEaBdZhzslBIUtvKFO8fwqrdtM5kDFofjwJnr3UzqixNkUb3PdZAQIpzWLU0T9HuiKENKG7FtKw3bdwo6/j9zH6VO83p0QnGg4p06c3qUOGWtFT/HBuMCA/8y6QJLJeb9Jer0g5k3UPIzCLfUbHSiJej/92ox4pLnGrgOkq1c09Yo7YbMCdHpQQ86nNtT1yOvGu0EvJbbVTc0KwrJJB0rQmoxYMn56McgfD9uP+deJlgGNHthElL1EnFlPIV6S3pG2s7LSn1TwX1EHSUVL4coECoibRrhRM5Lorw/JKvLvPHswEb6peunN4tZkb+yRmE7xKIgl+rP1bCWl3a6mioLODecDB1dnrmX1OBjStkrerPv0nTXLjZhldkZsq+PGW8Vqfp2R3vS/nJRIfVsQ19Mb2xIYgzz77oAy+gzIqQ+IQRC80sD3T2lh/7lXaz1GnaiEcVSIlZQrgLluoDZSZaTZ+B/P8YUb93no1tM4TvpugvXNtbo+wTyTkjdgr8HJJ3UQYlhOFT5jcGgaKBWtVBsTv+pxQvIyBcluPPVp5y6ep2yv1somJVZ/U3I0f1rW0fNUeqhSxJ3Q3v6sHyi4mnG73AONRBqlKLbeX0wmf8Fgs+GsDWKQmXuDIFnERfnMWg9pBk+L5Z/QDRU0YAue6SeP3UDxjKVTQeSUvMzz8PxoBW1Q0Y3T/8v4FSwmibWw0T9qiwA30+eCJA/vBVguBJ/w4A5p2jU/B8QZQOBVWG75PPs6EBG1gCexHmQnD5tGQfq/PqDH9MkkFCOiqlFtM/C9AZe2FTqZdnzZXJt87dkwDgZj25j0VJx5VjcxhpFkTC6aq2fNwpvizWOAtN2z2IUvfnV123KBlMf15Zb1zUUks0+gn41jCwIGzVIqUrRrW39yoyMdkHYyxrX45rRenF0NZl5CTDTUfhtX5L/qNdx71v2T+E5u3DTMTl5peqTw//hmFidht6S82bh8pjD6JWzDa+4XtJ+rwqR9VvdoeYl441xqJhcZ262KiXjJ64J0EhqQDp0WBPLy1kep5K/Uv0xKMIDr+o9RY64O2Ybm0Dj2d4+rWVIXitLYYM4chwSwALBw88HYJcezckpieEzZzL3zOSnegC2brQ8zIdLcBBH06dZpJv99clcYCWnWZri4EBAS/j2XRg8PD6zMlLu1tyOWhrBhE981jzovv9B1F7+MTCF62BrlZ9S5W1PLMvQunisUmItQ/o7XSam7ImlbF6/j2oFNobs8w9tJhfsg1YgVHiYBq1eEDecGh2MYn6FHv6tsh3NS7blqMVBwkkf9m0bQFC6EmZ/muMEAn0GZ5GA98r18NNmae3feNyL0GMmIyzICjocgYxsswz04Z+XeAabzmr4cDKl/Xk7sfcVI1lNk9mv+dNxQrH6Ri4hJy2H1eBtxI7O7l5RMIF4ayZYoF7Dmz7e5ExvCcYj9jWvt4XNPON6Tc4T//U4h+ynx8GD2lMBrl4EOxe36DrsLvllmHw54S8KJZzFDxxyW9vVDQMNsN5lRhGqIEJAW3NbuN9jIGLS/wMNuIpwQH+5ai+2HNyMxCrr2lJ05xrGmFfr6bbvoCl3xYnIS5X4y3vXgHeYLJ+aWz2pszowBjXjUzdg2wPY8e0w++ljBbPFq7SDMfqAkDtD0i4CcxE9GzXlybECXV0Cwje0YJrwaeL2Sio9+mJeiloRJyqZ9t8gsywRq4W1SZIuxOf8pnf+GNXWHmrpEyr4HFvjAzk7xtFkZAiMZGFccQNWw5Tb5Gzr9hNerA7JbTorI7vrcg96e+isSZ4qiHQUbgQVAT/iYxmMIkcf7PNJTrkBIuA3ULDuW+XsmzjYe3eHZ8H2gbv/KINoiggXXwRg3Pxbhn4vMxcTnUltZaY6O7r3+Wwwrqz6uZizq4hdcAmswuu1d4lgX4tMiXVDjqpFmz3KDYcaoWvQZJs71sLoIzX6shH7gC9NIHdNcbjUl0lS96yZzq40ZrWOAGBbNRNUPZvsV2DeB+UNib7IfsS9maLVNbm3wDflN4q5+7PEhHbzhdLRjFQF4nXppyL/m9hhYcbhaK9255KG8gVCxt1fXBSlLEjmJnxZi5XXNopaSx0GPyOmM0MxempvMgi2HtMdIJgEtr9dQvhb5b+n9RugRRNuLMRnZ5SCnK+fmVTpOmagfIrJbfxP0PwH5VyeezcFYzgsBQfAi15XAW7lO5tT8/0p7j5e79rZ2ejh851JdR+TE3IDEFhLHBzbC6lMct300rBUa44QXjNkIxs0S2qh9WEUV0gi+ZwqmtTsN9FJo3F3LH/XaSMvlBkFRn920L/gI1u45ALLLnKZ1zhgeG7dLxXIxrCdyLRxiD5ddIkwedflU77nWLFMVsJG5E68v5KU5rTZJwl6LTyRSOKVgV9yCMQqm4v8+5zqN9k+vI6jhVtTBEuXyp9AhkAwZSnMeo1+f/NTl62tt/djpchKqeuuA30Q+LInxVb/8Yv8ecDjB5zC78Xpe/Mk4iZJL/oQXgW1zKgHbtuJ9AUbQo/XHnoesu7tylFNYAyDF+rCW+jWPlcNOwr8O65qatWiPalXGbArbUqnk7I0XIgNxTr/5+22mmpmYYYTcHi9JxTAGT3MHdry/yFrIJTw4T4pNAu1JQiBEKTGpdRj2iN4of2aOtPI3xmVW8DDqWyH8jJW81ryMUsMw9/c8l22YSzR+rkr8iUrUb/3l7jniD0+yy4oBBdJG0Y9NA72IFTeFAj+gcNIfruoZvzSHKojDrs5otOq8bi7maoinvbwFYlGKSeIPK6Lh25ZTQDWuhJAPbY96aPsXU/J78BYKZZTQCGBptdKS/6KORfQKk6FcjdmOL+9xj6i+KYHv8ECHkSIaQaZdf2L1Gh3GgPeEFQScySsd+nt9ChlraD2nU+5Zi+nOHCW8xQD5DtBvdWkDGnk87mFWxiTGEUG945n7Vufg4cGr5eAErQL2YGHmrut5tvlNjuzAo4d+QEU3PhewdXpJVZ1wAWiFpNiuWrwl65fS7KXsD2JRdiTdYDpKVirkgdPh2xIzUev1/g8tGUFaNMcLp6ivDCRkaow/a0yaSSFikCZO8V0ybSo84Zl3qiXr5H7ym1k9MQ1+2A2utkw6DgTPWHYxu5qkhuI4q6UVBepVpsV2GorKyTMDr7D5BJN0yKR/S5YNiFDa2lqSYFsu5+CcZZvvLa1UtP07LaRHGfZ1fmQNe2EKZCEiG2yK1PsHLc+8WEhXut2EIM5XXdXytdOXcNcMnlQRH6hzMj/BxeEB4n/GrHBMSvDV58cx6YqEVpmQf1cR6PKP9zu8YncStcDTIQqc2YE7Lde4ipNwJmEaIm7j+UGh1qp+tAE58eblT/7GoOJulGkZNBvLG4HRu/Om2wP9mIUf/SsCgLX7CY9tFT4msMkUPqzbCM+B/CeOF/o8Gr5nzAB4k4ffHhYZJzV63GFT9HZEzCJyRJhk40zeCw8WHjNYxqcmn2qgQyBVl0spbcvrFbsh7QRqByzA8IyJCEaI8qK5SpE29nT2ZZSKng+lc3d3P1fJZ62iUvw+QZ0UjjaDdLqzGoapVoGIrx9msfeZVeapn95m2GSn/1CoB1cO3Iks2vObACd7BivOGGfAUq8rB3KMa8GfJGJ2dfctp9VtPWKrrl+Pc4Iyfmqa6Pp+F5t2MfNYilEul3tu8X8XX65esKYUTOPMgyEWeKMfSsW6tNllTeLB7btPbEjspaBEBp1mnJqzg0TCaV1ili9W3XYBG/bxT8Q8/Lj1zkOHYoN2iUEvU7mjlXXFTAn4hecXk2/XDSrglau34CM081KhsGpbed70mgEtPskcPiozunLoNpaPZYWHmKTCPmGbDQCXUSY7kk3UbPdR/yjRCKVwGF/gr1QMXWwrOLlqUa4VxlEDO40gD/CKfcjjU2JK7PkjxkkZPfiim9m2KVSl8XxE95RvRPL8rDnfDXYwt1ai9EkiWpOSYLc5vhCTHUV2x+JxIlhXWq0CDLZkECatAgr9b+48pcQBTn6MSCIHFB1GJ7YvQAEhaxC6+M6vQDu1Q21xH7BRzzdW6kJxqyjoOGJS1YuLmH9nNyfADBjD91xerR/ETAR6d6BtbibKdEbNLY8Qwzc+eUm9RyL6AJ/rLRONmr+imi/ODtrqmtsT5h7kWKHnl2DWJhPt/Su/kvF0YHknhQJmYVtOySbQ78S6cGDhcU/W2AAbGR1TuiVNdYIsSmzdBqNP0wjARlunLuZ06sH3eHLE/f1drAfQtD3MqJVKIvarbE0j1211oem2rLoWF8cSiNMGi0d4gGoRp/SzSw55j/LM+smg3YTh4curzL67RgcM7nq+CAgpWBWGMD5ffDNhtElWZ/jSP7agskWBVlzT05H3Z+C2ku7yW+HZK946gYLAqTyqqFiFoGXexKgXnegjS1HH/tzG9xMz9m+xVeQZuchkeTvsvCVG8ex6hPPuaD8j7aFrI7VpC+6/SSEhqAs4xZpBZIWR8+p6FXLbOlK9Cv1XdS8VU0a8N/CPNIy7310KgGezQIvjdAxa589Qq4RuKkBh7vIvAdu3S91dqLrFnLJNiHE62qoo0P5gjqo49W1ZvhZ/JaS6ODyFPpvIfY6xi4owNdPFz59qLQnKeA5Q+rkP/7yKY38UIehfOalQ//csDQ0tjfvBzxc6qMj7En6t6PKZf3U1x43ZYrVhHBDZ6L3jKEIAOENERASSeRQn2j9kJBcFhqCG/hU5HDRTDB+IKYRYFix2QmPxGyy7kXlD/p+yKbUfnrTFNIBswXl83ilmVNI6mEflcqu30nkxsGKsaeehkgAlcXAzVjtTXAteqNaV8tYfq7fzHuo3lRi58lJjMt2Xm1O+ytJzhly2xNjkMTV/ErE8fCzloAYXj45rzn6Um3yZf3FgEOtX+uLrMk6ITwGpItzPF4wXslCFhK9Y4WxT2ZjI9EMqwCN7qFoOUB/GG97wtc/tlgsZNUXp+x1b6uTsRABdcaTVF6Ow2cy29FMN7+er66IjLW/6iIFKMqBndJPfrcovBFLZ6TRUSSFq+DkjNpTxpMAt4eayDmbc2XC41uRwCVNIVWPNfzav5M7Qz+xvK0QhKMvCJKG+WiE4D+c9St/0Se5JPQ0TL3HvXz3p/OwlFIEWS9raeSYuob/feyugYayYk2QC7GvXswVNVTrGER0fDchoy3yzPvAdNA4RTCFZ8w2cbBGhWGU7TVhgiRGH64Q1dWTFqNo4BVpMySXspFe6LvQ3HDgyBcySB18napB+B8K8zqNTW6bLDZjLexup7vDywJWuGJ52M1XXtuOtDWHHEsmkMeaoj+Tk5Wl/OCpME5rZGK78q1qcLLhRrrfIeOWym0jyJV+5xEvGb3KklfK6TWpbJJx5LAftSHgzG2mJT13Rvl0spY9gUXtiYSsDio3H7E5kOD+OJVRzenJtu+7kT65Gk06I90X724tbGaksl6jRdauvws6YS7Js/t1J5QBer8cKo6W69StSFI7dndr8jW+RjyS7QNNnhkzXIldUQBRbwfDDOWvB8Gggp7kJSUeIhgPqivTO3DbFk5sedQxh1IyLo3fYQxdArBVKR/DDNiaVhw38gwqkvywMrx1vD+ECuWYroSIkNmtgO7Qi5a5m0lQfshFn8vLJvwOiHKo5cBcwrdIPE39cyOBF4EVUjjNQ4uKPA/3FG436dPbxQ1vCFlhpkFR45olavzT90h6GVsIQsSeuyfV6MVXCZfDv3H2CHI2G0dxICyg7QUt267v8J31l0TcI5TFlXDJEwhPqF7WanDZuajBC6SfSnY7VPxvxayJnrMQIw/8A44CHOMldM3/FTANHx4UTus68xsVY61NGvKBwr+OgUxSwpZczCsGHW+K4pvBpyw2V4fmepWBIfjPw57Naf74jBXu03OgnNivnPUc3owurOBguzZzVLoKBcvQqC1d/JRyD/RqkNqQaUEZ4yg58KgT5rc5K9JkoL/ZWB51lIJIkjldvWqaAlral70MBNc8yXXleXu/rgqt/4ruWwUyY/tVSM5inhVNE3f339q0ZrJa+fcAEfC/HDEbQT/AaysyxeO0O67rLQYFI+BCTL2FY9A5wNSFImKWtoOUnseMUPnvHJATWq1WpP/ePtM9OUgYuoFn7X+cjvqjtnJ93ns420VQBtuwH4TDpZyHDEpv4Zk9IPVIzeyN4tSemB8Mk4oSECR95JrCKSpXNcCQ+F1Vl8bQDaSO/8PsjnDg2+D/V2464ojdkJ7/6I2IAbEOE5DZU/WVYjrj3JWREvEtDaa93jjiQPCwh23TU3RmhcG9zXxCfYw2Sh27sxSPbKg+pV88UmZHAqZZ0Q9T/U/zLYZQV1jmUC3UR2ZfWMmIStOkeJoZhbcrBZpUNGaZz78NubrrdbMwNzLIBCSt4nbWp2uOMC5rkEDjMreyEPTAGVC9iWrTpA2DWy06HAjrbk5uxNA/GSbaR88QTwf7SK0RBtF7WRYTPiyLX8v8GrAmS4vgq+Clxl9FGapa26z4GknGWOlMwjcVUY3b1z00Z36y+2hNeUNFei+SP2fr/RGhyQ508FewMkEBJ5VGGoPvmXB9VpofcB0vqf92fsiS658UKNZ78H3nXa8sH9ZAZegzM+XX+bODDZgouQoxVKUZ98llofDpj84HXPEWhFaIATWs11zAwueD791SGS12ahcwainCF0kuEbR0A5Mx8ZqsHpocdfJ44hEz6pealZyXS5SX2XE2iJHMpdVI3s8aRGrG3CzWXqs7IrDWf7WXwbnSTo1yCKeHEml9nPFxWjgow0ZB9W4bZezwcnwbk8FpBlVUOt1m50lYpGVDwARe/AL1qBa0hqRc0DptDNsgPTR5/wGdv4gDKr/lJYuAuONUndEgfDobrxFl7w4Tbkea5B9L3MxtAfvp1V+d5adp18q4o+uL64h0Xf5ANZ94JCcax2Mj5eegob5KTzhrjPZOZ5qL0L/75saxHvMcbRQ2R7cZBv23xoQjN1JPHdGtxr5dRZ7EJcVXKcnpZpkqMiDCbMwT4GbUrUdIVeAsVVnDi1U96fo/UweM9LkMn/KBUpZb1dMebIUdDpobBtuNFW7UZOO4rRR+GLNa513VSsY1j9bzWFaOCKRpwClf1c+mLj3BTjUOwx+RLW3GENAJfWUzTvasXUaKYVMJ3XoNGnUZD8PKSKbpBGEGciLlBbF/EjSkIRPiMPxgGrXtxkMQ9DXKptT0j3Htdgy6FIs9uhKjklbMSDcg6p5XLEEOd47iIywiGuaNcE385BUmWWAZq7rvIR5UwdqYXjDL++YKoNvvkYsqW+0TtYN8yYSQV9mIDbKyE1HiLZxtHOwnc9lgPA8AYeH7m6AUa2lgKb7nAWwhiaMj89sQO2rDPBDmqtMETvzNy2nSP+YIVIa3ZD18ZvhZsB23cN7/5RzKG/Q2Ul72wjzsHo06y8EVGRGzb3sGsFOCbX+fQ0VuUQvRx5CI21cKScgvHT7RdleV6WNMeU/iJz62dpQFHtpYMwyQyobS52CPHHjVx92iEQJGUtsBx1kv5egz10ttP4IUfufDgGuXDt7iwFaZBiIXQawFaWS885X4y+3Q4+YlPZ8m97ul5mo4QVX6O5oaydgqjX3uK3GFWdvDxaQMySpkhOsJe6P9TNnTGpVKznaKNBy5mcTesZ26QgK5eqR7ftgXw+vhJUUYDzG4T3KGGZkDz51wsjnJx8Oz5fW8wIQyNDBLptopdAc85e0FIDjvaj2Jg1jiMmveKAIy3wWaex3piwqYd7vzrcJiN0YhYFTDWiBn0aJBdktu/OuXDMhQ2sCx2WEhHpOR7S7oa3GilExDfUrZo4FBp/Mj3culgXFOIv2LJV8SM6pt+5gq17rqAAfkhydJg3Hy1+5tWjgeCGJeGGqpNN+02gWwWb2gWEFCUMDCPhFUqFt1wDInd45O3iVfGKxWVCqLsByU0S7VAmjuoXgZFH+fhGaG/sq3NdIBU5rq/l5+8anFNCLp8Oi7MwxcmiCCKQXv22iIVaeMBvNfKJDcbWgaO5yZ1sJQmhHaM7StYoPhDBl5zl6gaLx1VI+y5gHdyFih/JS6jqotDUAXKJpa/28UB+OSW/Zyr3mt538i/zqAt6YLGQKw5c7JbWw+CrRTDmXOymGvrEwOtnNhPslwv4Ae51yr8W3fJorkZeo/9HWAJHC/ffooc4RrDBfrm/Xq4EZ8ovDGbyncjC8FK/Q7fZUqtpv9vF+cVA3I2T2JRjQIZ7u0V7a8dtgi6G3q5FpuTjq6VBEn2N5nA6QrxGRgtQDMjjFEcZLQ9mP3YFA2pGF5jBVmysguZwURu2AX4ycu6TeTPpMe6HNferKhFJwe5/gx9mSUcnrOjzjHZQDbraHv8kpsaoVj3jijQ63sIGNiwrw5xJguSXX8XlTgUlUrbxohoXUSUCRWQ3Wj1Rp3o1yMe8jDXRHVTiY0P1FnrB/dqjZXkO5Hbi/uaqCG5LGSALt+M4Q9wACTIuqpKd2+PPaaNMRnnwJHawunLefJ+YEOpX00uKOdd2S/x9CHqnL7/BVBYsLyRdG/r+Gju/2N5U3835X/qBxnuWMJ9LI8jy4sN2V/GiRV16GkPiT0v93qRoXw0jQPQf4tHEXA/IatKusXGoM3Tpw6kzdmmfdkyG63oo9GUCQY5jD+VB1hfm5kJXXXZnd10cfiaByk5oAzD6XX7MNwz1TsOuaM92IiwwEgGhUD3iQMplhqWcakDyf/ujxQZVMjZfUPsnMCzgFv5IlLAe0Uw+ZEbI92xrz0KCaPn5t29xHXd1aFH5JL/Lwj1BUswm4NFR1y5iTveRmmIkhCBvr3sDIFpASlQSMwM2KuwNSNZzlZcJNsouVuJrAPcZfVOl2PFe4Bm6xWSEg9jGBuRo5AK6MfwmdYeHKwWrz7WR3FgWyB/y4XkO4SNdTTQG6wbvK55JdMLQSoyJBNja6tp+lA/LMPIwbBNixD7Z3jqkfUrQubqFkAbGSKDV71W7lezWk5A0wEKRZi+gYX6I/knGGzUHxVhbde44+bz/aTShY6NeONFGu4V/GoAiYOIunst+bInNnF3+QPeBeWrLE+wPGj7/SgEuQu7ighBUMvbaX4zQjrTv5dF5GouMW9uKlMlgr8sXsoxLAMn2DiMYS1h0qlvKeCp3EOx9ZB67SdMdLLsvaoC4I726mcB/4REa2t/RL+YwP8uJIZli2ncmbVBvzylyVeNUCg0UMNgWy6YLM12TWRTel1QiogeaLCphy5pVncApCYGC4QVSckHEZzHqN6IWcTPJyxJ0D9/DscORPxvgy7U9SpLBQVH4br9meLkJWCtt6gCX2X5hJoNut8RUc/WHMRUYClN8SU5YWTjJjIxa3Bdn4dZcqBP2zO9yrwxsb9SJSTIKpEjN2B3yB7ohayPzoe4KN+UdzqxTzpvQmPUAM2smMt19ckee2xGpq8xl9dSWnuXdpgGetlTdrm3vAd4EZHQH1Ajl1Re1JqZ0CfNzwSMFGLwah19FC+fQDKtxLrcdYclE52Z0DeTU6O0amr+xioerasENX8JyXIclcGBhcNzjkDeQxv/6nRq2KF6J3CKBwr/lXnE9Iw8eJr2nE3Nd+xYOock6R5vmqeGBcSFKiHhT9pFUuI3F4BKUtyKkVEiwewzbQnSTb/Elxred6PWGIccXZg7ImdH2swqhRYGouEiRf9E+Y+bIli8qydrq6uPQRAqTHl1Lc6QX5cBkp4XHrPZwCANnb5SpvVcSvDHnSTFuaEXWNoMXmWCsIoL93Cd4KIpk4FDFLxmt+v2IIIKDVpYKER0MNRhWSv3v/jcysvTVMSSv6x5L0qQB0JlRAAMboqk3vEg9ulsuLyGnTig6G2F8QpIizMg71aMAzfS2ZZW9tBIOOHsxxA1xHWdO2v4QajzDZLL5oToffKKOj0qqsj1gxE2jABBe0uftlf4/1TclD+Sah07J/X8AWZlcOwZLCg+OavYwvhrrn7OrrTTbb8X3d9M+A7rmZHe9nFdz0Z/JR+ZZMLKeFPWFC1dcyfxjXBNPRlW8fD7d2h+bPfp28noHwSK+8hb2O9X1O/5PsoZ1bih1R5Vp23zctMB0eTtz287GohcWErnrdsPOJA3oKMxlnKemgEDBl2FfG3QL97IynjTcNjBWFobCo7Ox6J8IFWuGDsag85x29T8zhvDag5CsZms/30dGo0VOoG4vek0tVewHV7NhtWBE5uhyu7SN4OhEfUS9Qlkw2YiJ1HZ+t0AUYfuqZEE/DWmpah0wzAgi3N7agpzcKBOWTKp4rzndJUMsW3ACPUFL6PshCR83QacrPslNVU81z/SYZUhouKrOwBtj+PQfJnc9RvHCZA1gpd++tsxk45CTP3SRQ0/T4PMvwb+Ip5GI6bCfb6YnAfD8uxC7pCRTj/S+14w4z0idG72TOcViVaKaCPHGmusoHKzqXWt9XCVuKElzBFF/3XZzSjC6a6OByFft+QMt4mT6N9LKPs23Vh82BbEy7r7bYBeHCM+RBeLtNjtbmFHxM7Zuqdtz436/Uz1a6UTf6Q0hzbRTsdWlLsdb6wXUJaBbp2pr+DkUJqOKOT8T4vj2RszMxQ6L4A5iDcctaeakpFqfzrOIUBd57DQT58VpbfUzv/DTzQIyJmUzZ+v66Nr3czXFtB4fEfGePGTmkVfOIVl0C4CFNwlBzLNcXcL7n7rX7327C/J8jDqIbeg2IcM3bjXiOrEn05oo9d7DNUI+E6/ndZfrAjNqFrdxYIAi7NxEfPH5QU5gpsGxe9YIkLImluFO395PggWRCGWGXmDk2y83oH5mClZOHo7KEgh4/lusxcC1TuA7ScJkG/xyumykrX6yZzKZnQOJyRd/ZVfqOE4n9cHoFLiEjULF6w6cEy5ppffvowu7qOUnB2fHqVeozpssxVF7Lj4+WjfpxwbffXmmsxblBd2cPUV89YE1dp0XuegP0sRp2SKnvzwS2rsC9YVlCeKqVOGG6k5jevQeGBBLiIgmVQjf0aCQXXN4PuWQfuFA/HILIz79r2RZf2aWlD4zYq4+uSUMhJ0KlTERICMeT2vPN4MmImPeZQvP2UvZ6h9bA80biUSDCFwJ+I7ICgwISgm1nmlM2MkctjgwUStCgpjyfpJ8Xs0bdL1k5qPNiuGCcddUNQkTC0Dl+AVVLFCs2yqY5ue7PRMtWktM4ANkt5ZFmF7VqVqh/cLju/XPSlRS7K++84hc4kF8VQFbPv2C1CdX9T2kpNz5vorL1uUSoP4s5PyvfJ+HDhm7yGHb54CM0TaMdRm3T174MhkGGZWR/7HklYd3bAleCgmiw7e24hUlT8NkwSaqQFWPTk6DNsdORKr6cMyFFouxex+4CLqwfU9Vse5OP65mp3U7LyUButq7k7Qdruw1wqESV16iEFZyTovzCbpCHnlYjXn1KbS14wxM3CccJIQJi/1FQsdVCy/4du0Xwhpx4R7paHIqhjnyvwta5Nz/GOiH+ZddNpS4xSvVwOAP0yJf+IRfXKxTwj/my2Pk5SstnAcPOLvYq9QlDlw0I7R7dsIQS6JYKS6yYh1k2cu1FgGdaRR5LFSWCgU6bwWduBMywfsw9sDRUz05sKjwUlPhLHRNSka2YUb3ELCn5yH9znyZTCccR8MExLfQQ8AXhsZoGiKKMMq3ho7yeBpi/XJFORqKPnC/KZp5qH8CYEdvy0WLjZOkGLOynjqXpwCBcv6wGMz4cqU/askEYcD1R7uXWwGW97/Z6w3UhFQOK8TXm0BaiwRFKgyI9G5NEYgJzYgO4rT80VluPc0Zlmt8UFxp/j+w0RFYvzLsXXcddgIGB//vX+y90QUzkAczE3sad29CPMah5R7KM+Gb3yQunsgu4z3ZUYo2JkCvMtM4AsOn3HLdU6pOBjdSe/2cPvi7AIDHm2/mkPvEecjFIALpj/yi79dkodzHrNcXONUrhRynxFYqus3dPK//0UHPFMHnuW46Fk5MPymJoPlPhlrr6IweLqLYRRuVQq7IG1aOBU60L3v6owZOfbHNxtMjZ1s8YGfSVHFremlAknD82m+oqNgevEfYod7eeoivkSV7odnw8JJudKrS+J0mNZb6ox8+AOiaAgxvkFAMnchfGsPCDr4MhMEZ7XHv3SBQnb7+QemdKW6bHIvN0m9TI7v6n1wMKQ3IsKzBR7RVu6Gu3vIFnNDsXlaJ+AaLPqkBlt52B9FOVwN07TUXZxBmnBwncDxV9JfyxfHVgAh8A0vZwedKpbMLW27P6LQWWIzuRsTgSH05WiyGl3wUOcCX7T/UOiu7ucC7ZRCyGOUETjzKmGnVVPAyBnuAxQKXBztDX/77+fA9aMZYsAY/pK9zAw+q8YW8xbR1iVe87huYl9pJf/JDjn3zFCkmsqlS1DxE/bWCPfF3cLaRCu/lsCwY5ZGHgdNIW2tFZ72sxIdYHVVpWqVqwNz8nLJ31suZuD7yFMtp8FHkvWyyxeIliTVLhFyD2tWTk2jT/pq+CkM6Mdd8kfzbiGcREiqajtfZRA/fBe3DA5hung4BReIgZaDTXhaTgLBRO//jAXdhi450yni8NTkyTyWhVMg+rGuwD5ORNs7eOZ9wBzQPIshoMCuK/Dm9JJusL5IfkThYc/AMvYsIlqUBsgvzwiy8V2335Vj1wB5T8gRl4T/C2gHBznCrfXIrsCFi+NCMUFc3XSLFLKtQudcqI0QH5z+4EAntyDu9mPWGv1dav/5HM7jY9sGk993WyCYeS5xA7ftI6eKuuO4qcBSnyVYDW+s7ayb9bNVlbocSKQl0JleQD0oAZBBq6cq2HmCnk+rDnINvgcurEUPBDog5CmzR7kZKqHkgn5WjNDk1p8cN+SUjExNTiADHKmTqHHPd8B7J0noLPJfFQlXz+A0AB4xSGdh/01EjuBA7kLs2vsH5d+EKJQg90Wc8yM54sgrHwtM3l19cSlgjrkJ0614HVNKG0h/a3Lw3rNBf5CjSUJ5qwwWoJYuvVFSDQDNke7jlDBb3IOVybwW/2PeCBSt5e0Rrd2SXao4L3ZmmTxgaCnOL/gsXoJm/CPqr9UwDM+xHU9wZW34dlKJ2oXgHQr+9B588bWba7MMkIS3SUJcvXzo1MNtqfcUY0/l30YS+qFcYg1Y88keFM65UrXANIWFcq7v/wrzZ6F6B6o+5U2Eukrr+NHxSV2k+DOqBPYClS1OXdWlXHCpdTfS0UioSRGvZLnM9Nb6PVqYhDHJVYBWiU03SELK4CZIkSJuLsX/kqBywRo3MnS2mdekPoE0i7mB0/M6u8NXIiaetUSezy/Rsr0SiLy3jrZ9Fu6qgfmyNi1evL2j2c3ICh6pwHZeoGr8vFEhNXSDzFRNVCk/YULd0PBfNnxOZgvIJansVzIYk8u0llon/PPNkeekR0kZWqAiGDCs5fBsMf/omVCGwoSGI7zwakIFbEBQaiKYLJlMA7qGY3kLaKIK14nVujJecM6uWjGOGFYMRlg3smM8L3zlL0DVB7lRHFHKGs7KaDjxQ0VVIWYSUokbxo38OqE7lfTi1kJYWVPi7uC/wSFQRSDDJyC6ut5bpISwAg1CwQtHJ3URqkipvbFBGyOq6uZSSO0oKEQgqowQy0OfUVOdmyD0Rc4OyRej6vzlPGYL4SniW9FDgPzJw8GbUfzXbzMEjuvbPWI5IxWYM81OCWMjTD8gmc/19hA2NCyQcznXmo6TBmLTJyf4NHlcd1dEhFaDSJdRX5zOlSiWNOHKNi5QClQDncENoQROXf+AVhzrwso3HFWUpnnzXXk16H9MLsrGT/rVDIlfuI2Gjin3CEhkoEvWEVSULk6dns7I7/is6cFMoQjN3iBJn7uaTJhRqj3OOQRduD9tCHRLqjBXWnwxyod/w+GCGXG5b/bfShiQMEi94pLPjxOIpkgWrefiKU7swttiMbpKo7ofxLQ55g4aZEUMjZbefziMxTzawS7zv59s+emgqk4ZuF8mud2N2YeoEyzzbiSUoI4Uo0pG4OJPHcqV4fZaR/mgZrlPw0ydAS+s3KlOkK2niM8J9Byp5s4HutlG0mwAuC8LAoAhneYwj3Gu+5nDAi0vMHnzlohZSxFL2kHUYThz75+KfJMmt5qrWmThPCOE0rIqt/6IcYKb2NJF5j414hHky6/OPyf3l8tVUQY3JM01kz8vbTo+Mil
`pragma protect end_data_block
`pragma protect digest_block
f886a1e931b224b53c874598174c69f117eb592f16735793e90d574f47e5eb05
`pragma protect end_digest_block
`pragma protect end_protected
