`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
PNdF1sZ/nSA6flMtwsH+qouwdPhS53Yx0N2NFn0rQjU8RSkL5y/xxuhf98x0kf/8tNu08izU5TJbg+4IZd9bvUWYyEkMYpdwXrXdJe6j2yHxBHhDVzO4J6LADJLLA5fGKlQgVDXG5R10x0lSS5ISvSfVLOQ7c0u8nRf2VvR0Hz9xj9kBQ6k6Lc2LGUzbW9uI4FFaxBBOMGd4/4QBY5nJybh0GMfG33QjDNthxXm6c4hfajYzykekRkGoK20+rbLVa6p5G5/QxC+jfqVqZA6b9oAMCOZzdapWS6TDB8TclX+YtfnfJ+WlMDgu34CJEYLZTNrIOnHwl+nkDuX46JnrlkYN8eskdMEjNZTARETjEd0OejoJ4hznLRGSUcpG8OigmITKREsqUAcd1DfBB8r5PF2bhpG/C2hIvRL182tdUUCgLxX8wZ4mjbsSCaCWyBYqell5+03RzUJdexbgztCkAew8oAZo8o8PgOnyhT7xnIvhaFufTAAz/+1svoimNtrIGuxhGUf4XmgofRW6/VWRvAi2QrFE9PmgiS1nh+NE0JOFqmK6tnjkRBk60Q2VYZrDnYxNuL3RR3Yvpzg/G3UjqXzIfk4SQmXZOVVCC13YefnPakm1Km7YvqtTl3RpxPdsQvuYs6FjXeqWVpDFJSjeZbF2/ozq89F5LrleEEYvpKhnETgzDB5pXHpxOIMDiVtaao4Tq7eFfzwyjex0M0cCqTy7GprBafwp3u+xArBplQ3Or+3f0gcPKBl95BNUyEFxGo2WzYS6sCSRbSRGzqNUeYAZBUgkBzP9C1rEyBfzt6rWFfj49Xb2Sd9380aT8aqHSao/b1iATEdHC2G5X5SZ8MsbvOvZGOpTpjzPF55/uCnIHdADVK8NUBZbqejj7YcHVeDGR8meytfI1DosOG4d1VJMcPnsTpy3hAKnyCpam98JspzQlNfbIo+6dnUCDKsOWlmv03a8nyMF/D8eENqcyDWrF3um6h8vklLrE8pcArY6mDb0GCXFtH6PZc6EfvKAWGi9ZI6QPIaCr8gMyWaRPMMNO6OLQvIe7gcukW6B44RUVxHmlw6rXdagnhBLrab0/3C9ZQUbPXv60kMaBC49SdjYl50W3JugYsJUbPI/z37n351s6Szpjmh2+UYYdTaEZgTUe1wfBzQTJKY5MpgjjIgoQ985Ecc1H+6jBfbzjSUYGAqNYHFyaZBe6tRvMqBMtG+LzV+G4HJbJI/in/Ul/pwOqgKXJWVXg+0BuShZok8H/f0fMF21NuyI057i5N2AiqKTHnRJes0zPefOTFTRp5WI4rKYslvkIJ7OTnDA0yLDr4oFHK4Ybxg/hdHk+vB/wrkV1vVp6IonbLmFbBGTIwGiaHcSz0Xj3kRBSm/5PFTufBYPVw7TAOuWD84hgPFXgR+tvmQIQfpCUy0AnmTGPpFZcZK+/0iyrWg/TD9mJ38FOYBH64bRV8mKO3FFrzRyUr2TZl1y+Ktdeo+B73qcNW1ktD7mSTxpRPmo8tt24L+0uYLTi6gpjVQcltdaevggMPVSQd2HcBs4dmyhJpijdVi56rCoe6EF9VOHKp/Uy3mPWrn1VwnBYKpGckELw79sLL6ik5g+Y7tDCSPcWAGm1P7i9wvBufKlt3syeK2uxw0+rIiZv9QPWE0K6SGN4Xc5rylY0kdph4/ip1b7h3rkSjutJDMdT2F8G8K+Lp6XfHUSV0wqkNbGqliNfNS9PUZQlnOCJ86t2JwtQB9XITyX/mn3uE7A9NPljJmNgRCsk2Iufx/AT66zQsJj1W2eBR0WOrPui00CyJBSlv/DHzXXGsN95ul0bcbn30HOVONosFdHZ1ho27yU3FJE+er8fUXjy1uN/GGLJNg/iZ/rJ0eOSnjyFj5RdmTwYI3HUqMpUwJXCXLqdlXcD5K4FQQm0i3tQmZwzr0hSkeUhRyNal/R4lwSBwGUHqsvteuruOoz1kPdP0qxYRPNeQkrJwNQTmHT5VoSnKaO6jc5+7tK2EeGcrAGNMxejGhCjm2gFAfWKCN1000HmhAPULIVEP7DcEs1Sz5cpjhXs6ttWOizIQMdwSedK2dMjagE+G0jM1CYHaAHj6K9oEDmCxrExSGmcPojvIjd8WKauUeUKRTI+asTuXlk02OjwKjkvpsYFxpyGAL2hVDDLuMrdoasVuy6/VRIg5yGa6OjBiJwor0dXMyayfM0RuiVqaZztNRnEPmHcrHNo9fbT7RAGDfkXdDzEUukw/Y8uXR2Uka/cQ9lQcv75AObwnnRhZ41hK/CtKarehxZyz2ON6fQWZRgVnhEI0j0Qh23LTZCd7OtYROUz+GBLCLn3Egjz+QjvmQxhgjRxGCbzfXEcknP82JiHnOO72VTLj6up7VCApyYP1gWj1uAFZnuew9p3wNVdYTAGv7dzpFXXYcXSkwm2aRN4de/b/MrAHYonfaA6ajHmygdpZZ/50ckcI/yGGw0+/rSjyflDA54EhVgKMfd01O0GPydaineoAgPH/aNWAo3+Xl1Sn2EukbOHwRamr7QL6Wu54EPLS0974Vymdn3VIJk/OpGJZclkOvWo9mZPqHunbM7g5e4A16NO22ejhYnCkKtYyZQPmsOYL8JbbqMZopquKvjegDy6cMFoYMpAGecAdOCWbkrQKsZlV4ndL2gunkB7CyIoUXtCfb/fAy8pdDdc0zTWJ4ytGTiTOBHVpPDJwEDzFXq2yr2ug1nFUs1RdWHxGrMCWyv5QK4Prsz7SEQUe9NygwMtGsxhFbaenSxRIcCZDWvsQER8RmKcCtS0qh+xqSGMRloC5Au3aR8RwqpYasjtxH/oMup2/GDIK8LgZ2iaYjluE9gL+reevy9WrO+77PspSKy/UHNpC0IVnSPBQgA3roKP97lPEaB0N/Bqx3bOgXOVGbDFcbnE6AaQ4d9K2Rk3Q3DNIE0thDLArjifsA7IhAOZUJK4tpRu2aR9lfKx6on5n4iC1DlwcWlJCFEICZ/qbqARcZzXfXLIychtRMX+VDBCF5zIJxD105pUpafYdka1KuAKiRakLJ6wEjNH5bkxomwYY5FQL7x4rbWlYIIC+oFCC+gixzp1PqiS4rMNeLrdaqNyW3wN04sNA9tnQnf8gows0R37BDd3F7tUb6SSY++CHHWMDp7tCkrvcaMXijLbd17sTxLgKMouEEn9j6bMEzLzbAyBhTcNFnlL2uCfSW+NxXySTlWm0IwPbSZljP17fHUerNuzj4Rl3m9Sfu360nfHA35Vawa2DlulKnzjAyyx3b+SLdRk9gGOMpB3YRctgMnP2aA4IwOHWVu4mzyqERLdyi4ympNEOnqB57DWzq4kUhTVeb0sSLPNeexUw+XqZgCFEkXVLLodsqfMw7X8mSdU2dHsJ0RTZMKGLXqL9l4F2bPeB4C1WS/5jZHs2croeh/VBMwZCS0Gp78IG/vi3gcoPKNp7wfPZUQMiwOVziGGpTaGzq+QKBbbkCmvIN8rwMFiBB8hiOS7mqUshs1b81bm8jzw3Zm5iTpIZDZAJfQr+fzk3KvuEDvY3i187aN5YdxoPDSZuCf4FFDwgX0S+UlLvThKT5HMP79fbA+Dy1feFRcI70gydjzvh2FUk7m4vdIIyfvdFKmRx4UwdZOQ8LOZrHX+qYhG3c68SEiPLFDWpYElQLPQc2CH4+EMWf56g6xjDvmFOdXL6Igit2mlTxxXKmEXcEBMPKAXsgsgsveXwopIZ/w4SMavoMCec6KFt3jZ0zYemEMdKa5ZM9av3V0la7hetvltJ3Lk7q71/dPn/oMstezLsfXLSwcAJDf01gzCNt6dS5Qkv25cC+LPzItK8iH6Y9U7MEJZmXyAfTjIFVB2kzhCEd01+06HV1Yx6UhDt0wPS0sLQbg2As0mEDbAluy/X6k9nD0OKwax9FcHfGwUmnFfhcsjpukFJ+w2uUagAjS6oteOldBs8bogAlcJnUxfPfyPDM4Yr7Ej9ZLm1GuDncORYcs06iuotPEuMsgh78+EmsLbI5GQySpJI++onoOCsjM6KV55hZePoAiiUTXCbdSaUTP+uJcEfWA9bG8Kuxyl8hX64o+3/C4UG8dosERifYwI5Ok/giGy7GqkeiG+rTD6VZPkKcXG3ppF4wU+zr0EUKKInU3ssw2Cfx7+08c3ZnLFyJOYVfFm4f1Hmic1nPFRD0ZPiuonmelgvdVCm9kmFDkvY79EaCnqQmko+dHo8cygyQu4adn/j0Y2lwlMzxdohdLHYci1v2/b2Yo0rQMiBXHmYm2AYrv2pos22TXccCUwk9e7ghLOMA5gHLMxEDTCfgLFngnDu1dam80tYuk0TGthmYNufKXFzx1DfL22xot4j4KDJi6c0iW/WyV1jn6jAp5iF4uiX+bd+ZPmIi3B8BkSvFUiT+DJkuW2+UY0EwbJ0WJaWzBmuQ3Ipi2K9OXLe3LZJKUHYkAwCLc+89Lrqy6kXwO4Em8EY19bN4eRs62UAGVDsIvFK9a3QstsLSyZpD6KBWmL2/gN6bOc7nK+z/3SccN1g4eLGC2nqZs+WnLVT+SnLMb3fXJFFWfhp2CpiLnikuX2U2xehaQlCS3OL7KaiBmnp2/94ev3AUoyW34BgnzUvpyrbXSaf7kJI9dmcjCLOy9aLGylL5aDHRK1CKKxZL4P6pPsqLYDVqIOPBer3fChbZvgc1nEV35zkp+wQWahEw2tzIN/KeUh+74DsLByMLrLBYzNoap8wQ6GCmyBkAUZIQ8LK2pqC1CdPo2BgCIzhEGlloNVaCqcTTNe9uANGtX9P4WH6xsjKJb/mgDeHQIVKOfBPL4aqO9/0DU34BVTxcNHVx1a90crGDJTU1xoge54Zgea9wmgVAZT7Z4XZssUgNDZsuf27TJOiukE6zihycWk1MMNhN3XwjbP0PlAbM7kH58Syfk+uadtVOl9VSWb2rVyGMeUkhy4sKvG/5qUObCExnaYB/HM0M9jJRx7e9KHpyQS+YRy9iq19Jw+/sm203HjiEaRwXMfOFmLcBAkzhyAR2XkJJkcl1iwy8KqrqiLs4sRbxQChvtchYZQr8H+flEh1oFwIMj78Ld/SoyB6G6VZDaEr3tC5mrbFIkuNYChVi6/hbHyJP49GuXFR12Sn/NNENq4x5WSGSy1s9vgpZIbDPE2o+U/9gfND2urpmUN5WZKcmUTXFd4kRh+ZUPyCFE6khoyfI6zyO4j8S3LRNIQlr7VT+KieNShYKjXpIFy21GR1lHTvx/TQDN6xn9PjzNJAodbdWkQM8AilgERZD+vFw9366LmPRVC+FSS+W5FIiw2DIdN5UXXxMJgTLK6cPCTUkarADwuD8/uTWryeMZQtnj/AI184wny3vQ4JmeTbSJjnFY302q3Q4HLa1lNX58t8ybcXUeXYIJdukDhNEqbuITzf98FcnpGw4rZufJcPYlGDzvQ57nulpl+jinqz3yH0BLLJztssE3zzaT9KJqJsBwPqztIpG6CZxM7KPcPczg/JOBSaObql94ESC0pgKPMgS21iMD3aiWGEpypvSl8XXQPZPqWLF4R5+zFylkQHJjNEulK7cv0sHk7ctlbrtpW61ULGjiYVSfH42SYH1au8BfgQTBgt6Il63Frox3poflcvKhFChuA7GeE5y5LR8z72bZphOP5IW5634Cgh4UBs/82KSIBwQcie7M0Cl1WvdPzGU5NaGWkzMxOhDJxbO6NBU6zCnnNPmaXYghhVGMXcynG2ddYHqqKc/No6kuGvasA20zbw3YR6uqU47t3t4zO+dEWkmZeQOfK4MxRZu7RbXfyt+nun2FwspeEA1uZQ6gz7MsdupMA1JXOCsK0nq595jpIrodS4JWR+JhydGm+fEDTtToDH53BaFYbKWAH5FxzmimtrrNdVNpL6Cawj5DyZ+oScr+vdLK0ie783XOSEDy3pG0Jd47QaeJgAbDPRyud96Wy54VWld5UAnaQxpuv0FtdDhhlmcBC4FmeyrxTAJhb9+A1UlJbHiIhAJgIiOrLRmdEuGS8OUHpo0OekYjtJ2JDLeWFuhgm46kd9/jnBbRlhkJSOTmPnioSJMDR6pUCLT4E3BawdAcRfCc59+F0H5QS5bImW6X9gG71y9V9cIVxEFPsT66XPXK3LN9vN794rfOa2YPabDrpOYCHCCjZ4gXU6dIpXuSWZYYFwjbgMVMigZuy+gwxFHfJ76TcgnFJz0MeqD9w7S70ljEdPuU52jw3l1HI2iaqERMmCTYsRLfv1GLeCAqzmMNazGDvzfQYrSUZVstK1qAadWo2eW6ym3kSrcLrTQ/mopX8GG6azBlbUFheS0AbjrDpjIqMOM1IfiJOX//hHivIQoie3IQYkRGUzUYF0AFktTK51aN4HHY+DC2qHBJMjzlyVkJa8nDAAE0JCi6JT7tilsmzPfj4BSwwaKrDm4AQT/g/TbwMtw20pT0309i0WA1BUIBLovYHKUoFPggguOFb96FVtHrlGGNa4WPopK/NsMH+EV6Q1F5I97YGrBVKb06mSYuKECmSQz2tV3E8PekG1xcztMUFiSNlE96Js35xiXmgxaq47xPZZHaZ8UbvtOJRCeU4Rj24pOTaytYZQExBYKLlFY9gyabUdH35bLdOVfkctI5KThyhjSxYjcbf/iQClH7PshrP/G38VviFgTrWBfrcC+CYE1sew7dd8ptcd18AImHZGY1rlueJJfP5NxbnCfuei9xwcZ3THDD1xLIdTxW5YH6oP4yA8V4YZfKUyL8fxWo82rr9C/f2tcSuM6oe1kCy7zFVrCyl1v/R94U+UT/wvSszbzPDcvMhiQF4I9qZ/AT3zNEr6ITKaDEoHBVcPwfAE87nzySzpK9TXFbLixCkbrxKbs2+SeJn03t/MPSfbWuTll7tL25/hYp9I3wB3ZZlqtCaWl28CxLWd0LU6IxdK2Kwp2Aszo+WJWwbMQdqDEJef0Lhz3z03HxZLTpq1pkMMBRBZzQSCnBonAKczJGQHfhemGln1TT3EYm0OQ5JWGEDF25YTJm7a0q3ZUZKN+y1ZS7j8Z3W9A0GVBSX1KgNVjb6INvWe1HfL3ipmEvdIcR+BlMGnpcR340x7s+TxpXtlBzwJ+ohdS0ah7Jh8IZVSCC0pdvvdq4qhgJwr4/9oL2nbQ+vuYL0I796YB+IR1OdmQdFVWxkwOydgbQ00qntBJIdseqGha+eUzrYkusrjALD23Dhl8cA0C6rzReXeQI2vK0YmiGg1xcri+T+UfmnmDuV5VHm8GJuaF7875dRAOU8/K92hssIhtsPtuKCV+9sHt03/Re74aLwMvNFwalP23NAbm+/dS8x498B8QEUemuU3w4CaDr3mvlBX7sEvFDQA2Lr1sSv5j4NMqTkXgTDd7QttVZyHoOpnr3hldaV2wuA/Ss4hd2RajV1u6HhAGWfbgqDiNRsULR8SVSQaKwaLPvdfwa+pnuAlU5P+dzO4YKzXkBINgfArjt0a9H8LYpq87HMAznE2a5KZTDrD5mkwZDT2R9v3U33Z9+PFyAYDFxni1DBv7HcqSHqkRd1Y0ieeLcUZ8Cb6kLYUuYDEkvPyetd2sMuS/xdYcLVq7UuP7pyz1LXWajolqMnFvEDajxAu5taFMVS9rqQAphI7hrQJTIQArNAKjEJNwG9NmkgFVXz0UeERsz12/6LR0ABzWzCeJu+ktJa1727eTtQiUqnuqSbWcxFF+a0JFYMUXKtrUQrHU0cWnM53V/C2GL7ChMgj6AwDw/iXDax9nk7ld9bBND2NmZWGIFphFH1OMHKGtIkwqYr0CDaWg3hx+VG1RLEgQxsoXuzzabLJD8lEVSskIwiJROrMLHU7gXK+RmO09sehXOVTdwWsrza9U0v+sce/A4xAt0IF5NcBkGcuGh/nFxWVZiiP9v0YBbGGm+XKiEGoa3dcEqRN2fatr7gVjdFpcLjwKN45/tqnouH3gWlv99XTgxeLoGIdveAY0PpljFjpOimgzeYNzMRLVSMGHofUqNgei3/+95TNXrxKIlMUTMO3p5Li6ier4VlvnmhMtcr+qoFse6KaDfjDh17hQk01MLO9/xTFbMvwJPEe6r92xvVmZqPKzFWmLHSUSpO6cTgxyOXICNydrt+5+7NwxFgf3VAg6nTw5lPfFSwltnsmFSGTkAeO/LSBH8xwd0Sqg8RrzFKMt5g8K+NRWX/2SDObJREJVKBLsgFFqY/TWyxTbk9Of6Z3dAff4SRVPLYx2Ai6jf0eVAG1dEYW6kdeiEHC+HgwXyHLAMrNhGXAPMrh3jioDUl3hhyRg3+PNESlfkcBk85JShYDSz9xaxgCLNjpz36uRhEWk6eVuoZJLX+XInKPh4ZbiWjm3mD6zBGSy5xz4Iwd1GN9YeYNPlW9tGhjk+o9G1We3mHidxL3AV6Sakto5TBNXwdO6d6wrU8Oy+6tq3NJDLp8AcdzlvtrCRgPIoljaCl8yb2eivRNWFPBhxkkszRZaOEs5FD5yXxXaql255Ypk2c1PXc8PWUgXZOUX/0HG30uwfGqf89W+nVc4qkdi6nznvD34T5YzUxFrB4Za3yIZtH0H4WTHbDdUmipRro+n4QXpmef0JMlqeUA5LHP7J2uL8Xfl8lJyWs7GASxtnDQXm+Puy0RYtHjKlXK8W/18c7QpibzymfqEYm/tHlBtrxaKH1GghabH/7s7sleujLg5QB6Lx149c1DpH29ZLbkRB9fieIHick6g5TWGXJ8smUprEq3nMsbWFnehlmzNQMMYr11WBWFzaZUJpyFeINTRW75EO6kWBood4HDrrXZMnASQTZl4wfLcv3UP27EFnt3whcz1RFzJnUPMLKtwl8vjp5Qji7MbgKQs9ZnRc6KdbCfV7pCBfh69LOOkBUqKdkZsuxoJt4pdO2ANKE3F+sERPuQQ8b4tpQAmo+bzH49BLUB8+x8/IQWvKTG/BOi82OTPyvsUgm2oh0ZUjs6A1Y7Z7mPHwC6WlpVZeexIhaP31lUPXDUDWnAwmdVwudK5q83y3sTFbvh0BDbGE+qBdIp1gRl2qTT5BYcwgADeJfwP8ipZ5E5ag+DSzCrm1mo80uSz+slgaMIqZGfT+OPWyAxY1CPl8IOBfTWmhy775Mzn+vER7lyNPqhkswEPLC5xM+RvLjhgohglpVsq3lMw3ZyixtuAa5AWqQBBmXzcc+9pJuN8yu9Q9ZQlJsgQ5eS/jNVZ+0nyXJ5NYV+ivQAB3BieJ9YL0t+PzoVoS7pZK4GFv30OE8jt2A63eJcNbobStIgo43P/RQ6GWU87qM6oCl2VUebu9P8Gxjkn4g7tNv+xqsyE5rH78Qn+FZYLRkczmQ6dd7gCN78I8fIQxcfzG9qTKKX/4cLxirsuMIVq+LpkZtO8Ik19WbrVfAiVV02dpOv9c/8Gfo86TZxtyIVAqz0a0IRz+lfA0WCO5wazC9VrWbMRxwjFA11PKWekqgX7BZPwWCEiKGvQSrLnQg5lta47X08Pe4e9cpfcKzXOhwRwLNYgPWMRu5BZ01z9JMq86LOv9qfd8CVhv7u7HgApT49kd2GtM+9/BtmKJKXYhyUoICSc8xVWJKnqSUWhpubQ7FmUQ8+S/4JiGbEnac5ktaBEci97EnvxWJX00fmeTH+rD0ZVSPhbdRskesWvpmTx7FUoRX4T6Pmx1YgUMG+CbuHMWLVTFwMcNKqflsSmh4ESSTVEVFQ/Tmw99kMB0sRy2ziKqm5VfWrgXfrY/5/U0Nsaidmixl2uMoJp0J0Zoz6i5k5jXe7Od+xEa7py+IGAl5y1gkA0Lb93Lgtd/ulI2Ot015Me4d/rJT9Pgduw0iVoGKIgALX9AnPtSsdJrAEH2x6YewCbVw2b4kiuncxTtvQeU9DBpSuDIf0XW5MuYzV2dUAJ3qxXExxJwnJVDYYJ1fsgqgdlXN8R6E9kV5X3FB1PDF0sr7LyJ8gBzjftcbUTiDT+vXZHGFJfsQSCd3QtB8r0U/2V1HEq96MrPZOV9VL4=
`pragma protect end_data_block
`pragma protect digest_block
ce2d93fdb251b6845881c16f01798dfcaa5d82bdbedda36d1bcd401eba33c17b
`pragma protect end_digest_block
`pragma protect end_protected
