`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
PnIfgOl80noUFbjxULMjkLfib61Jh28/m74TpiZwwE1FFvfj/n4rCtQTCPG01R0jlLtUZ2F3aCLor31dOev1/xF8vP5cxyLbPTXzIsqIa8U2WH/JdpwmmrbnjuUjd6xWwlpJf/e1hVflmVRne/6i//c3VDp0mAKNsTEE+AU0kI/VnjEvwCCRMLG0p7orogGmlKwBmZCzBhCieMxg5XjzAaa/H1fjtATqFwtBZoL/15sS+hPF9+tZq1DXOjtx4MD5Ve56lt1EIPfghAGbTkEmM8qAJEiAFRdyj1zYMVTpUtZtCX+nNClpG25RuwRc+/VR0RovW4rQIeexvjiZ7UolHs5RsxTC49ZxbqRI9Ks+q3coqIp+pA6KlXmD/zkG04P5Sz8/phF2Orz/V6DKoCm76AhbqLmCC8rRRXqBoLuD5T9Q/XtS0dMiFgdqUIfaSmQgPaWOK0h3rquJ9lCSaIHoXYDTlaApFUCksK2PPQLrAnuhD5S0gYf7MjVbbHSv3Ecfj7/rzuIIzvppnvMEdLBXXi5Ze6DA4ZuaJ5P4ooPAJBN3hpMK7R0f1FBK2EABTYCRqwXGoi7cL/4ocTiYbX2EHVovoGTM9t2mhMNALzQoZyfpgS2lKDnGNMoHXyEkQACDhjoJ2CwbUr5ZGKQIs23Ttxum+c8l/XgxExDH533PvG+i+huxEZby1J8i9/SNUVF5Upg3QOvPGyYumcDFedfT2OsCcf7xFXZcVkeytumgv+VRoT3RlKjQK48gXt2ru1qn1BbIL246uzgFUmLeQeRbU678erfJtcvZ3s9n5UpNza5dGWn4r13r+hPVa9/oDkBHdUGa+gjUiZ4TVzxOZtn7a4CMlzK1LqqXbRSdQOByqBcMMXKdc3bDNWC0AYMoAj14ezl5h5Sbo4SbKjC64E9FPPmN95NtUTIovYQ1M85QHu/LXZZaFzDHn0BumqNG6j6AnTeLHHuZMaVMRB4SPFcXRZmUhx6ItUdi8/FMuBR5Hk5OqXwX4Sp9IbJfEHdeu+gJ3NKfR+Co+IA3VOcUophpz/8+QlsKrmGSZpZDO8ErNxVUPEriCs02e6tsP58eUj5mizSuGnRS3BbhJs9+Bpk6mLqlox+Fkv+7gGWmSl+oO/d2fxNlFIB84DfWa2vOL9OLGRmpxlAkOgZHVUUFBg8/NL4EJ5ZdzPWtbtSREMvDtkZ3G1/5rsh5kQFXGCwmVp7G4VTGySASKt9xlTCy500PQPgTJDpWKIS9pkYLQAn/hOep4wCmdFNbGUwv2ukA0ETCPabS9WLqpb0UtQr3geCjuLwa8wiZWft0CTDJB7RdYVjiZ+5m9YnS24oDVNqekzzWUKO59/PBiXYOtUHjzUmLJlPb6Pw8KnZaI+cA1Vz8T9Yfew8GFbocwjNk/TcKQbnX0jOuMdq9fJ7uLsyHDvUF1vSkCmM/rpya7F2o3OLmpLj0I13n0jwHf/Y2Q77AZSsBlkn3Y3JnB5e3k1808t8FqCtmu3AauUEqqnoJjRBaacWzMsBo7i2a5R+mcBpgLVi043NXV5jHdxVfxt/JLEU+DMprYGbK0VqG3KJGXDecUPthfRm8sfd68OWscEx5HsaLTAsqfTWwrvqE5n3edzuwQ7tvE0pQONmrRRkXUBEVUQ+yzeZlFOd8lztRJQzarIqcvpGG4ER0wgB2m9/Cu/UPzlmXYa4SPZ2XZE7+nBuvOfZOg0xFcjXvPrrbXjUkDIZIy19re4lvZmQ9wPJqwODp+OrkFOspf+0FBcqXv2Fu0ApSRc3IBAPozGvXWuoP/c41IsH5oUjr1cPWUaAhcaBpSuGfcUfS38wBsDci7qH2MtfSLBJwhJgyWeIXS4Qa4CfJMqPXUWm3nR3HpW10Em3K26o0TD8gc/g8Lp7hHPW1+WIksYSNeQwkLs1Hm1/VPnX9NEc5EjH9BCVYb3X+PEp8yRPBQch7vb8wHRFI82Xdo2XoS5XzJ62NxuBkOu/KtBYhWVd2my5EKoQMDWue5LfGbPo4a/O6lSbKF7ptsYs5beRr4DDhKDYs7AiWft1c1dlFGyQIgZrUxe+mtcO6TRMAi/VXbwcbCPTU5ILcjvPIXwxJJYZUBxml1GqdZs3RDqkXis8uWiB8mODm8CdB8jsdg4bgmeSkxTEIYBNjOeStaTu5WTXoHIyVyAo8D98xicylymYxLdXcZB3h8stYlttotznQOS3+Rh6tuDrF6fSvbo2aGQmlKhg42qKKsX0Se5F0fi0cPyE8Q0mL1Jn707kDWHPSzLkVS9fVPl3cE0d4OR39ZQob/JCauwf+ZdL4xg+mjDSXBh6MHNguDUw7vlaqoLlVQlrTdbYlRQhEVS1reZoyjgdP4S/Laz6FCFVTwClhHU6PGsEO7KXxzDXR/YG5ExItlXiu4PUKk2zT9WGNqL5hFG41wsbqz7z5CGErJ3jtwFuofSfFpShX2GhsEgj4uJMwMxvShnI8te4mt8AjB5HLaWISGbtLmPbxFSt9rFKoqF2Ca4yFJWhh/7tGOe4Go5IIiTf3fc4FWy6agH60eYp761a4gBQi9LpqQrlYvCBxkYOp2p71TdD/Em2xe7Cuu1Kb0syda7GO8UX4AEpXMI9eoQ5KLqKRRNj0A6T8oYMb58XWSAu6QysbpS6gKWcGuW4SayTuiZ4u8PGWrLc5gA+Xl0iKUtgynO5lcP+DlEQ/m/7vu/5pfOIrS7c/A8c2AD+TT3bcNT6ZBBIgyRPKIdlgfV83j4TVeNnJPf+Lu/m42jNebXW9eEcg6KoSy0gUr6D22Grbt+lsopzBZDDwxRAzhWrK+azJuTKnseCE8JINxpwdSvZ4AxSYystr0PrhZHBn3/Vh28QbVi5O15TTN6p6Q7VLRnXEPNTbzGn0TLUFeec0vqxclD40nJWuQQCEUlR44kdEFGIEnCq1MUWceh/RiAJo7NXsPA1zbWaH+7qiI+QVgycwArinrQIe9TStXCZTDa5IYr2QHm/NaygdFQ274Fg5TcmLi1Idr5tKmEhznEqyme4Yoo0A7W7AgWEBArYAtMEvU0uIntnrwRB0W6jSNByeoiecAD0j7NQ9JF+VVaNZrOWF+CyvV8p+UisENMvIitBtbWHIolIGIdbpEKm6QP4fOEWU+BRVITOAo6AhRsbTM0n+pE+Muqz9Fyu0kJKRJB4hFK4xjgvj2MIpE+UeMRb/QV9iwnt5+j0q7woeJ9BOclM/yFbxPjC1N1w7tsuf9SJ9R24//iDen8vXNKpclimEd5RsysDeci0K/DdO+0VoslKrU+i9pqnxO0paNvNu4AVs+pDA5LJiO3YHrW0q9GRVUJZ98hy2MIsI4q1m9iCRcudCpW/u1HTdKJsxLGK4mv0Xc6+/bJoPXIxj6ymzgRERP+17MXkVvzg6dui0Ikixp+ELYNTvUeaBPOLeT/MpWKpHr4YkqC5xY4vhScUXBL+6a2IEn9IvtLNzsVijvrFaRLwEkJn3z0dWG3wL6SAE/MU2OH8pwte8PuDWy2tybmrcUVHhIV5wl866olDgeiPlj5LD8qWuWSfle0veFO5JrnwNVXUmubDtw7BHWzvkcgVuGX6D2t7dM1sFHQmqLpiKTREBgifx0Fio2tz3YKEZmczh+/xvUNLfsYr2BXljH7hIkhJsKu/T/KW3quJ+zpR57d7X3RJ2PqwYGVZwCR8ZdM4y2BocuIrDOuPMChJnGxmDMijnn8WyYB/9lT1pxtHjk2qQQvNM0+bhODb925VIYkM1bEdY5lX9/8a4JjIeWsNO5b1kkg7RVeaC9GvI0BDlx84PL//1J9hhZ8TAlUguYF/dFWVyElROD85Ep9WehHXOjUYRZVgp2YANqurZCuSE9e/nm8ufo2OfktyQdQYhUcswEQeNgAXdjvmlr/QvSfEHa0DE93tz7VXDJr1C4o7fJjKkKmqjfA/XRlPnDChUMDpgEuVCgAKDSb1VcvsRF2pwyyTc0KVNB7rCsBzPkZchrbThXMxPSFQgDkK6t9qGd3p9NXkxrOddB+LKXIlAxq1V2bskM6hYcfotdi5i02Tpm3eLoolqbtJh/djYpW7L9vNq5tck0kiEWUboozwSkaVHc2O5U3E42fRQsk6ya1J0qXYXYewZzAMsR1mYgaBM9bQbrUap91Rcx3n3bb8HZ7h7Q3T7PWTO4RvUE4tt8FwnU0oRvCdlsweeFzvqcBJD2IOL8P+w7epGXIeVunxAzR3JebJWEJXx+P0PkNSsgYJyRcQEhmeg+Pw8nLYsXXYq7Q4dE5MyJfTG6Sp986YZvYmaWKtI0Is6mZbPr/JnjuOTfngD4HzBPjErbII9s+ljRNIbb0cygG+g0VD8Qy5wtZML09SjyPLoeJ2kRV4/z6vlVu31Btrgtmk+Sll7seFMb6ImAe3HT9Q7nsfzVKdZPya1lBKM9U85GLdUR9pNicy4TZ0lYajKaLygL9eMSKPkhSq3yWdCOetXaK1DaN+MbzuMZMkgDFcwhecUmVqiX6xtw/3h8TfiurEXWOJ1Aju3WrbZBF11R0/ThdbpvanQCrlQjfwvz8cRXL7+uU6NaarT0trwBoIbKbKlzS4vC+T8CvU0yX+KXRzavNWbXTWlnxhQe1HVGJkyAh8zat1ifR5se527CjdBDoBhQ9rLh70nDHLl7SrV1WaU2311AayCC720ttgYv2DKrxhdI5EF03RTckeESW3kt6WqkYExOoIIg9DDZcMwMiA22/dJfhDQ5nI6RDpypxxr9mwmA6Z/LsrAtHaffVWWZY2a985MeQc+zh2wfJz1rn79ete2WXC3hDJn9aq3Czyw8RxpkRoFcOsU1qzZ4EBiNlBOGeny5CR/GiG/9fiP2/irmQAVzipDRA0hV1zMK/IGQODkJ8g4VOZyqLIOnmaUqi4Ud7l7O5WLbGIe6lN8UePD5OnoE1aJy/R0OLyLZuSy3ePWuxdyGYPPp7fEmsld4twXUrOOTGQhI3iKiJo5rXCphf82Z2tdyruHjagrvYBPTVPRLBw/W3uZJ8rW9ck2iS4Kg5irl+f5Dl2nrl1FfVW6WlRu4L8wE+kKNGLRtPR2FDg/RbOwOetzLDyO+wsweK7s59vqjfS4Ygw105RDeXADBxEVtGP0VL+JARdZy9C9C9DEzBiU02jZ6uiPr6LvyRcMJY7tdqaA8FyPizxnvSlZ1EKqX4jLRiyxzm+Sf6EbxbnklH51TLjrEZrj92FlRSlf0d1a8KPB1ItBtTY6/RP4FCKvcic0cwb6mKiMf08c/EVO+1wloamVlBKi+KeRXx1KYzZCuzbeLQ2O+vi8DRnXNKMUh/03BAn5Pe5Qk7OIRd1+EFTaR6ws9Pln9yJ3O3uU3i2GBJvg09ZoPQKczSRjxg/QMqRFynJmiG0WJolnFMFH5B0fHd9KpzEmkx5i+QSNSlrxtmTUvwdQPQdPhS9bW6fXm97tmPrZqu2uG7l+jBAerTrXzD6FzO2K3iXVoKvARdSsCkvs5o2oJAbWwepHeF8tG42aAMNMItfCEVDKgD9Jvf+/IDFzZkrf1GT3DF0yJaSbv1PXp6oJSc1FSw+ndj5iekocVXTEVahhrxzOJZpxpwpFEafgxhFZkM0qvG6ZmXuszFerhYFkMfLxdkw7u2HBHT7LhsOHcDd/FS87U4gTX3NgBzmlbXbQg5cNrlfLbDkj/aeJiH2XIPbtsvlDz6RDLLo2i1gvobIAEbQAwzDdk0YNrgH6kZEc7VoGKtR/Cwl+pXmfFAE7tzIHuO4qO+CB4Grhayn0rvrcoBKwqBwEEE7hk5t/sCmzSjgLJpMZ84HFT10RPG2+h/AoY2/bLpaE/EWNSAgUnQxYBceTSwgdzH8TaSJMeJ612B7qxBKxIqOZh98ZeCtJngOVUGsXdSPRYYnyrmazhcbujPTAJ0DGFp2FIl2Mtrw/grExLj6LsXNsHp0KScWXuglDdA0CLpWh1KUjIJNmy/8EOPfs6Z9m5ZNWsDbQXy1WNIfQsUgCZkRpnhvHiIcjd2IrCoyleEfETkbG7PWKBOMZOveJeG7TN2uD22Z7GNdrlsY4FHXbOA53c5dZBh85D9s+MNuh4WFBO2fvFrKszxNs4hv0Fl5S/d3GWXdwN+ArUcgz0VzvNmz35YrSQAS5zJxROljsUitqJw4s+fTeqFPQDd0egdbB4/B/phxEEgVUE8uCP15s3GbBj8JgMa7hG8WOJ8c6N6ogKoFWwUssTuHeOQrtV3fu61pTIVZM043QOcVuN5Lw971fIpGxrim9vxJZwxrDR8sjcQjRNP8W2oBOp1v6RgYDR0TVbowtNEMhRn+8QucIfk77RrOEVhVHtpkZ21NVyA1eKqyBxw87ax6w3w6COL6yyDX4e9NmdOeMfsijOGnEZKKGNDZrDyrOjoWzX0di7J5zg2rs1S067g2tJreuGHJhW56jeNbReL9TVE5QleAVWrXyXZHV/57Ky+laB4qM5D7wGCqszuNRqFeSkPTAaXz11Vmw3IlV5g+GLSMVUrQ49KiRqOe8IgFC8JS/ZXRuvr9QBxJXPfSoh/DqXkfnFoegxzgAeMAz6sjbTWh7RKrf175rpQ9PpunfiRbzxUlahDmIMXOzImfeuFxVopfRe3fn0IZVs9oL5q9m/Y1xPktjJBUwFKwtT5ZSEuWH6PXBqiDiHj0UvcNAsvATHOdpoaIJ9/tNVlxrY6mL+LaZYzhQpvsMlg88jxp0dJ691iVnvmveN4s4OWO7OJyDA/E6GLT8Fjiike4H2CaqN0qnnVhM5Md4a8nXGffuE4TqkHwJt78vfBYJPY/PlL5Jt5TKPwHNfBnWhNVb1XY7XM0P/g/NmwyjxtNfUVNfBPg+HE5Rb7emRSnP5e7K5HtM3zMIppy8Z+sbWt5S+TOo71xJAZwb1Qk3gcmg6joJtB1XFfsfvCA45IUAsurA2ayQLwObsUKRqD8GMqEgfiZw85L5ykMroZyVyJSHb3lDhJ4ICCn0fzutk3M4sdH8846aUl0t9iY+Wrii4hYa8i7PhImoxLPVOzIC9vBK822Eb3/aBFiU9gIwlhjd4eNFCG0TPUxUdZ04uvnOQDqoB7jOmJULKdD0GhELhdVzVlHsEpDCX2ygbavAb+d9QmEoMs31o52E8pV14883NRYlOxv0m601YDn9PvEMBkScYHzfUiMzR4vJReQJd99w6q+ZJ0ScdOK5/FCQ0328dSl5erAUk+ZjqmWRTQHE7dheHl2VYVIA8x9eNeUjkfWhNO5RedJKuzL6gMWioONgvJfZe3vmP1UuqdgDJteYH2bSO3QH1qOm3KvVkpSdTnpqhOpJtQF0SX6junlO2eU44iWvV9hyr+rxMUZUB6rHVAqypmi7repa1mvZcyx4jDYTZPPY0twyKq8PYUyPEG2t7lq2rzVDLzcBCYTjrqW99WM2zhVk6rIOQdzYnLMw5BjqGl8sojY0mYJ355CTGYABjcsAI4VPgXaFET491Q/4gKInGnlmf/pqRlbHo8tmgi8yO4DUJB/ihlldiSsRFmX9FUG5k8AGnA4tBJeRMVAy4nft3OOy+jorvvXxxdU10YVJAA6TQZPwvdz3C1v95TbJyv+7hjpOCh0+xmpigOjEOBvqIa1OdbWTSR63TNvYTxc9nj6m15Yps5Yjme6LKquDDJ9MGHxXVB8/aHhHwsGntb67kfJbWSefyZ8+9IM1HN1CEA3RhKDH/Ase7xPcPvLIcr9q2GxfBg4x9uRReVjsyj1FKakuc3ClCg5SldUfcSkBkUUKgmHhSfbeGtwCw4pBjDSoZqKalwP+tbVRUNF/4G7Azo11lrie2T/ueD9Ivj+RdEukKJgz9ZuTJdn/YyNHuPY9qi+4qFkdVshCMcNOqBvmp67ZITHY/grcAHKt3Ya/LNMhh++L5Sh8Cw234Y9ulqLqyEy9F/Kle3hjVpjm3EK4vD+6fu0DAeNkIj5V2VqrXD5L++Es0h0N4b/NK7aKh15yoVjgK4DgYX6JRky+SCdMK//ppENoUjlWretGkBGeIWXUkKDcUGiDBXJoGd++kp2LvDpdFFQ9s2L4OB3jL/K+dV7q1VpM1x2C/pTsuhBy4/giAgHGo8TmekXw6n3a1uOAC5QZYcseDIlYNsffB5gOKO+97e5lifJEC77FT0miNEIPA9EYrwGsWZ5B3NPbkJU6u2w35zJl19511UkzTr6AKNFvkWnzZQaA8juBRtjCehhpDgUpDbDLgTvLA5VzI+HwzFeoDqqc88gzSKcYK7jPWgyK+Hp6bS0ECS/04A3NP2vcM/hPb4lxBkXkRKjTOXdb3pNJ5wUNNX9jXpQU+xDz2F9pdVqdKck8sZ0dsh1pqq082VxAjXLh4LFFG+mwfZbjMROfevmC+PQMVRZacl+OcGs61/6oU9ngFfijCnRvWAvHDZ+n5VN2SlWxpzww7TUM6TSBF4tlwwEdQggKqcQLGtwtMM7bDCFjQ4Tq7cwZtuJnQiae0UFn2ltmjfmA5LQl9y67kcoTqzjZslgtJWcESyt5/3s8SSnOpUGJAPhpc8eUD7RvVpxmlNB5Bwo+aBCfcI54VKNL26PRz0Aj1Dv/2ndcIsHJ4BuX1WShOwR5yvueV0E0eliZSqFzUNYJHHnv/9TVQZa0R2jf1Xlo1lMZur5+trsw3KBVtlhL1FiG/uCjbUqu6s5elFlMShvbe+y6AxeN2ZeEsjiH1gHJyFFmgh2Zdldvnu/hwZE8NgDbE6jeKROwH8Ffq5sfG2UlVpnFsxN1nRVF1nWFF1OY/PL5fX3ap2ka10nA1CSDUM3Z0PD1hFVc6/4sI5EOr5jRH0NNL5DwlCV47LQRNBk6QQ8VhC7CB9fhgbkDn0uttZnlF/4AqosiACWfp95bLwN/EAqaf/A80OBIOjYk+pkyp84eiKI1pFtOWwuw3aQa00nlWSZ/kfha/whSBQqUMhmB0pwdoXmMDg1oLbTbDLRsRO3IBmkdizl111t2Zpjp7HQSJXEBB1OqrDBLqdVYyfDfAPZ4Ab0CbZZ4SICnLZvvoFvN5GQyvEfhW5DRQYFadT+Ib4bco+jO9KfsgJRrH7a2oxN6xf5Aqv2hnc+BX6XKgJGg8izC0X9H7RIiufconoDl7jERu9LCWugGX7xVqBxHQsWzrkpWQSGeuejXcZIJftAVvYyYuqvMcFYcqLALW0Rkw7L9wzKax2iJZKZKm5IUIII79mzEabhSAvM4LMOs9ACMuXDZ/ReFs168vHu54C2/+gVV7iR7nX3/gVk8FId4V1G20fqiLgHJJi+CgxyGbQbp5OoPZ7aU3ZWJnug6eHagSO+6Wde5ZbbbEYliB9wkac8jGHpjqeNJ7WyOZgNtHy2pqpvXfXUq4HcSmJ9bM61/yo1b+hZXX9O35ae/Frx9B5gsd16wTgW/gXcu1LNXV1BtIusb6IVCIj81U1rKnFb4wAUZO0Ns6o6t1G+unJWhknv+iNTHj6+bXnD3393Q4fhgSbBoBYihSutkIdtOdkOSW9lW44LEQ3L/OnMKJ4aUDFK3TbZVKHxDvhe++V9fZwJT8BDQjxcR41bMNg6tIxZ+jALaJ2lVi0QN3ubYkEdJW7C5q156M0Nd38px5mVNrCK/FCkT4Leu+UI8CnmF2lrbg+vONgo+OvkojO6mTLRvpnzN/xW6UtDM7AnqW9VgLwYgtImUvdcIkVtzQicmi3V9aRvc7QSIoG2W3bjFZ4gB1tn/DOXexXNsG/ETA1j5TjkHc2YT+XBYTwq/2btvoHITyfgi/f8arzlg5XAnJOtsY0SFiWQcmFmUL0yAr/DOwCsDZWwI3lTUXN4FNIWlxOatGXKG8VeI5fJL5Jcly9epqah/x/V/fIlyFgM0i2GJA5c3bZjo5ARTskn8b95i128Sg5tOhXjqCu1VNfwK8+jRlOm5WLn3CfYfJ1BVfCHajJA6T2ubM/7HCgghtkJeMs9nFqDJlEVVFTu4RVOkQN6HMDwHwTF2X8r+i54bEOAlVU6iAoS3qgLNbXu/n8HSkclsrZusP6lYgLhgWtrmgE7xEUsFmBW+EtiZIYT7gO0PAgSrWg3bu3OrxSTiBiwX1mk28yL0+bAlFPbYpUs74VCRD+CLfEdSlzCWI56VVtY/BD7ljtYqqMFPRnE2biI/K7nbijoa6DUgfyMzaBUx95B44Js7+VfZJusLMpm8DHY//F6BFJPYzUfFcRpamqd/VpjLvOlHAMtjy026cu/ay/MuwewgYwRpeKyYwI/qEf2UjyEliLM/IApSd+zBCRapvq5pJnebMYh2wjdBXTks0fNQ+PluQFdKBoOE0USYWhYuaST4cmg+lJe8kqDK9sTFK0jGlUgEbJhAwfZ/gLOKce3k0T26UgRS0zc67X+r6UPq2kd77a5xTivSW/5l2n4MGl048jpzitF557W0lUJtsSZz3aE3jpY4fwWSrDnGzcU9W1esiKbymEW4RTtj6Py6JuUDWYBycXZ/VltDft8PvOnU21XUeEtt74LdZ2idcJVIs7RlxwgmfHB7vaKqnxnNHbnvKW/ojUiXjy/2dMLB2/QbF6KR4Gp5R0rhwaT2UYJIdNEdQh1Fovw9g+0bGm67qzHM26S8odeUFDztMl0HoxPM2Fw/EfsQIPm5NmbTy0J4YBCdmXLHk6S4sHc21wdVV9UWdcnsL01lxrHVvp89XiROyxeZjWHZrfEPiP6nnAHHPd7B5B9hdScs4aOv1lm+FHgMaLMAVIT7h5u2Y1mtk3qbP5tfXyFY5vjzTQ8yuDnOOl1+UiyQTSE3skMS0UqO6FTFsm9goJZNgSHnCI8CEunoBC51BmWVgf1OrufmVCsTakN3rLWEul3T8zli+FKaUvGkGSuTPgGo48qpiPIQ9cofUUewldfmHK/uaiN+/Z1R2IMo4rM+7mFMrfjMjguuLWD+kOk3N1xwUpS6kxc2Tjmn6rJe//TcrYZ2iBvjdGrPX4r6EojDrKXIjst6bVRPEFYfEtdMg65PnYy11oVJbIVSP1tOsRoYgOgV5F4aOGrJ+6SEw2XSiHNs4vXDpfpjc2xG5IeAthJGwrKhGmwxYQAfIG/vA0YFVTGK3Q2bNkjPIJ2Jd6Dg0KxGJkubpWGxfspACVh/UYjmQGyMG1ka9V64Cr7cClGbxtR76Mtq6URknEVqpRy6f3/WRKrOqZVOzbBGSuBbGH9YqMVSraKWNPT68LQET5y9ONzYr68nus9IjVI1mMuCan+A7WY46iyQ3A1encl39p8ND0t0C/nMJcm5qXRk6VDr1gaE89h8L31OyGAAHIO8j07qK5e8BaXM/ZEnBVfE7//xLzNpHiRAvXKdqGmymP4t3SusWVxaFeL8nGGLpmnF+xRuAvjRWPLg2lZgEmf7DpVzzEMppBnDyPnQRNeNApVC3gZjkgXeh92jREb++ZeOe6XPeACw8AAWO2ieDpbq7Ec9JpLNpMWfU9Zc9f6u03YMzSdwc5Elw26vDyD5pD9PRtP0Sq0DzYh/Qcr359hGAGjAlsCDBEE3VJ3Soausqcat/mqtvBzIkkvlaTExT6t5XS0Sy/RL3X4a+XM01amFPVzWl39lPtyyAgjftIJabvznzJijGm7LlutwfABmqQy/lcGoS/an0d01kkO4RcGxRDn5Bm0qTDocw9qCpYvMp16DK5snFlxs4fM372qdN/qAi0MRs2x+uETCfxhCh/nJrDZwMc3OnbQxVghY9MXJLpC5zHmfLz49VqzCWaK9eN894VYWtIpdlDDzEf2wDj+t3/lkzyPVgI/QlVBZhufVPG/WfLRngxD+nlRaWrr0AiQHS28Jtuwv+srxTDY4mRV2JzzTyCyTLyE2C2NAK20M4rLgZE7hzpdq3aF5GDLOQ2OnqOmy5gnJfqsz0hr8XRzw9zYjTNcSqYHqp0k5Gt+7K6nRDFo6pod2vQVkiB3HPu3kQrDMUEHkL/8PoCo00/t7lGXmHoR4ucByBpY0+ON2I4EsNSKyOBG6ciCVnOs9G1dQIHqSq23iZ7kboEGVFjyLZCkZ8BuJxrPXkrQZrk0S00ZYswAs86ftELkMb0IrFHgnwnabSjsUoSdT5Q54qZrrI2hwSbIzQf74rsJh/3X9YfdeZ2J/CFiT1gUArcDttsO6TKhH3VtjzsZlboVkU67/sakRtalZpknueHakh3YoWKr9mh/DEPcgbKiLf4GMCJPC655kYfQUkUDS/pQFXHDOcfC6cwHAi5cRsdgcD9jQCa/466FfiqMrSfNKOFU4UTlmoQR1kqQbs0hn1aaQyOVScXnoZtJwDF0E05I0Eqnvn5uN8nIveIcpFAzK4eI1LvgRz1AKN58zTWtND0M4dP6qb6vbmfhUwDyYkIZynMCM0FzcCYvQ1JLy/5wq6acYJSpeK9pFVX/K6Lm8YqbUnUKgFmQfaF0iBd4BusuhIqPtYWDq+hQFTLVJxiv/JRi9RwFb1YhHPhWpXTHhhXbXFOZFYsZtcgs5yboHPlDPekB93++aWL9ijEtcyncHq6/JpeyRCC3zvguQfqGaTzyI6Umy2PElPeKy4/ZyuVN7u0ZnViNeb9dkH174sq853AXvPLXg090u5Rnlnc9EiaRqARmGyQ67XCLbwGeOCRdY41FrByHbIrDd4U8Ou1cLHdqcHSwVa6PFm6sXjU4MHlCNQFsMAdkl4ynrs3D4nNj8U0jZbDjYG2GLYqGkH+mBJRoNL1s9Lr9dei/ek1woI3RLfvBaQsmyFz0QKcuyQIyObdyQ8EqCIBMug0x+A+TbyDygdtvQSUccACmzd/M9BnljzZiPFoZvaJedeOYQ32AOSIjh0C86xmHkMyeLj9Iu6xXNJTlVF4vQLfts6Lm2ExAK4Nh4Z6Kn2PsC1Fd34l7JMhDYTfSYg790r5jHnu1scrUUUPT7AQaWBbqVQbjYrwJyuWk7vFs0GEj7a8/V9lVu2nNK/Nkxi9+MOK6eKOZvi2EW+ozi3FKhKZ9jRAKxvzzumzvc/+68oMOEzZFpet6pW8Ln2SO4B8AtOQP9HDu1ZINuRW6bv42DZ3u8uwP4xsL5q2/Izq2YL9J+r5nNkRJ/WlCJZxik7h9kjxdmsrq/rMh1tgc/6grsh9gYGOECDS4QPjm8YRRqQdLtGcDrvCCN1O2EbvIQd2QMZBl790UIybgwQ/+2nudCmeO2HVA7bEf6KPN41LjdXGE4sOOnHL6jRT8YlmKaVMBewueTbVP0We0jRvvjHYFUN189D/U06P9o9JCr68+UP9SEQPnvMi0b6VoeKrqr4qcJbkNs9py/wHvUxJ0C3NDqCbPmYtthqvEPqn+dFqfxiCPlnlqy3T4A0avurIWAapI+BpCwt+NkCysgRufWkLfIcRhYJ7V/UlSJO3rtohvhV7oGVDYL29XYXSgDoNkIRg8UWiY9Du+nLeVMUlq3ztZ7Nf/gJaI4QE2bxfqo3afyk7nebBUX4d2dPWg4jX7RB17VN9SQWpWNfx+7IhiDcKilQy0tjSPSCTyl4PMzWVRRrAmhV+UFzJ/3nTTPkmhIb/5gzscItUYHzqio5cvSbY265UmACr0qy9xj+kbgOCSXHUNWsW3Mnpv4cMnTBl6/OAOJrSOe6k7jstM/pPT+InQv6E38SfOCr8F74dajVmawO+3tI4nD5s8NI65BKlyFYfit9Uy8Qqh3na2hgTUkoCMedxLOjI1gr8ycGeTtXX54KD2dcDR2DeKMOkfkt9mGueki8QEDjfWDT+147Nur/IBjVp+Pibfkd1c47ynytUFPkYVjkleMIv/0RKI8D2eekf7wzmYaRjYu0CL0F6aK+oZZDmVQ2Lk196EA7qAtM5EDuXrmVEEwHH3ilV8sERTVy0h5EKFtj2p9glSzy/uws/JmFj0sxUNhVplRvzFKjr7TdXpANXBUtgXK3dL715Qx0ObNHBgndfAHpyaVDVrS8348A4wND4rLhL83ALYv+/AYOM/SuiSjru+niwMNqcvlkIy+Vzh16vbw0DMl+UHF7GhbymKb40wgDmMmx+uFvE3SC1p5IIatkoQpk7djroJWULPE3wtM/ECh0q0yqUbDyBW4H7opDiWYGzlH2wRZkAWT0e4a1VW5zXvMCEfVnLPxxgmkQ9/JQm1XITIWuabQpaP8wLJecMTjOSes9yB9Mv4FdRi6CwhXTjtbLjgyXiap5t42/ClzooEDjqcMPTemf4LgVaPDJ/fziHjYkZu+PsCLBKxewYAFec92q002zHEydqJ09Iq9oYK/ymm+KF86GITPZeQs8FAZKrk=
`pragma protect end_data_block
`pragma protect digest_block
73a65f2d0b4ac122ff6329d617ce0d82931df82f1519522cc7ee3dd444b2cc76
`pragma protect end_digest_block
`pragma protect end_protected
