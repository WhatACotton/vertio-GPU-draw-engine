`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
kWzkU/tKoS3R+b5bkRiIL+yWC0kF47COfrZHO/rBU3qv/h3rsbb2yzXAIUAiXzEj7uLXyhTFTHt6z89sDdV1+B2lBXcObyKq5m3Mg10xuYya0MuWwfdvsam+yjynXq4a8KUIS1IZZeTJme7qaNVldVZTIi61bvo87J/AQ5t4KwF1KEJA/C0q/wfiSaH4GJkwll2tyD6LyFsaumcmOXVAT18z1H1BFW8A7bhH3XpoMhP3hC2Hvf6ik34TFgC0Z4BapcdDfp+cPohEiSq+c2ogQ2PvdZaDLDqIFjSMXF+JhLqkvT2u8NwxPx8Bl34tTuA+XkN+Xg1B/3/mTakaLI3CCklkXY3WDGGdpv+QzfO4PWtDWhDe3A7BkoGRF6TAgA6l0l9nfD9qNb4tc6sPq/7U17ZD1tBbvTQinfIyWHGA1mUlHbKky76ntol4hPXxK4TW5tr33YYxWZPLZJD/guLAcJ40qzXjskY8/vUIjpAu1p+r5vA538Nzm+hmrlSemRTF5h2ot3iFaW3yJ9jqERPDuEhuaB2ddo/k1AKBW7Uujz0+7m3zmIEa/pvpcul3a46tVtSwFidsLVUIsPseB07pOg4An0Lnk7DMe9SAwdv9mR7ix3KMpcLWAQ9hZ5k63FXCt7kS8JObemglFtXqFaND6dXqTaovGhBZv1T1YLYG+BaX8zAhAc9sFZlNEHyQJ6LsGpmflO3kHN6aojSwiBWC99rcrISLfQBQFSVqh3PAlvzdp0uOR/UAKtgwI4Oo380eqPe6yND1GoFfDh8DOf+ZI4PL7XqeGwyfM27mfKNvfEwRJ7LVUBJfmsZel1SIFlpS0Xn8n6tXC05DJvh/3PmkYwaog2nI1TtZYKMFMYt+vz85q7NcZIek2+qegIZ7Y4rjpuDm01pakDBj2mwsGcDIgrABTmv6AIAIsanjmdLeFQNveS00V45hsKGJxB9ACn0Fhbxe5QqoGah2TeRWgCSpwEz+xdTge7XrmidnZC+nlW7UsaE4pq3YgZJmxScuu+3YGthp3Vgt6FVdnJlQYkIwxlHEmaI/qeGi5pWwmSSZ3J33oXKANYqtySuCeEfcZ5xvSgkHx86lnnPSPSAYpGEJSsZnTi4FcqvDupxVljlE/JnFda7a4qI+2wHBruO02OQLkzJiopQHP/8uzuBxZfH2aPdpN65cOIICAsRE82hFXVnD10SdQCW1F/YyzM1zTQudbDg6CZK8upRnwtl8tAJ1SApzemwz7JXK04RItAdb6ibHPBcKZP9V0AW7rcMXwg8jHHWTdJLzEsVsB1HUwseh7vnh8ruadxuc2flDHJnNr7qohgXNlzXM5N8KboO32HCWRYmE9O4HQlp5Rn2XdRTVEKsYvKQzDJYnCUoeitPj+UBnyV9gyfI5RCAVbPcj7mhm9nHEQST9cYSEnFGcw4hcxiOnb2WDFW4QeiLx+2g08F95pMWpX46Msts8wNB+P+HF9dcgMrnYiO9tam3BlGFNko5cXYvpXhPOZMV8gdyor0/cEN2jrUMXX/XnnXDz7Er48c+5QYQ/bhObbZitDc9bDNoUk5EB54ZJp2kNeyrXwkJCQmOVD792GWOQFdwaG6hlqwyOFX3T2Uw6e4SvgX1iyOqy4ByR9Z2X3oDW7zqLE/QXfoGhkN7PMn33X2aIDCIldX576jU5fWjsh2ujJosglU32LMGOn661Xzqx6CG9KfgIYYwE1GIMYzJVLDLxmSIGthddkELepmq1qYMRpOaGNwbo4oH48mpUlj/QkHf0DnjxXZJLCT0kFhLdp2JLkuJQbxa5EqbFwWoJuMFOR3/dCuD423b37BGZZFSaA6k/afX+Myvy21YrDuCj+dVwMVOyEScu0y5KbVdzV8gOVQrRNaDYOzhubtk2byKi6CnBx1sFpWd2vIQbmOTOmQ27DXwGCovxHK6CsGctbIVr7XTvP6bs+jktXKvcrq8p5Mu+VBM59OysTjPSUh/l77zEw0iap9vHjX3FE5piBGGducsCFYHGvz8KU6E7rCaJM1qEXn5qkS++RScRpjgyq6oc8T2rGg6E3VbpIPtxWJ5Hd3ytgqW+sB9En2sCa17q+AqigYd+S0dnFzpGClxVn23bm+iPAkeLjeH1moV+b4ohIRNKFUDeYiQ23VR51C8g3vBh5FZoEb0sLmClNkSOSx4BVC1EaK2zqQDxNLqoXkamMWBthTX0By1FIO5WdACdxRM3WSCFhc0pZ6Iw3SWGCUQVQb1fJbH0egOC7LbP7ukyjw9AmXZ/u1LWPkMK6rzdfYPwWtIbrjVs55+xZQXKCOE7h0IWPXyNal/yXO0pEU3jii37BZ4f/sMPD87lght1fPpmIQkctaR2X7+HDTaIrySFrKPCY2DUqd/9VYuZA6Dc+K04xr/v3/WeMfV54oiGdhhGuKMk/oGGsrrEUAVEi2VAhsBTKWbDj+EhAPlVupJRv00FIBAftiOdu7hVdpkZrtSkD2SZ1DVtLxtYDNT/1XoqO/3sy/B5d66NAcnIaogdkwsUNA9IkmP7HpRxKTS29mFZToMlSOT5VZhj7T/D70FeiBo5re6XCx0qocewSOsF+Kn7+SQpEjUNxwJ1PpN4Vl6fNuorLLKBhkg4GfNPICz96kSR7P8cUgRXzIzTRch0taLKwNo8jqTTf021l2Hrn8ywJYUKYFiI5DyKoeC+tUW5P0ySKRs91s2ZJLIqO2bJBoLSDhXVZTdT9WOOIUmiyoyitHGFDkxpIQwFdvoqcaTjpBBPhLh4iXoCrfVQkZhVsdbYtyiKL7cmoHJzuCuYLbFJ42stE1liMWDqwvcCRVbxmCWXr4e9MKmGoCMayYFsf2M4kv4w6ho1rNXEiIO/FYilmBymu3YGkh3ZBbVVeYlRg6GwwdT6yD+Ani0hGzmcI6ylt3IZ7501VDTqmI0KgHBJC1vp2Z9rcDUNCcKdXLpPsD+g5EaT8UtEKKhBpj1g/L3tlg5CKrVJCYZ3tvJgJtAUC3sTSylsACFYeRKRm1jmx8myywwDaGVbCBeeLKMnCuvK5VMQUuiZGSYBUORc25xD5sfwLbrLYZMke8eROLCJyxccnpxS8Ih/Pb+i8bqTuM8O9yiYXauYXYHZYldEzQbpCeHo7iqaTdn7mhFP53HKxGNNkmmnsHmci8av+6NEzOfQd0AGfKCsA/2ay8v2lG0O4DvCzNf8yogDGgJNMTWn53GphOiWCVbit6W4C7d2ssdC+ZLPxjnQ2DmHv3o11MwgGnU88s/5nOEV40+S4WaRQECvENKA1Uq9lTYMYTxlHhaap8YuPMrySa0U6/1hXdNYz26FMBHE1XHL5vgx1i+Q3bSYZxaxppuq54vS17as1a8P5S8cLagxWe0ODOcbFV3+7QJQZcjXlwOxb3HAjmYaIOuwqORjNun+8IaW/v3a0u2mbIUdJywD/tZ3p7TdsakmTpWdt9hiBHjxs65TSPN91r3TCbSclHZmLvxJrSsIyHMbLQ3ToCuWeAJhAg0L7EuLQPDB10vwfM43VyAwe9WXDfYmIfc+bZR5b9rFFrKVf8xT/K88TVqXubEXFeRD9bKdJm3YFOtGQQOovOm4MYZv/Nh0poFpbkTASqAgjrVfnSi1i5U0AAWHtsgRkJ5e/EcKD1Dacx/53C3jPQhOPOep+88ylnAyUqqIgH0aAKrfpTN8uPoQZBpEy5VWwoj3LyRgV/9JPnsiFtcfBeojiClx/2mTr4NuFD53uxVFg7rsu3ON72l6fqkX7xqtV6883p4gDhsIVSveEJ+nUA9kUPO1YXynI2cyhdneQtMz9e4hvp0KMNCyRa9JszGSoRjTXp9IAL3BpPFet6Z58Q2jc+h9eZW9HV0D/AKSc7sOuGH4fOJiQZMVt42fQ9/eloL7ZdiyiD77aY3jCrXU5IBzo9/lriq5+V/bYYZVMST7Yik61dc1v2XNUYHusvdKxzelmAMJthyj3OH9uV7TSKFzWb4PGNWnU0ZwIvNuv00UhxYQfETuZOJfhD/B6KSz2LVFtHxWowLTK2ZqbDFb0wvjzG/fQ0+4M1Z4/dooNDdmIvqhfhVRXLvmgcARoq+4MS4bb2cLonQRL/KsNy0Q69gZddKzMy857Urp6EzkCF7XXe8yAZUVsy8Ddr+FKmt2gIZRO5tfIScCqVQa5DASuJlwnAX0DlC9N93ahW6cfYBwTqiCc0U7LS9w418N/Bpsb5bsvMcO8ALpASlYXZP1tG6uTm1kSKZxkg2Nron/LqSmgbSg7enp4psLGidxmtiDt91tj0AuzHL98WdM+5PuoKMPkfiQCUyeo6FPmiRuZVVT/JiY+KU+61MxCF9FZQyqfjsq6+vAUdIf4WfJ4JTpwD+PdjbscEclMJPTZJQVTRRtsDvRK2aNn2o7nDBBM+Wa7X57ejltK2HWABRipbizOwY3n6Px0N+qbKQeNrrkf7rM3AncYFHvQWV7Kzex7Zf7AcwNVtW3JFIIw/edbKm9QZjyM161N0pKILKWphrbHHureKkhCItnGyNypqQu6+S+OlUkRK79Fo6XpnT/1CIrPJ9hppwWK1dzhFqp2ImGatiHZ8nme5in3Fx2EKla9HQvjPCGWPv5Rb4BRdu3qGfBygPQWXJKP1W2aUqUiXM9veBlqPLRzJGe8QzqdK3+1nurqiJDmjAXq5Qfs2dGdknuqd9icKIf1+59QcS0AQdBLa1q7o37x6B1GTSsfAed5XWi4+XJZ2Q5ck91IH9axckrygz99zi6tsUmiFODgGcvhUFcGWxWv+bxvjN86wkDyz0Uc1VnA39E5WMhZ1HrenvGLqafGGc8Nh6ZdIGPypxxNsMADhaKP0QEq9/0hqukpywewEUhRFPA2Bkh2AaXXfRJZSvNnpH/H7WpSxk0RCI66T1M23NMr5RdEHYT9jTK7XV3WNkZW82xPvPXQLYNOrwNAK88j2fCCdFfoeF1qOt4vKUUDZbsHfSckVEtHkfi2ViPUAJa8Z6cn0qT6+sAulaKzpM8v8ez4BIjMEKchCgDSDHPSZPNuxkz3yuIueC3mz1peKrEFuR/2sMUQwEkJ6KAJFIF+miSMwiuyxF1PzMXzI1EKyquklXT+V7b9BGVuvKe+eVgUe7aonxgdwxOVGEgyM0KrqDlsewYkYiwxSXsRD4i2i0kniT0VnKVQyj49ISiSRxcQXWndT0ei3WoxFKDoYg8jgIG43VPcRHxebGI2wpw2l6UNvNhy/WFnn+RYaB3/4//7jJZQ13acVSGOcwfaz6nX8YZN7CNjZdFPCOPGIYTujyw7FEwDyOIO2uv1vctbOKZh0jtqYuGkgbHr6jXKz3q42bygqp/1eyukpxhONMlNprCXEix/JcHu4wScaqNO3QxtiwrEG9K1o5Zzw7BgJd2FMQX6an0+Zeup1i3CwiP0r54YVRdrm0C6/SWilhPBLB/iySTx913PGqiEIfw5Wzw5JVpQ01+KJxtbC7rToxAF6eiw7/5YBykLqBVMRRcFvPnQ7SY40pOMa57RoQD9tOfu91sJk5V6vut7nanFmr4RxcqSY064QS7jZVh78iYh0KvgYUUuvIr8WmAZzZXF1T8/PQteuOBs0DVnN0Mk2qeyEwvNBu8J4B7txtxTpyXrhUwjopTjVuakkfWye70ht4FeII3DacmaJ5K3UDjX4ShhMnGabFaBcgahhYGFI+paozAi8GrX2fvfl82P0zXayQwvLUrdIR1QI1vj1zEWIED3d4S1/E9lv1bO5GNQtxXLRmDrV94gQ0Pgj6OhGZ5t/y5kTr6n6YUIXp0xVJuVAxoTMVzgjKXuQa17Cjqk2qg+EBT0rLN1luIZvsnLJqccoz4minHTYR1EzzJBdZZkjn4k1jAWkHokjxc175PoBnUW4KysH5qcsJ7x0mpzeGgfnluRlVXGaXs+vGz+16SXWnQViZmX+yoZbMj3Voc5zOmLffOxV5lIc0Ksrt86tX/+Gd5jjSb3ib91/CJoTbuZ4fm92n+o8sdY63IZNKn0yZtVXqTxG/07siP85zBtYd9wA0nBiMGsQsEVKC740SxQG1mUEtjInOfof5icJ/XeiC4KCj3O2KSM2m6eEBdhUfFQIUpqQX2ki5jbYkrpgInLMMYwnSEaaBVqVlmCQbjgJLrU1pF9ZFAYTLV3Ts3dFInJrQGnlCGti0lkFNxScCsnOKjr4XVD1EJWWYQWlxzPYzNrP7kJ07A/jFzekZKMmU+iEwoAEPPdE9QFuD+vbKF1o3uTv9s219V8DQbquOwD3tKYmThlNsF9bk8NxJKwdRjf/bew5Mmbp217gX6PPvgpWva7rp5N0p2fz1HR/kk6UUhbFrpDXw60Z7rVZ7MOwzzhK6+ejPBtr7olwHkUYHBY44QTdqKXr2EbvIaKBJH2vtczduLVGw1l8MtYQHkr2KTjMVa7F0v/PwSlgzq41631ULxXBhrgfX+RrzRrKGO6qsBW3WbAXTokQYRDE5AXt+NKKSugrpNPmDf2N3BUS1i44wTSGpNZxmQ92Nqs/1j0oSF53YL19TbeVwITzhacupA1/8rb2DG4721/jfK+ij+bATeANQeUp1aa2rDJ9mLW1qceK2HlEdshGyYzRKsN2n89sqOAqgG6fxKe5s86mP5R9bPk755LBvHRzGEUGClZxuQlN0WLad0FJv8iYzL305bynSCrCPSZ9MiyyWGoZZE/ApXaKm7SDXw63ogCOZsVi6W+elEVP5xV29tVUV8dEiX0Hc9NZXVk3O6PvvycBieigRdJlWi1k5qZqozZTsr2XGZ5xHH3CsW4+ZfDd7gwTfCrueJwJqwjSzn49C1Qc1lFjqCyfHw0iHsXMFjQzgAtyhLuaii0tzVV2gIzfER2YhZ1J2kSbgROkjeHwiRD3lr+o67mz7IS1Kcp9FNcrz5odMORuiFXABhA1FvpTLzu/IGN1l1Xdnrqgt+zOff22nDWNTTNSaxJzHZ2cEVsLLQO6lsoqg+qBHBLf6yn0nS9OMrf3gNPXKcTM57ujbe5EEkkQJZWZNSRTElS/V4MtlKl0YDL33D/EcnAH4lMSLRSrrcMWQzeyU4VnoVscY73HH84APDZy8ZZ4iiWcPTtMFvZwpSDdzW+zNVaCxzvZ8ZuW2NEsFzVFNmFIhK0JX2zX9HIJsJce2lSMm7tCbXVctTTzBM/BJWFnDP6IWdpHRQMGeTxcqjN++NdprGDedcnZjGSAoGi9sj26A6e6pVmFaxQDFa2W9qo4FacKxNbKzJEevIqqNMnlPMIuiba8O9GBkRVylE0Dep3lNAKI+AZm0uLZtk8MZjVYf1zoJhYuyKs8m8yiJSYcpQkCFiEqOj3ukF5a4FfA1M1IdIJk6lbJaFQPP2K99JIvzM+TqKU+oTaEcKINwLs5SqVoqnu2eP2QRZ+955jzHM5Vsq/mXBrJ56e8VJ2O5iZ2A7GfELnq1/izpXt97HnhYRvPIkenbyBjm8e7uvklxf/9TQ24X92IdvKKgHEkzBSTu/LV14CRJhHaX5alrr/rOr3bOoejR6eOIOa7iJtdSkcHXxAPFk1Fx0zSoRj0D6VugymF7UMEtVHjRQg0U1CUwralW9us3wEQcfCa/Vq9k4XX6Kre50limakiM8Xd/lFqhvTGqwvzSfdb+VtUbASId9cA2qFKazHl1MPC8SLD5s5s3/wnGXQnDZABdenkOeFUMKQnvH40nYm+VooWl3fakkUDNhhd8CobiTel4wLPCi3RN5Ps78+fcSMF7D9nxXXSOI0Wu6Jhh4WpBsHWg31Ly1zXSMH4kJhuvZGEJCKLJacZndCmlg4tjw4IAL4VHeX20p+5nMsSY0YgQNxRENqWkNYgWWRwkquCoADbeQMz+4veIll681vHFmngengFgTgr2B6tkuFIq8SyZsFR/59pNDvZ/x4TRDDft4wXuQVUoi3y0PAxz1Dpi7m/R4daPz7c32b8bWwiRlnZKlC/b8rsxxrNEC+U2qQLsejxj6b3vO+zAEaEWL87LqDcQxnEnSgsYp3LV2CSrG8MDsDl8dfuaT7EC71+nSRG52yg/qBkNx3/94dJlKNQAWUW0eVY/uHCO2rwQOEqpbpXAGXEn8R5f3RBi0ivdxth7TV0FhKvqJNTrHN8EZCx9nZGXCOme9umDNisus/DqwP6BzjSR/w2sHz7tqjlLIUHjM0gTMtNw6Q8LDIjuEmWlOSYF/qfFW9Osr6GK7ZQHajS1efENOIPHf1O1VmLcLwnctav823jsBXhqDsWC+UbWCSn70p6s/n2v62V1xRvikAks9gZaBzUVNVuhmTwyFBEeT8wxgaOgM8lTFH5PDkePAPj6I88t7oE+qsnzu90I0/GAjyYSyRgw1u4aDk1+LYbsvXTR8gw9MBTqzDnDJ8/qf/1xQ7hwsnLUwEJldkD4qAy3mq6q2M0KSh14AJnVY+WWJTuRfajCer6bQltcx5QgOQBc8mJ5l2fXFRLODX6tNbCDYBX2hJB5S110s+9cqktLnV7ZI55J3T6K1RbiqmJqCjM2+w5XvGqwVLSt2+pL8TRq92yeV7G+UnOlEmuaC5IY3WemnILrNwpAyKe+IEp7w4NS8c9xK2zR/crkCONufIUM+D9I2WelcWoGv2JOaT2ltk/TUAiIuewF1Jl95HYJVoUCVxiMUINltxRCQBU+lqswwY8330U5JKHnH1saMqgmTckZ5ATnNmbVDItFwWm3XEIQyZD5bCL/fLMHEErJRaN998RsKonQDUiK78nmm77pdrUtzZ5rryiN44b3+9uMPCLekImPWyjsMXomNiS+g7Trfw/EI1N85Bfv9cyi3XXhSoVFce0W/+sxrzwXMdJ75tVYDlcJi5LJSvgFTgt+ifTfgR8yX0K8bpuVhTTqiLnt0c5TddDxDKhMlWKW2xKCtfd7Qq0bRswwXDpJ4Y4jQmdnNFoBf+03s4Vk908GNNfEtdcelTIig6rCof3VqC6P7UYu+/pIiVS7fsCCMu7EctYKfuxucSE/jUgmiiifPjVwjJGlxS4w+eKNkuu91mmBDzWPWMz0mlSWdIKXkbLLr4yoEICGd9JGsiDr+At4UjV0CUell32cj2pcTnzBiWznhrtBVgPIGoKTTpxSlLG9IfSgNhhvgib5uTAf9mji0QjxiTxjD/zRsdJBVqthDjBGeCw5WuPtynYpQywd1pZuUQBuWQsWxmKgM2c/KrdGR/7i2PCip1DxfxEVj6nBOA+l46KA0PaWLdEbmyETViLIPtJ/mFYfIPyfbsFOs+rfAQIlIWFTSfCs4z38Kpc47uP6CAfd2hlvu9K3aEZdGk/tM0+1MGfei1JmVZN1e0Q8cxf6Ot06O7tZIzvC9m+OckhAc+/XV7v4coTLCNUMUmcUQJlogkJKl/4TO0AI2F7UXZnr3GkJLGzPf+MeG9BtW0SKxKBAcQzh1pnKHFbHMbT56u9fpfQ9Fcq7JSFScNPchzlms+g6+kBzv9xsBgV+jkH4pQNuqMhQZVABL0mf9YlbEM5sPf82THcV2vrJ57xPk7XT7MH8YYKjxfAxQQuBC66nvN4n/sjr/o8NC1LCIBudivWClMRVMst8gt5Y6Ck18tv+qflGt94RuVmVwdBsnURYOPSYj+ShSQqGDYDJko2NWXNVaL+9L/CEezdOCWzyI0lTU19+l0HRBI0Z1OgcWXoo+y9P8302kcSckb+0iH5Dkenq5dodvZna8O3neXdXIg+Y11FQ4mj9FFtdqZwo1RwvLcSbNhh9Sl0qN1QMp8NcSvvUfWG8UUhHRVTtkNf4ySHfXcn8t1i1BHHFHfvPD7o6inJMEtrrOPxwzs8csmkWZlXd3fySiq2PVhrIeSUrZKl3N88RSEbRHla+ZNjqQvYcwgaDkNxHlbh2ypkYsEusiOCQ71isSoyTPS67oNRPGrWJhMR6hrJZG2S5E6c+M6nGtlknWrmePv3YrQmEa7qzizd8JtrLlVYZeuDwxZfmMcIwpsinapq8RdNFvnSeGEbU65VjtYpgd0phs53ULQ7LZ/M/wzsx6asc9J/qvaVWzT17avtBnLHu1E/cmy+PtJnfEDZ2NXRUSRb34uwTT+KpEs/+jrKI/BIQ8xNuA4sdXY1mA39jYXRQFGsUG9fNbTc+Lqhy+Vim8ZwX2EpJnDuqTKmtYJwbFBiQwSkY4TTlZbcM2FZU80pN7mxZ2nivz4TYLe79d/MCFwUVWp1TvWQyhnHj5FuG2r1ZbFaHZRc/x1D1P0ySmMc+1tQKGtoueXstjAsYossYPEC9ZPQt3v009tKG2rPilibOiaCFhuqgHNd/OiATvfpRaRp5q4LZ8IE4mP9xJjwprst+i5u5KySPFdm6SJZ4Q6l5dTfZT97MFDjJIlHEUFxhgMimpze6JWBllroaEzTssyRbqVErShTDL9eW650WbOso9z102IKiX8nB5KoK1dE+Yh3olhGmQgj5uft1fFsMpdpK24XeX70KAUsehud/MYfwzUiy3lRuyFwlMn+IofynBZkP18v7dtoCs/WQvZxJ7UGWCJCIfCkh1GkBCoi4W1Zgl4qyg047edwLVolMysxZPDivR6QdRy8lPR7nZcghpOlwVPXbT8StOjNkSwmtMdEEt0zG8ytETRkGfJ2ps2HhwJfV9raXyPQmGiheI6wku0c1MiSfLWLUbAYzL1vht/DM7VFcjtqGmoTjx3ocDAc8cvsLfUdaswAuptljXVHo59NXou6hMK7uLqo50oyIFOqqwL/P116hDdO735TIjQXXFZ+MY7OZJInY6PLuttkQ8hd0W5sHiCoKTN57DMaVBOSnc/TR43lyXzkyLo4+aqSnBTkz5lyfwqIYm1ww4yuTa16Fhv+CjC5Nxr+yn6H7ZYmxzBekEldTNUUlsIKjLda+8qDz+YA7WRREXgk3vAk/mm468N5OOz6RWCrop2t8vcDywCq8p3n2uQvo8f/1N8C7Tw/Y/KkNLe4Hyc9WaFwsfgAjuBSgWZGRnHQgNtpdoPbiQoJRwwgG6CC6Y1MvGwFNMD1a9HJ5/Iqr5Q2ngBTfXTIQDkce6IHopIYwFAy81ofZfJiByi+rBloc1oadG036SzoEy55NA1IWUSjsD2wwbTpe8n/a79jMf2hGAxw7bjN/0BFu3xAg6BAGpsMbMylCol37yYrpFcid0r7ANlG0YT4JW85t8mT4V9QfsdzWT4lLh4DzayUwT6HC/0UDrTTSjerO1/g37iqRxHDR6riR0AuvySMv/2U0Crc9dDjJDMLV2w0sJc7h2CMU/FotHP/N3WCLhJvo83A7C9PmNmp6nwmEpFJeZmtgRO9zFsNf0X3QYLl68Bx1ypU/ttlWBdl05tc3+xfCKlFEF8LX+MiFtpC9lmcXP2dmn60DLaffZolTrMQf92JVL8ux3HfNqTgZaaJIWWqq4hKxasWMOxtUI6XVLulQTTqEGNmGmIWNnH4MyXOXSDobS8S4Y/vKfP1zdbWrgnjvjnlQHfzL72vIpp3EUyK5CBaPN9n7lvimhOePD1v8DSov2QoTU8L2Hu5hw+dS0uOXG8pjQDNQe4QltsSGZd1hqJSK7VhmWnBgbV2pvHQVi31Qmbb9UiP651aYho8pi6QSd72W2RVOkAPb6+XzMvcD0Ke9ro2voMKHb9f0eQKBjuvC43QAWGcYkN50K5XIfxXNBTJtl+u6gF8Pb/D7kBtuXHPiyBuSO1AKsEViUcu+SlHZSVYQSlJKdJEwZpb2Es/Io83Kl64N6daUfpYtkSM5ybpdcruQmh0lgIK1bZhs8YVS8tTi9iyo3dAqngcaGv/evz0zVy6yvrkXYfjOJhsVWcFbuuIKiScKoLhsxCD0EYLuUqPNQZtPZ3/a9x/r7/va+vx/cwVVQPcyGSb+0wR4CI5RwHJnbDul0fhYw5M24Q/cemG2yfGXXADnuh9h0Pm6Y1Fvg2noeLsJosYbqfE8+FD/kwpK0pJ7jOmedW1cv+F3blW9UxtL4Cw7Pi6ur2VJ6mIJ/FFiwTc+ydMP928fwzSpnaUQ8MnUoJA/id5Mxaw7WyqkQM1IHHCZWNaOVsfGuyLo5jNEx5J+gV6hzsx2g8E4HaI06cEfDvha55VT0g5Hpw8lVQRz4p7+Chsu+oIFwHyCaMHNJDiOSTxJcuzR216PQOYp32eplivpfX+/xkIj9wWCqd+J69xujelnTjYsRNbceiikbpEbyLsKTaZdSp40xQlqVsB/Z5gs5D6nlmhrZ45ohv6Y4MyMsXWhCRQNhSl6xnf6pmufHityvDoEl+HLVEngQk9yNvg3oeTeaAg6zZCugDsYbuYX0DgSd92myJOImclutrCKaDr2nkUIF3mkl4Vx7CAUdCBFS0/Hu/AeIfQHzOah9hE9JA9nY4Xwofgpkg4sYVlld+0C7EWiD3s/PkPYtvaj03l/1nmaG5RnHNkJ5dGRy7eAwq0MwZKuDDT5xEpNvulMB2fR9rkv0BKhVcbuQMMnf5rnCTB5hEtL+LGuglDmWmM8Ehh1czlYuoF8dMtfH3lD6W1a3ce9meQkyo5LS4UYzkzHS78TiiNuI5RMwdjunAbFT+rw4fyyZQkjJpn3ALTmYyQ8hce2PqzcWLyVVsSm5vSnq8ESEJNSKjRUA5nR80FxF1pU3AwGgLEdpNBSlo7FLTmrKdGMNVtZMcvkKsDNTnbwZPxBa3M5/WH3EP6J9w+AjnAmDUT/tgtaXoR6ahW6Jhl3LRafPn527qoUbEE33iIGxUQH2gS3HTSagMPz2xUXyOj2PkfiFQxkKcscOpQMUGQ7Fxr5hFKg1CHfRJBTvEG/vVZ2PZn7uOSUD6kyfodBZLbrnNcVuY3gnje6Ze8TWvP6rDwfFhoWuiDRgDAQ2QULB0zRPzflkiLLXxBsH0Jbn0qzbYgPbNjuQoZJ6WXU46jGlOTvdDUK83nFqAp2Do5IXvsBV30TrXA5Aej4J+eBbjRVe6NtcrBJngaqOw7kJ4Veje8PzW2e8FqobvPyMi8JCWw8FYbhtB/M9RI/BgQtVqYonK0+1BTFNw3556V3BC9ssNRGDcVZ68mk9OAqQpQlMGomtrJpUfl2OUntvghQV9oiQ/DSLZzjNScUI5IebhP3MfFsCa9UA0QaXbsQYwwKdmJ+Mz+1XbL7bj0Rb1hH94scNx13CbZxK5CRS3coMGaVo5hOypwb1DjNwuHGbqWdxSb9mjDXBpR11ccW4s9m+bdOvm0HaZfZdTE9rXPLTnv1HKg3fIvGPpCggnzFwPcs5RSE5PENDtnC/BOyTTicl0ueydzDG/jvGZHZ3MEHB4Svc3lkNBX41ZVSYTyepgABOEjDQ14CDzZ8NDiYXed5S9v4IHhHMQ0KVGeN6O2AuX0E9UYS4/CEI+xszTIN8HWnXdIrDD5OhOwvm7fXG4C1dVeIZLXFsVc/z/FEBtAJNsoN6fBmYge0VDgb8VpX71mLxcLO0shmsGe827/nGz+gZSqbyGcgNvm9W34jwCi9BYZKly40Koa4haD363b7Plr7esDtTqPnCIjlELcYQOrY8cnGNmdcpjfWNBvC3eC37vaeNUkb33BJlsZkWmzKfLVYTcBMM0t7SJ2o6x5zHt7+jva/r8EqT7OJKhfGysUcQpn68tEKyaxoWCxLdAG58HQuVp4lpl/XfmMMx1bTueAjvQ2ByuYH+47L4TgInywEu4CB6tXPxoupkiAIhc9ZpQ/mqiPAxSj/zjeYyO8ZhVnwklA3N7GjrThLncE9fk1ZH4CrtyxTVrPL/sTTWQs110pY5ztC6fEydKY41AzcmYZmuE92Pdwj3N/XxZX+7lVqZahVJGdz2PUpYkMlawtXSkdlAn7azomBYam38GlVjTQQJSKMbgLHoNv3BnRNsjPJd7SmiGc1lo/6IEuK6cyFnde2ZlfXDaAWeF/XzfaleDfxUZLWmjY2dvo1+4rmTfq5l/2fsYmVAFIMePlcGDy/HTQINKYbYSxjF2mE90Fw97w9BtISyW33W/Jjk8bnK5WF1LzBDdl/68MuURxWYJbdP8piDlXMxVXEk4Tp3ks3reHisFBMde8fzhAjyFmGxkeSxmAiG036S+5L4+v53g5wf58wFE08itSj8Gwgcww0E60C0zXyXRCgdox+5x0shzCclgtTeO9niF1JFaoNmYA9NquW58/CtzkO6X+jWYaPrDheZV06zPCHyh3dqDOMzZQbzlUWldq3bl26ZdlTYVs6uyMHiXWhvOjSIU2X44CNP5tEkg1MiJ10XLLBIrd6FWWhrxKXNE4JQ+BObVCnPPVytstGv/krMspANeevV5iMK9ma61xgWy8Fx9uBJcR2Hs2u1qdo6y9l9LdNJi7Xr4BqaiY9Qr8gT1qoaCShhUXjPAE82xAntA5gnQu5gfHXv5l+YU3Fl8O4gYxkpePXYDfFqXdr0CfjGNgI22uvi30l+a+oyhpWJQKETCU4p/MTjzg/+03EEP5iMVbEVGbJEdiE29/1ykyccRArAlZkmulFL7ddMuTJjZwba3zaMq3+7gw7qDieqZbuV5h6ZNsffd8oj4mFN6GXV1qBbQKM0jJpa8YJzW4y9lQ6VBYyIgtvexVNxltUZDQ2lg1U9vmWBS/7WYqYFD9CuiCSBmR85JCkdXsay0WfbCHI9yn33i0zmzaNfW6ew+TYlP/PsMAbOuRjZG6ooiZkmmWCa8nflShYFfe7P8CPZvx+Xi8A23FqSQD80epURmCqwan/HAi7UnueSCAuqRNsWQmHzwD+vEsKhLXSjyKnI/dIjWS2jV7nbSuaXip3QuzVPXh3b0hPjykNizuv7JdWnnl7lWryX3fNBaFoA/TA1QhHFsl+ObQrnVBu7U9mlyljNln5DOXetkTXtki09/As6ygKLYgN9+sK3efEUwFhKLtJZsWTjugfzvYh2mN5Wl4bEpMkotu1HdZ50REs/AOTAyfYHf2ZHa179KDNGE3EGAthDCuqdMFl4dy+crhcFqzBptIJkox2U95bdu3KdeZu7qD0YNYUO5onIXkp+q/0rWSOi11+8L3rJDa4yR9wpokm4Vgp7GKa1AO82cCLl1KbMFWPkJ4tf8VjrQLHVgUW5QnK1NLWUhB4RRUEnAmij8cQl2lz6REBFbOiBN3gbmt1oHvP9nt7KBFLxQeXI9BKEAAWPoAQVjTLihN10T1J680aoDS1z/lBqUe9+brF1RRx0sUcRcaDUEKiQHjYmPUdRskVnDvBXeK6Xb7T4UrsukXmCSM4LEgHlHf+Ftlq7HxJYAplAbZjIZXKi7FyLL4XYlZx3bQnRhkPnDX78q3RliPS05RHP0JLCdIqsr4j1JhbY01D/fuPpWlG0km536t4lkY58bioBECNwhNDzaG8yplvLsufpCYUoLVo2wqD1bpU7XCkoGUWs7vzm5bZ6mJsTQixfOCBqztv40PngDwlzzn3APuHt/ADMlKMTL6gUW43/PBvYImmgUc3sPeZcaAFmKI2g0HQzSWbdWh4bVGU6fQBIOotfAe/GStU0IbRBSLiAzicQahYJVvCtEfyQvP9UegJ0bu3R97W2MQ9UoWF5cXFM6TUtpdqbGGYy3JaEg8MNyOPnC5/tLrqZEWptyztKAhyN2/Weva117aLF/0xlMjxyVRVkNUxPjdP8Z8gN6Yyb0IY7njxoNTYgkbJVCwS/dWiqqCr2Aa7khQPqP6BZxzZbGJ9SvBsPqP24JYpyKU5+n8nYUCYQc+Pk8cBXhLlB+MeCDqQALnUluZIX3CDQK9XQqeX+8hszGzw1wxGd8gw+6LXV+qi+pl15JkNXcZFmOp/p/XP+974awJn9VblN/EPp/weDqEsrV++4XvY5Y+MMAV5Q898BW9jHVlj2qSGcsm1/TmkuHeNrW9LWvAEHhtPlhHyQjvSe/cpGscWeJqL+rK/n3JZnpwNFhy4r4B2StwTm4sPOTRPeoqLKbuHsVy70QLHHmrsdgysi6V1cqfi7tMtdSSiTijXJ9zva0Op4xOusosS46ozN+HLpFxlK0vz26cu4EN3zkKzX1OoeSwUhscIk5/QlZ6w6676lRxEuijM7FyVp7uS5sn2JRvdsd5vMPlSK56ytCjQv1OEiiky5OuYnpwiTk/bHWxPke+YoYGpGPmh39Ofw68qoUowHGx4ezpZcTmz99Eyr4sV3Kf1lPEVwdL19wRypImVp8a8T6X3HdfZdoHzz6RhAsUJKzjEhQssQFL/3sbKtQeg1zLs8dITvy+ZZI7t9gJaEaYNGczHH8kF/UBWwSRkZB//2rMY7jh8SVBJbYzdLxoAY8ccTod/6YrIXgGBAWO3OwCq5uhjSJv3RWqdkDmSKNWfimHLkD+IvX04+xSp1eizID7+aQMIvI50KrXhxE+bkNkF5VFjekPF/ff2IJ4Pe9o4LdQHAUmsIDKf5f/3OhBbR93RnGeeUgrDETXewnMdKgsVFYyL/+1jyspE+m5hSGCIeCDimXIslOvBm+5DPNDB8EPzlpsPzMT7aUPhy+129lxRkdsVmOOzSPS0c8pxZmZGYH63g4p0wyXYfFc+wL00jT6ZHfEgkDurOBsvUwapNPMneFlZ/VUFd6Z/W1IIxRAp/cckVb58FXlHbRLKoQ7h2KPJVCjFPBQ4hcvtZmwqsZkw2JXhWqNdL88ZfP3jp7V+XF+7lrP8AUcvXcRKfmaT7CnuDS2WLywMcFrVGQ/FMG7KS07O739yxx20nItUCAFDWA51uBZrFJ1G6F4ShJ8EpGP2UCBYh5CtqOxaKilk2DvjnEgTK/BjsUJbAUg7T9hIJwL42+AoefeqmjTyXqXJlgP+Iu8tJ1ND7LnSIsrmXwVBFeAYs87p9rGni88P0zP9K4gJdLdZ1JLdE/ZjuqaKnhVsHgCHpe7lro8c7NgDDON3mV6/UapxRAbW+ND+wm47tX3qiGPKReYW76hQjwE7O920K0nTmiHykccDND4eoEyMqV4+N3iP2GN2v32gnCqL0+5HoXN1lY3YtKuaTw9a0tvlnaL3PQe2kZjdO/pC2Pm+czK0LUAxRO8deYgscxdHfmWciP82/e0L+T+hL/WKx5W7eH6FNb5Gy6NizDYvOlF5FMmM6w11hK9Wpvu0WkgB0kXlRje4+ONRDDvoEONai3Ekp0WB+GYTEedB+n/YNP1YlzPc24L7/R9NIscgyKtbiw/7peoTvYF9m3iHLw70mpU+9P6eK+z9DDWX4up023qfPHWzx4Itu2p4i7mMCbkGMdKOHaYNhr84WX9bJOXH5WyJurvNFqEZ0wS1VTQCaT9/dsHHv3tXcRx4abQ5G9Ljov7VBtxGrGz+T+iLEIf+KArFMwWgNKkDxGhZYxb8NTDiaACuj2qm0nmn6rK7Ly6Ym+RvLzOju+nGxDy8DP6G98i32xilRWCqd/EAja+vvwpiTrvrtcoPy6plHb/a+gUwWBSvgTBuxtyfMHoTPpkbRHszkpd4olv0AXXZONZyNH8WR77quJmyVCrzHnQboC/nmlxOObY0JvRLYAxRXiTz8nfnHw+hswsAP2M1+KotIS24WX5pM1rGkWltkjKvsWODmPyoAqIzfOTp5An0ZO6OZfZ6T/oRw1ZCWrJMPf5eYHjjbB0XeyfK9SKafoNjvHQMFzhONdb6ht1MzUAsX3xR6nTfjSDBJGqpLKxdAwcUW8/57oU1v5gHc2ppVYfUtZ4JDzEiapYjbwPw8+gWQcb7cTikMtdk5+9V6oooZFqO03OSD9PfNM5I/L87q195tVl/c/OlaQ8Uu2d/37NjNlYrPWhhykJ+cBXX7gqtKW0FSfnp3Ypjd0TigrHx/5pIsMJzzG5TNFwXOWEk5v13VEHmChUvW9RNfD2yWuCOZMol3jXEXv9CGqgMPPpYCj3DNlmpRh1YdCBb8wsvPuArPhhn0wVBcDybg24P3ePr5MInWUFW8KgaYgML9E/GDdx8pw+FiTqueV0/RcIPX9kgacNs0LhPRmQf+8zMBOEiVqotqqaSljANA4U1CP+vNwtYhGD1vGWqvrIOmueuUnCA34PQDqx1AIwuCmT+JW+mUEBwg0GWnFOM+YifkpaIO1DZu1XcdiAoM+hGpV8yuBlcYsRzTv2LRs7w53WPIaM5piFj5CepqznyLkYqBskbxBxds+nGiTO6qsucY5zu9FTi/3po7uefRPUMbRnLY0JX/DDzF0+o1t84Jerr7mRj9gyjxrka2fWbguoftAUI/SN0Ssfxq4t00UgM4uX9Lbydb0pFaQ+R1dwATNXggJnxMnjbbV1GB+rrDHT6fQ7Vao4kcxvab7kesgjzySVnH2D05J3UFfJNjhLMba4iOLynZ8hRtItOzYaCFn/EJEOwgn2PNrOlvDR6dWyZoPYDPbml5qt0am9EaJrgOfI1fKFCBtp2g/oleIX+uJgslOvIAVGqI7hdbk+Nd6eS64lks8tQYqlIcleqAEH/0UBOBSc4ljOTN7LwArJYCym4nUuVULO2+XFsvTJoRK3Lw+V+5UdNT85TW7h3c7zdd4QgMrKtKdHQWoe4hxzJOGw3QgrGT+KlJ0oXOU3a25wNY07GvjKA5hLFcpHqjCMTf8usPd/2mzBmnp3GyvigpeV+1e1FscnMRgCgujP96rb0RV+SS0nvV5mfpiab/2lBEPFvBXuuX1NRyfyc7Gb6zIYokmgEHPbvGmUesix0PTZ7oiId0nEJgDVTBrFURnyIkneJn7NgQj+RuVcdaF+nAa6gt4z6w/D93k8QEZg1Wuk2qMs/V0OeCU4kLEUimt6Dcua+F66E6LS547K1vKtXzYzS2Ye/kkziQhB4Hz6gbityNUbYC+JUcm/798XWLGJ99uK/41hY/qPsSuIwUQMAdWOMxXqHsgQYCT1mY666vfLtWDcl7B7o+KQwX7TF7qkl0RBIFXDvOQQ48QBZimgwtsG4RU2Db8m+YHi4guJbir0xKjpwikiXQo9JKHn6d+T4OvJNGAee/HKJ7dksYWEuEPlAHQIAxhUHZtkGa+0KlPjMicylGFCeGCAFdTy+Mp9GxvpNRJAnkznBfq5eMbRFeBJTJEHnouyk9ImWr77tRn+6qo+QadoEqMkXRd2t5vnouMV4H9y6Bb+BxQ3kXYBiFDLNZdzXSOXy/mMDjeL9D7MoPT9zKKXE8FOQpZH/MgQ0afysrZSOt4RtoM4ZUHT+U6ObiKSmC9BAo+TyrdmRgqGRjrdQa5ae8a5uEwd95N4MvKxhptJvdL+mWugcTSJb3+9GFSTH6AhVp8XesS9wITW5fV2Fa8UGbWiqv7WKGqqO9k5T3pVK64x2jSGGOceFKlO1NWj8NwRnzK+o0p6g4cMb6jxi+CiDMG16uuNof46876nbBF3ePOiXJnfKZfBPFjFgW++LQMGC+VkIHUaEnz7U/oEstOt+4Ob92pjcQkercvkbrGiDVVoANCUvnXm7F8FreRA4avYVwWzaR4M3s6S/ePzecg5w9VPOdT7ltfpRH5gWjowlH7vxpX+bNg6oCp+NkcBe3+b+WCGVRO3DqQpEfgV8ale20hsom2TecdNDA2zGxIb2JzIppfIh7PWy0Qp+nxSs8SB27CHcMW8IybN4NkqFVo6b3O1CsJAq0ri57uhQN9xQ4vOUEpMJ/q8m9K7mFCBuzWP7dY971rndgscHMTiqUejMGeBOvgA3BDOPSlmEkQWjB3an3rKEx6ap3LsM+FB79gC5ZDIszmRclUrzFT75ic6Cmksf6GEz9N2IUlJX6T/jz2YcJDucOV2/yTaUWp3ysAMudQUmmMbNM4NsUvwyatFykG3Ww+kyLjEBK3VHaMwZO6VKSkLx3Hseb7uspztc669TI+syfC8DOt0EEU5ULHfXFs8qFPa6blp4YLi2GYmXC5yvSEsTm8sR9Wzk2nWp6prHi8DgpXvubtmILG3bGanxFuwytCutOuctL6+mzCizNNsQUDVqPi4ytxFu0fVgpSb0kYIkxgpAQMOpXxBb1pj616J9E6mWDeOInYj9LSbuIal8B+E1dhlr0Bk4sGECmqyLLIMAKeo3AXRPzRiPfBStC9FIJmBJZ/YYRZ4wEFY0xl1Vz7p2i6ECTCupd8Td95Entm54WEWbN8SiHL1G8CX8FKzCkeO6N3+S3wJdeFteaG3SxcTJrGp5PuubLlI3yI8KhAtDf5Gqf18Yq7bXSuyojDFEmYOicXhmVfcGL/gdVbpQEkC0quGbK6n8Qt3qbhwocG7Pw+apgZqsK4m8FwP6lnY6KFjAYlV5oJo8HxWC+SJwMbZDESK/dyt1csqyVn5WL4tAyzuYJ3wzNMjydIVjqaTKfjlp5//3OgtV9LAeHHJdn8vhlOGTd2sJyrQNVugPHFEG8AiomsXYS8ia4QwsRVuTseDQwfdbhXSdtuuVt4iIo450V2axeRcTo21Mg/+/mYfqYMleRU4fcDyi2+9Gj1ivpU2NYo70Wbbb92VZB0WGNzAUY8yXkIkwYkV8kWGVHk9VIFIIoxvok37pz7MkgdCTL0Zzw3YmQ//d+y+0VLAaUuVdEC5BIX2AqedgXMudqxnMejwi5pCPFJSbGn10Lyl9KuDqeE6HpeZFY5mRs9hPBgZ0YWEpKvr6WpyzLGp3oPdLZG3HR4Nq3OxiLaKwTFF1M/fYiQ3uo0o950bS5fqCwOdVQDSUUX/3kr+XaoVrquqU2FdBq4M0Acz6yjV9GvJWFSSGOHoGTIYyq8238XwqAOMsHvdptaWyeHFj2kFvG1EgBQhZMyegVQVxHbAWq3suOtYZQPQi/ujApdH/wOkmCPS+XNGESCfpDu1NqPbntJ8hZvkx3q2c4KGP86oUW1OMsetpVIw8yR4euYTWxyhVWRLAqG02JiX5kywAo+qdsPYf5gPAJ9Z8YLYlnJLRf1Pp9KweI0Dbczsy+y10BP1fTCjmkdYby5J5EkSLyREoZruhaBH91AwCX324yAs/P2kdup3qhUwE/IR4OJiQE7F4DlhkYhMQglAxG9YFr53UPKIoOmmN/UNhVqyPeAW3zzM20hVZRspXxGWDolceNjuvkhQN2YE3iz8VFnBE8cYfJxIruFESB9mA1k/oSg6GrHloAxygoduemLt8RbRyHtkydSANOWzKJAHITdSMFDNNlsfD5UK8CGQ0LQ9Hj4JexXQWOz9tCB6YOe4wayr0wnGqUYFJvakK7gok5R11CHE+oIN+PqmJh1LgiYG1PJt4rKJbpRFgs2VFvmpQL0vzfK4plXupSAeOz6/wEMhd46o/Pg5N2IoR7hpk9D6kZwhxlDhEW0rpv1IpUj09SHeE1ZS1SYmmYk/mPuYH6VubMupQGvINTVVqs1yZf9ybp50aOhkXH9H8WDhRwRxJEF1Y4VQmDfmBUwF/Z7wKSkKo/ldeKR4Yk5j5VFxWlagMxtuDP1TkS3To63pHxsMMdtvmA2znqe67jPReLZKAeTmLEdttf3NKaPxs8YKtIHYT4OKq+vCL7u9XWKyGCWiWPc73BNDiWdlbILoD7vM1G6zAeq7JrIGkLcpw23bYtjG6fzLIqtdyQjeY9bDn0tS/lpS/1TC4f7cwrHWnJF+4nu9/HNtq2nBAGCD/RVsWj64mLEpdzKdYFzej9d8hHpGImL2FG9FeB29Grbc3Ynykd2jue/1RxKy3Zv1xoiRN0oF4X6O/teHi8ykFZ041W7k5mnGPJcJaMDJP2ackVRkvU+yooHUPtVLTse3iPAxY0oje/PDJLt31HB8rAM61+/hhKal5Ter1LFknpkH3ekM7ZO02L3jp1tU40Itqot05dkTLw7TsXHGGmgS6On9E+xtU7TapK+/StzMirBx85dBSbkZeBiBePTdglK9m+HrF+51F6cMr5Hd/KbYBToQa4e9mt+BDfiq8Y4bVYR22R+UsagdPJWZBP25NlIJ5Y+vWdWoR+2UlZYOUM5eQwx7acjtRAf1oQLPV5TLaufK5BsJTff0qW+pIG+RF09w3elQTrqK78mxtg1ZsAK3EBePhq1v99E8rcUD+Tv6pDCgcLImEFxdGUBO+cXqEyHNwejJUIYwXF1dzo7M2jCrkJXlI6awudWc92+ldrTedVURkIb73keZ8DkZOCt+JahxxqwH7gaBUzdwsPonM+49KSKritNZ4PHfryzWztUALL2ueDS6k/k/Pt7rSm4u2msXCqvWBFwfMvV7Bsm1wjpJu90qmNKCkstx5LLWuLhNmkbmviUNyvBG5Pn90yWMeBa1nXyp4KsOqHnafsOgVcExocqsDBU2ZieZ0rPEKHOM/XaISDm1xUDJzahOHXvHZ2VcsD/+csfMQSlfEVBJ+tmHPCu4uAQHE0CDolAlVyW58KptELqwWhVCGsPrlNJbqE7v2pqGEue83BpJZ3fT9oqh15/eVoglIdNjuIU2+jpBwBfOLBxJwoej8yX1L1gZGEm81i5Yys2oCo4yF2hCVdVkCday1CXKBLuNeLy2sf772+lXnJob8IwnOTzClAUJkRUmzpg3XjG7imaeQkmRCa2m3w6W8dfcqeM5TLOtGrAXLeV6GeuyakTDfAg4YBqkUjF/NShr8CT1F+iiOBzOGZ1VwU2HKw5MqJ5lQ49C4/urtJH8L0bB6oiHFrfj0aZ8eIke5XeG89wFBU1toOF8QUHZaMpHwiCVBdU2yA8WSW16eQVpqUCu1LvjqzxruOdokl/PRDyZz4FkXBI1PaBASj5iJfiPZJxfpyYULJyrWwyr1RcH3KWSgxD6nmMiEcOWL+PC6JnqyD/lPBv0LhzQMHfCWD96vRDAJhnP6gseUQE22T22+2ymPF3RK/xAMHzIjskx5ScIe/ENlGDS6Q51DQP7XoiaatY5sgW5XxOxgmNxpMChGFcd1EIly/rqui3SnyHf9E0DqPwRr6Io0N7O4sAYWx36RbQl2nY5uxMQRJt6mB7cOGchNgbwVmqc9jYtmR6FOO6mBA0HuHEL3hS+HoIaVT3VBAaVpkdbU3niXeWtK+WS7Se14jtsiS+oCc26OvLV1yX9oHvNPEHmETtyFjQcbCRkrmF3lVwdkh+5yb9a0zkKWUhP347+t2MJ/CGt51U7CsiVnFAtPm3MbS4L+JpVRXzxa9qHb7+BuDX0devmMb4QXUvZzyiKYBqWLyzTLz7OfAA88YcEKI3VYj0lv8uAnodoVDYJcZZG5/xHDfk79J/Rr/xdLUz8KWfUwHuOrnNj3iMc9PeREyzpRwUKKm0rGzZFUY1aaGdrSNKb2boWUwFzSPE65qiYY5hXI6q2ZLXyzgJWuJotbMVTggXUQJTcZSeMirFD+B6gZlFAOMbAswTzVYtkw2KdZWopdFZqwhvbovWAXbRvCH2+xy5sJ87iP4a5ibFY+qRlK2ifLk3lIsmBHHrMO/cyJlOeSs6gOcCP81vmQemji8csK3vkALyQH2drNQ2xo/b8CNTcFF0DHODyqJsOr9vM/BRyRAeSn60ul+vhEx/NlicThoOpnqm1nt2vEt4/eDnmXRon/XxY3EpSJ1P0nYo48kJudXRHuHROyJocW317Z1sM6V4Sn2bp8Br950WnD04XoqyC3ZOVNqFulas4EclYjn5dCUAvdc7Lq0cfZpeIfGCwAjMT1w2j8FXfOkM6eoVjK4nRkSWv2p69kb5D3HhlMSDb55ZshWl9DooWSrozf25Ob0rXpom6CNtQMAW8bAHPBZlfLCdoaqekWY8Az7kzeAtr9q3+7CG9zEO28Dz4Rvuq8fWmBL5EYT4sqC18fdWWgOgzpCZ+54ex6lWMzn5wH4kRWzgJnSzSf3mjAOycdvHvKh4WfUdVTthBy7IrSzpwhrGuezUfXo/Atq/3M0l7j1qJ2eubLsfnVnDMiHpXl4aF4lBQYLJ2x1h45KdEKW/KlGIOfLuX/+oV8OMADdUuORdkdJrLCn4KDbSIrgFym874yAvIv+OwXBSkjG6vrwnoFpPkg/axo609gk/Tmi3TgKZpv1EjjM9n0oMEvi5ZwKwOJkUhtw7hWxQIxA2x71R2Gi9laklLG++EIffC/xbsvoTaldyaK6KNDBi1tCdE5XF7K7uOV7jZzsercjeV4kZd2/yPV+daX35SRYpinxda6VzEGSpSqhwbBgdqPyKWAEe9anUJhmUXONsTva/5amnf63fCOUoHssOw/2EEAFVzXMEqXD+jh6rs+Y2vyj+S6jyrI0xyo96QL4JtbyFlHx9yhrhXyTvwAqzYt9xJySVoVSI0p7rzeS3GqvqBFiD97wmeOVXTADMIYlzmzrFPB0XC1lvdHWngHhAL9ZI8/iXM+FMpm5Bzd22EuCKnwoJpjvszggt0Hq7f6OOQcGML8S8ISO0VQxMQ/NyLWki8LwPFkBehmgx799vDXV41DxBA+PROb8CRafzgf2zgkG/zu9QCjDYCU7LvIOfSOuOVVbtFrz3eOLahOt05ajDJcJcCiIGSxb9SrRyClqC7g5E30xru7uQslBwGAmk5DtBAoSllvh8sBG8SaoXTO1lzRnYzeLjJMsx5gxo0S83RYRK9ajzCI4YD7I7JttzH3i/7cKr5y/XX4suiHnA/IoLqPMfZvwrEyx2i/Ef9VWbYf/zpK7t3rtyqcLF8qKzGCiTC0nqUpHxJHcjHWOfNjSBpUx4kTs81QcaZ3R4DH37KcGu6n9emIrlqxFiX/USx8UvYUhoedUf2Kx/5JChRPcLDcFKpe3j84ALYG2myitTCj2+dmzhF2N0WOq61wVKiBOgLwEKAi+aHGtC7KDrs+wBXF54psb8q+M9OxilqSiwDM3lhUSlo7pJnX3sxV15qcR1QNev6WvvudbvnduIALyuOEd8solVo57AAEIsZgJXEpYnpHokLf1snlcx189SZxfMWMmJZHvRS0dPZVQHimSVrE8b6vjnkmEmLEbLbdyYLRAx3OBnSyi4EXvsfLicYZ1EgcWpK8PzpAX52SHjtGWnfo4h9OTCIL4LzAYkTUf7qFZ5rEGMadhmFySaaB5uH3EYGlTc/ZxiS7vjqTNcfl/BCyic/jaM0kpy7uFbAfTaMa7Zfu+hjBmHtUS5+ph2aZj+JpH7vwkTdTMQUJk9Yz7M8X0wSUienhFkoaUv1PN4a9HzudfmFKZQQjq31zm43/uGZujupW0quWyqeomAaEAjMrsgGAEuhpOysm2zG6xmZo4pOEyG96UMaaoAdkc8GVjxHQ7wCxUfX08YtElORXcct3S0T5fCwimBoSDGGHjRayCOiGETUzkNy8unA9j+pzCU+Q8TVWqU+kHAgB+9W6diF5bgKWHOgBs8Ca9jx2QMd2JsGiVaS+kYHmJLmAFhrrOYonfB1kcKdi0WZcIgZGExRyTnAoLM18j8/uNZ1clD3FB23DB8ZfnzwqNRcG10A3S3RpDbJaLPM3Ydty2WVO3Vb6bYk1qqJlKa63RUrMhYvMMApb5O/G73V/VHEe92ZqCDJDsge3rMnV2LY6V1UMW1MK/OkcPF8PztQT19lFPCWKVP6lKPL9ouzp1V9MsoUKfALqgsQ+AgETgnCcsE5IBqueN8SQN4LNkM2R6gLkiGpq/TNUpYUgBU0JemXF5J814oib1608yvQPtIH6NTSZXOepPKBgD4gB527hTCerODnH2yhk1/43wk67LW8ncIekhnh6btMXl4G+AxEHSxDdulmrBV3BLbQCVGJU6MkiZQKsrS8uMZLmclfsBPRSxDRAUaCw8BhXvZ6t0JrWwhA7uX9P95/GZWyWAWDRMnffArclxVzt49OpM6OGZN3IukSugEIH4S9wT/I/a5qDNHfjiWWHBYVgs/RbKrTTCQvQVg1UXXarAiWauCgGt5qkKiww79nz/k3NDHcJTFisaP259+nNP9lj1DgBYJd8g5TOMyoYWmfBcwZk6B6qTKqCrcukr67FkkSv6t4+IZl8jXwoDS49yQ5g2A1NogUwd568tp/YMmwG00w+KrfBHdjtaV7XkR9VB9QNZ7qsya25J78DuPgUnfrKDNs7jPaB/E1FXbOLpdNQEh7d0auXT+AL7Lo9EoKHcYhepsHQeUnUIL74FMWVI36N/4rmiQbrB4xu58pCG1C9b/aUbbiZZZvrJ1lsagZbdBumM0i+DPe4tYmIqvIPiRa8DeqyfS52ahZSDL9Sl61bWddW4y23eD2VwQ8H2+oxw/dpoPGBlhBCKMhYM2jhXxNOJNtsOrxoaiqUHksAcsovcMgLxSnotzgJHWfP9oRMjEw0c1hYTnL5Rd4I5WKmUBW4Y30JqrRVIuL2OxW6656ZZBN06klKHbPySCZSmtDiMAaybovzx4NiujwUpjtXbX33D0FvPFeLbcpyLkJOtzvSzbB3cvZBSLdbQXzOujGwFn5s33CGHpcpzfu12A5wq9YnsjogX0tM8hWmbNuoQliurh8qDZ+RovzG0hUDMJmkDqVHOpYuWPcGHnxK5ixT2FTY8X6jMMLToJyZA2FVs/c5+y7PeSox8+a683Ns61R/xPwFzBvj10FnfTvO6Cj94diMSE+UMuMxpYuDts2lB7POiiy56UXWKQodfdwt1gVz9oBryIr/8nPh7pTtgGaWKqEzvYzEFRTP2Qw0X4Ivi8WFJsJVf5CP0czihuURTlLFJfSfgrATyMGLEv7byuVAjRQuFCP8peVIfx4rJZ4F1jFFoc2qgPjzJ/dQ94v01d/70DHRIjcI+wJldx/XF4NyiGSvqladNS58MtvVR36jFGchPagAztsXRW7uNW4u/5C8er3SPAvtbinl+F4erOGAte9ZuhYsPLqj/rOtf6weZjkV9V/sSfnOvSgPVuQSbi9qYLnA2CFksqp0igeK5c2/otxoPSB/3NRrudI9Xpo1es3RjCl12JjvmXx8JFu75KfjS9G7DO5SPQLXk5G+33uo/EOVmZEayRhBo475NwO5yZntERaTNrCZwr+EgQPEyl+GjV3r9jKmEBrRPsIwoXzIbVtUQ2BZxQx7GHuR/xinBnHDsuEoNJ1x96X1MVSSS7/Y8atccuXOjHSBxQHjnlT1DnavU3Dj3tZzpy7KeK1QKcGPnFyskaHit9ChfgZ2bOb6mor51sjH+1jvFd8qCX20ViRMZMl2aFVA2UAYVOLhkkIBPijL9Gk2/W/+gdV2vYtabXKxi0/Hmue0SNDSpiVs9/7iJp71/59zIPqB56ro5M21Goorx/I6TG3ZdnSFcn17Ss/MER14XeEm8pDVHG2s8HK7xVUJQEEZ8kebERtNR1rvsFByi2HFJ8n2fOV6/galQqWWuJMdYHKck5/b/wdVaX4s/EsIJ6dBKi2rGuHbAjI+TIshe8GCzWjLEnynPBEsgQ4G47Xiq1CIqAsKslBJrbuDF6e/Tdt9S4KI9QHZV7tRJSYFx/oHXoe0fhLsw3q+ECQ37pb9FBrx+YaFW56XDTjE8C/9L4LjPy73d2Ks16xdw5cGGetODYSLsXaQNd8Zk8NkRonXWbYlcDky2UnbN+ih63ZSsWvHAH/uR4HhWJNegi2+xCj9bmTEHpeJ6vjFI0NfowTP3lN1y71dR/LuPsydG3bs+vRQDYqzzDT+j3GX4x0GiQ/D49y32qzok0wPnzFO6gC+MRZnkHRam91VXfBhR0l+eWnhfVLBtEONObb/F9wrOEVWUgLv3jf+GNismnV/YRbVFXUMHCsd3DZcozq+/+RFWyvLvGwu+p9dz3xjiKH5hAZ4CnyrMkZD1JE3vtD5Fx8hpL4UiP2MJ0ve2MilTG/uP8VczHtbQoozgz2E48sJUy2WfwtTJp26rwCCv5Tkqvx9husMFrdEbL16OTPxevwoRRSwJczv5AyIF42ovazsmMtQQW5UBsLeSiimp+M9neiYJnPNEgJQtHbkuzxcS55BGVBASbREvNQVCJ7kGxIkMmqHnLSo62mvOg9MzolK0oyQuhciEONN6zchMXYisI0jJlCW37PkTo0ndomlJMI7LUPcf6qp8EqrVzdD21Nf4ne9JnLGTSTjjbVt4tZxvnUv8fUlcCWPLszhA1OmUiftUjNbzu9Yll5w/Ryz0jDjZivzZc6QxYZO1ZA8LXKPg+xwGu7wV4n7v6S+xnUJKo2V8W0oAb9bpVdKhhYODj+z198wIQw0RDqkTWOVHsbG7h83xzWAOf0VPIYzX1zAwg9rvTAQQ9d8pLJynYpGS146nTSCMyQKmxZwmyc2JelIh9OrFQ7zwe2AES612GwSI9P7n3QJMoiTpda4Bqk9kqXwbaIB0UOjk9QTvQc1aQ+yPYGzXeqcvvDgvZXrMdl4JZam7aOe4qJ+whLpxXcnaTw8Uf1yCMA+AlPAjtO+n1mJCnfXMHe0TFOFEdTt2NbgvsW3L6Vf/Mf2r/B7iXJghKn9mqPyHMNC4hyn6W32h9dXFPcfZ0IBvUu6QMg7d339w0y1804m0aX1ViP0jmztuXY8OnBajfHvIR2wx95KNPfakmrWOXaq7XgsBLii1nJlsqatvsgn09lWP/LZxC2rE4za0H5/ZYsVXrMX+wC6LsoD0sUVHyIyMlR0M4WyB6sAb0DVVhohfH5mRH61IQuZ7yaLRmoFDm0kIYVA+Mn/OyUFQ8Dgq4FKWq3u79YEaWGprlpmkYpMSO6oqcDOn8wuzy+xa8V+s/S/3uAHfUyasF9UHOKeIvjUBWoRsl2HjDVvUrJICTJxKwrQ1rbKYJ8q2FonTBY98lW5lHhb4nHXUhknzmnhTbKEuoKl6f11K4QIVej/vtEmifCp83WWOFBKVHCBXR4a9/gh5myClFqxAUQ5kSIdwEVZyjxSl8Th9EVM9CY0CaoxRiT7vkC93tCi0aBTEiDXFfad6dchplZTQJYTMSIMhjCXAF3iXM8EuB7v2P5SXfR5YxvXuMCcPYBcdg+p1biCCKpVDcNTrYuO6QMh69mbP6WFvqInG7+71UWK5iZCVDj9tOWAD4afa4yNY/IKmZzfyBUjLN4Zgunx2shmB/Q20/iSaqXK4hY4PphruqLKSn9/iaKoP6PAPYXTOcMWtgpD9/2Zs6lV9MZcdrh0fJ0PQYZC4h2+aYecyOjG/fD3AH85we1t0wNIAI2np38T5VkuRgkKROErjRB0iQX5IB9gL7PeVtL8c7oS8CU5XG2PeMSdzShjS3u6tu6bR2RaHPDnxh2pjbXDWcKsnExONaW9tQtOo3/EEgLXlyhn1B/YX3tmvqyDQAkQzb1qSirvkf3EpIJeCUd1eO1vqzIrsGAE9k1v/WAX7gXZ6s8RHYvztTbn45rgDt/Nz1JMuBRpCQX62txFWqp2qdClJ3ywYFT1y19yYO4M5DTmYvBaGcsMxPq5aL/s+dHcmvCIy2P6Ogl9RtXJ2u0IkBZI5GCwcyAG9Dl+xwQCpYjQl107Wmda0FAzqn3j6PhHQnAnT5868q8vG8GBVHj0ZsKOVT72nS3MrN3z8IrqP5EnUtzYgvmhLDoUTJmtVMzrWEycx5jbrKe5RF/DHp4tbgO99xCr08hVMlUfvENnxkSRdmvRWI0elfWXzAVB0notwrd/MTXuzL4XEcD4d54QUNac0t1qvNKMmRB0cy71Ls47yb03wFbpc1NDkKz9qIT1P92UE29qlPRTyE9lTcuOHCN95rI1BmPJRKlLRYwDeI/tWu5JbIE15TywXD2Zvuv2h9XiGj5Kq8h8jSknYHNceFcLQxp6stMY2J7e/lYz/2smBJMkFfAv5mkNk5JIPByW2kjch+B4Kg+Cmg78wmMUxyJ5ITK2yXtu3P7Dv7A5K/Z8xGGOaw2MXD1JHizBOdnuQ+33OoVhMJEU1W4pDKFrAcqUZ3vBpK6LyiVya0OZoyUhcl04kIMVt+8YaMa5o/pw4bYJYLfOqBICdxKA15o1hsgTTAmelDdu6oGMG0FbtpoXdSx40xrah6Nu84yjGOpRQsfZ7B1yr2hf0+8DjjVkQPFGxgjxVc8gJrpKyQ++IdYgFkBy5AZWff0NIRmUrNZnwWQFnBdfYQYBopO3GPb8a7gQkrvwCDhtd5ZdmolO5qOuGiQCMaWs+zc6cb66tNGjDHobhcZwJkhMVjrQIyTKh/3NfAHrTjjMVefdwNcCo5LAKLTx8TH4Wa13YgNBnYqRGVJ/DCqwOhPDpnNBgGVSJ8oXjGszlUA2dzyD6RKwieC8+NG4ONbf6flGO6n3giDGxT15msDhy1o+E7xqnylRBZJdIxQ4i13RKrYaAtYcH4hOLQrC1G/b3K0HTa4z6kwjm2qUPr6/b553CQjgooE9uS8sRX1RkkJ5Raq19PXsmBrSPvuUYYbceQg+t+dWIjXHNfx2PnI9k6VarpadoMlTzEbSzkuCs3g9PAyVgo79+2v34yOGmu0lvZxOF2LEWNhvFsl/CSj//XZSwPoU5wwIFEudKniV/vovQtP16MvP5YtgGXIb6kpE7QAH97vh4q7uzDIll80gPuV361n2hKz1L/a2NRiNCwUUBdRuElgykDvFiqESIetm35UAPAjCaai86PjtLE8owF4DYV9Frdax6mVfl2gDfRUoEBwsjpsmCybgmAdCOzmE64eFLJM5cpyKY22hQpbHInPW+r8bI2tnuKi/30mKqbXTWNoKmyVWCoKf3OYMl/lICPgaaHLd8gbeak4NlAPnH4oWCerEik27hD9rgi9DVM6hZP0ryZleaBUnBjsXxhxjpEspA8h8aZu7p0/DpWkj0Vi0eApiAEikv0gGb7IPcy5eiZ89VdWQCEXjiE1jUBJrAg1t3vJ93bNLLgBvkq/S8IpZCQMrRUKXVQf/US14GlMgmuNPtmTw+pKGkb+dstWdkXgmItOx7acVCz0gQrlPDQXG1SEXSe3DjP9orCDbgPa0VRjxu+qSKG5MkKKcglVcx39LnqZjmyn/w3dRFEOQBczJDWbydRq+W031Bnbr2i2B4EsQXF2Mt9SwSFxOlTQC4lZTlqsvz9Cm2cNWGs/RuvtAXtmWrIfnd9xtbaBDnIwf051ABVulXMpS56gJE2xndUDCBjurGGP4HDn5p4Jusu/nL3xeqLEnCgeX98c8nxqdSrxZD5wdrvUco6Kda6mI4TjkQKFkvIKL2cwkzX6/P8OFjm/4EsmUwgpS4UBf7Obc4QOh7A5xUgB05tXh0eX+A7Kp/D7loY5XCCG+rcdregYKu5/ErND57odwfA80VuClb0SdFKNajOB+FqMhOQgdwzyxPw919xRLm6tNMVGdj5vZvawqvoR/RhCqSwWk/fC9hAnefwF1HTLeN0kq7lGezLiriIRtFBftd09VRDtCmqZRlB39Bh2S1QO7CoJdyZTzjCU2PY+jDNpLLti/HAl59b5IQRU28/T4FlkcD+rf0njNrlGsQCNG7ROiDHZLBqWed5N2RSSnySSr7NdIF7pQB3ByOAlXC/BonNBgmqvgZWuDGN8tnJVgq7UZj7MZY82ylbep7CE+B0OIesBqCWWC8qQqxHQKavkGjfQIl9ePFLXyZyuD+h2gQyl0GTukrxw1nc3K7wMyut9lXXDDrRkrrZRLtP1esL9Vds9BQj/E0NE/rBlurxb0NweW+oZMnfRm5E1ZZqiCBOfDhQ5Gd3QWhneqfwSdgbGvv0Zlm1FbPt2nErWk0WwepbB9IwRWGAGdyLuWhZZ0nhyhSZkWlW0WWCdxSJ2JAnAzdDeQ2XXEWre2c5rM9N8In1UAOq1O0GusxHVzMs8om4Nk5V/fMPInxBoYOb0hgXlKH6aijpmz22Ve/GSRPCLReN+JyXhTir/lfk5NLFVDhB916aKp5QmTT0EWtlaPh5t5gqP7ImdSqSLaxVSJxAUcBn3JDEWu8E3iR85jDY6aZOfKqd8JgWpZm9LNLinfl3TcCNLX11jgwboz3RsLc2Fv5grBqadrC4Bn/tHlEVCiEarPTUg2xk7aLQtYYHJYZ09m/eJGf1GGIzM/29UynT815kTGarVyfUik9CIneFyhkuhi/VmYGQrP3twyWCOvY2Q1Rl3FbVBGspfVasIsOPEPj+svcgLtDZCSNuludM99YNyPEwSzTS3TNz8pE/U1CWLebF/q80CAFiXudsYeiipD0n7nKtO6NPYGCWpRgyF/lFZ/toPVlemmkwpOMpRtvceU34lhOCRXDbYXghIMPmkv9lJsIArVJsZGho0hEzi7gwXNQQ3GeAcXMei0n/Zhm5evQbGLEKyyFie9/MfdzA0SV20oB5ObExPq39Cpz3KDFvWd+QesibxeB2nuehekjbMvKwtzKCmGZA8cr/Zg0s74Ja4gRonmFTk73f1ERXvyCQCuXn31KRDYIHoybfapr3J1Vk6NUgFY6qI8RO2vhKkB0AGNw9CgTIn1BPM8gc7irMSz3gAeqb3k44Ry74j/2/f/Y6heWQEKzFmnJOexlp176+EWB09yVusvURRiCf9MwCJV6h6iCgmYJv7bwBeoGfKkcuEa40JRRdv3WrB1hIIvm8B7VXAwuCp7oGuz6FCu7e0BkqyBQYpGIjti7U2qJgIT4nMuTpxaC/M7RqKTENgE/AnxEmF49CZPr1sDTo2smtrSKGW8WOCRaJ15UjwAbNKmwmKzfTjeNscua/zxOM744TS6B0S67706j4NBMjzE+ngpqmVAnViPjCyJt3pgN2y5y2/TwNVVfxgmW0bWaH4q4IYNEqNMJSUddaAy5RXZxXvg2Cd+vGcRXkyZu6O+QDkmX2iMpPVqLvG4PMbN/5IOpSDEfLCH0K7HG56nhycTQenEBuFnAj4z6O+j1syedB048uqCOT3/HiqpFk0TS5LBGCuTSbSno13U/NTakhNwxZWEc76q7j4wAM2T2Ky3VW6v2jTe+Zs+DnI7gEXgnhq8X8E4oPyxzCMV/HnTCb/PYfxXvnQCKY37eiA8+7ui9kgdLacq7RewyrHP9khIYRWv7iIDoCxOQEgRFUix0t1+j+H3btwolaYe4JLMNYTTtAoCf3gjoJ62cdeJ2HPVlFdrX3I9V6QojH/HYH1m/FDUlLshuxuRE+FPlzxUKxR20g8pBaUHTsA4OIG6L8m2zz3OqXGM8+xFb8rRzP0wiCKkSNoxZITdD/ZmEYD0u6M2M+M/DgoALfXY+uy8mxdfh+/AggvLcldlx1DGwuHXahn+vWF1DsUpCX6lxaHL5HLGPFw4DRd9nRhPNL+A+0hW62BUiJHxen6mPgyQuQamWSRhRqoSWxJNO5PWCCRzBQYAm8QvrpYtLWg/yABBVHejX8SnuGC/YxXQtB05TxWFs6EtRzibKPucLIy1vczypPQPibaGGx0tEzsvLvuX8LYq9QwKZwmfcKeZ+Av9E0G+WbSKfdWVohyLb2H24JCRFVBWJWmTZEVlKIKATCYtWmZfTKoRNgnRoYB3Qvz3xfZrtiV28aqaGQpiQ6etD1Dp6SogJHzM5P4ailrkKdFJJ/JTXTZco1Epx6jhXxNZiLI2U0eVtO5lpeeaUATTrc0e5kJYZZdFO8OVOBTYlzhCumBPEPsKpn/vrCpsoII/VmSwqXRNPRyonDtvbXwwPxm16TLKHjXBEQBfv+EpIqLVfNyNkxx4SokECwo8nDikfhW/42LS1eWruZveiapmcAWlLatwinmsIG51AgMyWPgqYax5urbgPgWivp+w2htd+nG9dCGoxWT3CxMxnPR54jtcUhMi/BJp5iPlEsyAwDqMOYsf30yPxCKbwFj70GGJ95ZdjffwMRN9pRznootjKch2pTTvA6J7+fbeYw1DOKS5GDxRGDy1hr9AX+qlnQK6dmX93dIhL43pK/1gAkVeALkb3HvyiVGsXPNbkcEONIOP9jxN02RX3lCYDOZB5RP3/DlqgCAPanYEMEtM8MnbWEFoSv6H0nLmNx66gw6tm9bzC7uM30F7k2cxWRmg//bngvPNDq+DTcWclS8sfqn/m+YdmY+PAIAwRbAlHFuVJjrGuLsrZFOWlB2nqFwunh47IHphN645Zp9JLKi8I2FyrNEr41hZjp3HGUIT0hyfH+bOfGOTFgMHAu5XEvDfibJBhvtMF9VvWGrxW16af0xNWvqaKCVVFMme2e8rYVu7HH55v6AWewoaUmXmNqg42eL9tq71N3/qJ6WarMEpPdDUHch1F/Yop0Mr5foirKDnkl4UujB0tqPVLWINrcm6cNE2kfFqnss9DW4kljIKHzcgaLINcxC74CV8fgnkZ6RZBWMcgeUvDX1NVPxfUitCB3g1MFn1/PI29HOngWcNiK6fJHbfe+VHINFCx/txvmQz0WIxkEgeQmTInX5R0MLrtXQZVCE5jtugEQTiTeD1LVUmx2VdGhOHKo2O/xroXYMV2Cnzwrr/LL5g13TBAxeVLHEdoChyLtFPqRkAlCBsC0XwRkITVGsnjrtDh+Hlgw/5gW6V8CwCDJFDmB2ukNlNkVXqmg2vzrWpn54k19ffbCrcvdJ3y+oecmxJo2zkAXXGe6gOg74eQ97+NgQvBiclV1JnUDPmkyONVBtlBPSBEkKc3LvYWAGTCID3w0mDbxfk2LMbyFLLAJeHVG5dM/zjWhMogmWnZCVuhmNCMNQu7CjaLicT6pez25ThMkRQLxkyWUss4XpX3mX9OElJmcBQTZ8+zHIXIMd0PcnBVpOgzk+rA/yHuRUl3yve1y8RSEBghvh5Guy2ZFc8PfSlfRVETE3/meUi+l3SB50DbG/q8SUlSpKbefHa/rnYOij8264lIg7gl+/Jsgfcz/A5SaMuxy3U4kHmvMW7869I7FRIonnzO5g+FkaSe6DxAXA/M0GabZtGAZvA1dtwt340/cQGnYHjYmerMtBny1Pg2HZCvRW/S9jcxtw4cmainC7bnGY7YwzOVM40yi/xDxz4IrqQahF8OzcCZLYSjgnUVKKca7sGJHqN0A1lq240xu9/Xgv7I2sUW3g8MuMrPsM3hiOCLBw2OW+0/xzvS1lx0RBjsfwGwVEaR/gDq3rxYrc+bUFWnW8JnNeNufvTTUHWeE0BAqDg3EiQ7ZLfNa90Muxb15jAKsVlpndfDkBGdcqwvFS/8e8USKIfgvHAXDviHw+WoMiTycNBbS2/Ml1jAc0R9L0AzfufIb+O9x+LL+rTW2B23WOKBWNZxrdQRugSa0lHu6IwlxsQ3J0oFiw2m95cRqpKRGhVwAt+o/kAdNm5drZA9dc8a4wKb4f/kMS0IbUTDiLfi9DgoxEYogUclex2vueitfrY1QDFzhCvteGfpNXwiiscPFWg8PkMrG+L6joOtSe1myqDUPknfQT6e2u5XG4WVYOUaK3fIOFOIPDtBg0iSfEzIiETr5Xl1OkE0msXDImY4b0/8QqOSS7vVDmg5qy0lieQ5UuIQujhEkHkDkjKuUofydt9yomGHYqKVfNQ3rnSZuDq4zDpf/yiFlJJk3xRv/xrYixlcMj0iNUVH4RdYUZ+7Hkjl4hCO3GTL24cbIclOMyj6R0hwNeC63cQWv80oDE9Qn38nHR9/Ye1RTfdN9kdHvJXfgLFeIWQyVKVYacvfizBJWcjiEtnoeuYd1bID07AxOUPH9MnGD9CAtwgKlBoOYjIKEG1ZuReorVfQ2z++6Q0/+dKLZE+cP7cvSeQHhKj8RDnFig2DpH1O2Gt0L4iMXforn/cw0lgzctL5R1+63XPFpGm4dII7uSvyTP6fWaZcfw5KtHxOJBfV0UmCTag19gX2DQYQ0ltUNAMWFIIvTvcLsl9GKMsDF6EhD90GWXCaXRpajgN7D2JByyL8NMxSlCW/NWyROg9aIkh00edCsktkFQxqPE1S3oQulresXA1m6hh9GS7ZZGJm1hv6u8lsSExI+MUdUYKrAq8J4Tii8yDYlDh7Iy2KsoHvm0QxEE0DXiNaPEn2NpbToDh79hGcQl6vRgVH4c2buaoKmu+r/86IxJGFJoa6HT0YCYb9bn2bUk5OnPb1ti28clpac+nc641fTMZTnhtrcXXo8QRUWZgRNCuKz8PFI2si5VV+lSm5/q+iQi4lME6g25HUj2+DtvCg56Yg/ALbwYAa2Ze5xy3tk+jaNHQaVWxbYyT+ya92ri0QW3W4oxruKUmO+7lRc3LkHp9otBG745o8yVq4S8hgoqAkD1BbK+NYZzzHp5nfUOPMGXBQegfPtlFlFelm7inKltn08RNIJwx0Uw7Yyxb/ri+7dKtTqJC2fuQ3asYp2syX39/zmU1MUBhFLZBPy9VaxPpCjzr8fCKfQHWBrnslWkuwtqog8uMNvW3uQjKPfSljBC6yDHHYXK3EyNio2tSuki2HhVWlhOYcgYd3K3MuvHQGGHisdegpvF1+eTPwT25nMBEe5eGvTlfyVIq+MMxBBGInWHV2RXEoTEGqvOYulFR5xORb101VoIbsx2ehatEhPMvgKLjzxo5F+XMQbfRsqDaLHaZpmUw8mHqsMnWzu5zHOK2MeReXXKFF7EDLTug/cuoopkKlvHYX1eXe6nav+6MKE+LhrItW+IafWQ6mV6cAoCNtPa47zzCVh4kulHjUvKowYZYeffY2IQzYjcz4v4qkP4fMWV80PoSdafCWc8CH4Vazp9k2HZSzjdWy2vocC0cQAMqckhSWz10gtvM9evhQh10AuMm+2TTQcPBSwuuNKXmzPVnUfUbv0x45/wiYCR2EPaumsoPgZGelen5UZQI+s5OkyqmCDEQPdYYWNbuiL6T20EoSql31TmJkmE8MN/xdqB8c3pt0gYScIZd91dpH0u/ZB6JmsDSwI9ZLykA2RhU7vjwIALnZy4ZlLEOjlyA2z7DhW8DgTGrSDBtwX8X6F65Dq/MtxxuoLi+itwuxxXOl8GgPza0bQ6t0WG/Fhj/9+Y8K7aScT/4sI482G/O/yDjlweXXFq8y/pB5UzLxDg2YMgXkmrFIQ0RkPR93pjaKDBY/DM8ENzp4+mqD7twMv37sgXma1IxFbOWcwIf1Z0TgnmuX3mZgf9kAD+1twqBBxnAN6bXlwHHtKRjdEyBubIakPrcfU3YU1X9SgKkNC4zwfWkbQ0tqQO2s4E+4ojn1/guAPo3z4/msIeaJox6TGf2MuiJodid6FYB9hwai04VEXKZRztMjkt6ZEVlN9FcbF3PH377u9lt4hK0wF7o1HrviqNoMCSLLryaBuE5kHJKkGMkljfJph7DGtZU7GtF47XxPvKCfi67XrxjLEtIIKNxwYITlUPakgI7W140yVqQE3bclhWksm/VjBqK9VIm1DZBsktIUZ4ektKCiM5CBiybZOlR4k5sefU7HHptcMlamUB0Z2DOzzaNiY52xIQp/1V29hJ00gNY6JegJGysaFOIc5tgjRKlExwvnoCBAJY399CaF6puv+SVcrg64/wDrvEulai+TLIKvIc+5YUAAAx66ECiUf4gVoyQkTHKNVW04HzbTv3r4ytyS8kjovit6lr6CsJ9lprtpdCP1wXlaY5QmXigVM56GhHmsI9fK9/4qjCRc4KVPx4+c/poYMYMhx6hlhcyluXQ6rKckXUI5+bwOCcK7qASvjd1pDzmH2T09ST0sheYT6RsK9DVST+NzDagqi56O2BGddtgNYD750avNDOkR0MZc6YIHpD53vzHBW+m+aYHd32aJBoPED17ZDoffvdG/ClIT5mHSUV+I8fKNT7RNkNwvGik/xIDB8jn2IbrTlwahiNOtCs1cQtiiI34TkH9b59GDY0eUzrt6GsUXy4MFPsuti0fow1w8QNwwfej2KRxJZQVuTsCYwCUc48itEumk30ZmDVYOvhkqDHtDADcLilP1xf/g8qCws6OiT5cdQf4LIAH9CjWUzujxHH7Qwe7tzbF586LHwKUCywbjJFm0kFPVVFkGAi4ua/Bm2pnHAa2i7ZfCVGHq5tLTUHq7+JKEvY2229AmDOP4M91Rvtggq+lbckQcKgeaH49Kvfws/PeW79167GcSdWNbwd0Q3VdpN8HFC0DbUhRj9Hwv/+GKNUzMIO5PlI16yI6YxD3jHzF5jBHI9zj4DH6AMtRfbZNxM00PJgDWe8YP6c1JAUGMBHN/nMJZnybsuP05o49EozGZY1TvMYPogtKyJo1gep01M1iT4GX2v5609P7+PhOMnNJHRtbZ+Yijvmx0aeh6LvAWA/4BSh7iW/uUZGeR/BzQ2W4L2gRHTTJp2FOnLcpkFILi96w05WpN93vDyWdv2sjkGjWUScGQcUXC8XWjqtWyMYyGPH1MU9jpxgHwoqj5Qz1ffgGGIB9wYc8feUQG37qk8ItP1KabcoeoGq4bU8h03iuXp1HpqOdO4BbEzhT829IIzjAQLS6z4HFVRh6boJ75wz/CgnfFo4hlCvkGNLqj2D65dvgDKIY73dtMOFvXN9LpnxdOpESydpaLXJX1w8CKwzqyvx5H/hFYczx7k1apav2wMPd/WBVhKcDSwraiYUGBYbKBV1xqmM9HiLI51o/RL4+ktELQGpFdx1ilXCBcN3s1dClqVzivxde+6POLF+Tb61wV9mMlhWLZNVRQnnU98TBvS1ZMjUTjX/vrp7uss5oUMTclRfqiN07H+QTjvqXKuOLmoyS96JalDs4cvP1Q2Hi6RpuTJ+59zwgIZ4lNtKHw+Pygo7ODVvDffn3ixMxIyLUMAo3g72rBydXJsHYnFAGIIFEtgUAs+UCdkocd8Q+IdB96YLtEvv++YTxB5nKRFYZgAXkyj/7jF8i3p6f8xHRpLpOYcoT+Mb0tfW+c287ghZzrR/McdIVONwB69aswVOWpD+wn3PvFZ7G9BZkrAAv+EM/ezUQa7MwTI+asAIgqbxdw27HyWCJXNoqDmIqAjRjrK3MRoE9z1vR3tk2QoexUJP736ADXwu6AvqFkCFliZTZAVtCtyTotkh/oydnUHVHXIlFEqgpi9y3W655WVCZFIBDmCjT0/WROfSHFjkp7qhKf4AScVoYeyOgy3qhXEUtoQ1ORPJvoJARykW70WIFkdh7sl5a6MkXPxfW3Z8on7HvUoD32/GKceyM4zLmLCY8hlbLASq2PMXcQkcsPbIqAyFODEL5MdF2SZ0Mll0KwGptWRozmUP/aAPL1Jok0+sTeuw5oQOk+BuYABRXN17OAjALNm0Aeb3MMvlV2h4tG+Yj+SIzqG/Yo0QlxAVLxIu6QblhqwnWzHTjV19NB3jNyI/r7FZyEyf/7xOgL3wZoXR/24im0KiS7nnNMOjTBDruaksrYBJnNuNndCtJvj6NcKscuCkU/Okq1cpHFTeX6Tw6zGIdVZP8wh9CjtH/i/rtkXDwSW4AUNnOr1VrjJTDPrehV/aRE4sXMjb77isouQXaRJCk6Y6FWUkzKw+9VrmFVm5EbmEcgIKo/pwQhFKEEWq/JAz+8I+Vu2A8EtfvRMjtMIr8SgVkabXCepnOBtpj4NhHjBBRVMxt5d9et53CLhbccKlGxbOIFLhH0Gqje8b4GCjnuryzdBjKZ0S/boF9UHLsZDOpM9gdCKVMv/I57gfwGdvOkBonX9ou1lMwDoisWbLbs9McQEd4Jtk0/P+qmkc01G0PVJC8rvceRctqFbJh/emYHOX86Pg5NPRhEKcTXagXSLI39GXO45fI058vOEYKyyoLxLbNaOdu3ws9ys3Rl1nQ1wEfGJEMZAKb3Bf3nbrcdkU5eKTdmSu4dKcIqTBrrBWf0VHh0afVxl7snUlyBOwsYavhutXQNmc73SKwRBop6KsRUXFXWTtYTK7UPOJbc00UwG93u6m2t7Se35JHQbuvusnl/HjG+GhCy93BSKNvlIEr/UgAwwuoL6Jk10E5Eu1fAoWnkI3UNF9zc/2TnPyDEu0ctABLsiUf9HPNYo+Xnf8AHF8jAPxG+xmlFot0Q1NO9/iHtTeffyQNKzG5sHs721Kaci31nYEoRu3DQzEFWReyqTU1J87mVC1DhRAYTlbxxi0NgB9mbIPnb/N8+7c+Q81AJG5g/47f1gLCxU6iQlqs2YJxXuRYwPuNVRh1i1+NKwXreFXz1e47Fnfcqp7kdgAackwd830uZkQFR7XW+qTzKuYRNXZdbQssN5/yq/dCMCI7Wf16BF2xIkhkTwvxR927Mhv+T4Uon26mAxO+kn7dYAKFaJX0ebEpkSiEN4ymo9QiqIB5qQ2jtwz4+BF5BC58068S8P6b1rbpgY6dSp3F2XiMZtmUljMqn1bA1EGBby+Gpvzggogx1AEEPslfVTpyDu/LZWCfmFeamVfdicm2/5FvmgOwEgae0hfX+gdSZawJa9a02i7/7ZQ0VInvWtKdB4EqbFlV77gfGVSl7HjlFV5UVBiZ99UDNsgZcbZvxb9dLe4Gw6pz2uVXa6q/+byW0ScXFeTL9ElpAk62q36e9JaPnGUFp1T2mVnCDQ1yVErNXFuu6X5TFwd5LQmeG3gZ51xoGCJqUNx+zSSR8X6JZIpmS6R7qhkvnyCY5QM6qxLZTdtyJvgSTmQOiXLqXWBBt07U3YKkEPXglgXanysvs6CaauEv5FQWqiwlDhdBO9LzAYEbN3XWQgwL+lpCAMRZ2Bn08qxgL5+aPf+oo
`pragma protect end_data_block
`pragma protect digest_block
924aa2ea5227a084769c665c349fb364bf89c28d766b9a8016c8156df3ee7e4b
`pragma protect end_digest_block
`pragma protect end_protected
