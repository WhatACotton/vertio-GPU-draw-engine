`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
OQrkl8GKkW8ymWcK5rSs2V2mJloI2q8EZ6mRO2kdlVeIBHADu9HB+GEwHcKXN1WG8VLjJfU5Tuc4LtOMrzY1R4Zk5AriKDMAN/J/1S+2XUZrAGY/weGeesn+OZe7iD8X+2AXyfLGDAjHifvLtpFJrKC7sjjcnHowX0MtOwN/l8dPtHgnX8Lw5RLLPNSFCd7oy1sn3TP38u5a71I6XdYYdfdmZ3CTme/LbHIRk0R1GCObLPZuaN4NotGZ3EfylpUhJ+ADNG6z+OyuQoH7XJ8NMKrqvzT8UVaoHerWwmA67+RKGT6/shT412xjC1vSZ58kJO2mAhShgBJvR6zFzwkE7V+AJfbb4iPefdaEpCd88AM2w7y+ZXqOOoktKuBbdbiPsYdr4WHPISq8TPPO9YBIbBha72HJcNkQ0elqtfWvW8pwAaQoQOlB7t/chRQHJFDKWE6mP/nzqHJFMJLBGlTxpYAJvfS9r+FS6wu83m3fqn7JbxwuiFNTPjzoktlYvaP9BK2ZBIUxlm4CQMKGoMXQfTiXxOkQwCnjT4lvcrg9nSIYwQIZnpFz28u6wm/jXvrMxrE46cBJvqhrh+I0udO8gyQKcnuxyqM82wV0TRNUE8asjV+LHN2GMPBKVPkdhdyikiiWG/AxxhShSbzPt9NOB5SgmyuP9GZGOzLGK+yXTpcEZNwY08o9n+2J81KBRiEIW1N0ZuJ8BzW5gLVFMrC7qzKvEeEFqxdg7VnMBajUPEFjzE6YSrIUOVUqUs75hITSqnGKehRkyKM3griEX1mmwCXxfeyF7V63S6JAp4unj5RyUBFokHzwzr4kmVCnsX/vxue55T+oYSV5UqmhMFg1r6LPnHjOQXVbL9V6XeLCCrI1AhZxTgCxdrG/UVuRoRLGMB+J/v3o7fCpfFCsZ2KdJYb+h+Qy6L9gJu0Tm6uQyZkEzmnSokyiBpgtwTR6jEP2t3wOFi0+GFTlXziPnV8SBvw/n2yCl/5XVheMA3hqLi2owM2iWVMxT7c/707IAIx4TbMR+nCWOvllY+VmWfpto9GEB+abjJZpCjKyyg+mYLbNeuL7tMxOJDZiB7xMuYyHRKaF7yfadbof/jpFS9Cfoe5URS8urWkolO9eCRlnZB7cvuJ6CRCb6MoLx5cvkg6xZjCN9r/wn6Oqx0bVDJJxE3mnJCT3vBTQVBo0RT+PB4rVBOEa+2Y1LmR+p9qYko1usAVJPuy/crBtGpFBw8c+X/h8a+gKyfX4zTA6c6NCWkJ84wLjWfrdfIsvFEK4nx/T3a/yW5/pnbSU8+y8gr8WlDm7vzSjdmPWIkh+vmekdV38nKcbMYOZ4GLYxLhdPpB1KSkQ9Kj+fOD7IMJ8RFxHzu3gzhyvS1DXILWIvuO1WFxUHTqLS12tLk8E94ahMvn3aYKt/tPeDtjAJlSb3bmhY0olkDc4bQ7nDs0gDNyLGP99Y4yYWn+RGBCPEc9cMiewe2Tmx6oW7ZtpuiBaEulGKeV7nk9LPn4077BDnDGwJFtvvyoFtD7811QPlpiIlSfAyjSsDRRXiMaYtaY1YXWb9XeDOF5zmNA+W/+lk9/yv/aUl6HS7Xyp1m7loAMIabpdRlbcBwqy6KTFKw2kNNxdEuRUoE52sf7pxOPSSb2JhqJyHcu5gURCGA+Y2mXmneV8KXgx0pvoem58Kd9Ae7g+7e4aRKf+gJmBliAuhiJFpEugzFj7oUCA8pWSrE7MBaGZZDHbWGYumFuJJavRX7kYGDLg7sb/hdabez8eECM/dir05LCppJTWq3kLuO4yE+tFbfZxVjyjrjRtIyx3W96LpQ==
`pragma protect end_data_block
`pragma protect digest_block
f99291d373682cb02e3d4a78c7f8714a5446ed1fd947f4422e5397d564e79df4
`pragma protect end_digest_block
`pragma protect end_protected
