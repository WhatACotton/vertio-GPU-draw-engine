`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "bd232289599a8f8e7fa4b1762d95cd31"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
RPiktnterlNMmyZKTnvM2BmX+zwXSJmTJNOdr/1p0UHiS7UFVzJ6r+LPDF620yDZdFKHZhXKf7n3yezI1yh+M5TFJYBsYWK6BS1GmiKpwBhBfOAADBl+eGjsGRWT0DCXgV2f8V7vLYkcmMrfx64oxhiPy79jOY7ZSmplilSrEPOL5t+9o0f/mm6gI5bgUkDdxzzYKDLgP/A70//lf8cBYa1B6I7QQyyCnJe0C2goKWGQwNOBYt8SZQl9w6XGrkkqyWH6hf0XNo1Onqg2DGaDeZbHSYwO/8CH0b3jogKPyA12FybbYgQCxZwpOKLCZNFowOXcK5HArAwTjPdB3RM7vSI8Kz70YCqXV4BS8PBSc0SjhGbSz3hS4HQ/iB9ZiX5ewmnwy1sLZNzFatlFGyXhHI7MilRn19eOMWUwq4GEAOeAybT13HqhnSQvwvoA7ynlmg7xYM04oRtEpviglyqPv2ntWnACfKUbgJJa1+oL3ZWpwsConFPvCLaU5gbvqFHX6Z+W6wVz6UoOgAgGyd2nhthGNASdQNa+Y8MO+BvQKcNOKnN1pCV8OfK8xHy0/zNM4Ygm8qu9I3L1KaOpD/koZ1VYfdOeRAQSXKKfOrssR6pm99wlxRLfx8m0TGYJA4+WzrZtdImavVFlCLKcBzZIxw3GrTW9MDeKD+ZT2kTw4rsgkIMAFHHm/dNo3J3/L282CfAhmWjqrH513+ZoPinXad0bLeKbeCAQXFmPx98GQT1yDeQ1igG79pv5vzMhORNL6XpCopYHGI5Zz4g/hzCem3XYV4sJLOPQR9lHxOuuS5kwhL4VbnS3lrSTMK5VSPJZAy8X46sIeAux6b0I0Fy0+yNqzTpRHPkx1YRq0KV/kbMLTDnowyj+sdRqi3NiCd6v5OjwXd3+hjI/1jQbupy6G0v5bw1FBfEiB9U17IdsEdDps56EEA5dZMhzeSSu9q7u/hCyIeSdM+3wBKJOkoatcnaBwCK4V6LkSdeO+r1BPsvtFTwUSyR30ksKp7OkZBESaU2A+Heo9dx9tk9dEfTOguK28BevTsfTdMeflDBjWpL6m9KLYNEbcKA5XH2Q+ZS4qQ+xhMg+LXKaGIvb5lX0lvDQYpCE2bSg13KPWrCAQi576i69wTYeh463UGzxBsRsJXuCAxUNQ4iZ1IHwE+uGpia6+c5SI13iivl477qFhNAmJPR7i6JXFL0xib7Ai7uj0EeBMIP+KDUZPslBdtVKNT9GP3vOyxBzUAr2oaHCSNYnRvAy9GleDHo/R98enDLaDHyC3fgvPLra8PIzlBjh786LnV0QmMkZsDwZrCH3Irdy8PhJ87KluT/Ziz/LuNBZLO8uVVh/s5GNcfSK/FhjwPCBb5ZQdNvsUTmhu0fPnwmV4J/VmuTU3uHISQcSfoMZPY/OGSm2b3FbhjA21NS51kIiygr4atXHvHRmSVDu+TntABbya5kAlC/oul+XBlFg2fO1pn6dRQbLJ2/od71FI2fqFaKMgxU2xnRI21xQkdMkytaz7P4FlawzsaEsb6ISYgVt6t8SSAiH9vCQGLT+pEOzdzBu3+kw9jGThr+3qh4H9Soeaxs+sJ4XkA7KTX/677WvKslVaVaN7xRj12GsZYPL+llivNUXQLfWPle4+F4SRg91FKCIJO05kN2i4IkENQocbt8m4KzUyG+qpZGp91QjJZ6O++Fe6ExepVgFWzimRSmNH51VWeDifOzVxPFNKfB2e/7DXSk39j1qRBghuvtG8kWyvs8ubr6OruTDs7doFtU+UdtWQo2bEg3+dzeUHmy5xIZAEuZDmFxaxLoVceC5gbjKp9EBFJICZbe3nvVUCSwbfEnz0Sor3kXQ4TsJMZ2fvROrFw4R55W+9jsywjPI5GQh1hgTZl5Uggh3Yc8yFl6ozS1HERG/1ADbeFSVF+YrW2KJ6uyPeTeK03hU+z9DZfI8gsJDw1zUByR0CeXmvkWj+r8U3rjsKLDZeEocjRvjMF/BN3kCn9bW8CAmvb8zDsyJz0oQIDkKfMFKkO1ktcyt139cymokvlZDhoRzXGY6dVYNgEBw3CMWyoVn6Yvv3l2HYwJz7uhk39U8DCi4a3d2clqeYi6mPPBc5r+ideA2+4UfLmHpnjImgyL4PatTWNmZOZSD3Jb3poNQhZGVOo1H56ZAM8MCiobTqKCW9C6YgNU6MiZnOBap/fd3XhWUCQeOXLaSMfY/BjcrwOAp15AuBxstd2bnuSrwB2w4urPWiCD4GYKnnnivGegqs/GQchvmDqn+xEPv9L5pzBpJeTWYQ8gOkFY6dRSDudMmQsgrpEAAHuGkaZZnnLxjPjSWJQvkS26aLUoiNLV0HXMB06UGL2fLS4/5LD8iYYA94+xTE0ApQlqt24s+7vd7EpsFuwk1KCRgrNSoa/NYQe+7u82ViV/YAj1rfpezC7QvLA1r6o2Wl7eKUgKt9OPGFIA3r7l0CFQsNUvAl/dgzGG8vLwyuI+f4iTdBpRnlmZzr7U8aFCoss3RiQ90+hJpeRlfy0jb5vA2VxaCqDZUtXRlZIJKhfKfpDsytV+Y/Qjnr/9too5RQmf3oJnQDBdprOX2r1W0z9fdoW9NQnSEJVmzJTF1lfN9jH08SOjHb0sdbuyktG4BWZeF6USv7lK8XD+jEys2pz5+tJO9D4BbCxZmqWrgVNdJv9l3KmcYc0aypTe2I6++QEZcmytYZtt+kZlwgF7v6HNJ/KE7B0qDZMdOBFDvQ7wuDz4E7kSs++lJEI6XTaIfXRfzTKnfz/89LoYAysy6vzO7R7WDRX8lLLlp3oI5Jjbdmh7lWcsODJceE5y/ipvLBKX/snB+FYydKnrJoS9cDrk/apOymcfRAKEJstfYTy8vYAiVmDUF5ilTTGA4qafnZle9DByQzWkvqhwKI65NX5rgODAT7Yz2TtAHqI4tZQzvdiCesHFaVdZ49xY2D1FST6F7rbGT35qvex1L4c+hQoBwBBpRgDuyg5pdsXdwPANtIuewSwxb57SE7s1uKGbBTnY0EK3LYqDS84K+HP2jPjOS2gvRpf9Iz1T920ONpFDZphUGdPLaquy97EDCFkK3UIW3D6aVQhJ6RvFh5DAXUsEg00lb9VRPTRG/7PbaE8+jCvkQRuo6Lzy52EScJ9XMVKdUFJ+vaJMqZxfBH++dbJhuPAH/OwPUnA1OMoJPHmfTY2B0xYVfLSQCUb+h5PHfbWZl4G1PSG1ilSflg978W1KTr7JpCeT6qDrrIqUGCYgVVrSrlCS5hYVPxjMwGYqsOctqj+JmBesm3G1aaS0k0qlSOK6uYNuof6Qv40shcH6tBzcG46J1xrtgCCA7/blfDImFoyOP3M43UPGwJxNhbk7v7ykEEQtMV4TRM3d/XfrKUI6hPtwVbrj+OtG9RgqsIRsEidyoAvlogWPsPxqsvn8Bp4yh092z9AzrihIFgx2qTCDid0FkBW+H9J5IyallKkKt/3Yn0kdE5iFkCbMEvawd/Izp9dXv/ls=
`pragma protect end_data_block
`pragma protect digest_block
9e3f92ed3028c783efd5fbf34cc21db235bd860a3e8f86f01e7eea8300438d5b
`pragma protect end_digest_block
`pragma protect end_protected
