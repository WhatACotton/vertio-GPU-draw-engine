`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 15424)
`pragma protect data_block
jq8BQjV5gWoU6ZCTqUaB3uBZdpcyqKUX0WHs0ZwL8VLhvyRuVXHuQXGgGWrne59oX9gTNofFbvSH3iA4XaN9Zny5f+tWzrHPQ8bi83jWDdVdTD1KrCnuj6SwlqE4EDjAuro/nW3v5nB1/6NVktijtIUskGjKNXm1Is5eQFMVeofSFk59Wtfswkm2xGaqlKUh5HbcnJn68pV6Kpw690Pur6x/qqTEDNlGlk+44/NLBMsZkwgfYEchXK1ubwc9UlwE6XEDvKK0I+07ke08kGpqTQzdOyG4d18vce3oIZNeecC86lYvjvEvE629QMKHn7BzahlbiV+qJC75IVYH+Ng6rWbzNQ4OprcxkH1wQuI+H9NDwYrXF0801Sglwi7JCc2KoH32NOI/iTqFjAvyyMfQXJiS/7ZKUvh/c9blSXRwaZ5wo+6JKsDFnJJv8ScfRGK8EClFQtWUg8qCAJ8hevdT+WBt311NTl80Ayu+5yn6G3zld/yKqwKkmgfYwDR53AldDmxFp2A0mXChfAKR4fG9Ldyy8JtADw+BlAfTpnFKXAiNG6oDyRKEmDZZOPTSL++IT+BvT3L/IDyjgMkdVAPhpaSQDnGd/1n6QrOtwm2aVXs5H8vyS/HEy1m+AkxBt1w408Kvs0/oJXKb0RlqEITLJCB8/6nNWmH2bWbN/pEctVfCyx1ScSmOSX4OvMEMNJm9b97WDti4hUqznNgku1f8zkc81gP3BACgyNEIIeY+4mgJXb1KOkZL52M1l4scDMu4LKee2DUezmwZhb/ibqi/uf94txwqgQI190wMg4x65ORxNRWHTE4gIrlqKxZ7XG5gp8gxg7IiJ0kP8H0cXRHmB2IbDZv4Dg+jZs0MVTw1tJKJKQs+PQ8saZ9SsfDuWDsCHjOf0v1rk9dX8GFI4J/baERyhsAAFGGSiRGySJFgH2rWz8rYHNPuiYFGq3Y5RKiPrkgK6cX3xksULs9FqLOWdLYepoBLcJcvOpoYvTIeutwWcuxnxXMmz09n527fBS39lxONXUmP49PQQI1h6EqukZSL0ZttTCXy1xiLY99SMfon/myPgSZ2usFS9+p2cTOdErYu65Uxx+NGFoI2V6vCoqCbL05C01B5vuN1FlAfxKqh2liLDA/ieaC2f0s0CQmqdC7Ge0Ua6pTGv8Psi+t15p1phiUXFmsYVlvNVR0c+/QQBZykSHGc20YIY0p0PO8tqJhDWoKZPH4DzUAnX9bGnzc5ADV9y0kKqx0sYMyHiGH69Onp19WyUaaQ7t3RbFoT91DB7fH389jgW/+crQ/lU1zPnFhARd0bw9Ebn7dz5qU1Eo3vvQgzfsPC58ebUEIKAvAlpXV0aiaRCPUH/WMaU0IZ4e82c0BT1MKG77clttFkGeWdVdsq3FikXJ6DVCg1HHcrPUwYI4CNOzK2Z6TWpxJcHwCdirJrHBHyLQRql0JbqkDzlVPTB+YjbK/p1/RZqmn2NSOh2fi6zJvlvR7qejwQAzj1bG4v3aPCOfr1mZ62j5XjBvZ1lsVGc6n/cvURgoz02SbMejC93Js4m1bQW/Qo0Ro6lq+JVqg4//meuwedDkEe78UxLDBPwspV3qSExpD7vXzzVfvo50s/FmRIfBJXZ1ezTmp9rBE12x+Skpc9QFqtrsu5jO7hp2H5TMxHB3jGCoY/RNroVvk+J9EDmDfY2MS53bvgfVgqGw7+inE39H6zHdecPFnymDQpT2cpHass4rEkd068jC+gb5rSBBxNdDSt8wEI5j8aOxDUjX+TthIjGIMcMbdg3ZIvw6C9DMwVF2HMRtsx8CBA75yQ6gLPs6vGGK9AA3bmyV7pJ49rPFF1BV9Itv4OejLBpDctubWByvnxfGPSTT1X5LyoHSwjZsuwy56c3Blybzu74GAV1uvx4PmDnXZnU13+RjxeOvvLEcd8a6Cvt+ADI6W80mGmJHLcwYYeSwK+JQEyo+oCkBmyQqgQj1QIxKaHsl6zimn1jjqxKykJm+tJjIJaz4k8S/E/jU5pq0tZwpkC9MRuKzBfr0eaj6Twza+Td1XoO6hZruafS4tl9Lqnf83rtBccN1pOknWL5ieqHhPJEsKqZg024yzN7K7csJw7Geo/1ugbwVIZ9atcBLKWi6J2cugtHgctknqIZdBFEWDLT+qPqxzK1hTRIFYc3FDbZOZ+XnQstfgh+P9Enraakqa/hhSdHbc07ufLUpaDN2WJ6z98miSyBRX/GiFwZ7w+U+VCLmqE1JwIwhunnTvKl1k6m4ngCmw1b0wndG3feToTQSO+/NDgtzvm7W/vw0zFPHz9sWS0oQngD94zbJsBQ+vGQ/Rs+8rWzeKg0YEtbmb/p1aDOgS5o3mMsfAB2IJbPwiY6G+xLhLhx6EkNmCEgxKGg0k1rVLnfID23CuB38fuqJD3731aMotr7Z42sQXC7XnsZiNpMXJRQwZU2zrB182VBoAXdq578j5iKRL6XXOKnE2CBWoAOoxHyi+Lr8Pbfq8Spm6PWilwh+lTaKNjaTrtrk9pu+R4fEj4QPryhnZPwurLRI7wiw2JdjhK6SUUqzDm83VfDDf/5CylynI81i4sXBKwK4locOAooFJoolAbOKDA0i+VO0hbYHulf7cKwvFHJy0WC+LsU0mVWzwMxE37RMeaCgPenxVn78W315T3nHPTY4m9r7IZjXkoAmqFjaOM4tds35HiZ6V3yhdqV7wf8qLeMF3JBe15S3pKvGIK326+EKqf6zAPBNEsLu4VsSTSF/HGcwGwScKGRs/wQrT3WRbS3njz3jjU1quvbqLggbM/JctPHJy7QvB+qXW02OjIenY2JTrQPz5DxuNm7W5KSuYeIz5xKht30epUDHytoGnaS8Z/TFRPPcMGNrhcdA7+4E2wh2seR+abz3EW2J4WlgW+hXQXbxRec0FcA8tllXoXVchdDwOSCTPMwprCE13coG052mJR89ObHEO8jpaywTSG8CqYtpYYxOuUrIRcMil0RIp01YRaDPlYblOH0weXR2tWYpAPXlmB5xruwnU6J40OsU/NjqlkKoWfQUDm/t71DZNQbFPHD44mdjBIiCSoUaoRt51VMM3+Blxy9MebeFK8z4v+QR1BLdL3A34MHhoCU+rKCXGonHGGTfJw/PF6lxU2nFQuGw27UhO3r+Mba8md1n0lnxZG0WH0uuWNll73y4glUC5E64qCkU6wpH/hJ2poHUXc41Nvelik5Tx9dj6pIxJNJ8sl4x4l7uEJJQF73AHNUCR6QgkTHvxJUfsPKs/SeZ/i1L+hppQQGd4oKJ1JTxpuZLxaePjiQ2kLgrm4ffvd5RSSGT/sxbWbOaZ+AH5HEyJ1rFRxlexu8HeWcaDOahCXjmffvXXXmQmI9wq0cfkqSlU2tPuW3UFFIs1QgYkMvn36zZ9T8TSaF+GXv8oE20s+pjOaKub7AlPL8Km+rjAyDptw/8arNjQMiPhSBKYPyS1pVKKZ70/tiAjpz3f2KK5JUxRHyaxHyspCh325VJhCET+CotNGERdFYYPW15hArOKix6XbY1BTU78EoJbgkZXvGACgCBvBGal1Zn+3Zk7Tu4095SrdOCz1X5O49la73BcloqSXdiKqq34rLeiPIXP1F5vc3GGfU1M2lECpH1z3ULUkpvzgBEERqSzQP/8BaXfZ/h9NYXB/yKkLAohZp3JdFUYfcBU05tEvmPJKG9760QqpXyxBlCoF56fXAAmT7xe8XzLW+f/WWW6vGvN9dBEqTqR11RAaGN2ss4Rxqs01C/D85OoBzksR7cMpt+giZH8z/SThXVYyj8lDEC4e24vddgvJ//j0NgXyT9zgVdI2sWLv870I6pR7SxqM6Ykrpc0EHlsfpq0bcfq3Fs5h//HjmZX99MIEvXwVEwN+MWflK5p/cWAZeRKXe/1PoTBFZlWVi91j9S2CuSSCUyIAs5hD4Ludl4DehEMcHo2Sf+r1Xm3mjAA3tJy+Eyq6CzNc9hBZaIeCLY3HvqHC5wHYCXWqozEv61WYKJFOHRSwjt8jMfSlfH1shFnRXt7g0PQpdCWD8IbNcDnCbs4Ar8PztTFLKwYWF83DtAU25emym4bdZvmHzZLaXi0fzMwwYfMd+41/yX6zxc+qqTmhSLDj/OYygPpZ5tlElQ52r3tfV17r2b3793zZCYOCX8yGo+wNv/qCsREiYnmzzzdogGCnMgVDfwUqRV3czy+qH6oPIHj2e+Xx1bpKGCAucscHSmYnzpc8PBEpdCTeUSmmP4P4CFfR0lbOgiQMq1mlQ/FbgTPWO0tQhNGPcmUfWebi6upO0Y0SBzFmXqfLAXsk/6DJ33QadQ75TufibHHOPhCp/K4lM7Q14k5k7rkQjgkybsBZONYRXitO51CybOEICUPrvuKLDiY15dhACKD4RQ+nzBOX9zCWEIlPy3yfEgamewmzC5igpg7SuiSqN7cks6snHTqI6JHC5YF02xvipRoj2iTeEHJf4vicx4Z4A8oMv8TqWd1iPlqmp0xmhT9cZbO5gtIKbSgn3UxRa+PJUy1us48w5jZUps00mwn38zCKEv/fk4VluZ+ol9+f0J+QDm959dnSwb/klBZo5itfVWwQenbvYNXzGehasg3E81LTQ0+kRsHzGNjl2SUqv0p8wO7JNSfyMLhHsb9my8N+G9jU05SIAzD8//0EO60opB1Rz5DHzBuTcCfzG2zd8Uc+RoArtpOJfN0AW/GGBKIH6smCgv+/1B6yqdZT9rrjvkhEHDmxLAXuekFmm+auSHaEEahSW3iTzaNlzxJ2ZLKVKyQmD+KcDP/V0RHC+fEiY1LbqNyrio8Gmyl6fSmceVlhsCMIIc/hhH9gEs/lQONYF8hNVNYhLfMo748HMenQibtUGA9d0+xFzMxyzRKSQw9HyiGv5BhZGdgzGxbvnV3o8041yx65y4lpdVf/VxhjnE/htyRrYS3dSLScXVPzO5V1H9BnPlGGTrpXLSO4ncyuCgQ9JRANjAD/av5PCpU8Ce6Tl56Jq91iBVCYlMycmH1jylLr7Y5PvhkS1Y3xyFDONATNqyjbemXDlCV9zQluxhzwLmbU2TxPFafh0MpFGinJdw1x00cA88DvbMqggPD2fhkaEPJMuexN9rgeEmF/85oFCUnXbBF8mA/WVzRsQNTJbm1trcapiJlXx52M7oO0/1+MMrWAXr2pWJTEtG3vVpVvq8knhKL2MIwn2E0moHOXt7FyR87qXHR7j7itzUPnTbu6dFVSxxTJyxRVGaI8KMYr9WA6FGi7TIOgZv9nkswr6WlEjO2Np10N5ZMUxjvRUc6fY9UizR6M1fPeCyKR3GfEMwuH257GjUFKrUgHgRZTuA03GmnFW8EXOq8qAibOYxbG1rHQ7CEOKsD7exibVKElbCjjMlrtcx/TtyiPnMbTpjQr0h29nfQEg2JbzvghE5FmnkBATz7PCxrdbThlGGyiazKiIU/5Q170AsOu3SfSHWiRy1EhgKtrcv7ycBmBg37CrNr5VhAoVV28T91JY1fHnM+bD5WmGaCHG5uX+gKYNetUXXaiXbNlSPN/6dQz5Pq/NgDGxRI5vUioUCC2kCBeBwv7jTtsjbme5IlVfK8E0bi3KiL5x652XqUkniZ0LmgSZ0jwNURnqW18ElgIoi0z01TzC0s5sYUQJWUbFGoorLTM0af49cCW2jBI7sNLRsp6Dy8f5jFzIALLPsIQbF57Y9dx01tgWCUqvYXLF1AnQsELXQvBAR6J8RvaZo0mnRwtjnHclLEnyPlq410pSQl5QqLmoIYufTIGT+fmbeor0M/G84UAfq2G85g3xYyVmtpFWMooZ9KyMupzH+OaGSghDJihFZnJ2u+Hyf3WP7GXCFqFh2io1Mg9o2Oe9iu6fSQOhJZGfFrjfPkIteNlIqyZ2SzPQLZsxybFYFDM0aYhd0NSZ8hK2J5jq+DIA1QJ+80ob6DP8VDCtfCXzaC4ErNIYKHKNOQ4bjzyDtylOy/uxQv3cDCSjKbg9Ze6vJwwVKAFGjpIOMDXZij3nBPZRiWpTKkRLdWM7s/jf1DYdlwDhKOboe1qXMNjH2AEN0QG3UIHUhLTC035rXsdpadpDYRS/g4KsGxMyqcJVkob61Bfm0LL7vaO1qTSn/Zewiym4GMW4vpLicXaHlTb2lJ1hnyQWgSx+pcVF4wTM6WzLeEDjlzyHpyrooMWRhXLZnWd1QDw5v2sJwZ4aYn98IPnYZEsRHAmiJzudppwfw7ftzbWJnDFoQeEakX4TsQJFtdyHDxCkT2kIqOhRqrzT8CAfUvfn1ZXqtrroblAv9cpAq19xmqm4J9acl4b9LLFXn4cdG8uTYKTmVMIM0rqwAY9hfUw8VbmGemg7RyWK6g7Iv5Ls9jMeNoAgPporo1BZtxTWPPwaJshUQZfQ1SACbwMTUnS2rCqwuw3ZOs4GBqajKspHAlPRIQbczPGD/Yltm0gFPgXwcVwLRE9rVyjWoC0QCH1Vs/tHOCQOmp4ToDOA3K67j5YvsdMLjO84zFaKY96DYrky3mks1d9PHHIICSANJwNn/Ivau2qMTs0HDFWnWmmN4Ib0AYjXjNUNodzWa5bmDh+ruBk0inq7MRkJqe3Lx7xgJcuPT9RU78u/CiCvh7AnRouFTu7ECGPgSZG0yzw2iC4WOqBzCOycO7MWXFLNtxMNZJqaGg+Z8s6Od+EHU/lkHoXBgbQVqhDi2dLHSfPHPtUZ7zXtI1FSG58olc/rzieZxAul06A1NAfXZMWE7Ffkq+T6PjH8Hj3XdFgLpE1KqP70QMPCL/FlWXTwVJnMFixZilCbuO2jSb0eRKfw1gv6kJ7uShKVIbP5f26xmuFZrakO6ARz5eVeMN2KMuefBErRwQROQjN8EpSlaL1F1g5GgzH7bFt36/lDcTQyg6m3uuYHrclM5r+pQpVSQdmNEOle14RqTA1bVLn405COxs2ZgZ2IjBwVLGrrdogZlza7yjfsbEHB9gQi9nXO407TmBTDKJIlcYHgdxOEIYqskdW1s1RPQasNjrmCX1rwvdu1KJv3EezhMfvC6KCpEskUn8k/NTSrjtdzDqJOaUB12JiG3qU82i7nV6jldR8/ZLFaCHMGocutGfw9wUKF3yrESOYDcBr+G+q+2HjRmPv2beLblj3+Oz5p7PpczhH0NfA3xnsz+3vcZLXo0axbWDrdvydK+BU6p0LKHr7KCH4YZI5knsl27Koupzjndnkgi6Ji7ZyRaU1RwM4N8tYxX+lV981/UKHDZumj9mil5ihWwvSmVqAijbSB35yun6X/SUK+jInyJ5luKbYxFJgvzB4G/WuopRpmkTlhWBmj3t2iDz7AYY3LQAdbho1w0fgbxNZmu6ZMfTi+7B1UHDlBIAZHeD6hezJZRZeZuwpJuk8b/xz8c2gSFTPeG3hZZx8wXQFOKqwmJI1G+MLQrVMqnVqyJtXhw7Iag0n/h0bbUEGCk+0nc0mUvt+3gien/u9nluh3nt1Hjv2a0aiNz59jd1N5d+0MFwABkhQq06+oWH77v4to3daAuFG/W0EF8RXYq95Nm8ywc3LCYBqVpWz3bkMLPte89GTSEI38wMxd+QaANCP7zK9C5mZSccyACWJEEVUPFK/Mrycj5jchmPaxJzJVSpfyfIxQ6owSmTxtOIyuk4n5gINHXRc1Y7zx5QX5A82k0uA6f5Wpw8PYalVUlJzIBiCCe9ZF3pPNcVBEdNr47NpmTrdeHl4U3lQ3BnThuy9kIufwH57xT31s8s1vejPoa1jaAAlRUs4ZVl5frJILzklTjSb2zby++dwEYRWym5zGLNJE17UX1/bbhW7VIwkwx/XWYUFeRx5bjpmDYYK6/S3mFY8v61XIPVqvO5Bwa/UcBN1L0tZIYvEZvZEkfM2Wp6IU9EQgiTCWBCSl7Uhpgg+qFA8Sbn4W26PRpfB/kFtOp6eZjNtziZeCerb+fq+hBiM0tYaNHgt6rb9OulNiHM+qt2XPTEL6LEZtcz4SbeZKxNqBGrU/fokILX1leMNanYKenMYl9nAadiu9OTHOQnYawFtwUuS4dVVNUV4WsdDsa/oH4CR3QtpU0ScsSwH7hCCV/zDExUXHesMkRAJ9tESvTCegN6S98y/BeCfzsMFLEMD7PVXFGkS3HqlyM4yNETbcLQG7MkZ+BYPY4XAbTUKhzLN2xYgiPp+eJPIlDNYWRnZnUi8kGe6PZb+2N9wGVfO3M3y60M3gvxdOs248fpZ0ADbfpTeFLokAa/86qMcn9fPvNDwkgmk7eB0cN610hfmxkN0uDYRKtFw8fYB53apk618xbhsKocApwOpzidM1oIp5jyVXex2Wn6D+9i/rOuYI7GYT5DS6oeX1jI4lZBbSc03IR5KaWkGcQwYBp0AzdPik9+sae84euochA4zRisKCX273kDYACVYjdZOXbgUvVa2DOel54mPTClHHTVA5kH6d8zRqaNO4ZaVqt3Ky64LWBQAw/znhgiKj+kD+bKqIdCJ/zS7mZ1OOHRQsCWD4n1H3Zw+zf5pP7N4MBbhRFsIvezRAT2yaaglSI8nHkDTkGmBqCH+WrAZDfd0F2AYaNs93rCVWjaUvzqtGljdfBwXjxTacp0KkONx+0lcH+VN0kI8nZAK6jMmNNom9sufUrkIOuCZeCh+xDcOfx1eg8XO3Ko0tRlOLApvsgWhuy3//datuTBEiBRdSPOTfpAngUN4uSSCC47LCwKhShbwxRTbsd7S1K0NRR3P7bTI/Xer6coi4ysiufGye2sstuzv2p5M77l9f11grftd/r2L0F54XD3Dd148DvcZ6ZAqsuPJwHCtOhyP1UqS+4X0mPb4bxVxp/1+tD4jR25Q58S85N5I6TyCXfl7wUz4iyGCh8ZbiB6hIG6KZT/djZiV+ZXRhY6AsnnRvHr7sBvzw9AIEs52f0WwhGYm7LwPkpvj9ohzRwK8NT3qDPXioZMDHxJ+HdFsP5KI5d3SFpZaqNrh6XOho9DB3uAJFDUFLZB5DKG58LTPAqjuOno5efT3uYySghhgxYhnk6cyYijCg60d/UyLSrkBW/oHLWn8n0QbnNtAtUftTo9hAVPjEBh6itSNUhlKLOhYOKj52HIY9EB1p1VfI7rPR13vQA7vzgetx/xUFxzMflI8TKK/jLDtqPLZ0HeITwKRS3kXMCPP10K/o/TMdWquFlt5sytzT9Hty4gXdTP+NytLLDAYnsOFIMMrx1b21acdwHsDT6ISkQkohcLIsm7EfjacF7cePb1CC7eAY9WEYfDTJia4dEiVugAjsW7gPq4BD+LP03YI+58AXVrdQCFkTNXmo5H8+IGaUv9IoF41GdKyvs2SQBREOTpqgGMulqX5z2YI1xxNTVThT1miZ0DMkfcije/JW8FxTt0QVwpGeBpUN9l9iLOeJkWceth7rm20sQUYW+Y2DeDgL/x6SlwEkYVPAGmFm4MrOu+xrFKQTHdlIXJxwYW686GsM7nF4CmoJOaNdMgdSVCqlixZgCYpRZ3lT5pROB11p7JSo6LO9w7nM85xCCnB7U/MIdO0ravXR/RoTfJywSesKgVJ9wFzux3Dfpuu7/HAp6E6IDSCvAjjS9NzhxAYOu9FbEXiQV+aGzYCSlz7X7JXbXg9dkjuKb58MTtUJcLpsS0rU7+k9EIvnoFcZ3PJxsVA9TSFJsvcJRCZpaYytkvrihFzMw8QdFEmXRPHSDnKAW28E5mmGGBv26NnE3ZQdf0lwhyDL0TEVDtQAixd1kRJ6Xr8W3UVf+rpKf/wyi601g5wcoTbyUZPVsAg8q/9JgcTbaC6z5nqNbtFGY+i4f57krHIqxTAP4upFGAdub+ghif2zKZccmtKaNOCYs2ZhYpUPwdbgepREqJHb9s5U/qqkrS2cz5aiO2F9nuCuuZYrzWZBuYcoEbxR3fyAmViN4c6GpIlALcLgnkqDHPJzACvrHWojyOPVdtTe6cXzIJi7LV2rS9BGZnEhVBKEU4jV099MbcT+JS+rncKr/pNnhvXoEC2cXB1jtYZQYMjCb1s9eAdUtQRcH5tiJ6Ck8OjLl8ql4D9TVuqMbBQaykwfAoGv6ZRjY2HAqVJZo4seN4SG2STFzYaaQpFhPOPmFy+X7SZFfQkywkBNDPsdJIYB7N3fLy7bQJ8cxijYBAaQaK9YeA7JZocAGoJEIfbNHCC8eBZeEMMOGw7NDIPhdg8T+o9parMTrsKBXKQrrD2WuqXTPQk+WvYzsMV9mS5nbB+WnU9GFfBCyBeXgxLXxe+AjawCAAU8nBdJkuFyhGQtWOm129oFqYxKGWEQ9lpKmxcmntsaVsYxRqPvQnU79mmUcwHWPXTEveujwocd73K/Pi0StaMIS/iOZO0keoJkMBug/s/2fH0JJNc+iR+Q5Hh4o+n5ukZHZt5EnExyPLifGlAoh5mqK9qYRxTvXNZGahM2abGKUYepq0B8w9zgILnde/X66hu6xiMRpU9Ei4+vdxtYjt8dXsN2mW7dGGYS8NY5H7DVbaIEKbuiF6IdecsTWDlHrkwr16DUL1O/1tTvwbXknY5/C6CW7LgIlKS2dJSOkIjj2k4Xfo7xC1ycDAb9e1z53MMi9wNoEDWh9wX7NDYDcyAj0RZNYtnaPAmWYIJEs7tcaLmEACTOg2XZL67an5+rdZxna8axcsiCZ7FRVFhhLv9bgwXvEt8qzrCDlbhNiMEWBSsIZnfs76KnGKLfkFF1pK44qzrBfje88ZVnJVf686DP+2M96ReOGympyd9Zjmr92M7ny8/vIfv+AJXuKvSzlYPGZsZhwJwRmd8ODOwVFDtHZZTTQWxjSuAl7i5kMnDMC9wzJYDHhXvoFIqLoE7y3WAuTZfK3a6b2Tl/ICjek8pQyXyflzD5pKBDxxwTl+QQEItfjf1rJLx/kdvxrLExs5jJdTLUhygYqYRU4grIAh6ne9kSryzvUCbJJ4U7mwW7OO9q+hBLCag6FkmnEO9K37XAFKQlAxCTQB7h5BRmhwRUa2h531st15M+pH/NZbXbWjO63WDaLdgh7vrGshcEZncfvaxx4U0OPBvb2992HqdQ0RDYIDsadnh0gtUBD9L/r00JPMDIq+ZwFfewf5XBGMnj1B/NBv1rCsRSx3CS/4L5G3SoqeRAG09beD4ArsoZFN5HOeLNStZSUPNAh5AQTd4xW+Z7h7ftCQQXcnG3J5a1t/B1kDZ/rd3HyEKirzq28y2G6FBy4OLGghJr6gyAiP9sUNHOUYYLELdBav0U8++3sv//5W27O764sWGiiPvNzJPbAhJjT4g1N/i8c5QtMZRUoae+O/C8iBaFT5WFU6kUJ/fLnFBPDhrzL34+cGn1vlYUqSBMYYK5SL2smMNjaUghyIQmbqF5fL2KAmIYfnpJsbPeB7qiL0ljEZFHtAQrwFdCoW5qKxtyN5ChurWa0maqvmeHY7KV2MQmq7pdF/Zrgea8Ru/5Vwz/b91q3wj68uOSzpUjz8nFhWv3vnmgWIVu5sWjna/TzA1YkqdKTZcQi0RgiSLXhWG2DeMeUG+bIgjl4iytfGc+ctspQw1FHNLeWVBhTzx1ogjJHWRtATZbHbcJ9Lw6Wr6VImz6kWedRZjlMAFpgvSzmbdcPg1TSBMfKybkUujfN5pI5XZv/vvA5+80j/Be5613RSq19lgfTI5ZWQ7O4OCUprSA7wiw39VTbyEIvfkmftZGfl9fMUpCjmOPGQ0UWO1BcG+K/OMQgzK3kbHbsL2oyU4Oo/KMqBncduXuFysHsh8FMp8pC4WmYUAHaKi0E+CknvEW995NwbXbTD0y3CFkVZ+mY/rwDBrNDKbg7meHz2eJ/kp1Z/1F3wXYuOni+t2wVV6bIcfL1vD+72XuTiPXWHrhH5BqgQaUV4JAEdXVbQqnXjGhMFH0Xjj6oe+a2F/TTN7RxXR1F92MX5L1kpCUQ+cmepooYrTpBu4u4qK4M8GWVPILS/Nd/Vb9/DsykeRB7vT1R5/o0iJcY6bHvUO1o2gXBwXalyfGt0aJesPB1SuTfCDH/2eIR5SM9WP5V/VyD+NMPjNklNLlH0QScXOkhhgSJtleGEmzktR2h7oXgmi6fNp1PvKkMSQKdHMn4XfEmJVT15TQb8f8P+OSV2bIlCOUEzPNTSNKAop9tFRJE4l7kJswjF6JChAK/oA0V3qxUJoDaFyqNsyPWtcVM+aX/ACaUyqtSMPyRVDrV/0Hpp+0fjbe0ZFZ+d1T6Vp3muICLpX05d2zGkX0O8rdCttlGkzYwSsKi73yNG98XEIi/PIwn3ljx7q92LsgqF/PRUZWF2EKgXgQvQSrExJyTZ/1ODRjuxE0M70nSl/Tu9LMsT43dAK4quNM94wftmUYBNOzEmq6x5UMx93Dt/ti/Wq4LI5N6tFMz/Oc10keNB0KagNqyfXlf4M+ru0eR9CBUYfeOMRhcP7U8DcFKS2CXTtW7oOp57lhy2qIVYZnpGN8W8mzoHG9ltUK6WmHYXjgogwxUxGOjY+yR73hix9s4SsLkS3YtnwWwtaIk//63C1pGlWtEznWqR/MYnLJJGJGhmYLcCXavF9hbJuGtTiBcYh1g5K6MU6euTX3mUfpH/RwWIg2mQceHkWQEmsFhu+Hv5+UXt/0yO2Xno256LcNnfg3Nmi/NSwzo+nRF27lUH8tegbqAFEPmb4LM4AmBh6P0VTcDfy0S9E4nZ0QYzSB3m1yT4lZydSVT0A7N8pMd9/7uugeSRrFIDMAsKmx8S/M5daDumJGwBQaQxTbGxmQwkmMoV1qIeaTH8hentqYZjkfYFZbiIQjODpsVP1flXghOAusEXPQB0kjqAiqg/4heGpewBbEOjKofI8NC/95qBs4NlTl0kqE4zF7I2VcdUZPUwAsssTphQUZUMXmvHcRoPizQxbSyIvkQAuJPOT2YrDdAZSYQBBHMvugkYs4UdRMtpM/C7Yfeg4zlTvv9Ig3VioF5wAi9O35IgFk9mNYWwu5vCw93W1TwCVQ+YG3pVG14zpOYsIyG/kuTPXmkc3V8BiztUceLl19FwQ55jL8tGQAehnEYqtQZ6Vz2MxqetrLlG6amRNvnuwQ01Ecnuz5Ma1NQ7EJkYSeBrhmrMFvpjefsweJXmktAZ2WJqRAYA4gRIak4jMxwJ0Afx8HR3jv4qqffD35Afhsftz4t9nkzVkw6/bGOevHqZYE/kEVwXDE5AzENUkEdi9chaDK6hzn229MFWoLWR+5EJJMFRRKRCo4MjcBMTCSnWIqvxB9AdQR4VFR94edWkH6gVrEeunI05jCtHXyswxi397/Q4DImHOicK9iBGO+E+8OuxC7Ac9sXWlIPLMtrExbC2O7obVpfF86rCFoLCQnZE28UIq3apvD1ncf9Ewc4VOh2FypRf+mKrYEX42fx9qGmZ/wpXZqVtVMhg8Wl7f+NMfS/imSuZzFjGv3osWVTKcKbKytV3jYjiqbA17LMrKtVysvEalgj89l6A6VFbPAEV4OgQHc3KMbgu1ws6tI4MKf6NPctQl8L90W/GJQaBHK44HgQ3tRdT3ydxg6OyIvgzVNbJj3akHv+IXkhbX+ZkUIql1bUvaY9RvsATRU9z75fYe+8k+C2XmDK5D3sJC0Ogx+Yq5NatxbLS21rM1laqMo5b32qeOdD+mluOm9QviBlBcEEHDXj9DXdIw1byLgmcVoMyTML+j5okaHFUe8o/4fXwfdPbKmfTXZnZdhCacPux2c/97PTUHzR6E1F02lsEL5E+MfoZJwVXAWIaOBikNqHyV5/4IQKmkh9QVdETm8bXugXf0BOKPBK/azfwoNa0FYcxMBrZAESC+lXoE3dxwYdI1cYzkW5SOkBVi6IRf/CEQs4eG7ZmJ5jwn8O7DfpZirRpALRPGu/blMG/Pwcak778sY2bDl+Q4CzHZojLKSdjmzhUg1TCBp00GfbXDzbTzDem2a5a1Q+PIsKIjGrKyA7PGzNErh/5x0Gb46CPJ6K+phjvnZkZNk9bosW9u3e85XUZqe4KH4rMcTI2DDmA846XQ5FGIgh5KF5PGmgW96n/2/Pltu09gibwSK1vYazXWjOyA/Nfy6vWZJxI21yczFUZ43+Z9ama9O++fOHUAP2ac/sb+sWozYKNDu4NqkiNuxwwkw4dw2diwxMUg1EnMgSigw/5lk9h5xUK9gRGvAr/NjscKJ+TNN88+h6pWxXmgAYpEDItl99bJ7Lp78WGXaM8dQzFozSojtME97zh1eOXPtzDLX/AL9CxMWzbjQhAoKeX3sjyhkzMQbFcXz9MmZoiSO4adAdrVManDjiSkjO+GYxoDWbvfUfbAsJh/W8EBv+YpYhQzjmil8+ATYl24F2AlT66GFm07FSDtkJpysjusRovYCWhIlGVX5M/dUpTFFQRong40pMLlRDCnhA+E4rfERzuDkXVB2DowGmyNRK1ZplXilF2B/QFe9uSWdV7tBr2aIHVr3VLAEzCGaQqe95SKQhxdZYHQFNMTlOcy4tcctvCEi6z2MFVp8jIyQtdUSI7rYp6uROCNMoBlYb0fG2Kx+Zdiprwz0pEMO4YOoNlhjqoS0sip7p9Z6FpAOiBHcvMQjaT4pbam5Nq7l9aCKzCfO4EzU9/46Vlk9ErVYMHnYGX+RgfEtfkxXLaImL6UUyDyJ0XbcHaPpGU3QIB1XwGLVDPXYobXnifOsOjr3WaFL3Ph2axFyOQjcDFVpl0f41QsqT3omT0w1yBqKdJq2dHcjUAxSDhpwlwBwSTxGa9uFvs98ccqsBJ9TC4nt/qkp8Wf2bgunOtGV56ObmxPr9IFHl4nORBoe9zsLW+lVZTmiyUXbvN1DObt55URQO64AsJyWrzTfGHYwa/XZ5FduJ5OCnd7NF+7268PBa7oKEoRNO7uqNA3eTe+4TexyFlgMZRftK7dW7LXDesQKqqrsIpRLwriP6zI67NryQSpbs9InwnPKYDFbNRCdiQCzO0q9zrL8TaF/n7Eho3KnjEHkLt9LM+nKstF0PNkq/iMbyHxD/O1U1kCdLHngJt1ehTR+6PxyN+Tol3cJfu9591u7d25anYYTCFL9AQ1FP6va5iUf0/c7xURMldl/uikq+qwH6DKP9Z3yn7X/VuYkBEUpjY4AA0B/HUA4/cmQzBDFXlwLbZiA2wfKixMhl+2M2Idh0Sr5jj97cNjTzPJUp6jpAh2T67RtJfOIGdD9G3rsp6bW5U3nUFHBOQdk/mK1xM60GTiSi/KzQBFutoyqABNbKGuQw2eIUrp3g6K8Ac1IgvElIrF7+fh0A38pipN6sxBlCKYuAHo0zwELkUjEK7Fo+rDVLHYMS4Z7bb8OTm8D3k2hu0zQ/WfVG3J1RgjXjeWSObf9mnY01bBCDdhO0h8QX8s0T0gz9zDBekIyzbDaBwyMwWHjKsbG6z70Q7eRVWBjWJuCJIsBl4kthI95siIURLWei42EpSBH6xTpQF7YfLa2AoAjBKcirOcKMKFysOwYCg1zhZX+rhbgFMKJVP2x3ygYAIerDRPrmqfYT5SHyXh7Elnsope05nGX7GLOvK1Ck4m2CL6pi/FDfgJnSZDecj6GGDXWPW0LtpeTO2JuBCsFvDgcz9ZWvpjYPrHmGw1JX7yWG64kTapt7GI5u8usIEvmipXKglGycX+jRqNr9MQwnXbBjQf/xnBpCQCCLbdQHdD2uU8hyLF+z8ZGfmFphxcRL8tLmJlwdlna6xfvu4Qjdc1eNYCC/i2gkWGRw+JQtN3vcwLQ3YzOHJ/OeicCrXtNJ0QtSX6Iq1yvsvjRYJyZEdPvE52G80n4hVtiMXTKzYBhr5T5GKnNt5qROEJUAXrRRGKgdACf5XqtL6h/0t3cyJzoCD4MEikKzxRGwSFDeoQftu3aj9+DMoHz+vCSgLoBqbU4SC7jGxCUD41DZY8cGoyz8R0OPb4t70E3eYg7oUawRE3/16uzfkqZ7nmwMjxY3vxvCRROM1eJnhUQPj5paSeDp/HDiqmaiA4Z+4bL52fsDwLlRkd62PTfEN22+IA+KvISkHywenLULcKhrV9C5/4K23esmQpmtIn+iEez3b24AldzVYwjOQXDFgxCO0YAwQ8UQet3AmBCf4JzyhSLJzfZx59EB9H3rQXNY3EBzP8AXYBKW8TtW+iwqLLB/U2PQ76S5+fQsU7dqhEoJNlOGVP873ivCTrchMSfJJUw/WwnRrmuVUPHgsbKSf9tglKpQ8v9+gHoDVHiR0ooSW9j6RB2N/Er7illIpD1DjA1JFvwzKQUSQ676OH+U9m4hBeoY9bjB7Llu+6ib7g7JyzwPR91NVnzhOE3MG4vIJK27siFHdGhP+M3o04vyJ4btqirV6qnYagCktoZPEvneISsFUJMV2MPmK+o4pfQldo4Lq+yP1nw4OwMqM6y5ao0hS28CTED5lnP6Sn39E2JScM2tDvi/JbG2BRnHVnJmhhaahEf0dT2d4yaHEY2ywcy5Qwyf6251ZW+r11OQbHdgTgWD2DD5MLALYpJYpXAa7LJE5giEd+MATMY53f0+kAgVZPr+x1E9YzvREdXfuJIrnHmo1aOYmctSEW1mvndiHVt/PErjmUktEzki6MZx95vBmnwSZpNq0qU2+xlZrdNyQYN6zK+6O7FEwXN9ebSs/pHSbaE9WrRxCjmFPLBWke275RJxfjFkI+yUO2IhuPBvrHiwyPTOthz2lJdxJBjYRA7CluZMuVdPDDBLOFirsidxo2oOYIhXF20Wg0c7sCak8HbPQt+eyV9c+R3BV6efuDvZkfvyxk5eE7X73aWKHXv6RbtV+zL3Zy4ITT+KrJGF8wAE9CPEipTMASO4moPb9GX+vtmwXPNb7VQ1pCI8Cks6vfpwVpbKcGfWv48ena9zDI0aG0OubnVeotlFxit3GspKWLSrd4t1S6H1rKSfA+nlvUkrnMVls+B7Dylq3HSQnrZid5eOupxj3m/eGQaTu/T0qxaBYFIKXM0WTDdrCvjJXNp1rE/UZ0e3Z/iQlhahqwhpXz7JqlGYDj/1SO4/YJWRC/cTH7eg1e8wUdxe3v4ntCAvxnr2uPb6oYrUQ/74f1/ecC6dXAasHQK9/69uvqXY3fVsU4BiNhhiqjSDUbZiQ2tuLzQ5kmOvhGoydxcUaYFGzB2AfrMMvPCsvcWh+RtFuBqQghQ6ICiONOwdqtalLNkwYxDB1G50222V9Fj58rgN5lXTNFEW5lOXOhN0qCHZk2DfxRZze/MmpqRlxrF3IhD3AiKm8PkNLTyrE+NYU7qciHDxO8nyNGyNk8/OT5xagnN4lkQOkGLeWVE+NGsUzigRmSnGihBYidN1vo/CF9/LqMPMVILNLtAqtxN7bzrUvOCLqgdbtcWmEPnKRkY+BZRj2tzOzZvWNaE80TlNNxfVWpkPFkgxOJZZb3t5G+7TJIvz9ljIDLPA556bkLDxecC6oCNvzMPiBwwsXwLe/Xah6Y/+AQ/MqR7Z3/mMx97YnXffXeOMWaYlfK+6GpuAMiaaPGqQS/R3aCkMoLtdv1FA/orVdftSezLn6pJG8BxZfJG/HYZU2CVDox/RTzMxWkz6xK7IA1ZwAS4b9Up4dX8sCc+gYEEgMvuTmvoBsoTA3HdTdWa99HuNKORpai35SLTMwRjErO7RxRXBJ9xwxAc4zOC0KXO34lGrDgOEezIroQA24FZXvPL2elF2SdCAzOUIeUnyT6fYTCfzbBCaSMyQdb6syEID1Q+sQeL4/FGTOEc8Kh3MKCmpv7SmT7m7eqNPhyTrfy1bITucjxKD4vmSkBAyRzGlmvH14ViAiqDfLP/lvK5RAjbhwqaI221FmodU6hNmEQJXklP9UacWiiQsrXJOBz/gYnGCd/FIMeQRO5m00iFwjVKxoPPebatXyYNQssvkbEnti8GjBtFyfy8vjLpQ1U55uGzhj+Q++R0UFe94wcGbu3Qz2/T3rZ+QpdPrZ6i06jS8oMJJDzlI66GYaICD2CI0ekPdNJzlDF4nvS5Lf1Sn737XNWzO3Nc3Nce9ChLqmZ8WgvFPFVUkodXau8zVn//4fclPQegvtVB/pgWWGFCSL+g8jmGMntjX8K4i+pAcJWK9iwGbswxmRD0h2t1/H2sAIstDVAedQnX0daTSV0vS3wCO9hE92ed8J1nypiVe0c7A8jfgZXZ/3eaKS8ETEw9d+F3VanXwdRnuYQZjpvBnWY/wsiFfmVn2P1Jk7H2bWdM0E+GdX64K7pqFwHn87+9oP00JlcOOmhooOU35ivDm/gMU0U/As6LwR/3VXy90C666olgwFoRdSBAKzbQh/Yu3+k4xkaBmKaDIEgLi+E4vG7+3CNB6vxghSklj2fb5JLrmdgkII6aPbhqljYYSE4lt9KD+CnhlvWZZFYC8D76mei4Yis2IA5ygwWPWmV/2D7aDIVT/oFM7xwK/RwlUM6E7nH9rBT/J2vpM0vCG8fz6tmJXEgDaWToGKZOGo/Y2ijuIi7O3keqD09L2YxhfvWmIchR0b1ZBXGmVA3rjAF1w7YeWEFZ0LjbGNGvE8AOh+EflUX9XV/OaQw5VQxb+6IMU/rf0jKUsXzu5fAGZw33K6hRdozqjtn5ppEKdAn9T28DJwreSAbcgkuY2cXTWBPwaf6TlEQuquriUm+aPfLLFE5se+/humcRubq6U9XG+eEIG384SVfOgT6w3e8EOqaMMZqKSXCu9iYX/0msIHmw/+KoJD9H3m+woLsaR+mLBHjHec21AZy5x51XV+OjE6s4IWYM6xXebuG4hvVTeDoiHWMv7udSmI+99ISNiq6AGrEO1wszjidxNu2TTtGmEF708Ia0laQLR3W9oIGePQVFF42WWSH4FAqZVm8vaBWTpdwYT9Rxc2jeQugFD6Dt1FwyIREr3SiJpK+6nUzaISKxZH2EKwMCterfya3t3Ktgy17++lBnL+tl0ssgh2deBNQipt6pw0c5jQ8+Clqdhg4E4kgLeCxIrSfBDuE7PHqLSBmpPPzLtYwhvwg2wlqFBkhM/K7uX1K5rjVywwShHFMX+Kh8x8XC5njR6Dut9YrL8wZ0tnldRutDljcs+9Du1Yc9RVRCunUY/5aiZGl1HHTTCHrl9ceeChrnxIwW/LHRs780LHcWGVawo01fArtKQ6ziztePmhzNsMBapQNO2FVlq/cv9IQmTHV8zNnhWIWRzWz4kolFjVpuQsy4C+KzjNbhZu0+w/YmCpaYaHlh0w6V4fSSTflTq8s7Z0UgHULPotcwQHLfpICu0s1JpZ1L8Sg1iDZqSOwy8Xm+XgCGl0wf3v9/rebrFg01RAMP1CZpKUwEUNP1MfLttctIiNI9m7DZqQFl9pWB1ZYL6KSWhuhZ54zzvI5Avqo936UbYM7tHnvlHGRDO/3v86wOnQgPcAZQuC5LhqTUd6zwo+IZtUBB2jkFeat4VwjcTHdEArheG/qg7owLkna/Mq00K2+Au1a3LQ5PjA/rh760MTNNNwya0ZjX28mdKnaPXvepey7gw9e8kgXSWxN5kYchuSDnxGB78ApP1bqqOYvlmZjeKpVY0bTyUvie+1xAUc6r8EPvNx+eiqI5oLoEzAGeeAmUeMJTRYFcvKyBFxSoBsFH2f1xfpex0dVEj2f+eYyBRq2QrvzoAXmf39UgtnFFBzSGCywSQJ1n6tQ56l2gpzkMH5ssJ9+TuS64Ol639pSOMW89UC0ISks1AB+0CjaYqiZKxZeWl5JcB7bGXpvQPZ8tgXJsW5oh2/EsexoLYTG0sPlJodmSI1UZKCi1RtAhPanrScXaAmFv8Evnk1WYGiUf2gfQWa/fmdKR8oG28WFSfu4KbtpLU2rry3Bc6qlkyeK/zu6rF4bw0qQgmnbourkraZD1+LNK2yq3/g9p8CtoxB1jbkQ68D7hGSWPqCmajQKcH3zKCOSD4kRHSOKSO2X27nbSnNOcQDQ35LqmawDnjiSe75M8AUjQtrJzUoXYt+scWlZLdRmWy6TmPeFM5e1s1EhQxkjUYFTpwf/89JNdTLz87I1Reyml4fTbx74F33k1i+DkQY/u79xdfE2boIPMw25oHNG8O1yANyP1/M6NGlHgQgiiFbra1vH0o0KKIaoviywWgjI9E5sajvekubxvvT03QfvDosVMdcz88lLGUy5StNi4u5a+6QhAeUEqpzS2IBGfiItKsBsYxyCfgwR79Lb2mtJ8WFHcMsoJPBrGNm3PMFcMWJGax+Z1VGmZDfLRZ2+MCWUejl1krPpWJShnKIlZUlXn+Rtxqhu+hZ555mtUlMoRnwxgyYwOYJNZRS0d2Wkd0qvpXssdjV/+i54xEXEzrVgpjo6asSYSTdzsdtWPESClXcdRf29wdj15aXi456LYzcTRPAMjmmXPayBTkIA2YaEi9plExKpErRRZrnRAMtwZTdhWEySIx02YTnJlkB+SicWUOltycR7YNR7SCsiyTaRsM+wLZrBfRTtBI+zmZ0Rp/9K5ZU5dFvP9lMMWVAJ09KJ1cazFcgivwiBGyFvaR2He/GNH1LKEouccqOONpmCTntT6KTlwqaORKERzqg9m7dLovrymHNTpw68v8Qh6AasEWbsh4zUsUnEzKhmAIEbXsOk2l2HM6pJBH0VmK7wCYb57QfeoQYZyMM6gkMTbJo8n5OfpMt6qiNhks570zAxxsfZkLq7JKI=
`pragma protect end_data_block
`pragma protect digest_block
aa2348f23aa134e6a37a969a4ec2a95b46bca91a6862fe31cde8dde7046f6dc6
`pragma protect end_digest_block
`pragma protect end_protected
