`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
AkBYxf8jP/e9pgopotoS884Z3VFPAEZccoZsd9U0ZUIVx++xWgJMzcYc+uqoQEc8SXx16vgmenJ4gX3WdR9pFc3fyr/tQjdKW35Jc7/qLntJMGdmfOgWOVsTwlkfmyfYl+e+4yxYATbGlB++Hb+Po8exGgGm5UyTA1gzho1s5QoUi21i2p1k59D6MF+zuYDaBOTetHNeWeNvVBF4q0TtiqDaGxzl9n8eKTNJu/iyoj64FZVTo2xBj9m+MZnr5W3Rn7pKX+b28Ym9I6d8EtrF5tHVp8C6C0OQ/MJc3gFiCcQ5neg19TuzikSoVrByRGnkxuBWkQqR2BkkCHJw3J9jiYSUehvE6M+Y4B3o5lDqlF5kZvxIRGpPojuEscFmfwtBfPIinUfKv2r5bENzLsfhFKqBsfCPWeyPnVA5V9BQsTfBOHTXWEMfwlvKRtxszeRgIeNfZvEByGae/9iJ2cBkAEW/Kk2uKnO8tjKR7SkDF9FFjkfQGw/urTFi5IwHI3QrayuaDZnJa+hmj0wps0K+SwdUrpLvMHfj0QBMZ1ZNijb6gcaiF7i0DjEfcAGQfFf5UghxfnX+/iZWAIft0ywuLEyM1lrgwM0DhvHwiYCbflBtcuKU6nQkACd7jMH7V9BIFE+rW3QC0p3cdqiANwtfwNtmoqSRNvPbpHxvVw3+6zoouxFj4Z3MC1XcQr4Uai+lUFDNX+KO03oKXYvYHEKmI5Nf7BPiyEizSHV053N+N9gdbI4Vdcyat51lYQUufMqk9z/xV09aQoD5qE07JYedpB5FMxY728Qif0mHqOxXrLJAmabr6kgtfjH3uKWYcCvrF81dBW2LXey7su2fzrnYYNfgZPqacr4FB1GZm0XFSJ97UDAf1mRXk85MIoRPDe/PPMHmWsGXSrFyIrEcUZiIUMRQreXNilC3xyHrMn5VjdSpXxnlY/1HtaP4mnEbIvNYREI8cM+lqe02tzAbaKBG/0c88YpSBe58YeQE4P8WckBrN1MY0XvO933MEx0ud03aVMcV3rv01OOqBk4a7PtwdRF+Qmw2iQPu4n+K6Rm/oMAxKRKFMvc9xN2+V/BA2rPgjaj1tjZ70EP7PuKIdnaWQq4WABuCvzcR5cQRbHEpJX9WdBaug6zgixjif9sEr24GHkEPRnOs2bvLD+pxAqy3Ie2VvPc2yOp5s8X/WDJAPnUQcKYlJhIzyfJvBwB8kxf26KFXOIFaR7+hZU4fISXbrMwkpehBnj/syTqrILj6GS+WEYs4QJpFz8v2h3L1MKP4pJ2AK1owhvHgv31+wJtn1rmI8S37Jvcmqzsag/yjVDEmLth8AAtAFIQSN8JQGdCx7oByFj4izsxR6dz8z9NPLjHXz8QHw8o/MU2vnAkfyb3/bo5lwZ9sAfl95EE1vRoFxA9qWXX+kkz75tq+/BUNo834Aj50yDJVhAKPBuACir6XDGzjbiHG98dRaelnEbIqmMIFirEIj6jIEDHWKRjYhbu/vcQ0dYzcTZowYE5+sMxOXWNTa5Z07CiWPUasCTHcpnypXP/sP0NNMpY7Iez5PMXhGqWtyDwBLqYiATNxvKG+UmeC8LMT5RE7Xh4Xt/C6pIFSnQ2yGzMcbsMWQmlKAZuyVzu2Yf028bwfspKqY7WqMit5TV3HTKqTQ8euRG+nu3FgVw5nhxHHh1eDi3N9wuz1nm1ICCKJyupv+p+Y9VbAx/wDZ+CjkYQfHd5U5xfkARKdfR5TNlPHg7zJlFalwPhAjDuytylwp6+85yEEcUUV0gwnL5zUQeBTEaAt+qaMshiMrAzDw/YMcFq1pEC2L472ahNfhVBJ7xwucuGYNrMFQRx+6/0L9gxhnchKC7T9gA8y/n5lu3PGhEOqpSzgBvnlNRkUOEyTAEpNxLTzNqeI4h4SZz+6M2U5J6a97OKWk1Lxte68OsjHFBIkJLFIILS3Pq9smLjCnX6gojgWI15NPNpekW0wVvY9DhBUkPtq5GviZqzeDOnE8f6F5Ycni+ZQwPpyF77Gx40omLGRvk61/N4dOOmil4/MgFh8a2q2fU3Gsdk84W+yRsPTQcLlBcKySWGu96gtBWR5lauTfw3kCy1ZmGZc2B8sQ/qRn2foUpTilgk2dxGX+8cP2ktPDPuI7ASsMcxx2rsgwnJohvi7Tps4RchFaBs0+vbaoqizB8zpxW5ZcXxeJoIvEanrH3i+Szk29z6Fsxpp5CXktf+r1AmsCJ3SZy4oh0pFEtPk5P8WkNnI2DkjN3OonC4ArmyWb9zGkl5CbWkbQJN93VK043rxa3c6Pj+r4CpeTlipKKcJr/QhTIS992EuEaYAsXaLlJrEUBgkM3Tw5fq7WbJu16HqiZocRz1b18ctPT/TmHxncImMH30v4VhknwymYPsraxJ9IATlRK1pgm0yOhmXMComZem4WCjUiBP4uMRXl/mzQClQg+WZn9CMBpreSQUIkP5y+Gx7SQInKvmcqSb5KbqSzBcQ3ADxEKqL8Ou4K+visxndWHkngSk0rXiaXi1oen0Wgt4O04xWSYUFco8R/QTrjPZR8cOCqYz1H7o5NNN5bERO1DAHUfFiyqsQECTc01o8/hVFBWEwssDqLOD6o1r4pZQADv4FO9FPbcc/VKAbuIiXc4vq/LQnHoXVi1MJWkvuCX5n9d1kncDRbhVE9FWqLkhyY6Ag8zHwD6GZLrH2oOgl+xWJ3sx1rkkpwKCMOOwcmBKSDTbP3Usx4tb0gpNqMIQmZJtzjF3Cxdqy3CPWa4284dz8kMVUf8BI+rkidZYl8nZ31jVzq8Vns9pDvHI26D0Yc/NNqgkUDQmwjD+6oIyN1fuO8S5bElE9sYiwOj/uPUfi7fg5U/7TnlRdhUMMSdvbN+LzGdvAtTSIqam2b8zEQ6mz9oEpxUtjpfQyI9OYVUIqb7OUWjE3bIe3amOdw2ffenxRtca1CvjfkloksK92LZxp3fNSR85zGTmHw1Jh7WkAzKQHnchkqhCZT5dEaDbUPta3v6+l/B8qidTaHNMsG/6+Gk92pzCnIogPy/k0luP5aRO6tNY3tiHW5YOyS2B1q6RtiK2kBhlL/tXdf0IYBdYWNs3kwzXvkDQrI+Ryr46Y2CTjpVFCIaT8QgT4u+AGh88si1x6GfB/+Rl9NHrSr5HpJH1HDZRP8/KpGViDGLSmBIf6xiFZ2P/noibCzg+zZ4iforfMwjXPYW8vxUU0kJboDu2Kmo7BIF7amrnwVRnejS18yWLFbC49ZGjmsBmdWSBYa6U0Y5Ax8Um2vx+Dt3SHxVtRTBIKjTqRuPshFKY/AXMV3GqJTqtUpej30iCMeYJIL+3vAKPe6bYe2BSqK7RZTVtxhOMhtxHEeHSGLB14qORyA60q9cI+XNfExmoSRYUujBnbxhxmndeWOnoIWu9B6r/GH8tyQgjOXJeeCFreXRAR4GBHs1da9IPSV5IEtikimGcD375tcBp8xxgexpJKgydBUogMLKa+eTkgqGm76jPf3b4A0NJJZz+aKXrIwxSPd5tTas0SRac1ZFOv8RtsOALYIjzVeTTVQiB9i8tqMZDcA+5iGQuwBQU4FykNLXfEHFh1ZRMTpsgQ0QFWixr68CtzdoLZcW7zrDtiw7zu9B8kMLlduvmZOsaZSkGP2Hxot56UudZHK7a4hJVferG59mUQR2ae50Vi396MMyhHulbQawoY13VOhZF6ZQemuLhw6cIMMwyYUwnIcmrhhqBfBiqJ+nx0q9yHpwP2hb6vVnXfkBn2k8BIyaZ/SRUyLrEbn3OaF7L1N6lS80YaJdq+W0LX0ZnmqkcNxluqkD2lxpbn/X0lYPeyi9lRB7IaZXb0iAS/ZNuTBh2U5rTjsWuAFgnPM/xe8iUJdyjgGFPfy6zzfAj2RCV17PaPDxkEruruwZ/bsFasGjqf3IkRJMoLwBsthyPRcp5yCxzBrL0WrAU8DCqCuSkvdzHQ/YWThatn6CtLrH85hohWgmsG9422Fx5pw57HEskUuDaWOE5EO8URF4AZztY4+dzVb1f4kuLZ48n3E5fHmDzELeeD6E+KjZcKkG0p05sUO0yE2S8m7ko7i/jXgPvHkuuxA9wa40M/H8AHyhMWsj81HxJhOC5oXLZUnZtGT5LFcNZ2GWx2ZdMM2dQFjmYS7N0GXgO6yskagFye3wX6cha4Al7T3+50JWFd58BtBE6YQks5Rr7LHfh+DjYH4Ehi4okRUwylGozW6m5z8/NJisg0vQnCC29cO4BkDIEHb5UpJQDm2ZySo2vzgvIXIz71uQZJdVU7Qga0IZdALoambYVALVDbHfD4suxC9S+1z4fPE8tPlnL4SERCNX4W4WlMVbeDjSTobsFsVvEpIIXGj65nB+3B+TLwaiQHyRJLkUYztOjbBLHGXwBjYS1Iey2x79iYUyumN8/i2RPYLCvDfQICVIF2PLoiktz0WWvQJLg05JMCGJVOAamqpmAoS0tT+RO7NYy3vLIOd7vzmimGKx1x3zruSXim/EVElaHh56i5Mcvm4sOSMIvuByiHY2iGUIC9cGdU/MRwH180m95MhcyZFyTZ78j8lseeDuIqSnQDvpfIsgkITmsnJaXkowXQ7DaApBWpHx9PMiOzeM9NxnyRKA4E+1bconMVsIuXoEAj0okn02vf11kY3PptmudROKXiENuilWzr982c4hc3oItsxHMMglRNdYRf8fqcTfm14/I//IgkEKBHnGLjdgC/qQntHhp3SaGUlq6lUScSkR9GS7GSNf6UC48oibRup6ageP3hL7XFm7nA6eL0zJ8KOhkFOESF2CpqdFodAOpkaFdIBwB4HoOQ4S9NuRfRigZUhTZSfxylx4XNb2zYo+Xxjt2EAKmFqK2dlC3YUqEZOOIEfEVWVuH4iuEHbHeKcIAQ6/C1AhSRA3w+mBF+myV1svow8zFXjpIz2R+RNI87pxasq6vfd1Pvs7YbevilbjagRQjtDeG50BALhTk4stdIvvUozJ+s/MpFTsvSzO99O7uSp3TXOAi2Waakky6/InbJzH7OM3tz7vi7CQOzq1yIwqMO9nUESb1yEaLXFO6hAdFjCRuvUmH3r7jtnfNYnLJ7j4RkBRsrKjYUYa8SHDFKG51bibxUxyodp+1+K0HorLO4UwkbsIEc2gcIOwFzuGX5GvnQQmYy+49JOCjZOdvpwQrEf/yhHUIUlh1N79oWu9dZsLibf+bT1W9Wcmktmwv9jsMon/Us3huLAWShHO7uSIORIDb5UeV+7BJxaoU0c9oR7Nf20rxbEXTdukNHyv1Mvd0OlV2tl26gZ3rkB9slOqqAI0LzVd3Idzo2X4RBtKTsnPAQf/Pxx5vOlu3JGK72ywZqUfBbfutQMBJzm82uq+0oHtFBjqART94tAkBooHRc7jNhr6KYg/I/P3/t22AhLWBDBumNCSuP1wLenHf012ycuSCIs06uDH/mWm5Jg1s18E9+l1+PmVFJ9jIgXfmrYJvIsSbp5AANlmuByKTBFnkmZJQYZFkTZLTeNf1MgT5RuJv1/wnJP/LPY3ADChyCMWwp5JnlBd2hx+5h1ns57IkVK8jMn36m7s1a5iflK0t+L7ogD0w6ZnovCxuaYacUF3twxjybK1GKbWLpleqbtcORmMPCYZFQZku6e4BAs9BELF1jegjYoNnveV+fQpowa/aGq+AQHVKX2gMI4ERYucEeUiUGgNvp2Cxd6Ao2w7pRqIn0ftRxTcPZ+7f2AA7hPX5u8oGA19JD9qiKJ+gF6E1i8DDNsY6hTtTl2rGSc5pr7C9VkMcOMdgDG3VHXmsCHu4Q7FHGmrwGYqgXBGgqj+rSfhobdRa5UeWfZ5KEIRqH/fcOIi20JeaQOvUe5TOx1ote8z7bcAff+eyOLan1ef0+PMsHd/3u8MYQHJBIUret0Jkx6gdKMlyaKCA0EQEFy9EgWCP7ctdUvNaOnhL51V4xzA72ZRgONWGkL2Rekheovy8Ed141iUaxgFGC5dk6yqyL8LwNHZU4Z7dJqALknEKRjGrRo0NFiES7ySmk2qBpIBCs7fUpWhqoVLoeywfA2/yRlmMl9t82p5vc5gyb3XgMgLgUk1ULeyg0MUHPvTvHJMHgbfFfcUlHoYQhQ9d0L0DSZAZJ5XlY+DNa7aKZNtjpiZfRNZF9aeqSoxdov+8Jf6DL1Y0D7sChg+mU8AY0uKmxAByg+QDG9cfiIICgGIL0bSCkxuhdOocZyfQ6VyTiWv+MfRTmAXPgNZqBlIt5UA/0U3r+xyXifVW8zRyacz56p4ljpOxYCr4V86sjl3D8cDqYuFys/+7KFNuln14egfEae7Tg5dT3LuOmg8Xc4q9kyc3e1I7STSNil/QI4wOvzncd6k6adpD4Xcv8kfQn/VgfNGvJPc0RnYTnlq8RasqaYrpGG1A+fwibVIpc3BpePpWVCoS5/rGw4ivaUiIl/SQ9COLq4QyxxIxuQ8sACwfSBIdaq1c/u7bZopWVK8Bw8Ex42bzKz+/kS+w0M/dXCIg9Kr1yupzTQoZzfVDPEtuHZuMcF8iYCs34h9bmVwGsv5210iJJB93jtxVKsSSN5VQ/UQry1STI6FqSDxeyxgAAdWG6peHVDXc0sOHvLU7A/NtAeBUlNYv/Vxy8sCUqRQzWqqsiHOwASUB2gxz8DGOLsjUmzCu5Iqrv/XbcdWEwjrYk6AeDZEUCDVqNgfFCYyCFqAmDiciuJXkZpDgqZK7vkHUb7abxkohg8Fylrk8AIbq5d2HBRrQss/yd+tn3BkJBjzYpWwSbO2cvwKuiLwXoCxLRh8vfjLibiNkdzjUG59spGJzSb7XtOIp1PnLOt/8SepaeTe6gNEIilLjNUWp/551DIzDxiEuYLNvdfXAECv7g9kQhuRHjwzN0d7vaWpjrAlb8i9wQDY1Su33s2eX6ruJyk0IoS6bixUCDMWfMwhls1stelEXp4/v4FZIL6wcb+81o0mkPFMNUMbHiMKqTXQiIvb/C/KD8TamPt3GUzVHBJm50X65KXuJwpjpff/hYtQCxTG1XMUMPx/enkEzSZ+ktMhjkum2LX+dw+KKVfA2F88mc7xPGooc9RlF/IDkCJwkDkI079gjQjxb5NkIJIGLpN+Onyqlyq3RJ1wPv6fjgR89R5+ZWjRFZtdCUOqo6/x9/WIkJ85npuecQrLksoislMcsaLzbvkwyj2VrOi1RjNFPY384LTCQvHw5DYKfm2iFS/WbAkd7ND9Wq06PB2Nj3UsZOWJSvliQkVvFzH9W7BJnI4TPLOWoYGMalemRKchpkGd0xCGjYq+DGLBWXJ2lSYOZP8WMarV+vgpUEsFrK8GO7NPEEDljKZWtFh0+dFijBwXWb7rdQMCtzZf5LHo7GFJs/lYajfAta38xoGL0qtxhggtDO8cCd2ZL7VBKSyUFPq5k9hmpMOkxmfWLgAXsYmGbo80j4d0mnZg5hswfYhZEfjmDlWT7I6MV6jX0J40cYGgCRIxOdfp0QRhHkVUNU7BDYV5qfgUZiP8VgBi20nFkOswWFsfTRjEWDovEcEvGjy+PPX667EtBDbFRf+H2e/e401x1iat2faZwE7hvYX5MZOtw1m1Ib3uWJolggMLZTJdHeDKfujwNu2ag/qzQ07kNd4vtygCpsaZ6/Nw9extyMxYp93euFIvr1CLcKm/CA8WWT2prTKWTbbFgQtUWxQHWGbY6MI1jS33Zzj7Tyde2B3Ey0M93Ms3gDGocbi5rJrkd28NOCiAtuWwu2DTwSFUAeWH6KwUnuKS/2zTiB58DD8rf9Q0DbBihWCY/xRGwdJWYeDg/s5OJWWGbw5wADFwyD28p3wvwvWMCjFVTaxon6yYL7byQIja0wbyXH3xSwkQ4Fz/e42uArS4U8fy+zkXdK91pinyHwZ+5facNUGH5jOI7iUIcyaVNyM9rBHtK6JYxZnOLw4TA6e8A8flLl2ITh0RGlJCzzHBTRLRMQhjOOFDL5DwF/B1281p05v7u6YEfXQo3L4p1YA6jA6SJr3iVnmdYpxrCdz1sYn7WpzzisNJBupKWnBoEVKW6es26jPsO2khaMbOWj4Gak765hfUi4JMe6J/Q/Q2pG2RYSIUux2dzi2WPviwnjJj8oGHH5kzuqUs8wRjqUAPJP1JsKu8WZmxQnXId3BgkqPqE/ozYfmcrkV2e7dWqTXW3ekmEa5oea2Nw9GGIdu21Zcwgx1SXJosESH3sKtZ6pSwaILViatPOOlGkBt4IUR2hZ1VBELcYhcacpjN56/6dH2w873tCQDLgJgxNZ5CzwvAK0n6WzdDfF6E7F3emtihGyw/r8nhsm3rbFvgJRiwv6lanvotUlhO4N/6d2OhkTAm69C6mvadXBCXA9fR03jIRIe5xLgjESxXGpr9HZw/E0SMvqR+9E6tg+XTZfxh1jzCtbUHfeoYbBzC4gV3R7AFxTySnUHn3UXK8l2i75g4ZfwIOAzbjFrzSMyaevGiwb+KZMaH7HuzvZsXcOJaGiXYwiFrSFkLdwuDbYSJP2825P1u3E67AtJUic/lZSnHbhe/C9d9hDP8O2nc+TO3YVja6s5Rcbkg6iKrHkleKhdlpkeQTEWgDq3RV/j8lpug58azeGmd7RF06KX5Kw8iavVDDhfASdGXBdeBqgSkGitihxG2utQHB8dlhHn8gTiEGeV/npbynK4IA5Hdr2rK6VNbJIsQPFroKX2XyihJRwxaDy3T5w1Ztcw2G7ukqoKdMLYHpqJc1FLxOW/ePF1fDnI9VHSQI7fowCzuktIM+XBqZ8ZwgouwuN0Yp5AV17NLaGXOhSEYWcOA0ZcGL6hzYsN4YDYfcJqA8y22Mvjp2/Ytk3bwpToU6/lqRBIH2KFgDo1k7eF0vLGEZQ0rB1ByxfpF8qW39BTXK0eZj3YX0O+pIiPgcsewu4hga/rN7m5XAC2sGYWPQ1pEQZPPL5034MdvTaPOMV1YimqrsBdXyZO881ypgfb5dhU9p0uxvIJ3BRp3ZdfIIAFP6I0LxXUq1W2KUk5jXoA15iYaF5S4JzZPXv2HhvjOsE3lgrkvb6f6X/d57ZvTAHMKewBco29kxZ8XlS55JiGIbq6FRHio26niDFHiBU1tqwKiTnGiRoj1pXn2njvV/ftI2GkoY0BgruvEemwaiMVfdhUl/F1Bg+/xmaWW7jhqqcGJlrUh9gDgMZ0lsME8tIDL+DguUOUMPg+YoWGHEZGt6KdZl1CQCvf0alBzt5TIveEvfOZxr1DI3TXiWqT94pr7E77+a/yTIuyooxmTNLfRGD7up6dw/VeC2nnWDJQ3aW/aTY2MlOCduL1silZl7qKpdSq1N9UtTicbkPZcxYhy7ppqzLtAB0uusF9DSjz8CsjHCGAtlnctCCGkGPwl2U16vxi9qzG3ODYJqT2uTL8daD7mVR46OO4SeWkHoJuGd5PjawHytDWu/QFUNkmRFeq7N/aLwJE9z9jxsSpSI15t7n07CupApWm2E9BvNJ2ZPFoM5/mSWvGvmw+BR6f0KdLEPPLXKcJLQyhP33mQQbVJBdd1VqlbEIdhJJN89VpaPrCXOuTlv9/PdZ7LJuulqdN2rVHxXzkwBWObsI6AkK7ofrV54iBuvtV6aXDh3EiKodJSRXYZdnIvEMtI0RppTDfzykWhAENylG/6jOrLAMXcmDJMzBBgU1rfWT8IlhIm4Y9RLIOq3T1hdQg+pCFtD171iPz3jOVMShVgNUQX79nE3vKX/3qQn+4e8P/gVEJNK5s4NSr+GBpQM6nhDE9usZhdYeVtSPso2Dvvh8o73YX7NbrMPmkzVNs/3LXEq5QV7qCAOi8KUCajIBxSu+8BxqbqoK9Yka6m6NQCDiWPfughoE9nT2SCwyhPnBHyw6T2KxVR2bf7VOI56fOkyGoA+JEyBqV112u0KRn1LfMtihEn3+WqzHM0uBHzKPXHHBI7X5mnEWMtSxzyWmC15rgnkUa4NWiYvMHkeYZjC1Icn4AtUrXfIeyxF9UEUur2cqSqv8GLCoUUUrEzxuXuSeGsH5Id409DblEN+RQZ4eGgbMjz4B+jYkdZSGTGcO+6b9mFA7xyEJXmda4WdolJLNzrQ+qkxHCMmuOtmOTEIr8spkUnpO+5rsLoTtQvu6zmIMrUfinWHK+UbKH43+np6zsXsgsFCScVBvT1NZPT1rKTlxDqXejsoM3H4ftHhWCNcRRxrbwlJw0jc5vn4BvAZACm2oSF8Bbe2bWTloum8J4NeHwW3U5imdwr401zjvXYQ/WsRYsBh5bezj9KQXYpvbfcADfGxq7x7W3pi6Yev61AwEbPqsrryPBlWc3ieS+0D8tK0hBRN3yqE3B05Ox22m01qlgQakDHKyZFb15P/8hr4P+BiagqOrI125pWhg7ZOuCu337SdcqJ4ONZgmVxtum5Kow0WEpWGvbq1VVZPVrXNSEMvFsCmm5NUcbcFD0Um5i0Pn9Hw7cexhqE/mFH+ObRUAWcg4ltsmua7sF09+2fnpu02Mc4yZLfCe2TPcyMB+uikFUGhEfnnNLGJulIRfoWPdkXh+uVMwx807TA1UvbOqTfXOQhkVQwChRqfWiBdrxGksIM1lwc8grtfsk4kKM9M5Op5WmwM+rOJyKpAYvq0HO/lyfolvF9qCB7vYkplYBrfsVY0KC44BNaJVFpxf+FeOHxXl8UgECRXe2tWcbZFhecVzONlRCJGjsN7yebGMQ68BjTVh333uVhd74onGkn7n2njzpwpGcoLXokfTsdYFakBQsBdiG76S5A/JoXnDDoYISDZmGGCk4Ool4MjGzIB0GokYBqd45zroRnav8AhtlNjhlktmJ37z0zNC7vzbMWCY+rBy6mgENLXcQXvc6mR0bFfGRv+ylQJVVWw2ygXjayB1qofTozKPoLdLLrM6g4tfz8DYvHq+2gFtFm7qczLNUQa9kLFBhds+ofhOwZjhDyIuiYXtWGKY9qbu28Kmm1PWdxOfNCjKxgn0LwQIWMXBCtXald53FzCikWXbKyB9VtO5HduSUhMaVa0L3RQ+Bfj/6YzZeOrSkCe6dy5uw2v3VsE3nuF4fvvonln+PxrcVOJnkXI/CVrHBs8YNT/djbXVAmOQUAGwWp/FrfVUDDIK0kZpeGpBzR2qkipMsO6MD25uZkrwIwifabMne2cYYB78BTzAZsZUsILZZskBb2s1CBwk64f8AxV72NFknQEiTM6XOhsEQldKKkVmAg4KjXLnj+YWlbOTqp4R7XGJ7laklKDf8rWOjKYj2Ud4lfFL87HDUceJnov1AFAGgAocIGuRv566n8Wjlx/GfCtL8t3Itzl55Y9YjUU03av4mTk4zD2GkwbK5XgNTVLGJtvhJIzarBFMWhIS/WwG229rrdnnfP5FekcolSEZ8D+LuQJyN5AHxAws28Aw5y+xZdgwktwT9NUzQCABnHaoga928umMNd4TRdaAXnfD5/30jCf9hYf09m5re9Osm5G0gq4mnFUjfUZLXiWYG8LXYbaIii8kECH7OyxhSzJEG9Ru6mD9LyH/x5dvufjcm/54/P9aaBNHt+5p40OFKTbm8MseimM3l+Gm5GpfjEh+cbQuzCeSQuSV4RqU6Nhsm410D//1uplR8ykEhb9BdLcyIiqtQgTpYCM4osiJXX5C3Eug9Z7GrocUp7h0oM0tP1ZmiqUeZ1NIwADRZWSsio4Gy/qVRBeldgPus2dKhhfeI+wUSZjpS7jLNA2bPeAugVzxhtnPVhaXwVydTqfsFnZHabUeLDsWLfM3cQpzka32Lrtdb8ym5qsXTyOpEpTD1rgDdiKHZWgUKIm4ccE1V7c5lOlnOin/goEyRsReS1PmnfEW0SPUSLVWHzMLrBtVk5FEPfG8wKETiXF1NZo9i91eBMEl3ikL7BS2lOXrJZcW2rw9nqPF7Rkp8PKkSGoH281w7ihECVUIEVBNB2JgB0DMW58nystKWy6+jV8JOP+CAl4llWoXSjBWq/ZBFDC63q25P180VrwLX3fyDwSKYT8uCUPtu1qGDOtEDUSKPArkkAgOX/xmwy9faYDshurbhSoCQC6u8ssVlONaMbiR5mMU02xK+bvEn/BIHWgTCfCCE9XzjRBz3CFS3vGFYBd3rFXdKxoYd0LmKRwPjm4cOOcGn9OyGQdxMAlYhik8u/Y0bl3z4rnlx4GqeTaOxCDvJ8f14fYOjWR3Oecp/nJB5rKnu3LH/5guAOLvGRhSeXLyVVtkpZ5RkB/P/CGWEN0mcI3c9iu0O+6RDFltsrefbULMH1LagjdoOYi6M122CSqA7kHyDeeeamA+47ltOUGTOsTIQ6j/6k59H/C22x3wGpTahthy33b2GPqEEzst5vyT4ZMNFMMt2+GnDiAGyKKGPsSmSJWSp5a8Co5Je7FsFWKTIq66SFeR4osEvJqH5+j0RDK6V8OttMA6wWXBZuHnPet/6qBjt72EiXIj9AuCdXqVInwwED9niFhkmTFAzIHHNXoopAsaCvBD5gWxBII/uJfruF76JsAs47Y8TJK6tM5IGG5hv6nCOvkpb/sU+b04O2zLwE7Mg3VlXI2ha3kjZwBBDJvCCmNhOpZCULN/y8y/KC6vFvAF6VARYISemZbCFxVfXds4WxVrGyvHpoZhsvq8W8ngl229ZvDsj5SH1gJhJ9g8DEWTdMGC2JdMMDRrX72NoskoV6QiEZXJmS/deZw4GRkzybICkbyDxAcAaaxSMTMJW4LyCG+VdhAX+CZ4G1mtfdd6ivTEmhUF4VIKFZk1/r0Dv6AMYjatXDXsUjc5HdfaIfvNbZClig8eSHZ8Wu8RiSQMlGIluNTtU3vtBW+/AuTL5TSdafm3Yn+ubOQQtQYbD9H2JCy1DeYGPyzY4O4rnvJNUJs4owsCsMUUduPAyBqsgX4lGwz50tsYggrCVGuF//2bJB5mN2uLXMUXWq/7cm7rqVmnEcKJfOQGrdawQUMLpEe1d0pjS2ea7KdC8aHcznK+01hzu1q/61/cSlOQJuwUeKDozNwfrh3gKgv6uNcjwUr9MsFWEK8OeHyjjP9EOtLKa6n/S+4k8Cql9DF4+8cECsBp7uoxz6rZliPqInUUAj9KQIfyNeIaLRBuPNQ80vQb0P+bbYXOGaR+xkqOYj76m4D6UigwyVbcI73ahsC7X3be91eY4QkdJV3QcdvneBxx5o0D8sHfcLH/qQ7LTF5ZMc8XV3oJOL9YRbL5J4Z2aRz2Pi4tQCj9x1fpcY1FkWlZ4bQ7qT6mcamJU2YDp0ehnxv5TlZILueZq2Jb3kk2hiJBpfoVFip1n4gwy9O+gV+t0BsFd/JbEyahViu7YeXsemtcenXl02UjNNEQIzybxZFEGlIta4908A4+3FsiowiaAcC8o274x39AVoFOL2q217N+hIIhCt2srcK9jM9am8W/KCduYwzv/+7tckzGHM7L/IVzFMEQY3t7qA2DWAxW6oQdNFXxv0kLEoYT5rk8avDFSGbWqXHAq7kzjvGQaqJGfkwrCgfJyEE7QgA7O7ym2qa0tJgOxEJStwARSJfGLs5UkfwS5mnQuLKhda69OzNFewuXuCQoBAPYFyaD+LvQ+i9qgNl7jjOmK1Ot1JKIx0PtGReZ6CTqhwMvqCw4+dWQRm4mQO1IHsb3EMV9K76GUW0w+cNLPzAZiBxUJgO2Bk0hYCb5ZoTk42mNQQwcYbUmc+POx5kSP91FEr46JUTBgu7lQHfOSUbvCmJrr1rRhXMJzJaMHo5I2hU3TrATpUER2x80EA+FOqq/gZYLHiyPtT04234wdwOBnZsidf4P8xqppZyqzppm+eaiS92fDJvNkm9CRJRs2Z+rSbIGSFG2O12V/2sqZG77VlvMMETDtMWdf3DLmtceEYACc/nDmk+TwNkADUzZGWLM+5nnv/Zftr6PL18BYUxhiNvfFC9RNAzp3hBtkxmIAOFYOIMylWgyXYKEkzhIlLIPy2wwwczFluTC/6cdBNxT429YkCmK5QVC57YWPWrlBZ8Y4SK3bikPGJ6aNWR/12pkx0nSqhlqfN+wBJ/AhG01hCcttBS3V5H8OBaa9m1VQZGNlJfcd7UCHbIMPYi3UJHE4saKDCb4UCxhRKS79bUwjUn550Cuc65fiNtoMm1uZs03MCwZYV6BA2WWvaH5cOhmda1dROjXkkQ8KN1MjVZ2/8qXROGbJN46rhKIaK1PDnlqy/2ag/wQgTgruBFVn8z9dEVQJj2BTFo00EbX22dZjkPAe4ies3SXk484qyDCWnXrScxQ/3nGGZmBlHRvyqDDQIdEpmhPn2JoBFq4cAvmhEs9xCk0g+mj/NpjpZ+sOlRqX407V85xeYzYk7fHszHqASoJ7+1wQlHjtHYpe37A3yUZ171qzE7rHwkx4DzJesXIE6OgiQg2unSo2DTrkqE5jP47cuy7Fd7F/fVWCWs1vj1y7TPx/0LwNAkICHwk182ZGLwj/ZbwCkgqf/i6ZYLktdMs+SRAsJyjq9m7o0lsEK6m1ddf65vCPMRSdrYryuesKnAWVGydKOVd0jiqNPfDrUizDFYvrqZAo9XfWSzLcyxuorI4VHJzX36LfweScn0T0EU8wC1gBXQobTy+92nXr6br9IQUYhujLW41uoFkEHTxWZfiFxmu5qT+0t1ODlGje3mnj9+JikYhtvBCEaVVXZDpF3rdYtofMhRxpuZxETYcWNqUXjqjAN3XZp4X6kjnQfTaPmLCZxjyvbzy7DtwwlFWEgXecs9bv+jwnNKJNt3F3JgayalvO78KOffr9eDF9k+FJJ7mennweuEf+kJq+TII+gdEsJWePgnL3O0+JBBGfWL+IHKUOND/OJ4dNJjhRwjKU64IsqF3kX8+lPXxBnD14X4Rw2zIxez2n+WzEAFt/tMN5o3Xl0m/HykH9aeTqm1doL/jJxr6KokcTzbPJHKuZD/JXK44EPXKm/dZY3Z3H5Z/HMg82Yuml5BoiJMXHCuhTJBQeK0geZ36t0b6SKhKuTEFGjxhWRa8rIytoU+yYiP92ShWGgJ0qznI2qGX104P13al0/qp9ZeMSNKPum4iWckdFB12/6QrhwMlC00T+niUA3NBQTTAejzJpkGOMpVA1gDCfkheFfv9l3w121Id1n5qb0WZkT9vbgUjUALIauuGEfaOSoZJfNMOfXZdsdaOUXr5Zgnlw8zxd2SgVSzhJSP6L/XkfPb/6eRZRoSbFJo+dabrK6+nvucjMG5g68d0FMpmsSmUbM/BPTnd5uf7c6y1SQ1nimxhARdEDs+fK9NY7au/+lQctdy7UhMpQO543brPhur3ZRlzCd3tWZkyuOSIbYMozBEhlerI6GoKL17j3l6zkuVPPyMnZTFisIgoBQc7wVenDsgz67qloPxwteZ0tbE/YxOAiu3voEYYMZLzrwok8NoivZnjVToMKuvKRqZVNNWZXtTmEqUtnwFuBbUfwvY1icNE0VqUX9fMPrlI9jJvghY9qHxriWsHjRKz/Gl3a6pnKh/4YSFUeBj2XzoJT0SQTFmItB4UuxxLDOd4+gUQNQNvFJVkPpPW6idruntTE5MWH6BT+QULKX8u59sW+gJydDYeZ87yBWVr5PlUA1nXiPlKjYJ3ZuaflcK5qh0p2yiMj9124lXAGVb4m4Zamc47OX3EFUY/Wnu0ep9w6vbO2jgchWxptN+xHkcR/8iIEwNSWN5rKS4ReQLLhjxI1jMKCj39a+3cTHfGLEM15hi27AgGsCZMMSzPWf2n/sRufZA0g3Wm06x3geGkVGsTLo+9QCmdmF8=
`pragma protect end_data_block
`pragma protect digest_block
7d09ee5ce0d93c03f0b552b74d673ecdbde8c5a46fb2d554193c2f7ac2c8e22f
`pragma protect end_digest_block
`pragma protect end_protected
