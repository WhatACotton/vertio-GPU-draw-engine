`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
UTsEOXPEq97dTByCEempMnmEOhPfswcYyLpzbnPc4gfPVxsRt7fhSfwmMAxL2g5DhlWQqt5L1oZH0aA12hFuZKMzsQVfN1pAWTIM1HAOl4Kc26+VE7sGFotSvRg8IUNBbcBRxGxC522eQfJxxq3JesthAd5AY/oQ2rCO6ABMp+eVeXg+kStd4qRw8z6A7RW05xWUs/AonkpuP4/OT9WXw3XImG2mG04LhZ6z/YUpxt3duSrEHiDgGeZI+S5cX1fuHmm0+iFRfySd9/WnuaWexzF6hPr++5qoBe4kft7dum/SZ0zYepQJyfAF6qv5tHGi5PveJRdyEam9dv/n4uoVngs69RJPJ8lbWCZ7zWTzREPmsnDW5yoy2iQiX2PtrnBLWTCLCKIbAQ2NfirwUX0PsrwhOamIIi3dqjyyX7C+GIrP5Ubj1f2/SVFQ/r3dJxphoK780hKjSm3/CrHOvNEd/RyR/zNeyP4KUnRFL8/9HaGkqikgtVUNLDKD56m/fRYXzHFKVtIxPrS7PjrwOtTu9aALGYA7z2at+ACP5ijipVr7eeRlpDBBUedngpJhQ77uXfMsKLC8rlcF9I/wRsjA64h6agjdpqBAaxjnmolxoApI80E7LCzLeAsyDehqqK+ftXepubCS3vUW3jxIHriW88cHj0sHDMdIgG+dt+wkjhd8cO5Tmoxn2tdCq0oLQHG7GxP3GCEDO01t38zsQr7RhbFVR7TwFgHXS+gDON8UHwiWryCo7QZscf32xtrogvWM/ZDlOHu/R9aAI1qIXNBv5xRzlevZc2mwA5KI6A4uN2HWbiBUCb9VZthVjZm88kv6X8Rgya6OePK8ZrB7SC5QTR0YUgxCk7iJeOy6aBtQWEP9XWgtcUXPcd1amQSkmysxNxsA3pue4diUX7QFekszpcBN/Tc5I0nA1u5kY+Py7guGy/ELp77SKv9xHRtvQABmF289PsyHCH3XfREXlp58TP38q4lIAf+cASI8gcFRVxHn/RllKRliopvdwvPnrIIcl+NUu0NHrCNL9arhiz28sUb4eQUvcQGtxOAmrKfYymIMHkXifEqoZYqrCA3cxbfCkhwv9o6KSEhfxi7piaYJCQmwMXAyau8b43LkR6N5GM6ZMw+ekJNce7FGwwqj7RXSXSh6ndzCpbwp7XCn5IDpScGB5iqPcJbOOZCg9Y8bvM1HL5Beon0/cwnJ9xiriVEFYKQ3i34N9JCl/1A96j7VI8viJboIWmxD03H/XatzSVV/TR75oGSUfXOX7ZBhzg/Nl0iyPwB/SkAFatcv5NdRWgUUlk9Y/R9jlk+VCyEyFZdKJQfXoBs1D3Cd8Z7EPGK9fgpEjONveq053G8brcjFZGbF3shRGd975Q5fGcZGe2Y2rnczQWkof2sAMzc+fvibxQtou0BNtdv983+Qqkv7WtMa6D63IPojSUBWHwJlZeCrpY8UMISkRC134YGD1rEJ1IH4fPxjMjkvmFO78I0UUUmUhMGrK/vM6t/GiY3z76pB1Od54gW+3UIgmMBBQHnXbSLlFWGen8vvsOIr5Y/6tNwC94TxZ7KhWxkqFL53+SHq0vm4WtnHuFds8ZtrOsKindSJJwe6Bw5nhtG90sQW+N1gFPWYuxTViu8Db2CjpP699HUd1b4eMXqeLmiVPW9pimIvYtrw7h0itii0WWTlsl4jthopnXJLhr0GEY4GACOGIGzSMrtH8SUJLPZeABkggXuhIvPDk8eLhKFWvnDCgDHbNonDUxhzedJUdT1hPEt9Nyp/rMQVkt8+h1Nbbqbr/xIDh3NsmC1v6UK4xYQ9Hp5wXpav2fjU1vwMI8JVJk27eQ6JPWvAEnOFBQvB3Cb/YTFDT+R+/R33nk48nEPUAO7A8EWLepXJCIJoV7KVWhdEyxLtU+mc1KpqHwoVHs3PHHhtF8QWArwROgDgCgnnRF1IlhcwqHMKJeJ5O8+1a4oCAQ7qQa7PMzcq4+fMVAo4chPN+seZW9dFbJfFteDaww6q6ZrtvXq/qJIx0a8U/sqHtsCHIzTeC/T3wbHXo6C4aNcG60jpc1NX6F1ozybCPGaRq2ljEBhMtgHgErBZiZPln0tksbaxJySNOQ84DFxCN7ej08lu1j/FWijKnMomTVJHnp2TMso9FlBXTmARwaERYka3cyRNwpbMr8mO46lqAfSw1bJDC3pAaPgtJEz1Nrwtd5UuUI58j50Sw+ZDUnuZBn5wF3adWAbvcRo3z6Em83xMhHlCyDQi65qPxAF+VY0uMRzxGNZAdwoOmcXjaRFnPpOAjcT56FIKpEwaUPkXT/PjTDRnVuBzbX/cNdJwe8Zu+y8w+Qg3h/oa73XZUZwy6KCtaxG2MN3hDAh0uwfFeu8g6y2Bw0S4O677FlXOQujc1SbfUyFCmurhxlXpuxZtqJPltVtz9gPs+OI4aiwoAwgU+9MHi3RL2HUeDxnHxy/9BVACwr+/TIOmZkcG45kMI0bPxbb4ZdygnRz1RflUSxsVJOO09rqI9SQV23CUkztgvKUFJCl4XJLDKt21DWs9ZFYTMitmWAYX0lvqScC6Te7MoAYn9LNKQ1Dixf2n8PSSp8w+08EAMEeVCU+6Q/QnRbUK6HtyKJ+WpDH3rzV8cD2/L+6AGOpspUb6Ey39oJY/l/f47zxFCYdOngfUn4pqw+v9PVdqP3xwMZK6tq3RjTaqJQM2lHgEJf7LdKZBDCw7UybivVRhafuiH01xqAbc7354rcL9Va52CIMeI64DhB2GpYdnnDPrd+wrkH/tFLknmdZnN7VrIdrdwg9soVShRvNBFV6oDe8oAT1LZd2p+L+2iAK7T6PDUNKzFqfgXE9bkaVSysSE2crzrKsRwRTLA9+u6dMXJyh1Pr3yty9vPyxWmA0neaWFH9F4PgZhA69sXPNYgP1aDuuwTKfChVEmr4X/3WY0zda2YK1mCcEqPL5Bd/GrNjEQAhqllBwZaIK/s7IIOIQ/Jk/0iFMBeQJdLFmkVgHItckdTRyohBPuLb2nVg0tXuKrs9fk04A8kJkKFZa1K9Vk9rqZ/oZ8I0+tfwy5w6kL9c+GfdGo3uWIkO6GYrQqK4nGv841JEuQhV0vw6uMvcETxCr1Hmi1FQ87Fy3vFlc9TEffYWxiKG8uzHEpyA1kLJyMfil6Ey+c4kJZLyyLdxnVz98N2Uu6xV3RRIFb6r4JXsEMe6+C6AStOCX6BjUDm4ZN5Etd0KZnRInkF5YLSfTxu1VSdDCS51LKEPEecpGKYrMben85vAaIgLa05kPg/kWqz/Ri2YqRFU2dx+IkX/AvN+N0VmU/S7cY50ZDUOelFuulEkmK5jYKJBtv7NrPc9i0VMzLsht/7tU/4DY2uTtuWVnjofbwaM01Mdl1f8GFssMCGuMF/DV40cn0tH3T89r7lIPdwuZmH9a/PRoTeXK9Y+yYN9n1G3bqmpNxLkN2+MSXfMn7yIS+YPtkPYU+hRLNPsjpaVqfc1QCZSbeblJ9h/Au08vqkL+NAwdNIwkxVqhqyctZ+W9/0kxQeGOQrEUwlIMC+CK6gBvsqdEtmwCjy2mKrxd5XXOjZnCwpkXPY2umwAyXiTf1JAQWVlVoaS7s4QSU34tEgafNC890nsQb8Y5jRgpxC3xhYYWtztTjG2HqOVOUqPnCPEgiKk6CME+nwmmO+bRB/HopnqmzxuyxL2KDBC/XHUq2NrWhkvBp+V1X+NT1oRyj32FBFwBIS6h7ceCqC/QfEjEbgbGEUAg/Oo/v7TB9DBCuTtbTK4naFZUUIPOD5ShGu35YGI+vTn6I2E9oPbfLgZKISXFVEmIMBcvOW43orF9I9fJ2IGWKqLUU3qFpsO68pwqSGZLOlkvhKWwlSD8D/7qvfMO7HVLwwEhkW7RP87q3w7Wtu/PpUF4rwfWkOtKvl+UT+KB0xY/478axfPafx0882DSm6TU0cp9LjXVg+wvm8NzYzccYaPqGeIYdQxqM/48gTsX/kuXKTXcc/aGBjSE2+9RE+r7o/5gt4FoRuwQOxt05aumCf3DZpTKs5jZWQ83+zqtb7bzbr5TW3o9dU0G3Ms9QHUcuNOSSOcz80nM+8+zdKR141TxMbqqjT/bFzenlSoGYkmjxLsy4ZJ0/PJpZVKLTWJ/9yNjVxxF8biYe7fIo+YSPraxvRiuS9FivylManAJztB2WO2qwxODWjbfbjrR/UkOnVmU3bX8z+RSMA1WtQNDJOER0BCJ/P3w8a+HAFR211APX+hRf8tmIlIn/DyM+lf4MdinhnbRK33dEuEOMzt/tBT+g6jasIHxCr0fpnSsye7zol03Qq8k4lGoiPn5wPIqJfzTU1+Bw2X/50/AA19tJfzWVyrRlfBatpkVYoPmw5yaFMQ89jjCPguCw/pmcTboTX4d+AmnZZdm5NaHrLzDFUUzUl9jBn7usjXgNaxxPKbrb6CyBDLpBBPOgsomFcHr//ws7BB60I+EF71JaSnbROaclxm02pm5vW0OYCCyVtBHXewA/fmkHLiyvg9+FIaXqafUtcQ7ysNBgogDjH9f2+ol8Ae2BdIrCTH+XiSPWK/REKtCJXKSB3hs9/rAij5htj8hUY4oBIZ+YcCkPo8Z1/TDQ4VqZaMau4YDi/haI+F+FKy64XUNh7thx+07DJdxDrGQjokxZMDzBHcj1hSI3HaV8FkBk2nhIFeTQ34iSlzgBcQ6VmIWy4aLUgRQocsDSBGqPJ5NKUD/97D3UiukgvMJNlokGKINCHzVUtoovNkpqIKjEfhfHyShChkMHBFunCPg+6nJSYJbUTQsg1PY6Z0dgwb4CGznT+f41VDJc0wfcV0haOoVeOe98p6KT4xkk0OAtKCvTh9imtDMOrtOtB2kxKKay5TizwR4XMR3/0DWawClQkYej/tfLLNjroRkiUAy5pgDj02fsolfnSE0EwVSh5dPvzSQUs5a3/gn/HFpqPUrWWJoUxgtm1Lw3Zmx0w96n0sEZUSyqILte3VvBXJN/fWxpZxczoDAHPjvfioaDPxUaTmtBLT54Twr+TzQl4sYzziMa6cm1f5pguLhKx/nkpBKJ9usOPjbHClD+sxk5O3CLbkDjKDgweevueEB8Kw2TCX/KIveXRLFHdUXgKDzNms+2AYMWFLwZ8Qy4WQKv2G9RIwtWN0et7N8nRSQLi9bVE4bGwZDmzXCqZlqOoNoLLjGL/ZrZQxmJnR20gNbu++Zd5rVEtYfsWcj8wvFgxI87l61uo5k9LrepEN32sTULiwTE8R7c/TYm3K7X6ygTQQurlQ7fW7qOWkQICLRlZ2e26eOkyNZY+lb2T9FbM/Dhjvh/t9cxcfyVRCtwVteW8xqJlHg2E3k0GFMknv99fDwmEYzdE7x+u2LBZK0y+/2AYulJARF0Yc3HRWt6zPxihR/2ot2MtD3ZzkZ76DonfG8tBNntu1NqgbkQ5dOSf40rIgw3df+r/N6h0yjHg5rJMSaebGF1QKdPMDY1VDYQ2OUIId07K171f6N9Lj/pAVPyOzPvQmKnZqV5DEyjjLqecA7kl0ssAsI02eZDoaTpUKditq8FN6aHP95It13vTsjXwc8YRlP+VqfOk9p7YYOSZ1jRzDwm83oaNwEv/HLmXC0bnlsk7aMu62deien+TWiyTfEne/Y79012Dnn8gSYwFvWW01B7mAlJ+ZwwHv1KtmsS7zJ6RnFkyTDG7ADa6WavEKYs9qtCA48nmKyWJFEDp5NtIFizuqyAVCij+G7h0cPi6fHCE+MSIacE81v1hVPtYf9qIFCGCIgVWZ8lQd3mkxLpTbVEb2KKYz2uAcuExsy9DUNi2/5ct0vW5T35FCIOLEqVWloXrb079dwCMhvsIjF1uCuqhx0iscD5UXcYrFIDCw8LdACBnoUX3OmJiMQ6OKqS7l1D+UTErH2RL9EYfBpE+REGQns2vDkyrlOPt4hfXiWVJWNLM4NOukUtyGsLDFQCN+GlhixYez6D/su7BsEd2kmOaVTNm2ov4dJfXO/vW6ze/ka+K0QMZENKVc+bA2o9CI6pXgLpdevJg8cJP7REjZ2hgixPYDhdYwRitLbEhEXHmYoCX/1z9M1hZdbR66hWdGBkQzmXpRV3p9cWcKOiO3+pyGjPnyEulsROlqvAKbEnoq2VPsGyuDR7F1Eit6Iz1cNLDO2QG3EWAlwi00uw6iJoznBT4HHxdc7KKbv9IpudbnsgxRXpjx5p0uhC7hX7e7bEVVYDzqScLx3iOwNVDsOeuKMOrOwnXOrLF/yRfy8trPH5q/JP9YGuvdEmNv9MW+Uhig70y+2WBRfDVCSWx5Ebf3UbU4cAdQB8IdEa8+eawfmHqCU+mLc3DiqjlqvgnHH3f5ys4LhomOCGblk2RKByossHjSM7NKctZUwQ/SIro8rZPkJ/rRSulkCbgazRHsY+oznjvl5LkuYjc4TuVV7+Su72QKxl54CkkcMiU3pqrzCMeCpp/cPRhfKsU9pUGylPxr4w7NfY/kje0uoGlYmcHhD5C2vyR99J9lIYmMTfO6/+lITWkLL6Y+iZuxgcvEN9Jdj+trpJWa79UxdyMI1cO6QeS/3kz5xzcX+WNhcjZsBCXnZ54Bg3gFKGyJl0qY3dYQvsnuUSxekDbGXOaSimo7smCv32zcNaPIZ6/MXfx9TbhO5KxcWP2DGwQPqJQclX4Jh+bjI8lXCDv6XyWESFbkAu+UKNZca8oNJo9kZeRddOmDnQj764vsphSrzBa0AkncrlbkKLOKQQ4xd6jBfQWg==
`pragma protect end_data_block
`pragma protect digest_block
251f7fc5b1f25ac0335085b431c7359dc50a6fe645aa9fbd25938a80a9ab149a
`pragma protect end_digest_block
`pragma protect end_protected
