`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "dc6cb4e2e63b50c3661660de404d2797"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
1X2n7P7bJr8lVEbywqoLt0hHgixWIn+nzJ+CX/hNtp0weOme6tnQqqebQDa01wOxMPSAqYFYtAI2hsV0Zqa2qW9ta57t3M6Q7BbsfBkQ0pgy7uO3oWL2GQPecyMLSnexDQ+dc3aEIjCbO3MDORpbGVejs4f9PUU7iMEg9cYFV9qaPkmsl08PFupaJ0jGB99QOzafCfaLXBVNU9muv9f545FdVu9ENhmjuB797AKEA994LlTZxlvf3MyinZGUCdbbuHpH6cXOXYs9snSfRT0x1S/nkVrexXWCXw5EKvkGTeNdw+RImrkYOaXI7a9/U3bvLYYFhCSe3QhmSLkTR8X81Dicwcnb+RZ/ftJ9HB6h1WXeeemUBApkhfU42ucR2G5BwBEZaZKmzPNWdQtNLOb25cQTc4Q2Q2grsYg0AeFkBnzpHX1UzOjNbo4A2hNHwp0EyAAE2eUNLTj2yeUls8i9f6xlGbCRmmNNIH4Nh/xDUx0BhPhv2ksMtkW5QRMfLjc7ruzqJhdDDrUus6opDMXra8rju0qCPVBIN47+ELwkUoEAjlvMw++K2IQc0fkyb7pLee6/OIcVQzNDY4MB+bpyzm5+lpsGMUBz5I+n2NDOACiJJpKQiSGhLHkteGRZ91gXpIs/bTZQQfSyWze9s75TV64O1/7J9lRQg6Caas5UfaUmPQAcmlBQ64MHmKrLP4oGvIzyjBnIqGkybFZkm0H8HzUOjWV+rOBqMQOln0Jm8K5QBp8Qpg1l1+xVZjMjAT0nrhu85cvtyiPs9gxOELy9T9R9xjIEJ+0A7WzSCF6huXVKbfCOmtuAT2Vnb3YxjoxhsY7KCeoszVcpaKoDeRhES62LbPQs9MjbhTCq8R4Rg3qNw0hnCh2Rb1kGA5/7gbzP6A0VI5TCaPibzXVger2RBL2lzGqqskDbnQT/h/gA7OnSojhOjr3qr4dYT8jspKpBwYFoPcY+qPHys2/gRm2+tszH0nJ3ednxblG+kZm5Drf/LjV5kl8JBO3uaheBq7YqMpofZ2LhPZG+/9Ihwlxi1NAr2kD+m+z1EG4cBrlewGOhR3D+k+tg6jbe+9F4GOYntoBWYEMHkMwc4z2BgDYKkesryaA5hgcBkTIt5bxKc3K3kcEn8ZP3IvEcHxFOWfVqNj/UnyYv92o9qruYsyQwV+UbgzAo9IwtYacYKwNXKQczU+Ukd8XpFj5XgQfWmjV7npcPfslf576jyzCJt1q/+lutrg8FqDNj57f+tX+hEENASipt61B/7vPfhA44NzJhoeB4s66SUzSAMbLkdiGJldnEwVW8soeQnBriuTovNVcUJYrriIWhqdtEKTby99DcAAPPSm/Og4pDxMgOK/xz1qOIi/KQrbv0y5SuNcDvjBMKpkf8xeg4OH69hmbNS59PQvFFgPK/FLkzcIq9P59CKV4Y/sMS9sxQlux7FS3PWJFp/24PbRHvbJIQhGlvQ/KUA08JoOVBPNZUz/UusPR3lJY+i4CYjXuUB41pAWX4QA1e1K/zRZZHTaJSEw79gcSef89Q/D5Is/atTNwZ7e9CS+WkM62An8O9YIS9cyvnbIdHXruZkfXSjbEQDniNoOgyCjsS+LWjwh+kemHeOZA4UAg51r1nV/5BNsxOrchW0FoipG3+3qJ0jVjzF2YWR+1S0k/O0evUlMIEUd81dz6Z2+lhQzwmIkIlTuU7NR+40je5fjq0mEEPGUXEHryxzFNPz/SmqeBfqVGgtZQ0PGGlfovNaIab+UJ+OCmOx90+3M08CcrNAYH4qjstOODQ/TUXV18tOxIur66CvldtFhQsOhqH800KnD+bzCfXXyQ8yZdfmlYKnT36UBtOnJ7SxnJU1amRyOQwa3R4EHlshZ062Zs00GnmYxOHhILgblJ8PzaL8vy6J9tDzp4yY615XpiMAa1nIhh1bsYIA/W/3wMziwz2OpGY3NUW8kXCNDzb8/l3ZRn7ecTeljbpSQWF/pMM1W1llexePTbOruGB2bN2amkcNv1C5xINbptwBcRpuM1VpAUOahpFTRReNnKbfhI45WFyy+nGSit/egWtioNNYyMoq14QwyMGn5Od2tlrEyi7UYdSCrxMYUTvcmmr3XlaeMkHzTksPcE3slWfpHs6zrBx/8WFRzy8gC+ltXiqFXShnl5fu308Rg8YrGgHvv+M7myXRDb/VAOgzoCr/GUJYGPXhcl2xI0FuaSiEmLCYHe6bunKtVGrDRuTTq8GgFaVZA9z1zJek+mKB1O9ZPaltAIVNaaIgoelBcmnHd8bGczOoZoCX+KQMlJOxFOAvI/qfJGGEHra3xsfP6TK42ivHBWyGKVeiC4FMZCTznfs0hyFCygXbW9XK4NztYTsJFfZnAu+LAPBV2IC/6m3RVKXm5fC55oVVGipjIBFzkSkKG9tTpCxJYbfy3NeFeKRp5Gi+KTkvc0M7PhQNERGsbTr00l9VhNRb1iAByug2YcpYitmMZiJsIG0OB+RKgoZiR1f7qmxbagd5qNjRHRbLg2QMXLAjulExTWSsnNvW91pNZpQkgg/dt7dxK+dnOWie6qMd+0U2j8wtB1HhOga8y2rYm6jZx9cebvY2bq116O1x9v88jc+MxLItgvreoKcFTL62pJM7ALCXMCewLkuceDvDpJINhbRmmlZPl3PRI2bih5sxW6yIxoCud8Cdf4/BLGcVKsflmp/Q4Q/KNbtgdB15n7a5nILEJmZIHjey4Fi8OnvTDC66CwAhvLfFgon5yiXNqmqtBHsWsGUu4mHboX1p6V08YlZrrqaLuvutslJexdpVhtF5RbtAHMOzDEKKXHFqtlGGEkoDtGLVz3t4L6tXzy0njkIrZUEmILoTswlTcJLcFch2pX06YpMzxXexueHhf90dSbjqugpZ7/+To/2z+jc4HmerEVe8ZsDhzYkm0J23sKMD3GRJPPVf2Nup4S7P9xtyKMqC7/ZHzXnykZU8hxiRZvSntbAVZ3J44n7knVN7Npe4Ky3BvMRaMtaQKgq/g1DBi+Kr6I0tHE1wMEhMjxqtJlrHhf7SgjH69t3gyfrKhQOrtceQU6mjnIUDWHvdzGCyKCeYiaudYW5N1inT6bfgBxS9t+3MeJjr2MJ4L93SqDuqVqinL4cyRdBkWq3rF3silt0Rx+IPzJ99z3hMmeqQuQtaHDdTmBqWk3ISqCmQ1Osp1ifKwQreio70BCwKn+hiRxydXng+EJQmD/Y/JRFCgMhPgWD2Pfn5pm1GqJFJG/bb4+FFgDtl7gsK2vZ3TnPfHuFMzi9MDNjq2GDxs283VAQ7pi45YUcpgVuUPoLrIKgp7finmiwHGvqvh5VOcb0MCqhV+DY7xpPkCKeTsyTGeffsitXvpel4Dn9f/PmeIKVX+oB695khnXczvnG4Z+OkwnxFzm+jKWLhO26nOjGTP6KJCSW2INp9DIH6x4M/L9nxFbGv12gUi9qj+isd34oW1/TOs/w9M54jVf3YTXO9QvYRyx7/IKeH+DTT6lKYHk25cMsThXrTmqZtxaq/UeXpAlCKPtP4RCx0evDaga1dwSRG4qbYLgwpxgaQfr5BOQ65G7UcIOI4hyklhDeH/K6hbNvosFQh38kvfavscFIs08649oiwdfxJ5t/dZmOTWtHUX4iMDWg4YIhLGQbEOYdNdGUpA1jqPbKzkZPZn4hCu0pueRog33KB9NN+h5K9fLAI3umxEH0QBcUj+qg343EF4is5uj4abmLsrvTNWAlBK1dhV0bFIUXzA6icSS0ufsc5JsT/G+bHsUYbTYyaVSqPppEtqghN/53wXXcX2a1as+p5xGLOURiyM1Bj8OmX4g371eHGHCFAjSadz3HFZzFop+AZNrMZ7uZYiyrjemrJ1Ie9CFRjAelcCrdZLUFD+EQbXWQv0Cu8Dl1u/cGKVkr/ybZU5TtGmDd3otFx1z3fDr4LpVFDwLZuYHsYzU9X15U/ydHC/bqHzRnDhd/mNrWFMuGwwTAryFk4uzB0q4Nmw4PBzOoOtMaARBbDvARCRkGTQzSgoCUaaK/m+R4uju4atUxDHdXE4msiSNTddjgR2JH/f0dX9LhT6GOwDMmZ5G46+GylJyyd8GikwybNj6i38SUnUI8HZ9luVJkOO2Oz14mX3XwUzM6H0eD4iNVfLeYlsqSqPTYII/ZH5oIMzJ+vudnpa3YwVcyuGkTQHhyfO9Yf2Rjyf1SvXSY6ZyZPKsKFGzBDSKoOYtIqyPFXm8FeKQAQ2tAV64tLYmBUJh5JKoD36Y7m/CTruHkdoUALffLgMDz9SWZeOCZXS3Yjp68UKg66Dkirn+6NjBKsmVydN1hWEOBr+LWeInT6vXbZUwGkOzdTaG5JGZ5macc9jQQSSHSJECqDBymfCY+8pjOB+onCEMta8CyQkyKNkaVjAMqVFw7jZQwmrTNrpCXI61cKPMvCTwkllCPcKaqX/KV8GZZJVyRgQ5eF2S+5YEiDnecjQ+90J6KH5sj5E7Fs8brn0Nh+wn28W6dK/fG5BQ291yF2razNCnroo6ZcaSiiIEJ7Sv+TO7FImDp0MsshoH8Ws4rX86iZUGTYCNo8HoZ6X+CQYvOJ4eHJUPGsbB7lgEibdsPBZS9HxmZGSJv+9pAzj2En9PbVXlqLDlBFVEk0Ij2CR/OzsxSHBWeOu+XHBJH6CvU1mytMc4TRKAEDH63nYZAFXiIZ6ETxVltxEc4Eg2ooSWWmBA7j3u4RgJAD+Lv0VhBO/TyF2PQBj7C4B4eqpKZa3HLOHh0c6qcfdQjkBb0aKK5/109OP3ZYNMyep5nFsSCiHEdD9pOaciPCVbaCAdc2LLju3X+3D8ETpbgZJRaqbOYUTJSldvjWBH64IOg1SRPtFCUvCWUjgx07qmAStXdgCoIgEJUs/a9rRYPu1ns25FXq2rho/5qCX/WgDh/YE50aX2G4yb8tQWGNwX7RslWQoDOF3r3j93N3lRvqTL1ZDihjIN1ARUcLp6QoZnTkXgDij88KuWb2wohO3Lhh/qZuayBldrZV9SS9El0nLkqPZwer1p1pVp7x6pFeP/4kPpj3FCbuI4on33e7DNbOm9FlJXVhqMISjyOTeBtC5qou0E78XL0vF29HB+L011UvAGjm3IofMgozOwRLqMpHOuciiJBfbWS5OyNAL9Q1ZS15zSaYEV1xCC9JMR5BDBbLPEh8L+kabpE4Lp6h8fpDDAS4FrsbcZAXzeLHP23zVgaFKKlXpd6wymnRNex7p/TIwBz7S9ez1o/SqAJQMJWztfw4F/YjCypQHrp4BqAEY4brwpaq1iTcLc2iHRqdHhFcZ7y/0Sb3SzDS9TmOHGBrt1UZmM/Gzmyzue9+1Wj7ekTmkyMNiKQ9TcTZuZLLm2mqfhLQr2i//wV/GSPuiHd57Du3U9YAY/CdV9HgpYa8MxbuaW2tGN848P4YhL5Yd6A+ev0lT+UkQhZx03EB5CaVauyRJQ8kuuWKQoFZYeF4Z80zopKN9oWKj54iXMq5GTsuLO9924rHZwG6Wy9lg1cuBMwIhE3s66KaI8Hz061qp7Lh3mgMHBNrbrYovFnkmsgNPzkU3SM5RI+Cm/cZxwFdEWznr+AaHREvMGImjqerR8aTMZFtusjDFv3Vo16TbpiCEfgIEMA+FLeylIeV3uk+p4rg7ADG+kEinuxlVZp1Y+C/CfT3pytdakKDLdKuJz12+aEJvtOwnZlijYJwot58eKYEtoaQCBbDWK8AhFpAmb8udhCvKwotI61QettvWpuo3KFC3VOY3K/9pNfaPMOxh0385ISsz9DNUm/2zwJjWIo4UEGZBPJrsDEwxjZEXWfRCNN0XFc7vn//RSTKtGxS1lKQdqPVoH4zMou+zTUNRhlo6o315zqLpoV2prZzP8zbPqY7Ap6VWTC/PxtoBgmjpeJd8QmuSZL9po5vThlRi4cqdZcCjuX09C2e2EZFMbjF60VxArnbDf4y057ME0VoGn1Hy5I2aUtpf8WcxnL6hUN12oKm4sHL6UqJrLpWp8kR4VxZcfccpKzO+4DlHp0ZmewDMaEYYx+yDOaNSCSOwMBHYvDqQ99AVqAoSJBlKnw2ZMY34Wc5bZpYVbbZWUcu0Zfes3omqlw/Q1nRDav2XEI0sm1upUUiP7/q+oIUg2FwV8Eiy62fdGQ7vR11+3d9ww1CQTG2H7xocVMdNe/mwnm3j8GiS3W1NABabsBlqovY1ZTy4f8h50YcPNdHcjmSvhAdruV8/dUY4N2Pg4cHaZoL2t7d5hCJQlQH9tfhgKXrHPje8VjWGDu2I92MILFNeDTFjMXsKtW4wWVKihWS4tiCcM1CpRvIZlX4iQ9E8mVCRHVEwvIWBSCtHTXDd5AKBnRGPDBIoKckp5WBRPL8F7x080Y+ivPTuFampDmDveKwFGwPPydQm+5ucordSUDjziw8ALav3Gnl1fRz5kug5kenEUw91mTx1FTutWsK6bfuUeuTq76fm0Q6ZtqjdqDuFJZ0ipvBPHn3CoV3nv/WTmXjruda3Q9OvogkfbSfZr0nVqD60roXXU/yVBum0SrvkHGz/px2qJzIufHAiBu8SALAv7cjjEVwuzw3MH58DWpYaQTV9jT5/GgHN8BX+LneJrNQO/hjOchN3ovqR8hxCsZDYq10+n/bDPBY0nZLnQ3cV2J4zUkaEriaUp78+06sEmemnMCfc8qQBoPpxfL/X2m3112JHcnToyxqEgV3CTAHnP7W5FP5iuAeV4RAOnCKnjgzJ6gF2/z4B07xqYTkQ8l6Nyi0GyOSdYfhc7tn2JHvzpaxtdfTY+gNqyefcQTac72u/qdR5v96efZ30X9IfO6hv2VMa/RJvks3nICXo+/GLeQUjlw0FtcK2GIejtIuEobGwhPCK5grG8wKaEBUnPuB2L2e7RuPwc5cj4KSgMZOetrTYOTGoAkFBT5IVePewLxprI0cnz0WaabNVFDyvGN70BaplChUy2u0vi5wU23D93o3DRsKlTQdi7jkDVIzZ+lUEU9DR8vo3bFeJ2OQ08kYvmHQCOl4pGc4UVqw7qcmH/LlIdgK5gqjAjtocDBGCt/MQRahG7J6D7FWXLLqAVupr1Z4mV6gWk78VrwutoNGD/XomyCIzOydXvLLOCsXn6PscQke0fzhLcwjq9JMur7Y12EhazoOQXeXD1elCSAXY73hxRNcolTv1oW9BUYOM0Tm6gtfiqlS1ddHVg5yLXoIUZ3OHT+FNJWC6cw8fNe95wZ6lvxgQq9CJNyZlXGanznSAKKn41gogdws6+6d8BKp/nOMk7MAKWVzTNlKwzYPgCrlYqIWnI+cuyG0wZyVA0gfwYoYKfFd4GDXk5v1k1VVa985R2vXOq5ihY7L03+qAtab+XC/wphEciST0aGKa3Mop/zu9YkhgoeWC7qIZmsg5q7vd6whdC4i0MiTfOKNRzlwqB/UTSX6nAUKrB1jHduBXfza1lwS9Ys5ifqauDJdom7vgVjBLtFpUq90ikVwer0TyKw/AQGInklA0qAt5kigFHKoMwpJgc8v/6hODSGxr7xFL3L5LalNkv02M1wf5KR4aAz3TeCBFbywDq4Z4ZhcLNJeRuBXO9U1u7WbEeWE3fHZH3RWmUZszOSSCBbf52zXoxzHhR4wlZC0ss648sT1S0XPygIejnJUOo1G28a13qYz3cE8mw3qvNNmlsbGWvjBXyQWRKe10A3CC2GC9NAxiqW60h1LStRoEOgIIg4/ug6l43tN6gD8Ie2YRF6F50mWCgBqlzbG4IaaAPWsGSFttxUIBlUm+roYGrBmuBQRR8qDjRf3otphgAQdsen7/Jrg2xDQzhhQ3ZncMwVrvJ/zBbH5a+gTIPLwicd0J1hmq3WgU2kUksd+DJyr+HSYBTYI4lbv2T4YjcdDfwpplEYFmCZjZaYEPQIfihyL2kZnHQd+bFHXZ2zPPQH9z5O6DoluEIqB203nXI0DBJYOD5EqvnwXy48PdYNTVjoEa3NFywimoPZ8UkVWCBfUVxps5If+RosDL2OKASymNL9iNkewYBT6wGMd3I45PhcCkDDmiXVwKfzlZXcuBHr9/UX5xe8FWzNAEN3NxScC1HKAD93GP/Mne9dZoilg9qbB9HOhtBclaQ08xprHPnINB+gaEbhP3UXKIlYseJcji++OAgv6XwtbSN7YsLJ5k1/m82m+RGGfsn+J+W/W/G5jciw/WXqs3s2UcODrb9zhhZBa2MVR25/A547FgWCy78okvZ0zwe5me3Ww2Wc64Ne7t4agP1q7YOqIvARd+/VioigfgNHtWG+XEfEaBWhBoPlSKLEtIstIO7dQLZod/Z1r0oM1qNFIRVTNQgEQylsPqkIyKVSyjWdjsrTOra0/sxOkUk+YQncF+xMYSmkHyDlPEtifPdyT2n2geQBOEi+8pOhO0U5ZwA/Bz+Ojmo+oBjU1XP2LqDSNnKAEwNqtEF+LckvPF4KZk7Ic34Nl0a5ngINwuhIrbaOQ5+VSp4lxgenMUmJE7EVwu3nwaiDzZs7W7+T9vPrdkOw7X6p/uApDvEwCOES6QSoXSrl0HUVEI4Gi4j8z9OV2Ui7MSO4YnQKGAfNaO1N5CjAqee19CBRpWyyWxOqhklsV2i9pNGjBGklGm6Ux6uTpQHdgOBlcfRxeA+neshSZFOqItWc7G3EFObP5f+4CNoQe0wUo2A9/HDsNZLYb3ln6WQU/+f+ndFGX9B+vyNiy18AuNpyl0FMULRi3nCoZtKLuX73BDfKMPbn4LFQO6TROvIvagMMWLqYlpdExZEl3jzuJDhAF5zxAxEN4W6qzOrisijw3b3z/uFZDNlHhg16Mu8ePrDJnQZVvjnSSbYpKV3O+1XNxf203jwAKgdpuxXKb+PHXkf1N2TUaq8xDWo3GajUARJguWwnEYi6BzOuze6K6lhbYdJA35nCXz04SRl52lMb8AEU24Jr/j4iJLfAxw9YcVUEl6GGYkdiBzLFQAE6nsTapEc41ahIuWOpbfJLtlYFk6aRz/DnTE54uvnji/pkdFSOG1Nzu3MzlsDmfpx97SZ67ltQYblpsnbVZDi7EIOJPOWK8x1J8PlAQTWIt81bFvftHU1xCZpxBlAugH6coR0/xm+YAg7PAZ5JqqFA7fnnnQhqJLmYELKUHXoTphMIwPcr7vzyRwuM68V2MbzmovMqEcudoz3fC8I+qoyJb50itDxIewmila/Chihg6S+SCP+K4k1hh101OH5dv2tx0Tn7Nprjop5pnLNFDJOj94SGi83aLu5vbl+ME0y2bnGj9vsrd/oGGHImF0V+qtIkIgI0xO8s1m7i2esJx7YvkSFDL0LKqHTNGV6dHjxGOqA1QzhrN+LGqbFxUw3oXL99f04IgMrZfgKbTCiT3w7nGYxFNnvCeedt813ehDuKoJxBQpQQ4tawIUC+Yew//AR5oiT3A7d3+6bgN7bktW16nnLJSytuD7mZqaXC0Z1iZ0M9qPsYROtudK2Y45XstIC/AyPQNdNFAe8ND7F9lhZiZaXeHr/NAOrnyuHvWa7+T3YbReVV2DEriBbsfi8QcmUUw0t+oBohk6w6ZYGZUYfR0GNNBZZ3Dn8uRYG/ZluPrppQk2yBdt4OxX5Ahpw9pDj3ZIBGeNnMhN4NFZY9Lyr428AlWMAb9+TYHyWDClbSkJADe1W/gRjsiv8wPEwKDz/vOJjqyqCqAFp2CDMXv9oLLueGWxWuhEs73eLN6QttOKYEPA3heK+Eu8woZ6HGTxFLgByqOdvGVa3uyRfZdqwc25ZDKHzKTFBnTNKOnFf7GrU4g1saOl1uCWwwCFW4ajAhnqs+hMBcAR5N3VMAXXaY4OuO2xWcd+YcLJ9GtADHGyjyJ3C0OYcU7Eu0ciS6/BtQCMXs7v2+XIqdFcUNj5x6BPlZ9oyStFJGy0v9DyE0iTzRZK+peHVqpnW1PU5q2tma0MS5sM9QhEGh/vFew8eQ9otQUe3PIrid9pbbNkH7kKazjXnJuoFOHTvBzJaqkP3xsM+qjc+IB6uSzGm5xlCMFdvweN3DSMsSoRFUlDku1AvnWXmY4INALqN+aUFbqTEWFDhi/ELW+gGiI5wU7uUOdLFF05Les7de16/PQ7PlStXNyxtbD+186UPM1NVIzyc9ffQAA4AqWME9yLbINTrgG0bx8J4qehjuZX10L0tvOgF9gE0any6sF3vsstcY6tsK959FhbdKDceW1KNDUhZrYvH+yQyW95hq99aahbKSUG7WLTBu7N4Y0RwmM7YZ8OfrTxm1JamJqEVUAUN51s8Fvizd44eH5Qh36ElH8Wtte8DL8GtK4nXr6WTyALkDRzWHD93U4wCeOlRo15+KZSHnJo6DAJ4fu02yBsxXlLO4mVB5CXvMw1VD/ugq9/k2NoLI4Ul+mtXy/ogMDeqldYkv2bRlbXDJmv241v5SG/LL8i/beZqff+n//8h41REqrvhwiFA+UfFDN/SR5EXeqUSv7ggcYcB8LTBMNR/K4Hrm/QWQP0RFwKmrC0NBfq1DHpTAsvTPRK45MAvjOiLmhJ+glQxbybdEa2PNN9mLMLz69cbue4Jfd2bGtSDYn5FX0FNGK6Ggz+KZrs7zGeswUKCzVJP6C+uL6rFF2BNS9jspMJcY8jEsJFuDOLFGDveOtadBnsvGupNEiPwpUOl2SXNO+bI+Dbmc0UUoPH7wzoXyc2e4E1lQ617eiqPYjc4BpZPX1utCn2N5LIZM1cqbIB3KDVgnPrg2N9fKoMyYULOe8lRsBBIi7z5J8cy2Vlg3ZpfHAU0nJr6k2vsk2ctes0+tEO8a7IsSS/BHX4efLFgg8j5pJz0KYqf6Kb0rxf00k5C8mIlDSiEMmdm6VV6vpJ/nkqJ52oTZXJBBOlSHKuNERlwxHEBg2eHgE9L1rus0qUCX2DhNxy0i+pfgNfdEHnOTcwKX+ptFGPHNcULlEc0JnEzHo422sG9XLRND7qvUeHChE6ku9B7Wyu+lIn5gtevKm5e6jtrHX+MoBOqZufdwmhuWVuo9Bd+n8Am7jlh9bnWsRT99yiOahHr9qutJ3gaAZPLzoOdXeoC/cvWNITh95acHYabX5DHKIgrca1c6wzMbUFHKpIjsjLVJ2tXttVZ1Bvk4lU560dSFzAdlJlumjzNvS/yxJravR+tvDyueN5oChR691o/tBXu7xbWxD9UrNx8dp+arkVq6uA0vMM8amzmB+aCtWbBp1jnH34LKzZVMgejRQR2HhNp0cQ5y+/KiU7ky0GtFm0ck+oloNuK0NA5AT964MrPXmzsdyuDKc4OMznbVCY8KObL1fuq9msYvXUk8fjOCCS+gnAWBeRT14rd4Ydj2iJYEMu439fIplIpyRfsJxsmJMzF7zYmUIgwORVWOAQOrduJty+bxR91JPgU/cWTadiMuGethGYqmIlJu9WzyvBnIMRvXyAZgGYy8AGAqywuAf94FTZcKL2f1qFKe57+DZySo6BjyeERjh+dcWHLO/CZZ05Tyj4vhjkaFqbodoOHS+nzscYTuVwiPWyJ60nKQQJkdDAY/W+vpWLEhRo6NJWwRextuC3PiZIMaJL6pqbtlAv9sym9g0JEexHOHRjXojLjpkdXBNlP1zRG3qpazht6Zw9FXPWY9dZcLlz92+WiHu8xMQkZZgJN68Yk0loE5Qgz7JvpVMdkfXOtWNIGkw3LroA7y0TcVsIhrBnRZ9ykvMwYR5wzDq65ZyRTvpMpqldt4oy3gIm5+oHg2tyXqKXD41VymnP0hIn/dPrphFbf7SV/jIm8KBFp75yOi65qukIB/wUBurC8QCK/ncuikC8/NKRWhBh5bZ88uK1gP9diFtcQgNPyKTWBOqd8JuJJCw0c5ByGKM6EsBuipApKlp2lucjb5vV4NSXtAw8sN2nhAD5vzjPruNtKtJdQXMcRXHRUtnnNroXxeXkdnhzzZhQqMLhtXYB69oot93+XpLpZsLGN7vl0zJbj+XE6yD2WxlEisujFWUC9GOZd3glfSLdTua8GmuCnfBI/4Dq45wGOQvn1ED25DaFYZQTVouCdQ24vuQCROIEB79KKbiGKxeon9Wyqe9JUGC8qcSiwWkdTAKHzascdbfGTiQbbcKIsP3h2eD2FBf0qQoob4RhE7bC4OcM3JBPjBZGS8NdbQf7IgPnVbEOJr26Ejxnps02M/6TCMgh61eUZWPVwY0WMCxPNgNpu2N+otqz/8b2OpUSIvcYddryiBLBYpWOurOcs5inufwUdiyO1QYpHM6ddjlFmf+bhQVtRrZ3B48LnApBwvBo4FNQcjgMeyXDyQPr7Jp1BBcTvljsPViPk4ZDjNmYFzits39Drrnw7rD/lvnBUM74U0xsaOgBM6JaNW3X8838bC+I8FQEnNwp5+L4jLpxNceckK2g/n9hWgIJrwucKFsQ2AoFCF1ENeA1ubPdoVlwU4k/z8jNUugbjEr4hgkka5NrmOkx0+1CXHbA2k2dV8pIKZ+IqMMea8s0M70IuuLAyPj+ntoeXjokTP09rE/SiFZ7OtpJW6e2Tp1dZm2AhjqNGAZqS9pPIpTDxA8KyrbSnoQ86KbLCAqPZN3QrBiWyIDRq2dneYNPEgvq7A18DVU99mdq735/O1AgKe2mZmOFdlkuoSm8Gk9bWZCTHxVknxxmOSPqiWMdjK4Wj8U4DjHYF2VNhjgSy5XALkk892U/JWoNOnXbUzlekI/isCvd4UKBISDEx4Wv93Hs1+c+6c4NFsfms8OG7K9jvchg2su0s5h+FopOM0k47WzGBdab6lRdeorhxXNAH1KnXqctDgMUZ4/ZaFjuq2Dkbj+NnPoxh9Jk5g4ny5IcBs8bQ4C1eSWqOraN6jpJsGLCaCg8CPyXrxaE1MSQC8A3Yyo3/oXpzARIZDdItDuG7BEwllyZtQ90blrVVjTO2Y9xen3A6D0tj3WN+EELfQ4VzSKZYW1hQfutDAcpGXvWsNHoLg61YTd7w7cISE4yyBUAOVqqNa1kLcSIRp+pKtj1PIFV+i53xQ2gSKSFSJuEozuRfyYXzmloadlsL7/i2fa9dmIgZUHzW/RcoLvyeHJ3OaIYpyh8hROInZPUGHNLNU0QpkLMsUFM+isI50f5IvYBAx+0ueXTc+UQ5ACoKG9NPZ/zkN0/4AcgWGBTnu2odlSSZqMBbT86NmIandGQqtClZk4lqAPCtZ+dwO8dH2bCLMN52ldDBOGIauNb5b4v2sGmr24VrU9/5Zk6jQThDYDzSQPlAX7Q7gp5rixDUAYuypMQNCfeT0ElviCKYUaImFxBrvLw3MePT2Ai1rUV19+rVdsUhOX0PSnHHidn+8Bd9cUcVIbHL3JJz42/HQOqP35qLYRuy3t5o1/K6lnSmg1ZJqhfdgm8YxtKiq9KMpu38cIkE7FqQyQZQc+qKbyugIkPEWVKUtOUm8DuuRMaJdhVLx+rUUPNavr7N8Wl6gL9wF4jMFT7Gw0YnnayTu2ZQmLbw/R0TmSK7/lzkUjqnFRU+IT9IBfaeXOrM1ijuBlNK6SlhSm25/mQ6BTILafJ7ifdClQkbmACRE6wgBPRzqKViNXbRZMRTqg5h8oi0X+gKMGx1SdcLz/HMBpYBYi4rZMwnWc8RPablTPUBM2lsxx+Dg8nOICyN5HF/800X7EqqpCC+Q0gFdfge4bNM30R2Oj84k5qb0TDVYxbk6W/PqvOoI/aajV3SX0Vclb0qbehyDp20tJNi7eogITZKh+uvjum8eZJdwTOSmTZwCrHJCLzj+PES1oFyGNhKKyrI7++HlMfHCze2IIPeq0cPKrfsnWLS87jEzP2kVUQROXz1kN0ZlllLSzyw0npfsf4JDVm2IR3ZXj5QmYa3/wAq6VRqoS7ex5AJvGsXRGu20JXNKkCag+5OT5LjtP4u9Hbxf1cBuWmdp/jYEZPnOfCuYJNpcIZ4hTAvIXk4fX8XSQG8cWqE8NvbcL3pctKKLj89oCwo+XUBCrvjKa36kB46qqRaQNk5neb9Jy3wyRjhJARFCswVeOhs/RYJOaqFH7MpljrwMUben8Ky5NKL4qTKG1MWPai8gqe6GNz+1VjHpfXlCJCfhe7jfGS72yjxYiwsX6gPWszAxWboHqxoFhm0GcoSI6kADMAB3Mu+mahggFSPVWY7Xs2s6a/wkesPRom1mzJ9yjIXfTULW6pTEdj+PPa3GSQXKfjhHwoFlvPyDXS1Ng9vRpbIhFE6xKwpHkNb19UZwl8bnBWA=
`pragma protect end_data_block
`pragma protect digest_block
80ec3a19c3793d1edd6ecf333d5e7939039eb576bbb54641e11188cf2d0085d4
`pragma protect end_digest_block
`pragma protect end_protected
