`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
HyUMV/wuiEQLI3eK6F3md7FOxUCR9OhOklHdh5gxX5ckP/zHcln13LR6nbwqyfO74FXeitzWKKI+r1m6iXzmEoSVkvG/M6qsDtPk0VwogsdJNEDrOc7YtyGd6Q7n0ZSdfDynkgnXUEh5SSt9M+560WkSghgx5shZzamq5mxWxkQ3PvoCaaEoD5YOJcUPfoMrdE0B+OgHasUDUv5BJlK1rJ5BLRemKMc3whT+uwt1VQZKfRJu3Uv/NBK61TkcZZxo+WQbCcs/KHON7viCiOXheErt9sZB+/T5RX4SuX0mlvQoIzH1O1UINPEBF5tLCWfpOiJ53gF/AXdk1ZvS7AsHfGj0hszK6Q4ANpsX3QQjfp3iABN5aD1D2Dt7ogw14vHMLUK1LgqyIJC7qCgdPJlH5B0j7DV1amIi+x1n0vmIRbDWzKJJhozmh6nHT+1mfGm2LcXZfTKD0QktFGfsUGQmq03aq8IIn8jW/yn504PUBbW/OOSPlU96kjZWJ08SE56Hy4xUsSJ1/4rNVs10+Zw8c80/+NTXeMdVuxJ6QjNi8K+YRA8AHz+d5JX96Zh2KTMucDz/zvafIa/wL8Bq4TgCbMYqO8WAS45y8kuTmXgutGtFHwt/UxtVMJXtBF19qFknTq9nNJD4yjaHBBk1NfTiR3ih3Us6wrZPnkX8N5uJBjABhgcOmxS5Ic36PklbiBxrQmRGAiUhmA4bX6DPYoLjVraJe4qVkagFe9vdiFR+hbP6wuBVSVUy584jKALVD8P47+2NXnYvVTg5nCEGd2vVqkQoaE2l0kxMnyS82iMq32Ido7Pzfvy/QwW+6aVl7VfCMXvYLNivFLoGLUzavwj7mjOZwJB5tGqmfcF0XeK5v875Uml5nOaKx3Szjt3P9+KvSdYvZEa217pqC5ksIJbIjVGStDKabUUk4zNqKu4aVTpQnVFJSFqNg0DFYpEkQV98zv9UpnbP2jSFaZO0ErMVwoXFSegxptmGs4+k25z5BubZcKcUMgJrDO/rWlx44gY3Qr2AKRNecQxqlaB0V31Hm08AOxuwarKck8Qsb/QSEUZXzjLnS0KnEm1Y8lGYaKXrO9EsHdRImhn4y1vQ3mWvYm9892YNb7v9elHZY/j+mNdBsul4exYkgvva5568jR4m06qkESuia+ueQmgbBF2QuTMmiSVFjI3Mxzw/uSKtfOCZM9btoDNYGov+AQm8rZ5efJMl6XqGC/zQG9IPefC5w0IFnrXdA57jNKKcZDXfZBacogEkpGgXFdSOThozjvRtIX/6Ltwq8usf9DkMENbQsYtv0s4ujmUZgq1UuIMZH5VwPvY41LBvIHXUj8v4NcXuOtrGwKreMdqMgdEsmnehAcZ4f1HUKyd/eMRrmQxT682wqjNkiSzTi/w4qX71LQgMnj0PZ1x1xn4jvbv4ZLZAu1aghGleNoN3rb9w2oS8xMo+JHr44qSmxf4WDM8QZvxI2CQmIZt0ufRirvxkoCWBuUZQ9eLXtulPV2iBrKDi4esN0REkDkym25DC0JUvrGhK4ZWEchYvHth7HrEb8Qt0jZ59sxNpxZSaDvcUYLUPqDbYOJnYO18HtT0BfD5mdavQ4+ehO/88SLi7JA7bYdCEP7v9Nm1dn/Hq+JUsGVR4sUTRYA1xswVdk378djXRfNuSM2tCdC7OruKBlXB/Y4hJp6L4tjCQLInJ6tGXdVTSwvGH4YEYxn1qZnYpWL8wrIFC60/6MS2hAgqa4FhyxJGNQEcXr3CV67mK8ViX1v6rFY3+j6/IafyX+a22KeE8cPRG9yk3JWa5vS0bvSaj8rgCb5yNko/xHKboR8ad7EaTocpnsz/5K+7V9yWTrsQ4aTCi7tnEThW2zPm44NZO8rdz14UIo3Txrl/rK6fMcF0hT2gMAzj4qQwZXxjItsj3zvL1MdteACNQdWFoPCD1e6X8vxxDJlnZjjZMjIZRZlE/m+5z9I7gDPQMpb8QDPioYbcIioi4EOVkmjOOvHqhWMijFPfL9+4z3pG+EAj+mSjpB3d+LQbWpzrKjq5ddpMTvEf/sfWzrDa+hgln/mGo7imRLsdfO/j3D+9WWtTbrOaWQzGSY4WYWVfkjNxz5cKS/+jmtRE9zxaOaM8ar8zxFa+/bSW3K5AM6iHQgPVteuJbL9iyqJXbbkH4FDMt32agc0OPZE4XtlMqHI/Z8Rlw6kRffqnzD7zi20SY5Qcsmoqgi19G0XcAjnJsLkUucvzSs43RwGpc04LxHRzBAbSKPLxiUlQHRdq2OP1uUgz/w8qsa5jOpcUDUOj7kewwHCndmuWh6UTeOjO2o92cABgenU+Hi8b/Mao32/nWXBKKBHgS34GJYMftxJDZg1ZQL3FN/qwylYcWcxKNRZX7CfbpKiPqNMnoq8c+GOMuP8JzJcZk+BEGxDTAMs650jBh7TUyLcLe7Y93t57xPApg5zL2x36jGvgRTkwdivTUEguWpvbZuwT5V8QdUlH9t69nEmmQmPcauVZtKVCgiWbxFkVBcZ51KkQX3x9GsONKF5MVe3zF/10cLy3pcA7/HsU+LppA3CjzRCgAbl9MaRURP924FbRWRqREmGe1wkgttXvcjd9SCo+Yh8hloBql7bbA5JoXSsJKlT0VO9/5TneH5ycKveXWi3hx0EPMA5AEni39PozOkGb/XUfjQQw4+v2SGrwzuBTbWM2/gSkQ29LfNl4zmIF10DtAURgHCDOJBxImLEZzoQsTVSH6XQ59LdwZyG/4ClzeiEfUrnJrynCKFLsLHD2MkC2D/fmUCL010RQB4v6GSSLstlLYej3RMUc5KMvad2UejLrNpprTcOfwAkEyf/hJ/FyVUYLT9wPiFYRavoGA/eYDPFET0ke6+SJ55nfjocxy0s6ZG2Q2uoUfdydGA/czXRGZwQQme7y5eleeTAgo/sy3Hv0Uup2McNHKvQ+CwEIJQKc66AzykeVtYWVvr+nds/c93MmN85leVuw51aX4PeUL8zNyM+x5eIEfmV1aVYEEpKsT+gpbUsyt6h9QHSvnHLuv0Ay48c6aobjU59YwJOYwety2qkx1YOw3jorxsylqzu0VjT5f7mEW2d3wpjMrX7Xy+B22u4TA+01c5XJvhYDq8WkOe1S3M+OCRgQiWL8kCby5msU/+VGhOCzm/XkFXZ1OvPzlQOf+TTYWrADvIMwUa+vpezdnkJqKm+wjZg3Tge/3VeOwiTs+M2QY/LY3tCfqwVPFzdU20TUdAJqDTL2q4zM2albsdLBJHGsW+cauwb/tejkrgFFAh1/UX9gAjmEUxzBWlZE01tAtaZtWu4FQwiH2uTCAuZ+aaxvkosbAlhVNfz1ea3kl/DVPwVhZWJCMr+ZychP1zoUOIBIATvDaqq9oZ+SY8fObgAsAQeD3vl+bM5bUh1F/IPKsaWFZIwfR42vyGMf359n7aTqSYzah1VP521M7YnEaCKuwUdsoVoJQBCzfF5pIyEb4ApR4JWUabJW7pPgC07NixQex29on13H1l12NejiOHfzdZ7Pe+cB/hsPnV8sIzpsK5021L/VoKTUztpSn3gy3VSGZSIpqPlMPIPjMvxAzmGp1C2MTHJe5f09q93HJuMx5asOc5rbR3gjRXVPxGkuAhnjjqON4QcJeIJaGVh8t3zpHLWjtRhPUA+M1y0rqcl6eqMn1HgxZFX+aIgmfNGeadghAv5X2xdxtBgrcOr84qt1fz68NP7uqwQTbM3w/RhF4g0B7UhQK9yYXAQb5Eksp6bcPciCoRwspWfeDQVkHk5ZMscOJZvgLxp2Jp0DUrxXoMyCn2zZ1PKSNc7oMLUXnWhUDzZfScloIpNkr3dVrPCYfbk0wmm4MDkpKMJBh6s0J0jSmaW7+D+OMg2p4wCBx9RQ13RRAz3RL0d+jZdRdL4naZcTyRdIq6/N/ZbaXeF7WV3wjLRdmWhSsAeb6TEIrwv5OkgIIRr6T+BfPlLj1Q49cc7v0PR5fVPOfVsBqH12clK7AAWZodvw6UWkgM/u7fXB3nVfGDOAtV/Wobz/ND/FMqGsCHSwAP+6P8OcQywA+OSWvxJ6sP7D8Cz1IdXrrRd82eNRkNDtglfRL1mKt9xZTbYVzuKxzNKxrtaQh7zXgcW4nEWBm9ivYQ+SuEkWAcJ4APWPvAV8Z54z1h10pH5YujZl7wqT6f/xlKYKJOtY43A7yZdcschaXxd44/AsEgqaiNTEfQ+hUznyg5JO/+d+RzRuWh8834cr0tFTsEjxx7LBBK/kM3GnzkSLYb7pdNAayD6cnGwvQYNXlikc5MmVExpeigDrSTEVFZevbFJ4gEVkphTbOjGkp0iwAnXGOKOei44uWCU/b13qVQ6Bi4pCNwGGIgBYv07VZcjQb+vFMlMbibe06Zk5V0EfKI3pcXQi1DX8GQiJwWp42fjgotq0HXGM4Bu9GBeuC1OwR50GENAuuVkmuhhO77wPN5jJ24yKDDOSCKO4BUoU8S1yNteo9KDU+9WukTsfXBEYpAGc88CJVNctdO8EsUIZ/Ci5u0uTotWW4Xh8LWJCRW5tL+uIBUtwq44fEN37ON58VZejJKOkwXKhp6v97dNkem3eSIkxHtJaFzvWHybWeV8BoOv06+U2xIXfRepCJ+oasqCZSuJ7ljONgJdoPvOIxyvTWMIiBpK6VQ+7plKzYKW+/rUeYqWkS3x/IiJQlJ7lM23/a8ImhH40rrP71fHdUmGjNg/R8VArFGthg4/TU/6Ohkqz3okMmO6dFnn11V8O2iqy7qP+QY+3OlLzrZt27cFMiwGBCFz7Byn7ACyhouNNqB6SVh4y8RVImLX7/ky8ZfH1veheDz7ReolxDKOs6KlKec8EF61k9r97Jqy7JqV2dJHUeKhBzzQrvrylFWVR+2thYZup9HrW3zD7niQ7tppz9sJ0ECTeC+v/DNgIgGAPugOaCGcUyZJ9/5rZulrUOcIkX7dbMZzvd4LXF7a7R2WHpi2gzUN52vIm5WJEM7u2RchYdjK3NlrcdAGendvDNXLkhNSM+XV6hx26W8IWhShepC2ugjjoI1qYeW6FqYRgYIWZXT8CTszrFGc6jqur+DLsMfPp0yU5h/OpeCl7ph44gxvLZRpJviYxRMNUeXTgueWtALPLSy6carbGFV8qloVNTNFCRk51IvxUDjQlu9yLmskmsz+YltRuJn1RDARbPOoQWH0MUy6d2lA7bqJKB2SAYwULe0NhglFPE2r/ubcVsqALdAEkzhAGRQs1XX2CBkAv+iPnJEpyxGVKSuFjpT3ACQWQVX7xS47fllnKPB8lo/FrI+b9apiBO8u8taSjjdfsdM3tyCHlwiUyTFwWUJw70TX6Kw5Jhsr4yr7s6jct6kpail+vl82o6vzfSjSVPTSc4JxdzgnRC9L0ZmFIYYTlCIIegcqng7nxTMF3jshTRAKr4Uh8e+seT4IukN5vFypprjKhTelegSHe5x2DCPP7nZVgmLk3/ZWbomX3z9fLDKRQG5XKcbL77HHbQ+emHj0D5j1NWUPHjfSYhooWiJXY1SLBMqQv9G/2LjSZKXE7DkJ09fhgokMmy/LPfxgxTj3Njpi76V9VuxoZdycUBLH5CJxaVEU9aC4ALRbHtmp/qzEEY6lBHODcEM019/tHiY3t8ykfNTRPU37FSU92C/vf3tB+Sq6ynK92xxqz0jP+YebX35cQqUOONnK8udZqoGdJMMhm7NuDiz9sdToA/0CPSRhvydPTa2ACMk9TwWwY7YHFOkMby4U7rY5Cl63diTx33kmewaeM0ECgLtAFQk599jIDWiX9MNf7LJasZ/j5d6oXrzRVGxUSldZklRuZxDJmHUVNPxqq4G5k0yEl1vK1D9VWMIYEzLa1xUxZYGKJBOQZPZuf/VtkI99rteyn1O6QO5uaBW7pJH2SZL5ORsWPK8yzKZp2tY4oeZh5BMyazJp4lQWG9dWr1MlgYqj/msvs2lUiUqEI6LE5u0vhKujgeGdaoSqPP6EAg085k8IbgV8HWRL0qSKTEkWKPuyAsbTWBkrFzdmuHen+ZlFae2ZHgvsgTC/GnZC9to6M3E6WNB8CCbsc4Qfx+IeaMfR5DwIFo5noE97neMcdL9yVMouJlvW60p6eiaBAwzZLOdY7tId2wFVJvFgCLeyBiyo6qqCwvORf9QPRlyP/3waoT9odirkX/70+4aHQiis7Ht7zujdwZxqip8VmrOfKLworotglGLTAgeF2bHzS4jNmMroBNksoUff0RQiM+Wv/IuNLNHCrt2dNl79kzQPWIchRCfEYMM7gu3iefQqWO4PXRgBDiLwntKjBOG+Uq86cL6QFglVgphP6nFNAAgJVFoNJDV023bbaNx2WgHAtqPavUBq3MY6zxmLgQYzrYyrIlOS5DoPLer9iqdGhTmOFjkKDj6mkREI1ArEVvZ/BybKTRnbfL3xEV0Q6DeAbq4Px0RNzs894ILAhWj9GmYJ4/FOv1kcrA4Mwh2cBNq4RQEKMQRd24oFqNHyoRNPBl1pRbWftl6vvy/jsZqla/URWH91o7XxqOjyNFQ+i64ml+z21wrYuxzjTgN6UcTc8PewlMsqXEav5ckaTzxO+prq8hcJVeJPxu2XWcSkPQl5wyov24Cb3cOsqhgT4lNqT+o1NeLwXaZAfhFMoMQMmoKJ1EqYcwa71bp7pyrFpHH3i/kxZd0IpZuJpGWIC8SrpK+0CdM5Jr7vnSISU7kD7gxw+KuECU2xTpeZxUwhPt21HrbsK62h0gUw0jwDuhiaqmIB3vXN6WAMdNOyNqDBFDYFkynH05MtaZmwHBpA3e7f+vfoyp8qpwrUp2DrvXZaGhuD6Dy6m6ew/SjSqgYTi98GXCa8junx6OyxCHFMLVSdLKzTgWPHIIEwR45mUHTrhQQI6llqpoFyPuJ7xHdvnJkzO3ZLjw8ueHMMJxebAiwfIDuLnO7ZajvbTUK313woS34mpYZiuwxLWz5+U5z/wW0mJosP+t8F10Hnz20DpIdQGg4nj0oIfJSP3IfoD+KojCCAhLV1kNgrHdCgonedV6XMnaI7LrQR/6ARgZb8p3e8X+TqkbEq2o+tRx0ruU6LnulZ5PKWsFP6m7s35U8XHCV6g1Gp01aiIGO9wjWwlm5m9OOKSVZWPc2NpZ8jVIT+k8gCWZv3JKaaEJ038XU3G+LclHXtgUPvWUxHTANi3Bf0vzumwD6PXF2YsSJAIYtdIePM3r0umbeRsCzgYKerPHVrwjUfZJQLv0ig2KPIiwEqtmcxq+qdNlsOif5SS6tM7bVRbpxX4VNZiGNwapUUBAsbJUvAGzBLKt7BLODVAyFDrhIkWFBIZ9LOljfvS+lusbchbc650EkNlXDTqg9+sUSEKL5iUFB8yGFTye5bko5cE5yYZp+cYbnBrCWISS6TPG6o0ch0aFq1wwASGf9jH/sAxQJahSgCCaRFQunSxa1zamb2/aKu4J6k+ri6o3ZWHUSQ/F4ajHw9hL0hpYCmM03oINlShSGKzCVTeJRuTYGn+ehGDHzj4rHuZMXRvKeBHjamtx0189A04qKreuCmaqeeCAEXTSf8mjG2VQUCsNIyAExLyqf2aBAuGGYA7ZY39/Y8QCz7p4epgEAxCTqJNAcLyDh3pq17YUlsF1SYRNzrbdyYCRTMPHGVyz3TvMDTLiqin9SspOhtgQmLkRkb+TC4Rb2jpVy7bXQfcEYLQ5oHPQ91hNokOP9+VYaEJN6/gwu7a6AGI2SnZQNySxrkmoFmOzrPp8IHqmMpp+VSmmU+utFvf0cr0SnogmoUSHznRQAbRMPcoTOC591f2LccUQqswjLDzQHXoypSOKOcuTMGvh5lyERgzFbGXZIJIEohLZGUbu/0kPyoD7Rgnij5qCC34YLc4ix+zAfNfGOmfxcBJPN6Aha2HtU0SFMyq+9vBuEnaOSL8sjO2UVjp5xI/9D4/QdnbPBwZbivDcbXk759QWkQc9U36sZVpODVwrWwTjnsIiKGDYAXp0Bn9YTBQprD3HlmJOhKBHva3wHYYSbD718EkGGBXl0wCf0xElr+KildiWe2mYco0LEcV38Olf7RFIe09froYUU5FNRU5EGXM2frw/FK+50tkE911FgRH4kYpLN/4X2wl+LAsm1i1ZdB4EDesuBZTzjFBJSbMN8x/wZZLclF8qwajcrMmytG+3/YcsGiFLP5hYu2xyMj/MIRVBj59WdbTa7QyU4ntofZCAlXPkZDFzB/TtJPA7wUiY9l0aiGbZL7o4098dX+o1t8PRw00OmSP5vnQRkfAwYFLRbrZbiv2l2/x45o5/E0Md7KXoHx4AlKtJHn/8nm63hnunEVT8is69CRvhUazIX2rBpp0eA/xYbSFAZ61kA3rxNSOL/aHKjOrV7YkCKfUlACW3YY7qiphQW4CTc4ZsYy1H39Esi90H0LOrrObe2eAQVS5cStftRAeWIHcKixkDSb8Bn0xVYtlDnnUJRhNCQaMMa/e3lAx8EWDZ3RHuk3VX0hkEcuJVCP2IcBwjrLqrnNjaYL9qcNyQYITtA/jkS5mnFdqwLhwBcwBV0pvzQ1g0KWdswClXJfHzk1U8tGgtplPooD34u/AJSaE491goAImNTPRRhvg+bOpqGt/omcNgRoQFuYX+Pr4oZ2wUU1koQyX1xjMgJPOfSRRZDHvdyll+KAhoE3F/6B8H6y2s3rBwYVjKvkYBH8AXdEb+PYav0++/aouL3fkCfUjaIuQidpF+nVOIWod6B4rYPZRRzxwMEt3hzkxdw9Nc2YTGYDBrtfQx2rEkx16XR450xKxXlBBLV64fyCc+WSXDLS6E5t2d3W8u1jgGM3qu0neO8pbA5kORj4ovDmmEzEyihfBKcUvrcFLvHqG0xchpQ2n92tc4t1GnjuERHnUFPrC7VrA1GKMYw9SdsJt4RsKXcjlQEyibPycwOX93YecFF8LhVn6qpi3fVXBZFJJQ4h3wMCK84Xfu1JFbMHVFxuWhyJ5asOwIHrlTNcCLdWcryn+wsBqbZNXzl9PP5klu2wAp0R8iqWSghAQwoGKRkOv+icqVCjOuo2lNA8BjD7H4SY3r5HB/16WzTjZ1O6PqiEaYuba4yBVeY/ufpWWiZ/0F3SZlYZMnfHWTImsKojSa/FInygq5Vr77M8EFoqTrwNYgMj1H7TcE82v5VpwGRhWzZ/st+OKZ3IsX6svBkV97pdO3lZ8ouOTWtCX7kMEAHdzjRZrRyJjg99uMQ5rJ4B3Sq/o+eAeeMtY83fEd2s1eq9CnZNKkuvzgo3WkKnFXX0+SfC60MXR8mZNSlT3ETADsNnwpN4rhPeRjL7iGAWZeigTV86O+VN2MWHkRwBuRtf08gGVszMsVaLjYSXV6fMem+gA1C8BXsSjmcROX7vOsSfwB/Xe1wIdmxe9ihsY6r3X0POJsAMaAUGPj1seyn/Wk9bgRLij5RTBFRM/2AtoE6ghkJrmBUeG3bPKtDl7JrsClKMk+03+UfNom/gAvLuZWvy1uuPuiX1EDNIj1hpi0GmCbC+xv+bkl7oOtWtpsgkZW24pvJn5wLSn+lJELB8u8iC+iApubDYmgXHxuAyAjT0XzyqkXlc6v8JFwEDlv4bjwNqRfEJa11WoEgNclg/0huVJNxq7x2n9B1KiqhcoznLi4lYFMAT3PDpbN0/OanItZ1NepqPL2QK9mXz+GaJqwGA13T2Y6m8dwQPdFiAb4xnRAokYKjrt5AsYN25UsmWdOqjh4mGupIcPe3JvsMM4xGZI1f+vbW2+vg8rI1nWSCNzpkgJ7AERaVrL0KTVpiqxyymJ9ceYo26MQ9VBwh0wPA51iRQssQGVgbeLvCSmoOscNj++BOY8l86haDF4QZ8SZhO4krMjfH8MjSMVjIFnSyM8mUEasmDk+E/+yuuDqtOLtXIBQ1LPboLMHUMCtJV9rum7mFdOaxm0DGSUJI6X+2lulDF6Xfmg2evGRawAFiZ0I9VK2a07U8eKdsomzxKRhi4MBX61acvjfbbiXDcFi7AgDWnlCnmsE5S90nuTiidQCTKt8ersm7SeoUjfUw6lpDeCLRDaICVxndGxw9LTwyGAU1SKXMIjxBtYKU0iKLpM8cpWWYajr85j87BGutC0iED5SY+XI7cEpFAFji97NBhJnpgl2FVtX7/DZivgaa9wIxzwqKBWSiczP5NEfZaJZ9DIDLVqniqIgfJOCuZwVtmnO7Pkquj8ADFu5BoOKKoAqwGDJGUGrzrFMV/cNxo2arJnvUEsXD77TMRJHi9O5UtsAZVRKHiRQbtF2BADDniuVI7vAYOCYMFkQujsTok7b1P6c9k1nqBbCcLpZf3Y+6B58Wbso0hjAvHWsqcioEMMd7Y/f7Q1phoWq4gO7W74/NfwSwwHoyO3dacWnWiKNe0VtVg+LXWTFS4q0lpTVda3bVtlwxkgtEQQT12Ai7nCwY8hN+Nv1td16yuoj//YeCOycU82Yzu1KpmImKwy/Jf0+Gp3hJYCtz5XpekrvVkqwcKB7boq4Z1zOHnThakih3tO/63vg/GUbP05oX2xVcP1KpR6mXbPw7IvqhHi6fSgKTsEWbEVbF9JBpf5f6zBAS2pOb9uvaJsVxZKx/lFjLE4hhZq/VO+u/pDHKvuAPG/7CqUc0ISulLa/53vk3nLkkS6Aa1v9yHEtkrG96MpbWd9ZFi+REZVgW+FSu9xxAgS9ZnRM9NRJz8pgOKXjxt2XfIqN2lZ7/tBajAXuHdGrZTFH4RZJaKkjTRCokeDAoqjLos/dwJg/hzUnDII0koID5EKvif+VbBD8Hwr2n9c351NJ/mKvGCMTzLAbUtRnGa2dSzMnSowyvmK9gHM06m7d8CYoaaHHq4Vm3cfsVNdFmDveWMvKgEQYGkB1O5TJOf7OsA6XrOg3xpaU+Rn4mZM7PsIV+QayxUFmPl5Uu9aU5xtC7QtDdCz3x662CueGNSfuR4fdB31EdpdbFWeovHJNZrWKIy3iC+tEgQxTlOH8y3w0I3mEcl//GTES41pTOCpTnXbWIPD4zpyiiJlUXbErx0qmZaF0IXjbXgCgMrzXUMkupJyyge9xBOYer0xOFgYxfu8KnivvspkKC67HFPyd6gm2gEv5vS31o2XYKMxuXlk6UHSW3y5DsbDgKP0eWLr5MenmXXG2fFaujvSRHv4X0b36ZIokbsbHBsDuusR4vhZ7AiVyGK68GqwMk50TcD92b8f9oeh17qrH/uMVXDtLAtyQvh9TKsyDZEdS8c6hw3PMPAbSy/8e6ReJOvvXQyKIb2ZvYK8i7bM2nanYKFRamcWY1pBW+bXp1dATjtk8SG2mwktW3chXZccI+JL5ggASbbcs1PVqxJ+O68Z7Q420aDdYbOD3RVUrJE0be1b92o+VYBfJGKZwJVdPHTWc8KEMB2mHQcP+XOfijPcLr9nHzHxXf3uh4Bvl0IxlVXyL4QZ6ZH5nPJcpdWNx4TieeEkzTqIaT9BBmePel4bPiEx1XSSRi7CM4ArPrdf7DlJt0Ch1DyufdJqzihz0VqeuVE6gx6YE1wtI0J5v07Wf3q7eSiA7f2BsekrK1z4dXSF0NPqpYYrnD2Oe3J4cH9wzkqhU1wHRrQCaP4WwUC2f6UkP2ppuTLWFyQmrtllWWqCFL0pDK2eQUp8y7BtJ25y5pISJmP4qZTvMdtjpqiQT3ont1C7L8JGGwq9q7VlHc2JD2ZX6+IhLeFCMpHQ1CelU2KJ2N+SVKuuC3rY/0tSYMSGARhPikmpAL8ykBaHM4Z58oCwapq/PhZgI/gtXcH2Dqu7bhi98ue6es66DC7b92w2doj9a7QrGCjBNPqZ3PRbyyjkNq3xOguJtCDXvA0Rox6Ii7mPqazVthWzUZyWHhBAgf4p7M/dIH5JqB699SrqyiR0ycAxyEM0AOPjVvt1qx6DsZ7Y3aORLQ5ImAbMmJdRDWYI0pr8jSCj9E5PYAshuZC97lSWpxpN0DXHLpwEqXFcd4RVmhgWcd9dUfDMIWY482LLn3xGK6dCEAWjSxUHtNBHjmhBQ3EbGSQzj6fXqqL66mwYDceR5vAbuGgfvOalxwEEoTZVMrMBMz3rJWtT5l0GmDcmxpyFMG7n0LAj1gwbqNQOqxkiU+MEG4b00SkPcbZVQZn36+u8p6kvhzMF9XyALUwe4ST/pdy7HPMkuI8gzs9QvjuE77s1IImjfI8Uei+VYy5gqTWjVXm6C6Kaa+0ndLAYa+myPWOdg/zKKDQWG7SK9lzD4dWrNieUHT7IyhspnWYwf3/fgvgZSRx4sPbFe8B5amGkeYAOjZLC1tBUJMDnmcQBfxfR6H+QtDJQhPaJpEWTGS36SwNmJEjmLvcK/TsT3q1Z2Zko7ig7ADfIRL1sFOS6+6E3K8D4ObwgXE9PA1B3SkAThmG5ln7GpH1CgcPadqZ/ZdYbW6ItjIeZ1g+AYD+0+UjkiVe68L3eqjLbEyFxaJaBeQwQ33bzBAJEBa/5knl44JhyvzgSP9MbuaKUTG6036asiD4TnF2QeosiLw9ek3bwfX1by3pfJZBs5WNSwe/4BmAd71NAcjQIf+eUtVNTPUJ4y816jFbch/hLfWZ31MrLIOilAjPXNXAbtWdrFEbH38KYkR71pbIIbawkTq6UwD7qzpM+J5K4Dtx1Bk1rxfdeUgg/gBNgCTCOqvVDqxvUhAvzvTiEzFXE8+E99HFPym0tTq2+tCCUkYmW28Pt4zXZ+5pwAcCCHSk+9Ik2qo895kSHwx7XReCeQnxR7ElrsQrYbkjFFCQKTVU7oUf7Yfk5Ozsm03kOPcS5K8UwkS0PDg2mYkifsR/Xv3jdEzfF7a2eHaxcpf8y4Z1XB02VQTT7ItgQkuknKLlIAJq2XbSUJ6Wwt+xp55j0j3tJ0g5tEObU4EZ5rxr+44aGDUNRC7WzNm1ZUVJ/6lZADc1ouNz16dq1MxSmJC7Z8ZqeeLBd29dzVnMuao9XT+xwZX3SxWeQqDyct8gmRZPQ0TZBG9pNBOACFF14Lw9e5NJ2XUXcLAvhmoosdXf7VAQFv+grOIhyCHdftrmz1i/UpA3KCK+iUut8C2hegQFO22kMlPPA4GDhlvbJKoXvZo5QJcnt19xcST7EQ/5W1ENkj9Obv7Dl6NYzX7/ml3fdl652VOpmyRvbEh9uxzG9nMjE8spHZEj0XQneZ4DnB3KKrvHn6LCR6OePtlwzDnEXm1FL/KZqy97CcBSpg18eGOuhQf67vdR8bQ7+biuARISGUnRH8JMQi5weuat9Jsq9uPjg+XCbsSDtpTM3wutQrszWTllzgDcyfVqsCN4b0mxhmfFHVuCC0ABx4yHvQ30ApBnewoKYrA3H1u78eyznQnRZJjKarcEymgttmJFTEI42Dk0HeqXXDEpM/p4Nld+IlRJ1bZaSIrNi9FjzhecaYGG4UDmMnb+zwGcvlZRZbam/S7HFhJKk4rwhadX4ocVWrN3Paii+lFref+Yg8/F6n7wFD8LfxtfT7AsFYwbcX5VEe326lalYA+ARmNAzw+cvMrYTYpPvUCJ+9FGIDrTnYw0xYWUx4fxIoIkKUXDZAba/TL1IJkwTjleraUlzcijZCyRuYaYTXJvUABJhDExqXw95q9K1C+mJlHIvXGUzF6oVMRh5ts/toVIVJpMHLNYP4qCiYwArjaCIyXXABT0xnNX0xSiiq05Op9snGlNvmLgxys+RNMddhmnO9njSTAliH2qQVG03iko49LnGxc/rwiXtF0K1vNcHvsOT0JBx/f/0s0zCTAlKLTDqt2sadwAALKIRSBaVJUNnHfGy1dvk7l397OSDKFTNFk7mEFn/qLTXBzkFjh5T9frIuZWbJCStJ5xL7QbsstrTy5RTMQvknhBRHXdMWqstUyaZeqvXy0FwaAWOF7cxZU6C1/zWvoGGZlf23Cn0NPdDupPI85D+d0vkpEb+9b73Ey3c3wZ0eCm5dYFuukp2Kqs7FD20KGV1HhXpPZxJ3MGzCdNHWIafe7LVetcTN15ekGMpPoptuXnsXF76WEzyWkcCmT018iWp0hdhT2JFZwx4EA0kg44RTf7kwJWk0di2IpqMvU0cvBy2mT86kE/9kRbRjZ70uiR6eFMXBvG+yciduayxSsDeoi4K3XWIr5Zo56yudbeXsxFZPcbIr5nZKgc7xevmb313a3fTGF95MmFj9FBZH4VpDORJrMfr/X02aPI9Fx65l6ZXjp9BpeVyFQ8RqoEc1AbHGc4uIBWVfBzmZptPVNCzBi4RgEWORD1dn5slNX6PGr+i98uQTUAWjgw6QmTZ7FtO06IboqAhrjg7hbOYuhWyBjkvudSDlybC0K/yxF+gnNKRYxHWnpRYuJOEx59syjzudn9pXUtxlGq1gTHPTOAO415AE2UBxNPmjXSGPVugvzTrUj+PsUWQRgJTiWdDPyJTCNoGrHgzjGJ6yeYx25HX9k+2zoIl3VG/zY6ScdKNg0qnxK5uYe89fzBii7995bJWdXWgNmw1xBCLcoQ7soaBTiKbJ05j7Sg9s+n72XoTPA/jLVfoJtD/ficjkVmYv+7PhB6eJLeLpP8pJ4Bse9fzX2/jJU+E5X04o7+lzI5W3vBzQ6YR0gS+KIYN8qS7Q9c6liYH5Ul2wTIB3jd9Pg4mcRsnF5kGIWx//urEmUsGviMhALR36nQlqnYyJ2v93wxgTD5e9oQb3f8PAft+8dxgj+9xGwH8+F07dHoJKltYjOfmhMf9bBQHBW360UKqvVX3OGMoTJc3ANS5D6YUVVvU+ZT7hK53mMHSs4454Z/0cHepphk/w1/oRLV6YceIYjlyQmVyHQ2RrG+ANplLfcdtSQSSczHjcp7HJZ76i/SWIkLtc92KWOgGt1jJmeed11xsWZ2WejPikFtzD9iAMzALzChCSPgcZ9Ji5X/DIzKra6+taNuuKRM1A04Z82uyCbXKZ1Z6ulXjVKEQlkcws+7CirxLCYR9kPk/LvAHtHv+t8iKTbkM0PIBhbMzpRllpCBBl2VYhfXTJxrVmwFjVf7vz2g+K/nu99GG27Svv+NpNO48/WNwRy1r4NR4y/c7S17X13M6EEyticX/iwzLuseAvJt/EJG7nko0tlZzaz0HLLYngP5RMwjYbyON5hvVmOHgGYHWXwQ4AacGMNeeQVddOIlBEOw9GPOrBHYohesxZ3/BDTj2jOKAApWhttCW32fvojNf0OupmRY18jQFvzptv9o1+VpO9TizkHkKIl4LJ0iYJqpWvsAe5JvydO548S37hmc7nLMAqjwFjxbi1HDao/04KXEusPopB2dagkMqFG92fEyEpMmGS4m1JI01WAoxis8Zi4+68LiFrza2JBD9kDV7Jwy/Ipwfmv9jELIxE9OuOCtz4ue6AbaIAwAikgxHijN55BzmrY3BtoPl3v0GVvXENFwBC1mFGL0HvN9WqBOq3bMgPT/3Wx5m2ey9FTHtLUSlhn+0qyVXiA4hTKZHJRJ001JqMnfVFXPwMwS/4ga3o7xR411jteAjXDyzXxM68OkxayF8Uh4xWmqEulu+wXXB49ao37SHkantdJFYzVBznOxtwxj77QI8sh1RORvK/bSH0BcpuKrfP6NGbF36HbJEs+39yRw1o+xgXF/9kAeOXqC+fwMHaSJ02aPgeKU7lRi6BkOVVDKHQlK/rGW7v8tqATxJFRg8zDLDgvMhGN9JSBQ6Iqh9kgKUstRx0uwk86FYK8Ujm4iUQ1AvUkXQo+x1IsDh6jiUUeyAp3ZX3KAypUL3485nwFCjocm9TZKranxdI8a+9EV7+6aC9J2/Uap2eoZbSr/NkRr6MX+MzwJ8FSqD/BdyEN8frUk4+h006vyqs06VwzASkmFIIYd4T/8L8xWPkIYiIXrDdh4jkcmu+yMDeIa3GHwoJIKlo4tZW2pIonA4tL7Mhro3uIoTCH3wi7jxJkOH8vjlIQ3OKzdMIA27jYGXv9K12woHYmEo=
`pragma protect end_data_block
`pragma protect digest_block
e04e2ad2a9d0dcb359ba78fd5b025d0a7f5532ceab959ae55b8a3e8e722f5bf4
`pragma protect end_digest_block
`pragma protect end_protected
