`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1359)
`pragma protect data_block
E8XKxHb5OCsyUWDn2GsdN4it4MXqwQJyjcjKakn9U5YOaFD2S0QQ9/o/ITRwgseriaDfhY3xvb/sH6QeHIugCA6Luvl8Dydg+Erpj28/swsvyNcELXHt6ZIADlZNXLoMfnx1Pt5v4qrARpokJ3Lkv8F5y74dLamrfvP2F7RxloSJVNEyWEzIdJgjyYwgmR7RHlrQd0mY/dVQ1js7tZabJ9FCCHAC4Z4BqS5DYXdB7MAwkLMUeWM3f/ty12hTT65jddLu0jEES5JG0ewxcKAdQF28GYQO1guYv2D3qHzIqh57GZY52jegNcfkZXSX44jp9UFVAtHdSp5prIJmT30VecxH1qT5zNE2fmwVEBl2i8CxXyr1LgBbN/WQY2PVX4TEPEaP0G/mUrJHOtMZAs9HyLfqYYTKgVjCE5ivmWcQ54LpwqpFk0pGrZia83zZpd2cBL8ss4gzzQQ5eyWU25XXWGHkUSTFG/AQ0x0fQn5dhM3TWwrOCHjKk3TMzUJaty/o3xpZ8XKlljnG0ZbkU5ft3sGH2CyrxUeMzOdkmceCbg1WSiJklHDUnZ4c1yvt96k83082MYlhb6leofZDdJT+aGRKGPt1RWlbTDuEw/Hk+dmH4vrU6ixiZ1cJ1kXSs0LSHtqgGr1fuX+2ZI9ynK9mkp7T/CvGl+GStFYYZTRpTrvLnU1Jdevy1xQCa6Ti1xGqaHQerlL34WAWjU5rOXY9fkEZNupR4Rax3L+fvH42j1z2zXn6MCCRdINBfWR6nnVwAFi7jGlAgs5MeOu+mA2le2byQNERI3tIFe0evik6yWr1R7Jvzv8qBM/daTdhsvjmIACOIKpL0YwjgInBxcJ3UymAOvlruazYdysad2vplFUYUweLETfgT0fjbp+06uQ23zLN04iGi43BG6vO8jknueJxN6JtMFoCI+9Jothe4TZguRpXFH3+m8mL0TDKdnykhL1fAuKOKI0W6UHw+g5HZ4u+5pyOeAPqHBuHp2Ibuxq3znmBPFB0dQNy0PIDDzzcnWcdhHTAlC5y0zlQZ/w2CPi8Z0fnOjOg03PE0DGOY4FlqC5BMKKWzUjgJglAsQBBwLiLcsFtaOLfwHPKyrotQxIEv1cJ2P9lMt0yCc2fAhCey0rzH3tqnKhMEPr44yY7OKBm0h4BtDodyYkhwRCCvecOgkYifnSaLp5swOu1GFGqzXaVg1K+OJL1CC2NU7ilHGm+1sS9OpZW0pNAdfRRForGUC6hEgeU7piF80tteZk35EtXzS90BddbpyPcPB1npmvLQQDXDcomsOAhttAjCbtc16u3ah8uiQInlC/7c611dKMSEln+pQO1TwlJjuVJp+V8oy/2etshFXTP82mSKjsoslxIoqPFeCOmLpGhjv94QpCtNpZkqXSpIpUkRtYcv5bVMM5MMWYIVdgiL3yzOK6ut2DJpgAaddWBZhlT6Od8mISTUN2KpL8J+oB3vnJSPsg5vvtN8nNcM5jo3AXTUe0DWvf2pCMusCGjtK/V7BDVnkHncYwCiQNISHAlS07lusNoBRlDzt3DL5D4UVcpEpxBaeNp6KiazyHrUlDSKKTzXL5BHJuBXNqQ3z+VX0SqPtpk3cXWaTyG5w4A32MLyCZO3T1SgtIJmZKlbiNW83PcuhHuDsyq27A15Fp8lwOWPXYlrl29mmufNMu5ggNbRZFz7xvbUWNwFC+vorJBO5rnllbkyadQthZ3Dbw5d9l8qjEA+THRvkbKDC5iNiPZBoGfyPr7k07ndm05ce8Cq8hVDletmKEMolRct5NMJlqYYyBtUTAxlOKBjklT00IgNw==
`pragma protect end_data_block
`pragma protect digest_block
94a5dca005b8e1d786757561061ac1de1bc2ba9f18c784d7be2afd44dcde8244
`pragma protect end_digest_block
`pragma protect end_protected
