`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 5041)
`pragma protect data_block
SBR9yGhYo4RzDVY4kFw7FFoLrwl1GrB4FlFV4M/T8Y61GY6TCZT0PUmkse8XZSBtJDXHcczwDLqbu1ZxKV0QkpFrGaTwjDR7b/YGYxRi6rjok1/t8NI/elYkxZIosNmvAGLNuHD1CJTTB/MPpODtEojOZRfT82X+yBIEqA6RxpxHmqevgX/FJtiCl/jXlGaFighDJYCnNVV0RY8gp1EX5icD17PkUNm0q4tCukzHBoH+PryyXzhnfgv7fQyz8cYmJWORGPceChpRUWK4NSEMhpfeeo7IjJTtpXkXxHCIhGWNKP6Znt9CU7x3yDASUwUNFBao+EmimS+/B2ub4HjyyEgNrd5TWELRYBvcER064xfdcGZaECpdvseGd7hhe3nI7j6S3KkZkLG+2jLtGoE7SULkrc+ychjp7NUJ01toGJ4nTiUihsazeyqCTOhXwJNJAIT5UBy2IeaibkX7cf4HgNAUTpalh4LLi1QW++Loh2h6CNLixw4ONeAYk1CEOKMxtAkNGtIhRaRu29M90wk25u8Z8OpzPUPprip49EIIZ63ti7K9lNQX3cOrgJIR+NfDKEAcRgJzzbUAE4/LlkmUJiZRd61vKpXdBJm3/dci+Yhv5uaHWDv0G1sWzaIk+hQ1RndbeP08Gndg2DTE8oAqnYOfHBFZS1ogdU8bbPEAiFG0fGp31re8qNbC0D19jpLs0OArPU7xk2n/s/kWrxKpe9c86vqmb5lJdfW4iFfIP05KlhrXJjjExVHgF9yH9mLispcxDlucO7VLVocDPpM7vFtGoW8yk5IxvH3SQk12G1+zv5NU2dZwMmkghaypm89rIWE0A3ucWoEmU5iVazlx1Oy5NzHELq0w+1xXpSQc2vMXGQFKxwRBxxCxBiz9Sqf08PzBBEwdFdEX8Cy3J5czQvZM4R0EJpLBLiPlnKGnXqEiL24R/z0Ps2fH/w02tNdtvhIMOHHHBuCOKOPHCpGJ/vZurRvwM/Uu10ZcjGLoDLmo6Gk/xL9xoCG6uGQ/JrAAUwKHuwzu/vFsBOfblIo5mN6OD9Ut1GV1xivxAobwANJsw4Wuyx3OGha2sshBzOEKes3CJdPSN0PxmcKqdFobYJFYTfOK/Vh21JjtsDtseWSMVpFhejeup2pS8chSFJSY3YC4cXDREHn4ZCBWfsdNTBUHKIb2eUb5OcwUBWPmHcVbbyOSTi+lFirWb5xHzdLFraOVQIk+UVYDeQJH5WGouSmcFUkNMbpM+GF4wKbB209UF6IEnOOljNrtCDBvH4v2RLWLrmXVR9giBF9e4mHPdzFR0IckX+R5dyYGwZRaIDWflGyKjBjs9v4oiuwPRzkpJZ16119y9PUCEZfiHiCskqs9zWl945ThnV5WW+I8gzeWD5bYPRbXPFzycxohJYftbBmUGj6eDWianWjg90aAgRH2mMK//D4EjmKFYCbwR0dfRo5Eo09y5Gsu3XnLY+iveCjp94CHEBlQN21oLrPWuOTetQzOYwhH125R/r1hWJtVB5p20MfBnq2/kXVKg9qFIA0ohjufBpuDGcBuuBtmnRLtaR3GK3+zEyc9FY/oYxO0qfYRqT8du3AHwyjWKDpqtu5EPx3EbDXneKRbfo/a/QqJkrp5g6x+sw9zvZt6RrlSHtBto+xwwHQYNBNCp5+rps+XZZsx9EedY9ojDlJ8F20nQDeGDPrK19gZ9N3ZdA4V/8fbz7FVgsaLnHYXR0t5xTptuDsKrb26pfQHyFSNbpxVxrIsKgOM0H6ZV0lf3bT84iyNKVXLCrkS7t7LCpuAh4pRYxPoTekmC4vWyAJCTVkszsinvMysr77j7pvcrQ5FNSVOBnut2AKhiOHPKEtuke8NrniEIeKrJUkn/ib4bt+DE3d3zreOaeAxHI+Zm96ehnAYLVsnx6d2t8qzZl/PMZJOdB03m5Xjpr5hndd8deQgSxri6+krPHe92juL8C0tvnGyzGPlPwqL0gK8Di+YUTYxH+zJK2N2qk8pfzVFNNp+6L7z2qHPdagMgCRPAExSlGihx+SInMd1nbYyj5ChAe4jAlWLC3fFlzoqXWMEWzJJqodrFrUib1y4RZb5vW+56ojcQ/YiMWAmNTbSxX5VobQcpXBdPazFz0C+8QugBEmFvIhZgY/TPorvwZeYNx/QSXLTlzBAgKb6v9dPCYMBZ46H+wRjq7i/cMnvbpOt/AbxqgUGUmR7qdwvdvz0z73REU8S0l3GnoxnZgsm0A0BWYb2qVHC+I47mPej4HRs+dUep7uuu3C9JArcPGINluyAWYodHEaf47iIfZbjDN96Wj/Q+8TwQhZs2uFMvt+G9e3Daf7iKIb2yr4Si0OwXqYVstmMskJcHwvf0HtXNiL12QZnQ5oX5Vh3OSHwB3hnBy+UOX6KTc92Er/tzyAHAClbVDHNa+D0rGYPC7uXGBtC9ZEzVudvTWjCvr6AyajEQHpZ4+yebjU1wHlPnsSbTkGFiyOCwdeCzRP+MYcELxvfQiIeGkyJbCbjOJ7G62vy7I8rPbmwG8UZf9n5UGj2WeDiNQri1NlVB5YPBLM5tJaDNjGJ1Olz+bCVDsuiIGESRn00gfS/w4wHRQUYRjwISyfdEGxCeWcIsXvet7ZVne4wD/NBS4xAarMeeXpv6AjcfAIO+zC3LFq35EuKDGcvteeGhrzk+xBvtqG8FE/h2G4M58uY79O7z0SN6AI5a8r/J0O3XKuxTquEypEvpjTqiDJeNRxz1KeI6BlqKseMUqRs08ycRJHCzGDhhb+Gf0ydmyHQs4QDs2/RqjZjMv7yS/rqweYzKSV0UbLZsAdIULQ/cvcgblwONW+e+xkPVCBOwU3QpJdQqpiSlQwVSmhZP4XG+OSrH/SXtoPgXZCJEoDI4ieHu5R5RryU6aBgbpIQAnHF8Ir54eMRSaO15OXCjDMwXrcakOh7Va6H9tMWSDLIujbid34x+Kx0lTu2L0giy/SgqBuVXFifvgpTPYVuuf1xnniuW+aqA0+Ol8+BFT84ZOx9K3pehTuu5t2yrk/SN8p32GCxoR6GaSZz2AsU+qI7HZE2I6lmSRGHgotnM48rHBqcrVC/LYwnfCKmPtFp5/M4zmVnB1ejAtSal9e5nIHbJACAo+LkxRxF6L5hZGgLHKzibBNChjYjA3moDMPua2EB+yNOygVsCL8MJ3MfMspuGO7GVSAX2sWRM2iMejyXBMTqEgvyJ5aahIBScW8K5bbOvoTY+uZBx/WCH/UudW9PQv/xAfbcYuYOUJELnwnORUrzLPqvHq2Ytoehjreqh/j3PEywDSSXi9+nCvQl6iodxh0yIzf8/0HWjBYVgmiGZjBubeqVGETF5OKkJ2mv6AEySKcov7k/KpS0A/2+NEGKlkxrc4+UXLYSCTnDxyHg3WM8i0gzORHP8v3iKJ/KGF9CGUqsfDAjtN5ebiAEG2wXYyZ4Ycxx3y9Sw15YpaPDjKDtILQlfbF526PEUGqyG6+CHKjGyBH+GofdQAq5Avxi7Ju8Bm+7ebSDY7+/IULgKt+H/lyepd6Fqf4dU1jwKlRIsIKV3ZNEjJrx4UC6Pu6xMeeKZMkwBqLtkfsuPiRjuWsF4QRH9AZE82W5Cc3yL99L46siDJu95/xUWAFLcrx9OHP0hlP6OVy74ujeoP7cyVGQqsvo/h6HaRlPMGCtq8USWfYlIJn/7ETPsgni4bvSjql1SJmvglM3LeCLv53CKaSOWtnRz5BtDKZhOQZFZlTtlSSX99T8IxHhbiQ1Y93PE2zTarBQ+qR6z5MOiVx1ORYdhzfF6eS0BEWy7ijenJueNvjCG0EdryTjpX7mc66r09e0269nXnPIL6aFM8j69GYL4Pc9dfxQx+znx9h+VTFOWOrYgYyy/gvZcG3IMEmlEVetlDvQUZCR8plEae7K4edxdl2tmUp3bp6ftOziyKeLOBV0wCGCUYnKJi295UWaL3F9H81jWNQOAUO+pA26F2272StIKf6+nlNA+J9BxNyxPGhNHbO3Bv6DasUfPLjRD121IHk3eLEBi9HR2iguOtRQzqWlgZBSj6YpPnrOMCUH+ni4kUb/1pxbV5I/THJd+IasmkT3ZBuVTkmg/s5yPFvKiEmMUPeHkl4VbQoj7Ziw9sxIBVUtsP7yA/gMpz85OzrqInuqZfqN4h5Z5yfTL6njCyH2AVx+K1htK6ghO/JrlrQCagVHssB/Aeb2mHXXHVMEOSNWOpPpwBUUrg55tKss57/jJvnLjl1V4QUOXFWFqlGG4kKDGp/DXflD99WTMir2pFoZZ73GaP5YzO+H6BDj2DoOZL7BjaO/sumJeuwmpL2M0SqcS789N2CUERWIlmn+6gcfB26ensdWUVBifGIyRD8JTXz8iSU/7tKJG1ezjC11dRmC93YVVAYaL8cx8fFXa9SEq2T5Y9Czp04awRU5jArt3307P0AUOx3Q7Mx2Q75d1msnkxRHvn0bFoMGg33OKnK9tSCjYzwfNe+bGkpkzrggpC1sYhWTb7/JBsnz9Sj2CcTSe4bpFRfwOqp5k38zBH4z6KRwjoJCEA1Iw4eTbesQDTrzIqupolPXe3jmHvkxpD1/CQRc5OIZp+n2H1nCAOAjqCXdcmvLn3PbhULGVDt5ygzC2KdTCzviNxEnU6m3W4wNyXwK+WKCSaDs/v+cRhSPVMdAlL53O+uZ2M/TrZWjcH92zD5IAc6n2SH1lRdpLv2AvVUA182l+2F3Wnw/hSIqbcJGf+xWbVxN5imMWR+di4tcuS1P2ktoCwNO0EDJ6SYVfnGvm7XZJorWyhlKUDOhJ9rFSTPm89cNp7/JiSxHA+Bgxb6hfu3PsJiHAiR8NlDoyF3+bUxfuZqIx4PXsc1yc2WDqHbqzG9KWPkzCJEZYb2hVUrGMlaqEchy+VnVKzSlhaxVpN9IDY0z/Kg0UE61nb3mB8oawRKpRy2wT3On8xu2XlIWR5Bj57vX4btE6l66n3nV4bw9e1/aSfs7nwjm7OOWSAkzrhjW3GopNsfhooO/us3LOW/G211ZCFXkTw8l/1teFvmgj8o4CO2L+htP9qVfoP2WY25Q3YDf+qHUJZ/rQkJNsIsHpe5bqA+r0XRcz3pCTmkiaOqfPETeVt2LuoUS3gV2/asvF2KlgHVxKMIZp5R4XXRp0lraYdSrg0uGWLREZP7+X84MzU+uwJXjcaatKszduklh6AqA17x0mGR8PyOJmKK12+s/07yaoO2p4l5I7wEVrymwVTWCbyu5kEyfhYxX0eMNrCKOBMhNzTlkocnfBQCHxrNfctDyXjYuHOIH0rSs/CQCqJw8aJTwpTKp8w7qiYYMHrS4gq/KG3QxLCMo4yjwZKnnS0N3v3lnvaVF83UM+13KTvEw3e2NGbmFOovtSg+KBwml63b68TybMNj6ehjK0V6rX9hgjgCUj63CfM/yldshMMgoAd5F47uG1yg1tP9C2Vd/xJPFprCbjXLOEn6ll6ZOT0r5G1zXMGlxBTGHzJj6s4JmjQ/rrsp9fSOIx7cGJte9zddP+8W5bynVmsK8+x6ZTK74XrWt8hhvbfLYKWxGyzqc7s3D7GnzRSFM9Sw632/Ianr1R+SICoyI9CG3VYdg9ILhRVywNuM/Vd++xAK7RL7bPiYDMwB/iO2WbU6hu6Pw+1WlBGW3iDmbuoUWxSOSnV+s9NDyoQd2x0ry1S0jdMSzEjWM6Iuna7c2nZMHfpjBcYE/oRHw59if6Clt56Fl7St5At98qJp3spWdUfJk2saSYGznes48yAj0Q4q987pe9xKv8b1dKozGgriDTuSgIOGhfg0azAzIg30j177vZk60nqAlCTDbFKqK4jYXDWbUZ+S2gmwzoTBD1RD00zaqNxaGRhb1pv3XFsZPfOVV4z1tXJgodPkY1Iyd7Ph3MdTLpjByXFzzydt4f8IAsIvvaUwF483u3wt4ArZbLrhJJR4Yx/xO4EgFzue/KDZ0IOLN4w/VnC7+YeQPpGEfk1DuTGGH2HzPumhM8JWFLOnIDs+d4dDUgvxwv78rt6OZQ9mhB3Enn0xcfvJimro/5iprRImEqF8Nzeq1O+fhsZpUnhI7bWpHpdQlENCCpYOeqyh8tzBBgIfTRz1R/27eVpBJDJAX0p04mCZbgf5y+vJq2gFNZLXn4kkvau36uv0tqMWA/8FaMQf41soIE/sULiw5uiXlmFD5hAiDtfUuvjCPjWCUAaHyWk6GG8N6Kprypi3z2J7hQQxTm6w6ZENzAVCvfH7p3K6/GAr5Qo6VaJcpYXRf5MqrPVRs+lLsAuUoEDUrWARljQ61amf4nEmpX2ZtzH0q99bjZnsbaNWTfiCY83ivqmuQzJ1axzyNnh7AY4z7bNkI17ZR+aTEoUJeav2ZTpxiOPIKX9bnOE7FyNM4cLO1sKVM8l8ezR4inLEFh0MgnZPMxChPb8KskWPKNHfzEmbl2fQgHM2D8YEbT+VWLVCeQDBZ7Ontk4DhioZwZJN2U/eX2r1bkA5WhVxAV2R9jnk5nwj/9yeSzwLWyh/1+rv7N/lxf4sAxjgqedzR8qzHIKn1wg0VT7GA8udkP7wQ2PfUf6pd6f/nSbMRnsfnE7XzudK0dejDHFGpmybmb16xTx6jKEFzLv9fZEpdaOijFsQlliRnrQCbevkQ/4wAoMmwNI3nH1OUoe6hTIKcW+nTUXbXm7pW1yg8bC4Kr62ES4snPaSchlH4paC3zJeDhSRwWcpGe9tlGdHhzADi2sBSLsYYx6G1R6rVvZ7Ikg==
`pragma protect end_data_block
`pragma protect digest_block
fcc71dc61b71d4a812bcb698192ff10542a2e430655752fd7f9809c94b0b0845
`pragma protect end_digest_block
`pragma protect end_protected
