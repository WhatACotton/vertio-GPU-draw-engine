`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
vWzmtr/o1yKJPM9d8p/yFVMuz426rlP6bD6AhnRn/xNxX9AOSbWvnXY+FeKYZv0/CfSs9r53z+a4lNNCHQZSDpCI6iJ/zNWuG3abIfB303pRqjjh4xJtVBS24gj5TWDrBZJcG6Tq2BFEKiFUFM+ov/cBJmk8ZTMbzOJwpGB8RcSowobSQbwGUwjTcEDfe6CxPP/CJ6rMPE1EgVUys0XCwrfK8hXXZJCQeoy9R9XlY8IkQTBsectUJI/m/JedhA+eweNDHNAfJ/iml72AQsud/1DVUusISqBiPN2L9u/WhFnfq5AFuHbY4EbRq/hhgxMbNV6ftGADj2JZIj8vFKSpXBuVhJY1SzJaEUWtuNH9cgSDOjyL1sD3aFyZvyDQcf60IRVwislK/h1uljY+efn7JUpoiUjMKgYfhFspsfAZ4/hpWtS7TUlCYT3my5wMXP2467zkms+QxsfwmJyLicxYOrgXE/y6SEfwet0w374m/sF+yp/NfYqaDo2bKuLt+eNPD4umd30Z9kx93mm68HWyPH5EskzZS/K+7cD7kvZ1NoPendMYYV2p+tTtxjFUObnln1ehITadHjDN1st4QCp5ZgBaaUU6mgHEJksvY2hAq96yiIGWAFzHFs7+2+e5VSN5MvjtR29hlvdoGCYGU27Ehjx5Pbq1PwyqaL2Mk1AyybT1QcECpaorAWIuy3J+ygTDDXTMGUAcAqmXRDhfsUtCK/ZP61sDTUxxJDyn6dgRSA2hHDKOTLT9mbaAql0yj1a7agaD51QUGJESzx/miBu+V5ohtIIjxCWk3W1DBkjmfm5iYTXdxdjkhxx43PAk/o64WGIbAjZT9n78fzgxnrpg76RBXHfWUyBZTnfzbPzyDLFOKjKSVsmFFQOZp0zSZ+haostoYaAfySi17ZA3QgI+9NPt3skdJPrgGJV5GSV7nyCb0SvKw5/WU866pRcSrVjPk0dP09MEkFzgM3OFUGo+BtYsbPieyBjB7jDPNfRZawZ1KcPBNDkRKTG6kkUyK3/G/t3rPjLEf3yNraHT6wkL5PAKjhiV27sVrUROY8jx3noRghHQ5+McStoym78+QOC9L15qrj07HcRgTXFrI+fQogXWK6oJaZ+4AgGsLJ6DpzLqs38lgCAjUVZQyiDuGtmXBe1i6zMfHuerLymrbyhg0F8A3rsdwpjSX2kd8bMq8qAJcwzhbyziByTyL7KLgjPp60tsKO3EqIBjkoCTSmtkQQshQ/XOAkMBEN1JmiSaPOY2bWrF8z8y6f2ngDisSpRIIzbmD2OCZ3n/b8tk5lPawGSsyb/JnHj9bMG5moxzVK62Uh7L+5k1TyZ58/+R6IFt7veXc/0Hi9fiomHbdc1npsu0IsWbxOJA4tAsimSe+K66hQ0BttElsZPR6SaxNqBnG65jK+S4TvtqDVa2Nzt9rlw3/JAR23k9zvO1fyWIbZaBAjqDOh0o10FVtr2iuoqj/bu8uqqoa28OyYPxhCMR7VheUGMYL56Dw6JYlxuQVCVc4i5Dznnrs9ZljMjfzNp9EQTXVAF7nMgSubFlh+w2mgaR9VDBRDRKy5Q2lHzNNZ20vhfsPH5SG56Es4+vu5wmgMc7m8DoKxJCL06F2klHNmrVVXNdViy12vm0C8k0mqOcxxKHLFQup0Qg+lsGL9gaYdfsfJTayvSFKkaHBCxX25uH3rzHDV3ZT+qo7OmOKDem4UTZGxY1q+aC8HJ3BcaqQpvugR7JOfSG/LuctcuI3g5OuhorlxmEv75IYiHykLeLF6WGraHRc4+LF+5goeAzxU6rRv9Hq4OfV0Vul5NBPbgp64b+LC2pXi+gA8lLHC2b/snPgoQgQSFxaAsClQyWnpVUZbxZqauYDIY9dpKpF5/dxYnDoo3ffiq203gxEsaLcq5XxZHvf6/1QYe2kleCay4lp8/Kr/Qo/QQLc243PD3gSmRt9uYJDO1RhhEXNWi7kp0+K+PmhpjvYgBnOT77XOWqpe1oHXbJuDA14lDGn+TptCP8opgEPIOzBRfTtJQpKeBPwPkIadpS3M/tpwkG69nobAzp+hGFx5Dw5/TCrP8S+01eiyWo+ZUXFmfV52ss0AJQ8EUmgjePHjmBgVGZ5AA1I+JQte2mzPQ2BDgIhdBlg079TnHvsyq9dOxZBROH7yPClmpaFAHjh2K4hTL0PTPrEPz2dcwrbh0d7SW5HuGWuWOK2lsuCuV4x/GmUQ62F62iWhxNVf+QglPrWAwjE/yE5OKzD1sdbIbKbQsyE4DTO2QIojZ/LWlalg5RecWMZ+fKqnfMcElXouqwrCuiTBFe5z5dQOP+JApCKCwFlN87R4HRAgJT0g45a5L25DCQ0eoie5gQQAHPck6EQ0XQ7Chiva3zbafU172RUMJJJDum7t0ztMsDKX28VP3Jurisc918bhM0+qGVABlLHmTzQrKn1DVIy9LrUBesIVrD4a9D6dIlS1WkItx5n1Hm/9VkMOI1qdJFUqD0tdINXsnHfSUx03EaQXs64KLPRB/gF7UdsDVms7DPCsa+jzTaA4ueyMb9EzqgD9YHIktDOjhey+hc0Z16/C/DRyaljxfLKxQYC/cyROXNcAWsQ4LzNlKyb3WBSTPasdc7NKu02ECinCPuEyo/0raHGxEKQHsC/TooEmJ3QWWmujWZIB56la50eGpV14OvYyWeJuQJCGxHukLzoJyJ3yEazCGvbMJPOSOvRbt25ilYlXpe8gNH0uzfOcif24VyfgJ0WiyGwdnSi8VMsPISltInDr51HxGsFHaxDBpgtFjHzEXRQ14TmyOqfuS1JgrPKyUMVNmX9qwHe6t226PHSFPE7sbjkqxlRBoLTcpokTwrvtF/qTne9k4uxK/53QoVYxC9235RwGp2imMfJRlcTc0uY39C8W2Msp6nGfTDWgMYa4x3OluegaaUp3dv8oEbvXYDOUYJQYEzEvEQGcJH8TOHUmkLYfTKrwLiuc8ndbqsVzxWaTfxBvhqZPTnvhi26CCwNHlLbi+kmRjwRwKcfW9Egh7A5vW8PRHBmT0Etcpr7GorgMRgsfpEQVdoBeK54w3OtTAquVYR+osu1JVDovfkg51BURUhlQKggmDKjRpTleKfd6j4JguMEDdBOjkuQHSZGgJC/Bysp7MpuvfDlUpTK1skwZbefCl0tOp7tczNY2ixZnMrGTvTHyCrhETeo860v3GSySIZd9XiAUyrlqJWvBNTu64nbUtgl21pukTQIT37IOswLySY1M3TJe1sEtaUSYt6T1ikhQq5gHlPTfbDefTkwO/OzFl6qGr9DLoEMnEUsehKQJixupcBtB3Z7szrHkH5WV0ozQ95nidIL37MnTq7mMrHa3velB23njLGSq8HopVKfGRAqRExGtGoxyIJ6sW+8bXp62p/BZNuDMnGTy6TNBSTY2qaH6LNBOV4nHVIB9F5IzJRMrCLJpRFEk/9zpKvod6o9nY/vX9bIYLlOC8OixPxIVeEESanZnp93+bKBGNfZbLw+re0K5a1CTDqz1/F0PYVH4VtSGPkQD5qaYYPLvxK2/Ql0V4CyFZiIlshG5CtX1KoXPTnjCAzakg4tr558RNUho4ELLsPCXhy60XUkI/+LkyoitCYOHvcnP/snDuB/81taU5T+z/1Qmn7T4LdWtfmhfaHXwrhj+ZCBM/1cLpiwxVF5iTHhnMkeaoY8tiuHRtySbc+WVMJHSGsukU1k3wXFPeOrdJzYD1b7zuQhkLGHDPmXw1Aa/64mfinvk7doQGSArGteBbE6XkABlW1z0Nia/sJppbVdkobtFybCEINvlRIOy6m6HR83DL6nmUjEBKvK3SFO8GpyUmSuPwR8nZK1IMfz0HiB8wFM0ypYKtfQt+AXZGVcG40ZckERnEWj7qPapzFNwTg3ATU4hbdFCN05AqWLE88BEAdUdoneEKkRNf0bxMYNa8nnQkSKCgCZlMbb9BCMD45lQz4LBkOxCUomwp0DaetKL1RbjrOI84sJd9z41/jkavGRtEs2k8dZ8WDIyyW3wrIS9pPsACJaVNatv6/2UzzsI4JK11uefh6n+H0QKMUYXZBfFXVRpeJDNjZQ8jWD9PzwIIJuZI3xNRAVrKSCJqJJmi83cColdpEHCnDntk6utUhXm2d5nkBUaVOEGaWciaFo53wwV5gI9UgstAui6Qk824oi6u8zT9w1kSTA2qOaMe8Vu2JARqJYPC51FqFfja5PKlI3r2UQGxglxX2rRXgi12T0XKiE0crDekAXrAFN1lv35owqzwUPwFVjNakRDZySpCa6Eb2Q1IC0GLUvH6/iy9CZg9PPUlO35juzX+6+uFVEc7VVksy3uTVIQUlhf2l9rZi6G4lC6JCwXVu3QEHi8N+HkpTGzlg11obcrimuEApou/g1QdNmXyfW17CEKYRcdvLLa7n/jDJ0GFFYVLQs7BJn1OOtkdr+22sqWkYsLEK5Lcxgpz3HN2/XbMg46O7wXYP9qVICuCJOAjXvGPYDUcvduE0HfeELTDDe4ftGFmG3ZJy49WEvYoDSzZSD0U9D+/IgDS4/dqalJTSaey+L4TCI7pG2zpM/Y51eB4Hagk0irYiLz9b+vqUaK6j4O173F9djIg3ZVQVmKWSS21uDHSJ/sEy6PL1J49Sv2MLi8HjfXGwEBdgq45+iSafHktNco4bejwBYu9+OuRe1LqmCHZz/RcuxNCol1QN9XMq9UnRYgG3gA809DE13nrDI/n4LnAh3RYfhK0zRTzQs+84p4taac7QnGmCmJKGC5OHGwhLq+g38YuV7OLd5JZXRU+wwbQ/YS3wuMpBtZ2WIY1H/52KMtU4rPXbjS4C/Vfw8s8T4qbQPPNj+O8wdIa63uJ4Yp7ioMfcsALfAQoUkGquZflw66G/jfc1RVD+nhR/vXO+H7JvomLSVpM2JZYWu1U5HHrJzcwGCWX+DfZbDilgX86eLT31Z2Dwih1pDJgGJ1qeJ01208RsZV6b8ers9lO3BsXsORldqmg0Bt0LnaAZClbEO+v7LFqct0O0Awaag8IYHX+Pmx06aNJz5kORw1so4UPq4kcTSogR0/ukDhFptufifbZ/7ePm2Oo+AUErUYonPxwG2qQvYxWVkl0bu7x3SaQ6bVArE2MBs2FbVveohn8l96uwyY1ZRQV12F46Aa+lzyiqJS5Y8h3RdPYidNNTuXX+OkuPtumDGCEe3AgYBlGSWuaSHIa0zIf1JWw0KGkPZguOs7y5bspLJzQePGdsUDuAO1QTVEr4XzCJ9OQ8BpiB4xpfj99o2O7AiCIULvfsj6xgaPeatCWUIvLqZ+75tnhXLllfH5XwKywVTRwZYVKxh6bJB/BltcFXXxWR9pT7yrwZK0tuGq3xRQDq+r6auWozOd/85xusI2GGdbRQ6iPqT6Eav00Jl3/sET88gbKfQ+HCHDBFesfHnmDfAAiMLMCjLXNu8vOMhVxj/wv5mD8qHA7Y2Emam+Lmx1Vp7gchNIzGALQ1HfJPwj1gZOvin1xACx1/ieyB6ASfLZglEUtSuk4bwjLXe5U00MiM5Usr7LSERt6l7GdSsljZpJO67QDOCO0NZhZrqnC9tzz+dLnFMU3KjTXziINyWB5LrWejcIGKSArzX6c/nA4Js5qeC4yBUNwca2cWyzRpGrtTmh8Z4Tz8b1NR90/zWoyC80bHb7mJEb3GVJfHpfoizip68LMARkFO6CskZTCvXDlpssMzs6A9LVHe60ked17xWkpQCSShAAH4+XotNkNUUzNVCnec2FJOvdNqW8wi3rtAzWXp0sdzg9OO49bfGEIukG1uAj8b417NieHaasoO9H3EtDMRXqqEUgVtVXl/tQi/OFkokYDB8Msj3LrI2kUtClcQ769CdRMaXhkWhb2PnR4pLEkkrRyR8YyC1RjF/JQJEXMQ4brOVaBFxwg9m4kvanM76r4oXtmiW6eHJ303xQxQcftylynmlyHqZQT8TiUq1L0FLp4tx45gTjpfVlXsdLUe8FwaGnBgcoGFu0HqTSvsmkKL/zZa0WusCI/DmgsMTvO5m7mrcl9gQXeASdbCnaO4x0FH+OX8mkemHl8al7890yH+J2qbrXT6iBQsQ+KRnP6z6ozUsLUM2W6BnyCEz8iDOXvJVLZWdhn/DQ/6rteHwGywn8dAkZ1eDT5RofBsi7I39yv91urGZhPJMkYA+kPYNeH5QEGYyBsjZEiHiAllVTPoiZvwjc4rHLRNhnG8cA01+eQcIkKM8JKdcQYznlcEfehsS7udzv/7GgRShxe0bgrd/C2wS0APPmjujI2KQQEFisOmnALR7OE2hyNg8EqFyuhWKgzhZ0SJsNV47c/al4zLDXeH2uCwv9b5sVaxW0RN39PxjLc5jVvidli6uZkfU9u24640bfFoy5fFONA7KqrgeT6IcMRka/RFhC6z0Fsl0WiGKLfo89t68Lc3gj0AJBJoDMlY5SqmODnmlw5DQOmGCrkYLm6ASeYskS5CgPMy4DnVz9esmi0eXUjcVgqEk5G9EnuJiEk6kfQJLu8F7lj225ty3E5ilyO66AGbkP89gmg19v1Xh4VXKpJ85szrdN+WUgVCuW3PgIVJbrQUNbJHQccE3PQa+j5Jex7B/xgPv/iG4guiJiNhz6G3usRs6LglG/vKThqfDca5zRCtuWyGkLkYsT9j6ouXbZqYVipCG77BhW36SF/Qq2/mG2AQ4hD1yL+nMeSBQiS3DmNZbEP0bkDk20ZoZ+b/Xvm8h3IciSNFfA60EgLuNcgGXlIKiOF55LaJDr2C9HCEnmWqe4aJRXYBtBU2fcCdOiLUSLAPy2QMpT1rRvOD5KtbWVRncE+WsBGsN/Pv4QWI93KWSrvSQMoc8sJdhis79oEiPT+YYplH0no7UCsl10WZ5J5aSrLOqx01T8MMR4P7WcLxc+FVjiz97f5wbMdOlMrGJ2ru6j4oR5Br5n20IyljD+oNQTvglBNFY+atg4j4N4HSEdPqFPlvmtOgJUPoExzdFIfkpCEv69Gig/DexKn6wFQWgmrxqzP4uyEH6oXPnLvxujuOg/Fa4Ti6g3zqzNwUolfi01VvOFBOGFLVzFkw+jYgPuMevCZjBhX7BUpWfgWB0UCaM4/ZnlOyNZTfUEbBqFmsAZLaZFOcHJh2rlp5uV46dNB+fhxGF+FD1Ut11ISXosvMbejMGtyHDHS3ITXNtaJ7uxxAUn5PsIuumfXY423kndvY1QLGeutkFGx7YzTS/Erykas0NbCSiqmtq+93urzoVr/ZO/UgI+ExGNhvsfRAYY20HuGruqCy/yC3eV7qwCHtgvWUMhqoAwqw8stf+r73iDorDKuttABNqNi+5pXsR3E4jVqM5k8D6mue4JGQwLPSUZtAiKoocAYypi1I3PFlskHhEySgNXnkjyqYuKi2G8Nb+m3FN92EyQNaH9kgbhGb8Mkm7E2xKlrJZUNLWkKm1+VW1i7hsgmQaKlkqPdY5U0a1LwSecvZFxOFDJdAvLglHqHSw5wip97zDJcXmkGNd6QH9ergEbkhxRtTJn10Ja3aQnX7BkyJuqPMc/2HVNnh01I6iqN4GFJaXjjJUgA6My80G6DCsNmhV3TIERYx6d+IpK5Zb9h1qXxgzM8cjtiGq6Pf63Bv93BfCDTBSY4Hc3P/unuLbzSWD/pohuC5gjNkWKi6K/1ECjzL95v78iWEvvRS043XbzUijzkVZD6uxAm33+4cR4HDLd6oT27bC0b3hfhI1DMcgNpWdrtsB+nyVaqHW6174vtzrUyT0mJZlrdd8ru5AYcTvC4QT99xabY8rLexEHT+arY7cdMIV4iJa1n2VbdI/wYW2id3EZ54hu8z2DxkyMNzRHWinu+VQ4tL/djB1QloCckE9WxMk+BMrr3VzIrg64xuKO8oxxd2MF+iD4wpExOYQelbYOPwBNYiOYHrUK99omNcCZBBAbLbNpTHi6wdM7UlP+ash1rxeepuA+BsIZa4uCYUABRfqNowZpuEvnGtPUIBC2j8rR7HC1z+mByDfwfKy3Ir+DfYpi+d1apnKLETqjunudUJkjeUT32y5Q4xsW/Yn8QDrua4KZKhgB36fiGkxZjUDeQh9f6DEhhpWWnvTfpxUqKEKxnsOfeujdT35I2rDpdBFDoWAHVDSJ0yFpiyDqoCFnv9FmPw68egz9U7vBBIYu4KwFieGjDfF2/cN9tL9EeVaK35ylsbVIpqxshMFO1ZQYFNGOSuKXeqsxMaX4kx/S/zmaqIn8M9cL79KHgLeotSZzJwYIk5wva+V8lfqHrz7qHVA2mStGNoLsYLyfI1vdzRWrZTrifbE3Hj01c9D8uIT9D2ANsTwKUF4v8n6gGVqAINe4HAdJAhnNZKrSFpUVdJfY0p+nEziGLhGNYGLl/YPAxyPmQYj9VifbqLL6R8UxCLiyMDICmVwe09hRCD3yqWmsIgWiCjT/I3znjekdtJuYWNg5yiYSjHjmmkQmPzQO9ZSJYJT6vLMlZIfVn9j6x1ptLV6ptBajqOjvD90SNM/J1DvjKhPKuQxH8wGG/5SWPqfU7gPlCUKOmMpJzLp+qXnfxBsjS1UO5ZolVlgHr4AMGuAVLjGr7dXK9Dv3VgtpTGVP4HxOkSkkGnTpltCE5Hyo+KgIQEuHnse2g6zN2Oo7TYeZa7Kaor4AiEwgWsfRYUMrnFreXxnczFoQIKaR0z6Syek4hZP0uT7usu3mfoXX4Gh5iW8lcQ8QrYEzJErKHMpdVRhwkG5qN6lx2YJoeB+1tPn5lCGRvQZCjt0o7QHrfNaYRQTk4qAM2hUOmEMC+hryAd4kd2Gk0tls39q8C79S9glxBuTMmoUgFeY90BMqeWEdwd3Xjip5FY6racHyvjboGrdzJafBWVLChJTfUPcnkG/jXwNLNrrMT7RFjIoRMBoU0PElVk9CQimjXat/MWY5C0jIOYjYw0nUjbOfrpkvicuRiSvqALf4G2ejxu7mjnMvgQka5TpRrxhjNefVPAM3WRDqyQOw/1TK6BO1G53fqUaUOuP/b/DkexbFMxmNajBmLA/2Yj1MtoLEdoLFAWBNYdTUzYVq41tvbnQIdXk4NavuhJ1T/k3tI/yaeHxYyo7SV9BeygA50Ppmqt4gY8Iriuthcvu8fphviRw2Kj4KLloQbHW73E4MWvHCiDr+m3aREH5VwZTCJe8ZgnQKaPZeMR8/eDvyJBuM1d8bfJI/KQnQrGNhbiFCW9eA9r6AGTtCQ2J1z/rTQcTkq9ULJPv3jj0IgdBZC2c47UXDXzzZ3Qpf8WZwuQqUwFGcS15F3m7EU1DdnMCrE6fKQV9tQsa5ib+LTmlMqp+tmBtN50mlBIV9sGuBJiQRa63U8lmdI5TKvmMzVngGsfvhwpeD+pFjK+Pmc8Oc3CN0xoXscO04Q61ffFAXWwGn1sOl1r8cxwelnpkrCjobWcEhSz4qhQ09U4w86sI/OVw7xaeMZ7cm1ez+dnl2CcAprRfBQDV5av2r4T60LJZzHB+XG3tp53FIyw0ppcjj9jYnBJH51MZf41a+1r4IQRfx5yXoo6EUhLd+1pOWrKJPYiXNopoBqxeB3VFBvHVgvbBsfcgwAYGSDTUbxbS1ZZwz+Kc1ZJ3xlW0LZcmmQ0ndGG2iuzESCQs+T5bSkMHroNhYhhFExyDL1caj0ThvhCGiLh6Paea2a1El/KJ/P8qdRFwmkX+5JG5PauLKBLoJsbfOtYDneWR7cTH23hJ5oU2ZjG1pMTQMyPs0mdKAOJpfVzN+2W0gnP6Krhcb1njaMJ9X+FyooPYw2D4NBMHASgbl1FWfUhE9lXFeMB967C5lzxifIrJQmdS3L2tWAYWXU3IxNy84nKaoW/UXN4HyAzsQ2uhkR8M/oA1NpZm6lhPA60g+0FDkJxxVLgss23+3UbrcABOfoq52XHslnkFWgf5tg2Y1XHO4omr5ksaoZlkvJTylrNKL49pVuL2IeCRnAfAs7mrf4+Y7uGugT4Wu9AdfCJsQubp7kEWXhdk4DpWW5AqX0a/zhUtpunDnoBQqPjwEeVn4IynTWcY2++QdKy6Q3i85lGbSg1uZHE9dZ3r6MiNvYbmvEGgQPfx199iOmHZxYsyjcfSCFB7TAFL9SCyaPAOAoZpOWxxJuU9oMoPr9EBQMX5fxYfl7gFdz4Hw2sSU2aa/fNgwltHFHUnLsU7Bja6B2yzMryZNXdCiDgQx17IhttCHihxBXOF/4BqtlxMEt+vmRiKMIDjNIK4J5NB1JIKGFn2VdLX7XFiGVoA9wkQGx3ubsKPcjyrUwScDFBGdd3dRSXRec3Do6Tu24ETj8r613MrofnTrzyETfSWKWY1PxsKtQfZsNE4tCGkeQjYGJWMtwYQ4cqEVWROLZGR12Wn+NCQ92FbFej9P22ZYZFngRTabriPbE+WBvYQS2wVfFSmYgZBNptMYadEzeCvGhu4ImkpJkimkrhHr+2Y1cfpGnHIXb2XVT5T6/GhaNqYqGYFbEwktgh6dJYl/XCppOUfaIMQ8OFnQcYwwbG01QY47NdmsUwKjfWXCnX+pre91ZojoqSL8J5nth1unJ2oZYGnCTjbiALVeB1U1gF5EMjsS4mpwIiABurx9qqHXe4DiE2FzGHvvCTXYd4pNcpWB3xo/vhiBs0tpl+RCfjhkojFsu9i3itfsvb9qmAQ5EK/yLQutc/sr8tDb8mr2/rppnXkb9Gr+6Zzg0rR/TaDbaT+y2X13ypwWR6kjc2+k7Zp/DucYZI2OaM08LpZYYv+tNAC7PI580Iqu5wio9ejGNSu5xH+73xxpiAHJhyY1SzLXugQ+Mv2kic42WUdWihwXNiVymCB3kgYQr13Xzrj1ids+8jJ1kCnY+hRzbnTuWoPmeopTjX+nZdzW5Y2C9ttuSWRFsowoeXRL3CC/lPTqdrwpOlnqedBwSh3gsBj4K+mOtUuQ9U70NRgjAz5twfnAKg97HBKOLhVDNvQSyZn4DrHuLE7abYY5Q0Eebwqg4ALY4Lh6KGA1HgFgOwKUfv8VocjKkIN7L9NYAs4KMtWLh7Tpv9z22qgaJX8TYQ/n6B+qBwHWFLWzRjLOYI90rnanapoCIj7neVSY5R+Alvyudhvh13AHz9xwWx4BPwscAVFXt6kuc47s9Ex+QhKRSPTo+iXrhYrvVK6yvkvy8ALW9GB/tGhKCjciAPfS1NvvYQ434jDBMPIERoU4C33CbJbUxXQmpeG0+kh+SWLvWX3ksP4fvqnml63JsKCp9D3LibAQIttpxgc0l0MKX2OGwMKANPVJC3cGq2GfTX1ETEXqUlO8DhdvrX1GIZV0iLjU8vxPrgMKFA4ePoV/PJhfTc0nZ3BhC8vFcVmH9DeABueTkd8MUlZTKTDoisMmAgMmMePFPBCq04IAiOwAdoOzmO+0YxTScmAQK4HN2PD8zpwvFoHKB66HDTePBIh1Dz9ClG/ADrz/rD7oXfmR0WzULF+Sz/wRmxsbWsE/WPcR3NRFzGhwEvWx8/tj6qB6kUku6O0WdFRvwLMjw56LAr0wQbcAYdxyyvZtZiVKz2kNrfkaJK/+zFq3quqOwURjVAzxLWJhoMwOXJDEWsxOoYUkeK8ycNGFBcscEvbhhnsGp+a5D+1TlTTtLFVA1XqKBR6+IPLglpAkQtIBr0WEoil6UZq263K0islO3TvQ3cWnLLg7CQ0hbd/5l85nfq9Os/qNGBsDn7ZM+pVCxffF+4aXwFCQekmMMe+Q4TdPuM+bOZmPrAvUUmVSuiTms/IZvNJZ0hjeUBzqOz1XHLCG0bHCtQPTigMhuvTOULshCTRvpuEk0fcpLVT9v/nFO3pP1mAnXaZZ1idLSqXZjMLl0JmQ2y/U28H6QCCtcdvOOAgosmBrEvaRpcgYZdgIzfTQPJQsikFcMQOMoQTFcdT8CNrBCid9dvD3bexM3yYSk+R28SGhFI/6kgUbPHyX/InzYTrfx3VKAnkzJ2MK6+kOvMbzUbEKjrA8OOvKrxIpd0UpVsA26URIkvkE2LJxKizQzzulq8otq9kXujFWDd+6gsXl6fnN3bGpIIo4002mBnOqnFBfqcE5wYCtWazo4bLm6Odxwd1g0GLXdDhdW9ozb8GSeLTO1FhIjMZQNOPHtAYjfMkTn/PsNEHm/zG19MFA/7fbGR0uOK8GynevG01EdIMrRvDJrvTiVGa7PyKsYrbNmPuMyFoowZZNqQQCK1z6PEjIZk2D2IBGqRw4kt2Ar2KlgetKGyC5aLD0VNx2NtFxklfm9aVoHJyCBvip2QZRWZ/rptT+4kJ/4ahVLw0bBmrT9ubN5eD/TVAeMLU9moLoXoqteVhBPSrxbq95Dbcf7TB/0b9XFAsn8cwhfZBfnP9b+Cpsf1n/rzcPW1SfVCMrVDP0TLdAOUtczUOKT5mBKTLNnDOZQfUlAvctJgKgaNZOLl8S827ZgzvmR9cjhJXPpPpXuBEdzInb9qfQIHcwU77+0KpB6IQMtdQdpW3beLSlJV9C52KWQJqX1FMlA4sYhL3plqOYJppk9UhN8j6wXLDZqrHwctnvxxjVwty9eBNUOoyScXpkXh4jLJvobRJ9UYzPQ9tspFrf87OT1+AJu95+YMIMnhkKnYUYD8oJzqIcDfXKUoqkc3G0kqymZ+C2Sl9VFHetPuu+RLgJviWnd9WsmNGyl59IfE286cgpIdvlD/AvE9W85mBnjCBmQx4GUY2upoPngWLIRU0K0glsieWF6sFOQg26yK90mrD6yrnZJ5EwVKrr5qVATO0p8lvYh/Ly9obKw+LGtMopBupKfOwkSsfn3TJtGxORPSjpE3vGFhh7zqAHOGHIh3OdEp0sHFkZR0s19i/Nw5Ebgdw3zLDCWP9uuTJf3vRtfoC0EEtNh7oTRtmM0AkB/h/b1/kEs6wsniLPjkvgOXrumcTUV9OUxittsxFGl5MGPtkkkw5R3N511sVe13ybKbvPtFXKKvQUFpl6mQQpZCFR94E2DU6/pqvXbgL+jZCsN+F1srs5+OzVVALb3xq4YgsAkbd35O00CLSvvGssY5/b3lvm3N5R8qN1wJAAegHDLip5bQXUTxy+cFhx2FkyJ+JyWXWbRWURfz/GnkSB/dCFoyFBSl1tSZvx3HyXAARN6Umh2Co1vPuR3K88coWs5Iky5g6LoI2Z5L+7wtOM8ksM2o+a8HhPZJ6olKctpv8FUEDJH0tG4OU8iT3qaiSsMPQsIBQn1I5Z6qLoxSZQeBfSstXSQxJ+/Di89BCBVJcM4JQ9if84qfSAvmNcyr0VQF5zm/b5XgOehLdV/C6YIbB4y1veVGESHoBFgt9TaZkmczJ6u4a1tGxSP9cvHBXdUqoltjvbZ6FExUOVLv9sBykdXSIEIpjFM1L71M6F1NrSHJKGAmFJZNKShHMaN75TI823d07c3jTcfo64RubTatLtObdqjz5ORe+JeV0L5xjyZy9qU+26zgqx00/HFNfz/5Lof2P1Xc5llgy8cTNIFRC0jv3+YFHf3dY8kdnZynh6SN5SUVbWgd5KTq/QMExz3wh8OSbebSkdKV90kcG/wKOFbaIYhgqBtE/ipou3L93dW6bLi9lQuVc7LadmshPnLnMuGZuaGOj3VdP42powTf3eWKy7JJhB4oyyDUH9vLxPWJQ6x1nugftOlB5tIMlVoXIg1o0P4sFlzllu4Asyj7CQjQN8uwzKBNzQEP+L/b/bgy9CSVHqHsspRE01Q5bJk6b11uo9je+xpuxzUko54P+9LgsM4XcJwyAyo/oea0SAd1+bS4vymt6xFEBi+BrA3CK1hjcHLB8EqWU7pU+vBMkq1w956yu8pdz+1YQDd1OEo0jLin9KcQNrbmTov3SAiA752xUYVV2dj3VI7AYeq8QRHdTT9D7WfCoGrv7vj9SsQGiub67nnaGYI/Dycc5fulIiwQfkOI6z04+muJMzp66guSvKNYJ4jy3ptgSmniBZjQ6YosHDvDqXsLeSvwt6V/bSsCaCBw2X9R8xyKrlovqCyUn6SrVNa/qEZq+7C9IjGrJ5OeU7r+29q1jft/CEmtIawqM+17Fm4NRLkQ8UcPYoBXiK7ziorlXoYhRXg6IgZoJx87XbiUgYFSK/3MxS1UBzgGvmirVfLwkDkOoFawvRip4rr2sj/gr33zcAABVwnoOgQN9KpV6RdmYRnVGxxfHjCGNO3VQOWxBpe7D4hBLXJSljg//NZ9HahsEc6t6b0czvdw+xTJ9dIhYQjVBeOEkfwDpj+3wVyLaWNpcOhrgn1PaXm+L3++2/2raSysJdEWoWcRCWDZ3as2M745NYySgtdl7UHLqF+kABGsW22/YCeXhd1nJvOIQGn6tlCXOz3Oysmj9oJxCFM/AVdZVgFAagRCC2/W+MPbBRgDpgVDstow4fV95I9DXktTPnCNKfnIEoipYNgy8QS5is8gxRc3Koj0IKGvgc98JTaT0sPNSqWDLY5JbBIVeIuBf7RT/aeuGoBz0rjU+1dFtJ12M60hmWKtGAntPERFCFhs9A0vZ90a43PwOOOTrv8zjWBaIpJEuBMyu+DFPDYW/RUC2YTz1XxYPb3+imzIX4fUm2BEFh+xQSC17kkqFqzmxxwWJ+qIz1EWfR9rLPICt9h5StT4QHACuOB4PA9OoKnzAA6ejxlDQ9epXHFJRF93AzBF2qMezX94CQvrrNJiZptFuuILhaLMEgBzcHBkLuyOaDoiB2JAG60zskf6bM2/FZK+1fvZeh/RkeopDT/EXs8qRPsBaEFdO3ygOLBfLhZB5KSS01kbz4fTzbCrUOPXAD4e3sEm8PNFBlIWi+OEOrrdU3n/GcEjG5Sk6mTY5Ar1k0hIAZzXFiJRhiDwIANEHfy3lLZCRVt9QjCzK7hZQpFwj7+mXFXUs2gOSqCwrSLxbGLDwFNsMEOdfhyGjXcwA/WbaW8ZV62HPVDetXcSdjtBsTc4Z0sdlFc2aBN7XSjZ6oTGACE5wCSmmJdpTDN9+a54ogjnCwpbrXQB6P2vpjLokhec4PbREQLLgAM6Kepp+7lJezIEb6iaR4k82ZWmecAhoxgu4gMoxT+EIF4Syv4CrqL3BC2PnAVq5aDBA4vCFm357XP9llZO9h8O0sqc1DPf0hScFtQeGpqYO6YC5WpeBmvIZD8mMZ8OjPZiviFKfVojQAjD13pYZ5284Nyvlr+DFfBcrFm/LzrZqFLuc4Nc09OKKe0FJa9t1UPOt729IcVWvXUl2lEI1KdlJpdSeDKCBhMU8cAOcceJYA2DYjvg0UYkEfrHUSLMyqcOzGX5Bt7BMt2RS/2FwE8Z1NhjVnBWcwhGXnlfUKYsspoxEa1PvrF3KNLtzcRoMr0Xt+na7fJfFLy4BVuHLibbwn6mFFCgwkCqBvSHrlWxp8jawfyWQhZsXehgGr9QX5YD4/lwljCUZT097qqCBsFcG4Nys38rKa2/57eQez2KxS66vjo0CRc/9kpysHYOVE1NK3Yf3T2heP/ijs4RzgkeD0XuxgVuMsOtsn/8eEkSxMN0in/Wbk0TwRmNG5NlzWo3Zo8TrRkhwBRDvzBlwT2Heelr5i2rqld8mCaL9oUX3oS1+PckdRO+h330U+Bp6pSkYj5vkziFTsQgW3n8G/OvuqaKmyBQuSbttMX4Z1/AIJGKysfg+xGg+iT9puNu8IZVZlDSUK8KlPbj7iz2cjEgcLnXcFXND39lIDoBtKMB2bEtNo0Eq2RZ7Sw/37gXNBEK3MvyMSLQmN4/RlIRgQeg3lkqZ44MEtDp8fAFKKwPOWYRvBEW3fZLqv1vl/2nRSqP0NVSmUEyCWiKZlSSpbvMmkvOcMkfZgAXNuAK6jdDY5FKzPDcZ3pOk5Gjov4GH0lHxjazBZoGFOyWFB+fKBySSkd/QED3PP2uMI8UCQF6ovS1vWUAVI6rTIwa9Fyfn68nIs2SPQSGP8jeebiO/2o/enSKa/3H4A9AvWX+joa9JJo0bkepTBU2/BPDtjdWWF69kZWwK6rfC+w60Z9WS8aK1ZzPfyGsX6WYCL+7tXNsnwsFk9Kh5geQGUEDr3JK44W4V1SYq6RrbH940AnzOqolq+EY+JiBXpN9NkJvH3v9ML8kwFKIivE4NcEuSobjGGlX8NTF51h6HWnGwBzAci1BuKbdexX/arHgF6x9tua1TOxf8g28/j4Uwpmb2ck3o82QVZIT1STVXmqe47VUUOc1AFGY+9l6/3xE/dj9Flrfgr37QTdqCmFZzN3KrtMCy5YZHhyuFhF2pXOPylD6Aw913J9BMbdE3ZyKGhxUEEjk4mSz3JzQZQ4pvrLuR/k/i4ayAuHeqXz4d0LU2thX/RUQ1LQyzZHTbbiDtJeflGTrP6Kh5rbbt6D+r8o5RJRa8Uk9m29EP0XTwSQtGtdSt0QLgfnHkJYxWLYunz5rUVVe41AiPs59B2BRg4WBMuwxk7HlRDTq4RuyJugKjffkLawb+Nb7hwaU78aaEHlSCzxj3k7Ki0wvxQ65hGKbCuonwxwdZoRvGBp4Dr06jts0CdXRitgCs/ZJpW2bnycuPkKKiO+V/UnfJ2h128Cwx+NKAhQc2aX9Grj26Jkvr94cIi1+hRhmme3Qs87wXzyrakwgJMKLXrkbxGFtsvkD9DzuQsRGs0OCFqbmc94pxLt3xEhO0WnkZwngX6PLiZIVmkXNyj2A34pc9oCsE5hINd386qQFKtd0cHKrFFHYTKdM4M6xsCXK4wJfJD36xMkOz3U4qRlQEVIAN5JqZzP/+AHHd/vwsrEfAy+h6mZxWUq7owQSp7VKQVKelG/rTvIlZ4fcjrkOZE+N0ncID1kTVlhtFAvMAk7e+yWZxLa/Nfa1P/0b8Rwx1qL4Nc3fRJ59QW5E3qJ5TjF8xZLe18A1ylXd3604CYcAnfcjL8IOLPk5Mae7JPEo0mdfSlKWDliIkAmoSxp/ZqvEb7WqMo/mf5rvK9/DLrn9OsclxuB5mTyaldBlj4L5mX5g7OMZAmZuosa/RmTsMe3icukAsmXNyPfHq+734zjjpx8KApaN9thGJ47kg4qM7NkNZu80yv4KTBAq/yz8XNsmmASNaAcRYPle0QR7i2XvOD2P2XIXHfbeRlKOEVFn2nAhZR97vcepsYUPkJai6XFrn+7Q/kBRkc1N2I1ZYG8fs997yrJ+e+j5RRtK/UrW3BiaXsytrkBiqe0L/aGwoIbdZVqUFu94ON6A5p5OVtOWdj7Pm2JI7Cr2RobKHaafNx1fynFne4IEsnpAISW4DucrYFCthUi7LMZY2pf0elrexzq55Tk+EWhtJG89p/tHSzVKnnxy2IQdBEsGz1CF3kVIRMm0LSvdEIXidt7moKIEAa4T2cEuBgX1yteA2ISrvG3psWUVMLwd/TzxSoWHaaVyqVMsYePCbhCTPUTzsYgYz+pCDvAIOI6wk+Giox2FRiyer9degXQ7T7CDzZ5Lk8kWiH+qzyi2idOfjYrtp0Yim7eOQdiJ+LkQkexRLuzdZ4UP9LFn9y5izM82uhI3l9g2q3S+JRKNdEfQRbfyuxdcSghvYRhaGmosDZkvUum1naI9D7QXMNntGYmMVZ9f2jJMSn1l7aLUr2xgZZcCBYWSA8IXCc3gAAg7beBwGYqfwdTWIyvdoPD8WjYH9BSSwPtgStSpomCb4c6AHS/hWdooUCuLod7NHu6IdDspnm/PzrwZc8nRlL311fX1I+8T+PBEbRDW/vN6UxDYPl0yubVR37o+Je75/Q0yAKFWNbum6FRkhem30Hh7kTvoDLcCMxGIIyYG8osXSTKsTNRO7dgyzgVhFm35Qp55QsbENtwapvpI11s3OUcTs+VDdibTq7Y7o1RR9bFhv72vuwwLG9ffOIQGh19Gs/BnbG3zPKApgiJTWW5UIYd2XopGKx/RkG9Mp1FIZiP2EJLXF3sxCr1KtXbpgk3Gr7n/8/Hksq7es8tiItXgX/muv2JU4zJIWf8HNW/gGwIMT4q/LiO1+L5ongx0aCaStYrLZDqNWEGcWycU8QCJQcjNFqF/+gixJvPUXIc3CFVgo4RQsC1TNMWqNyC3BeDm500DR/bW6zJNY0WdquVAsyPlyGL4tnUjf5Tp5UagwoJsYiZO3zmh6wSevnjfluPGy64lKT5RYZ+mD6JgixjZoolOUH3J1LOZH6YzhUggPjU18scnBUk0MqAp96kpuGFoY3d84veCQFQcyybpWDO0bwIRoYVMNUxSMXJ58yY23AHLbBeUN3lz8GMDGDB3dla9+xIIrUEr8mpYcB/uizZTKrSbFCjmqo5+MxocLHC3VAHRqInD+Az6kPWGa3W+78GpSW/ws7lv0/1ufRJ31FTldVwwqt2yNNdivR7t7fHSi/cNGOMfw5FVcKOFTPb3JDV/WCn/j9f8DBQ+Iqvnlq0cgxFq2tzhd6Peh1BSaQ0m2ICAqEskxZ9uwI20QLAQ3XcUEMp4okHq0vKNTQHnZogqk2wQ/TSmaj29EvZcYk0g/QdtWUAFQ80ZVr85nmhN90sNSO92ilgGTNLNGGojYNFa90wDS8G2ESLyjuDFAn9qzXIm29I6J8xf1pIr1lxKq0R8TWtw4CAwJInFvoagfZF/U+goZPzQNEiL6jdKSUQOeKQ+dWBeLtfzgUJXJun+z8d5ve8ODBh9+FpQd3mUn7InFNh2n2qpch0CCOreOsGp1qVRQVICG3kT/hnA77Q+eiss8s8BLD2u+ZhGipXbtuWvjj85ci1v5JNB90d31iyBiYcsUyAJqH1PHyZk8BZ8jhkIKEmCMmCgK+bPDorvUHt/0v2lt5zRhWJZRhD0RzqYMcIIIypfNL13+VwGY35msrEA0lKOHNsW1aDoM8gPjg+aoj9zMPsDDIptaLDQuL3imJ1yGbvrkH3rEi1QNfW8+Jyiq2NHGoUZIXY24Fq9TKQ3hUXNamp0Ndy7hndm3wdTTrKxKrWzHeXucqCqv2huN0ETJkHj0f8tbwHVnGnbISsoglxyRhrN3MkOBe366/J/QW3NDSyqh9ROBsBz9r5DetWS4jFyQ7LoozRQh249UIDdmBjs0T2Yr3EWhy4gVt6zYO6BgFVz3QZm0O5C5+knPPJjxIuKiFx3WoFwFibJr5MK02Gbq4AHTFDcjgP07hDvCpD+kTbYtjd1x9N7Liz3JeOjLUJtjXHxyvr2iZ5AquQU/PMjIXe5c/osPGrnYVm2wSui4alKEBAD2p0PPr1rXRs1RId2E7U7YJXA5AaS7ZvnVGJgeWbLYsTOQg/xC3wPAD2GeB/TJCEyioECdFi7U1VKtPKspvxb20fjh5nK6hBRxK2kxp46NwJZFdPycT7aVQnPgAB6GEA/4wPZ5h617o5zaG0DSOA3Dl+R4cmRqO4pcRBpqpTqBnMvu8gJ0pc0mKecmUAhB48Ney5EOnqgDo5cgYzAOWVjqn5AN/r+litLcIXAnergYyRJ9mniXIhaJU8Xv0PNjp1jcU3zYkdA3HrwJuGi4t5fzb8JZXw6H7t77xyN+w6eFz9N5mN6yam3lZ0ghOgrYid/T78oi3a+qYcG/vCuFemgXzg6ynqp3UbjElDwFyrTrLvUn7PhJf47vvDvE5tl0ni9NLxqPdRQ7cB3NGY9iJD2v2Ccw2fRRo6Hc8eAEVJs8PI6GZUv28m9G9Ej24jDAmzDtjxHfFqfoHe8eTBs4oTiifZVxv1xHyWhhAA3eoUizfS5JoawVfBTryMwX4Te9wKfI4g9QI7MPw/q50rQzBqTV1jj3krDkujfoS4TqRS4Ud+TxxV00lLGOnjUsk3jU00DJV2DbvSLG/JwekpGYLLDZM5su0sqMYfEs/H4XWuxAhqKFgjR/+8PF/FoSX0+nycR7tWPmbEYNXNvhD2AtIiFyEnCi1g8KmotL9zb2Kc/RgopinUQMKRN1Uksl3dRKh35NuhFXoc7VUhtFKlvoB/7lxjwF1KsO/kpcnWZ5KWMNBhBrQ+m9+X16ZtrKwCMYUWEU4MwHZjnuiTt4Wqgt/ujPwbN5scjwTaMYW7MHuJWWOG6Jz+1bbDWjro+3n82fVEksXi3I3Htuu39qTTSN19vF4n8uj4EzysqbhoCLtnTU8Vc83Zctu5xSt/q1oh34CpFJzCifA5FM6hZEBH/Z0zlGfM9RskoQD/HZsYmYme055i9vMKz5lCEfbqO9ghDN9UpCMEx/V8kjrfQHbrcD2TQ71vi4qSuIcuTiFTk4cg6tMa9qohqFu2U3FuJqntNEGrOB8SSXPIlV/ZOCoRc3ds95OaGYXtEllPGeMclCaJ7uHAOpr5djrIq+vBahD7yTXpMKz7ikYNCQAozAa1jQ/DgIngv+gMVv2cOT5kvn953BlRy9aG6X9+WNXgtmLUHnS4BOLjt7jhzf/zryWzi33XSZjAyEGzxQyclKiR5151RCUqNaxPTEX+Og0uzCwAs162luVkZ6xzPHcGYC8V9DNZH7EAbGkbXxAAyN64QOBvKg42oTXohvElcTWqdt4NKA7JRVSFV0TcC2E2X3yb2geiaPNE/loUP8gP5Du7a70Ais7stV51HPLSB11LvxoJ8q962GNRFbV0cIBUv9HWRmmdNXya0rA29JMh3tzFEuDXJGuqbY8kuNAVbmTtno8cVZTH7Yw/Oa4+jsgNSFuMBTkzNOxmqaY5h8zpER+X5bs4Qcg45Fnb1EVUQuipPhrWA3dSIRLsRy4RguXXsZTWnoL8G6tCPKOrpvjuGxisU/3x/EHFrHD1+4Xk0knoNWy+hyGT1Fsr8eg4cHxwLjXBO+XkBkIUTUe4YVMIxmMTBfSg+CHXiFAKOtsm4KzZbVlqiNiQ13Y3F2EMHtMUNv7646h4xu2w6gEK4Z/qKgC5/F9rSTUx25QbyaIRr+go3tnQmHhqnMyjkWoFcFIyl9A39wBY9G8+yS5QwB5oUvvsg/whCRXEMxYDpgrBReQOzkmq3gTiJDjOkjS1C0TRJGWUssJDQYZ/O/LS8eMEH3evxrvjLmcEfYKStkefAqWUVtFZRfgp3vgukdFjUrhv8w0BdFjxaAMsv+Lf1X5pelflqEGdTgIIE3ZJPYIV8/lKvY2fjZ4loXpPwt8VZt/Vpt+iBluFSJtYqMz9I9sy649YOG2ia/QiTokcznsbV/hcnfNzUzJPdyk81UAiP1whtr+dzyaSYSn/EAklH9Un9J+XJK0oaVIuTrkfDbW0dABa5EAKGGc06kPaXmYGBNtxHGR0aUHcQP6LeEDhaxqxixynTXW+bvzFz6L/DtKydHKihLHoahc2wIb1K3CRKUM85E3ZUTXKNZX7j7inXCwIwQKhEZuFtJCkejLuhctJd2aofRAJnNpn4az1bZ3Nio7pHiLcjTD9jaRauRMKLt2yN9PUY70JOmFrEoDUQll20WroUGinOTIEhn43zsLT7Zf2SgoBdKDQ6sdpynb25aJmH3vboGyzRXnNLEFi+dnTSwOVUX/emePRqM7veRTiOUPN8kVZNFCBZFpibBh0uAH6S4x65DemAw8sa2wH6MVl/GodHcet1lWL2/xG2aDqVhK5t6YFQsK4z4TlJo5esrPznsezSAQkxjVv0Y+sVVHMRD/kz1f4xvSYE42j/+A+SzrQ5XfEUhm73+nJAxmDJscVHKs07UuPmoY1/Kx/cOkNmnfFJSdGBkTgpZYFpqHy76+5bEJ0jgJM26qXh3/Mu3WdiVgvk45e7vV3vy2F9hPIWaCq1pC+yUMbCuXCyYk3UBWRig4dkb8BgAneqvviWf5Oa8pcaAW08Z2bSEHJVGOXGvvQ5sq3nkgeDwpZ5ik+yFfYlkMXKTjaByTnlMAnvf1yxi0VrAyvHJBdXrbHHkpCuUw/+s2X0/2TZr+240Wg6QDzT3t6qOEYQDd39V3K73uS+RzzAAvhvfztfmJ73JIxk9Bv+hNsdvaS/8jttEGMkgYq23KBvdq0SYvHlcS3Y90ayI12kQGFYuVcKScFvloJdsKJWALHh4L4F2u2lVlt8oVFY3G83KoOH+N3g8KBV2EOQRDKq732n0K8qp07htCJmoVkI+CpJeQLIibQ0NgdknbOQbwwlAHgsRDOkz1s7bJAIFuYp5J2o3Gcn8OW8wj9ghasZNoCxdRflaBpzqy/tcTbQKsaceXhlgawExbYEIA82cmZTf9Ys4Pvs0uvR+3t25YRpD4NP18xqrg3aRe8RvdkZLTxpRTVCUYPJ9IGBB+lpe4f3Ap1KoXEdV4kvnPVZI+tKfADJRAAvmfONkow0RIt8Vq2ZSDJXyb3YnfRCUZpJ6YKN3tPvx+c7EBGIk5fDlskxr4pbRFMJmr2nTCOoGpP51wkuoLUY6O/jcb89ubUsVsiCzF/azIeqgz5yD9kORPeGwSutTMDjBlw/dwkD8uzWniVo5mucYkX4JTgKH3caTfoPPyIifxueLBYgidV9Qjebt7dqP0YsUwjJYSSzyaMD5aNe3fWo0zKbXsXqMP4K9IFCXMkufsHhtSPmU1gAqQBAIyLkQ2dt3iCFM/KNNlvwCGLjxhZzrIPcV5q5epTQREfnvPTqpIUdDGeI4cWCNOpmksYi8qU/fkkUspHbAkwPGR4K5/EeaMOV84NEAJfUNSO4y4Dr/E0hOW+7LBNdZe6Z0fSLYu7MP7OGq1J2ZKXJx0dVzIs0xn0/ugDfsP19hQSkPfkJqbLeZxUZvhiN0r50k64e6V8MszQEBmKrkXbrHaGxh2WKkqnMw/TZ1b/fWwhCHeYLeEXTyX/CppiQO3QWeTJWj61qVWWPTAiLyFnnXhf5V4kq0h4tnj65xrc7aecrViQnUlaB5//uHP9OUzsswYMVFI3uXaa0GlPCWT+5IDUz7Ihm5YU05eC0d3R4H8olaan7JjmVACL0hzVckKe2EryCP1buhCw+OY3loAIqkNIbXlu79Mwlcluwn+0YMVbRnTDbtZKp1FPR7OZqZ33qNxDvkoZq10zQ4K9UyKAZtNTxD5r2M79Sc9Lzp6RAJGEnnAd+F0kQS4U8d8DLSAqXG9r4w4oNG58xK+6uGaF8ZIKuoco2Zfc8xkA8h+jzaTYuJc68TEtELlVQK72D1NiJS0vaUjXzh74ZVFAwNOwClVBYKytmSntLUkbFhRPZ8nvMwgcaFwlsMN/wZHneY8YtAOpLaEzeDes3nHQDT81RmHRuwzkRWey0dOeeKKL8qJ/Swu6+riMW0jMzPznaPOcLNqCEoTunOlihCpSXPJksrmIu660+4G5sfc8H+XgDVYORFx3HCvvzVnI6mIrrLxc/j9WEMCgkqBi7so4XPNMdx/w4IpdltP0GrubipQTVKmViStvXrV/3MoR5MHwyl7TNAwNsTx/gv+0M/kD+WsuFFtoRnzxmF250u2cE/fu6/wpiabsNpluW2XO4HKK3hS+o5iobaHJ4WrY/2mG3rWt72f6dSyvMgHkTd7zteCYZSBW3uf9rREb7JOy3s3ZbmZqaCh/qAZg1NSAMULldZCvC798UKdFox4WB/Ew+oDWCV3OZ3JMybwm7M+AcKGFl1fzdfRaFtWOxKD2A5x9zZ+UxubXPIkCbW72A9T/oyjR2/6WvZH1n6P1OsTAeCUXJRikHZF5QgkgWOwxCFDu4KizoywWr4TZLw0RymsUsKHfAek5NEHUeCbAkXb2niu3Aqwi62wpY24yYJ0kLNo7YYi/2x1aMiSnzIcPKEX9v4nrXqL7+XVNRYpKrnOxBTb/U7/tmzR5hRylmBqA7ygdtXJgZCaHz61nSr7grJB+zXeaIlfu2Npiy6z/dlWUkAwVyv73DQeYdGr9bGwTPD/xI603NBrpJvuV0h0vDnwfKPADbKru3aQMgWzLF8b5FeWTlgZ92OdTuXHuqnhaMY3GOTZ4QSq/x9bNaHAfpdovOVE3rSg8BcRZDgy50L+IsR1KLWmw65MzTfaI6SAQ71G73Kh50QJbSjEcogOVlcrQy7C0v2yuOcNUjJzR/SeGJapQbTuSOhVIpvueSfa7IbwQr8+1tqDuaR4+gw4Q4fKAsXHiBo2lB6XIu+NWUWH6JTxDCYjsByTPLbKO8XVTsGy8RhpL/WGZBlYOUalgyxnOhVhFawgF36fbuYgsAULMfpm81CkyigeUJc1gKg4F2OvIfr6CzCYdjFFxnIsN9zvdxNhdXtAsQE3HajGUWQLQx1oG7mFaJfbH5COu0urMv22HTZvDXEo5vKpXEFI+BDLHHubZqmwrXvW216TpiK/I5m9oQEXL8AYswkTU2eP2UI7WTYpn4cqrVtW0jnZODeSqGS70Sru4/LgA1MgyctUvcBfP7sDzjfOmGc8mB+ap3hodfN8KuZN+L5aZeSToKCz6Q+RN9LDDJ2ABfm1p+p5ezECXqasbe5FX+wg445YQpEXadCjMFEmuOK2yzy+J9taTSWTTU5H/JJFEVEXErgJBp1027YyZkorr0VXz3uO4jmtci/yBmJar400/nAQSKBtcRJ/6a31Uv+fc3OG1msAOk+V4fdRp+6EDsWnz2DuhEjPcFqWtDnm3ssRISL7XP/HbRgVJvxSrbSCspzx1pPIln/udBbTM6phtN1HqKdU1DHQlpjHgmFws7RDOkIoZhwhZlz6z+JuXdK+eXR/um6DfPYVe90pQX05N7RqqI2u5Gao3v4i7HTTqxbK6H+dweMAWxuHLu2+jYF5F4J2g8NtbjvrxNBhlwv7ocJQrmboihuEmtI0iiybxXnA1fexHBwNG5EM5GVvO6pQeghyZOgtOWKOobDAJDxbDVvJZtnJz/aHga4i9d5T1KzwdZ/de10v7S5969xTqj3bkEcfoVFCpCKcmugJdMMEVW6kFfBGGW1ypF4haroiRIz3GoIBLmxGkEzi1z/GSVGHy9a00fOoqCmQfx7lMuxbUJRiHAqyo5hVoHf2Ygk/YZndKPUiSh4XZpabujBnFQyp1d5pg486mYPnMRRLh4zxwHJwzW1qJ8NlVDySHP+V4aXemm53ul91NPXRRcALD8bunONwhS/gLm5LGY6C5iKrS7ao/JxtdZhCdA7t/UkNyppSdj8zrtFGM/XcJA5ecVv6Hl00BFPl66fVDrdv8zph2jR1sueat8tmfSiWylv+STSGu3dkLGQ8981QIQP06lT18fz64HVl6ew/0frRycJ4P1niC5NaZdq+8TONtvTGfZpw4yskqja2nSu4fYuIVVzPFH4xMV7eHVcV/MD5eKRt2r+60TgvuqQd0qbW0l/zbKt7uwmgUrf8SOdfkwKSDIonRW3gkm/IzKn8QXe5eAYHLfTk+NmwcoKYjWiHHNA3BW963ARYbPUmmW6OSdAsiFuzzyf0thp2SeJFXt9FV/STiUivQirmCITMZok7cUM1sxcu1faB56sKBkHBfC+OnH2qDLPRIzIpFNfCTfIrLPqXcXdSA251jd7Nsighb7Imz6fTFMkEDEtXDonmTAdwKPtQCwS1oH0CcxlYyKu58lC3wAQinSbDvU4cnOHtNHlo0c/jbqif9+PbwX7Rbf2HzGVOk2dNksCrkFKTmJUbeVX+C8CF4eEYKRfD0OnyYlTbigEOg1IH9wJhYNXdRyE4D/ItJg7bDXgI2LvGGyPosLl2o7Mrp9FZIqgyAgFuRoEp0luO1BlhK3mpnwX7HO4u+rUcY4XNv1OHIh/vPJZGYq1FzrSRlEPpDjZ5ChnlD7UFLCNgxQZgbTrpcbObpi7OPpASlq7cBYIiG0964T3lus2oA/IzEMFftWE30XVDSC3GOCbbmk4cBwOHj6cjiheVVIVZYNfojwiytFHKmPIz5C8nsD1eCRwNDGMK4tIBJRvIM2x1TSsirN0PQwYKwB6zpxXKZHF0PmfMOoE2ITnrY0NfySqf59ps1yuQKtGmnDC/I2QqcwTTLAZpyqyLLqU6Qp0hI8r+8zi87wUCtN5Y9PCF0hrqZa6575uwrJO6Nn9RnnAX0tF+Ad19JEvzYxn5C1xSsFpqyK0eGqLZ0snpGVi7WoVF4PqRchoX+twoEeDvIxguv4Agql2Aa32/iKroO7FhczIaCxFwLYF/WEe5oxRF6CJBn6p6qCp8EP05EUVeX0krKtFHW9T/FqGeExs5soKcruYRBrg7xCijapskMMm01h27Ppu/4LwRbVGfwM2TOlKoA3HxFySbmpBX7okd9GeRHGsn7JE+BxiOsRPcYpOPR122YVlZiKrPk9TyE/RaOg73YO/xUmD2nvHPlUKQQE0JIGXK++c5ST9bVuIzWzrt3kM8KXSiBd1nVzXj9etdUDbmjd0LFb7S3HANStDHQ9c32xZJU4u53xRBjjq7xXEatspfVTfpGOWYSJQEKcUP3HKV+T7s4wKwI+DC03uBDgzgSh8jVtQwJqRn4OKynJ1lsDFOhS+ZpPYIWieqMJkkMTFVY5gdPEwFKxwj++HaG28KnjNvMqNw8WdqpwVkb4j9IKsAZ7ZrggSvfMuAXGI4GxQrCVwuF3Bn6Xqu8ALuY6Qhxn/GH+Sj64QO3+m90kaFCbCjN5ZdhGTS8qGrsp1dQaTRZMhVJgQ9bqPOjDBGKrYcSBBJQScZ18mdMe3lfCCOaC8u/f3fIRN+Nw1RSYgUHuUgy6oyaCvrHaR0QR1mwd1VaGu2DHcwP+M97+/3uizN77AhJIpvRnKPhACOumIht48NIyA6gktCoBcSADbs4DdzSgf3d7yCActGU/cBfKEMXKnqMAfXUxoncxk8w39NySTF5+Wt9GJlkz5pKWuI1zQRgJCgGcIMQFeL2Gb+h5kyyDOEjxMVZxkauIk2B9D/j/L7fh48VdRvWZXJeXaOH0QZINcpvY7siOCpz+rWM7H2lcIZ61WisDZCsdNwz4xBDSmSUz964zPMHhRkNT1SF1V/6pPYsiOL3aKtC3iZ/yaIw/CXImpn0aI9GZPk3VbBVjHlOCyGN6yPBX1NIVw8GDCCPBISoGRyyMNdsdV2zDWniKcBeVoCk82zYlmj3h7aV8x9hDlnAQFLDB3ZK+bywhzJZZqN+3QWj2c2BoxcXka3Cd8qJPTsz3zJhLEChXlPCE55b9GgzNVf0iDlDJxFjUEJOg5FAcg9MfGgJAubyH11ocZcuBVLXWs7FOnauXW6i9djFgdudM9pbbKa9zpoCtTISLbfaUI/LUIXYsZ1vtHrCnp93jiUA7MXqsXPSyRtH+Agtl39lhvKup3SZXpWTJdpO4lW6rVcBzj8NKm0GVeoeJQqKgpDLUD7Tj9IPTxWHO9V+z3it+xqsKD1UBKoqDG4PCgBChecs67+TMeCHIyGy6YZZPlUaMyHEg9/GCkHQTcbOUe1cyBXvW+mKCduU9QWr3M5k/FrPRVsizGqQvccGxcQgvzjAGm9DSQOj9QALR3ZZjPEuGNUZlSbCqbabMA6hO0KB1qhg1B8agh18WkGsreXsOUxk5TqcTMSxINsXdUi7FdCnpq1EYg+3C+br1WOZVSxZrWP6Z8cjhLez+MBmjvAdMTPNML82JC/631Hub9MGi9IKEpJXi5/9W+52+Bb0MqNjm/O6sw/qoD0LAI+gBT6iST6LbYMEhmk2v4N3VyzFle8mLPuxnplsNPv9LSI6dUAVhF5GVhSiuPwhg8E7SZU0GFO8aSVvvZ3b6NRf9OVlO+o+NIPDfvOLHDdrRdvIVHe/QFTlBocFFrsTuVuOPD/TJC72NnsZimnmoOsliebhaPNMbJVd0T21Ya8hHfWPzBmZuwSn3UAujXJU2Zw4ohtFif9vG2gsptWznfGv8h/AKwLnlTXGT+ZxRbLNOQDoI597NlynSmG2pKQ9vBjZyJ5zLEiHuA6JVcoBzJ6mBoKSyS4Kp0KQ+Rj+bQkJj6WEJFBc839VvkpgvZUyOjd+NnUf7fsor9YYzyUHYVdrvIZt3tOxVqvq9MWDYFakrPco6biZcG49IRZcFKyH8ujvbUoVC0zaiZLRcQ41hywuKhbNy+IreSYvIXKQxqDxczm3TsR9YwiMzm62yXKX/3c5KSL2SO0gI9EszyAKgY2yDetPvr4jZPBwjwkjSsLHhjqw8w2Ab6ba1gIHb8hT3BVjE0Julf+1I4d4Mc15Izy5gkUzw6D5jJOzOcKk9/qEe05kJF1Wjq94P6k7XoNeBqjJ/+eMAv6gNTg4NocU2sm7mxl9cF8HVHXgPzH7KeCX9K84LXHasiNyNIGttd+9fAokmE5CgiEE9numjrny/EASZspnAjAhxaPLPN1XgHJ/WykYgKPeYfpkT+r/sRIjN7yZq0AaxH6M8z8MUs6LGkXMd1TFwPrL1LPCJGAuMs66HSNy0sgPLQmnLjh60s8KvTyltIDXalPl9Wm4M7AO72vDLQLi4WuH6bXLBIsTcS7REsYySeO6B+3hwPn+SUAL7k1pS+h59yCSLmoT1YU5Xp8BV6yL4TQfNXNqn1i+KjoqDWaIPT/p4KfYzckFz8iGBz8LSr66xybAqshtGZMCmShbgY0QxTgWnsLXccLI4/TbUpxAk61p7T++ruu10tjVNFxwTr3Gjm/q6QZPkk7DQmrusrWc4UASWav4XpFatAl7ESNnKTfcJhgOwOKtv/7lVfCbjyE4Ou1hAR20OjrYJeTdUSUNrvhP3WC7BIm0n6RQDhb5Y7da0AaTV+DK06KKtG+NKtS9881baYuywgIL0Unp5YOFvu+2Tg5vr+Zq2dma9OPbtcxvkHJPbUM3TT+gaL73cxMPbgx8/pwlCFrFdGeDyRg5FLZ8QAGPLImlNTxANMPG6rsBPtNvU7d7t9sBBBEk7ZknK5XeSEQEFOiwPCJ1znPkSUQ4RjnGBYduFfCTxva3evF5VErkXMW90EN4JozASh4frvdJmqW/6i1qayNnGTQ34z2R2QB7sYsC6Pexl5LRqwvYpZIglWzuMJOqPvMxe6ZE/Ek5/yarB5mPT3p+yCNkH7rstMqx5YZQ6ujxbhYVHizNKpIvOwxA3OLPnBZkA/MWbaz5VjTuUjo3azegl+hy0IgRjsdc8Mf8BSf+9ag9KZsxFhm/9OR3T2kBgr6QVcL9EWCAYdP8DqZTg2KLuEBgnzqqfJg0DIaKefOIMRJ0uw7RxCKDnSkwnktwnP5PGMZED4hjd7TVuETjH7zCgvaKpv0ZndXxejVtZA4djLl4POM2uPDaaqaflZQoj+MP9HybB6bB2I6hr04dGImlumIvr4dHNqXiiH+TwSStbKYmqXsqrr8PpCnvhoBtDMW9OMBjiYDiZlhg2e54jtVWu9/tFSULAOpCY7npUoJTUKJIAlKexiDCPOyXMdh5mPpMYWRXU2e9WXEA9xSqcoaxdfJGm6LaqaUU5yDKE1KbDziR7yhsEqppx55I544TrGWcqYof9GiWcufdiawP4MBwzKVIgvsS48Ri6qpnA1nEL9Cp2g5YEN5JKwlkDPOWVy4OmIBIxZPvSWchl0RXE14gnuloY5x/UKPwh0a69qZu6JydCITVCm6UR1/WOuWQyrwhHt0unYHSPw4Z0YkLFvPnnBrhrwVA0vpuaaRbDYhDmNY/EWnTzDb6LQSmeZWcd2M0LtP2woYqpEuaGkjPgt3xlpMOYDMjhCMLc2hXl3InSA/9sTteps6d+z38LqgcFmUDpRnMDhsNYEEQnP6R9vpDFCBHzdGd1YaxaE+Kk+8EdLdyYPmea5Mds8UvLGTK9mESTu3sXMocGuCZALeUb45Aed326bauXUfnEvih5N5k34OmnHHPRtd9chYWo1W8hAxbEOBn70RU4FivYKN5F/1kRl+qx/rwiq7VhclHWtLvowRJT/CIoH3QKIkEM3difYyepTjAbgWreDp+YnZkxRczd8HHSyrQGUwIAuyJ0DFrHWYcSofJorZA3g9cXH0a1oQ8y1B94kV3C9elYi+yyFxAxp45oJ3IVCZ6ZGf/xofRAn/n3dlZB22RaVqpb5b1Ezo6nO3dCnzO6Kd1eBlrlkm3XdNzgpNPbeqk0R94+b0SZGHiO5jlu51dKX9XhCOldoDhTOWk1PPVRkWU6ksKU/fp6o0j5mcF1dzmba/caDoe4hPAzy9MSxAf0b1+VN8F2SOLSbukaN2MC1qvoWr9mp8j21D8PpHRNEYg8oNzB2KxenSQzny02z1AaOw2DWHVnFWbQAV40unFPebQWoeGISb0CqpnSC31WwtlrGkWUQzzDaHfYoGvHITpjvGQVzUeEpsQUlTTdrYumS4aq8P9G1yUXAblwKzzhviJXNMnvVfayCMKaxxLTK6RookotLrW1bHgg8yq/OilKWVcMBHdIkBQgR4fu+5jDvUBFtnINUeSmiCA8KpG2X7O4ICBYYT3dc+pPM6pKabLyd4N0x5sR+I5SleyWeWuTjNQUmZMInHmqmK/sy00Lpg1V1LmQBWpUzkAVtXclmIRqjUDtDrhkPFErRUogVuNUAZ8N6J44pAhkAqANL+EKE9qKY96O46pSMs79ty0ruucHsRkSzWWXO10r6SvApUArdA21PSt/htaLIJaULBvCmdry8dlBDkB+H8Mf7kzuDOHgEyfsIS1KwY7+0fgGL4UDsAv48ZbTTEP4G7TXdgXw32S+ZU3LXURHKPIUcAW/0UWXP7SW5ICe7A+QE8pOCir7mr38RvHbLP4btoYAsoFFoMOjS56adnvvrsF26YESyS/Q+hbK/R2pJxqZzLH9U2JFY0EztWkIkEAQ88jKNwIchf4BDx/iYQ474QMHE9YGgKlfGBLIR8Cg6MvsQMgcyyluZuq71vYx5xraxtFtBCER6HnbOofu9fXJU3VKqZwkcwMgSeWyTn+dHuHXfKBVFI8qs7nFZZ/x21yvUAEg5Z9KGBidtyzqHMGNWIlszvf+BAfPN2EGaaSAGlz1p9mRm4LqbUjsLtY1GZ4foysHbANOii1QY3ZVTAh91LgG01EIg/UwCZ462KC4o4DBN6NbsQfbwy8SZ0CW+AvqoiHd5y7fyr7GD0co9oUr1Cm9GhNZY6V/j/pmu/9/NLRZmo5uff+3l8cv46dSj/bQJincsrhYtyU3GxXLXJleH1xBBMrTjcY4YykMja+NNLDoseszxIlVqKIgkabVWtYsqdubKnlq/hbZPtrTWYhSwTzpKCREXas5rZdCrYXDvbRyeimCGxDqvGn9iyOvYfJ3wmJYpae3GcVeWRrii31L2lGEnMwCZqL0wWliXP8dAaEqgy5UTEi1QRgb1As5kt3Oj8zBcJ2V1hK1zQ8/mXGBNGznwaP7v53V9eJpnNxEdB0pmU9/xlHi+e7m0uCwN16nM9O+qwd2a2dv13vhj9k/DSihjziGPnbamM91ZCZKqNH84M2qzd8xBvmElltX2JyN/GCeBK8V8i6T25tS/oIT1kK5JYFMua0Oy7uyaA8osegUf4wo5dDFSNht2VYiBrKkeelUdTtpItErVTRBMaGfUQv/G463tL3c/hJ9SFGhj3Dpxxv4PyHoSphNtmTUYVNUAcWjtqQObLmm0SHGQaQHupz/ORwz/OPzhitVxeS9D2zux4OHKFaEGfZs7pevD9TzyuW8LfYACnBokGSX2wkZbYkzYnmZI40ndpGrg2zxzx3u9yr2I9vR4ApMJJi4h0I0o1opcYhZFcxPmqps+QRkpcl5ZutEGuoXNeWndcIk9QdV9Kq+WPI6o0NMIvgvW8gSaLG9LR9aYHhVeHJ0hpgtyq9pmMz6OxY7Xyq95T3/vx+MzMRA3Rs+KDMsrytvBvqUGiq0T+IJk35ADypmRYVRDDqjldNmuK6uYDur0VvQUZuNPk2B6DR0xh32Qvuvyd+BvEHFd6QCVwnUSnRdJvVWEfhE5TDAys5T5ZfYrT2FH68pdNS91+znBVxeXQWZQfGs7yeM3u0bTUkrIsKGUFr01as1BcRr9E/RVOmVvMsGR0beVb7opGnI6LDML9lvypfWNtOnXbzgkdKf9Hfavh81JKzOhP5nZnLlsbK88zGyil+pzpwkvzmfHs6ObTEMXVeB2iKXvTcJ/kXlNXtm25WRnACbn9wI80KuAruHe1aXRogdRfa3H0FG/ZZYfKhetlBc7CMmxwOyh19p1OttSs/pOipETqSWQ3DdFQAMlFYhJ9gLTmCNmrWK/obj8DZColIGsQ1jCjIeykslAIOmc7xZf0DkOPXYtGxvaBPi0Wki5apHd/mX9F75xhaGzgfRsRIQyZzLf0whXx/XesxN0FOi1Tp/n/1MWGg8hGQuknt0VUT7WqiuWvSlvw0gH6wJvWaW4Gp36u8J+1lxxFkZldFh0h/dlqpsjl2HifS0H8HY9AwlGxet1J70BzsHqEZcnkPJlN5xQ9NPthvoKaqLsnQ+WNMOgnPa579Z5LdLDe+Degi1cRYrf2MBwVtAaRT2DtL6mN6At6uTWOMFIajQQK304Uh4BIexMT8aHHxrZQdBZpiChRBn7/StELQEoDazgBjnbwwBABNer6H5HOxUZg3J3hkaVrL5SYuPulrGeJpSNbachWXqvfPEquSolQGID+JDrtkYgOzuilXYrkLvFsHen5shex+UbJvvu3BrOK1aiZqH2ImOYvsCINU8cNCU5sSpi9Tq0Z8uQGux9Z52SebN2d62OCaNkVRiumOTvRKMdQctWkO0a5rM7omaRFxHpWyOc7r/c/QHjDJIv/Gz/TyvtqwKw+KEUI4X3aHjWenQ9FH80y9C2bnx+YJHS/V/KFABBvB++yHVLN7FtdrsiL4s/7ZGl8B3bZrzTxZi8D4p7iFxtpyWyaz6zipg2lduYLU7LRYpKZ65bD1RhQ8L451ihpkWYQdB9QiwoIv5I2gY4pdmUP+8GM/ozxTuZrZ4c/v6JKSgrKF5PjRIaui32EoAnWx6iySdqu2iPrsb92g/i7AGvO84CWumenIJZhUl2ND83NI+ARl0PR1nfvU7FqjgU3et73KEkPVRkeUopRuRWhZdNbXCldDo/uaykaeDqVkOgKGTXrpfackvkn6QQ0e4Sb/MHzyKaAqCFY3ig36rMF7AVX807N/j5HWytHu9CkLEcNlu+XOAKSYPd68cvwmNG+TXWJnIaRq6FDke1UlNyS7zDvS320/OdhmWtaPmveOK+8p//x7kkdbDqCE9SKC551rE/h8ocB2qU+Mrq+UvQGLuojwOJ1MhIdEiizSeqGmBR82vjRg5NFAxh265MciSndmMHaU/bSCbcDjLnmZk/MYnQCeBx83zzv5bbwGMwnP6frvGgHYyqfxxrEO7LfnCixmoh8vdrl/Jgm6iA86gp72ANkd3kiV2CA9Rb2QmsobFSouXq/ke0GnL+19a9QYqov0g+Ky2/SerCZFkHlGB3LRg44IsY/fvB0dqdXrPcjjXw1VCs0U3rIffoOeXXn3ZP/MbZ+GdEQpJqpPDJhmQAavHCiyPZkhLzBDgjEK+cZuVv15f31D91EtDQ9MHU+6U6HEm30KoU47ofmMRul/5IK76DWqhVlR2YYHYYQgD4W6Uz+Si9LgNL+PzACfJceg/gjAfPQn5vZpLRj41/DoqPpMy0qM+jFazSJ181UknBC9ZAWI0HSOGTAej/bXzgWPo8eDNMfMyPPgloMNgIYea2j47f6c01nW9b1n5hNvVyZ/qnRbtcyro46Ceaq8HORXItJgHcM5XC2K1SgGK/9y3dQqoB1m00UmgQONbH/Kai5HIuP0vj+833gD9EZMw3uysI9Gn23SwxeakKDwHAYqYkpBv7U9ywN6YXmLA8uTAoxTjGZ+rfm+Ea+mNPNq2woLrPRcxPle6aLra7k9poQyKYQr6vsOaN2XUuq3BZsCv8H9v+fOt3PJ3eirInz2QixRNYmFoUENVBaRqn2x+R78tCeZyXHjPuc94S5HuOrRUxnMdAR3zoF0eCvJCcHSPm1uWKVGVFUPI8DmO1seHC9pakemNrWEK/kAIXWTSy8O2582zjiXgAn7up+QQopI0yqPweT52GqZEtA+fdV+EnIKk5wxy+H79KrVwmpiY8t2RmfHiQlUy+xKRZilmVpjXfczNp7/rArA+J8UBI552RPY5t3Z+8jJTxo+pAxW+8QIZQQIqmRj74Bl8gdftrsk67eJT+bx23CqBinQgVyYIWO9f3JsR521T6myEZMvobhexmYgknMmtlaTqOWJtwIZVtrChClGXlEFQkQzwfPAAgdzjgwpCltxm+JsNvPdEOAHGHoplDqJB6ZPxPPs52Omrn0ikrOJlxSl5tosUoGY5vXkQd8aU0NAbxxDHqzBayQ1BfOyRM0n1RFORZ5wqP5B0WY6C3SdWj2KgSzk6dJf4Sd4HutMzawc/yQVrfDjZEn1fmXbbYhtOwTOOiQn9cQnyhCQoZYNGDh1NfIfyBXkgXkna4cUvnQXy4GXdYfRWvGYd1OG85j2Auaq0erU5LQJqYVbz1jTs4djfyXDYfH5WkbhW+roI9ClsFXU1FN68zhezmvJGLjkqfHUG0Yy8RTZVoIcqzLQQTLb8peLPHrVdD3qPe8+lu+VUQy5mCxzyqx9NTnAPaUEjsRrHSKa5nHq3YCGo09/wAOmx3chen1zil+uDfRwJn6YvC31hvfkCcjAZOqBeUd5+H0dhGkkQs7G0mEu0neLDhDqwZSq2H3YqdTXMpdRYv4BxS7zc2EEfbcHmJZS0dDYjRbi9q3Pog5vov1Sm/zPwBUAPBe1GNCS+wo8XLH95JcDJm9N9WWFqror1ZLsXp2HfGM76lpaLTeXXA3/BwKK4Zq/a+Qwl6QJjRlsElbTjxptdCJkZhmPUJ9kQFxUdRHimmLGKxeSnY0b4y/aG+2WhinXFATGZ48taU4RBjJnUrLwhduFHCdgJAiDqWLP6Zq5pgyOx/Z7pZ8n743wUk4ZH3ynUdd0lv/G7uQmaKcgyHy/CLwycRErGQh6OwZZRMSfiH4El4ffCuXBDda53PEF9xAL3RUO/FozPxucntaHxmZSrURBmyFKvGUFU86K+08/B/+JSV3YVg1OtFJX+HnUvuy4WUyDNZiYv/0yVMw/hCcOH3Yx2jDK8Np9aGO8nKDeb9zFTfSarXXzqI6jGaYm+hLOZsAyBJgWs+AHoIoEuNszyda5nmkfxxM6DAB1rtVWwgLafLkK7kV6HFCtBaBbI2CuJiiEGDkyb6QJgaff983Kfd5Ehd0HKY3hj7WZtT0jkwQgcroMw5v55ePy77sxGpFAypzMlrWJkH8bU5nGyMyVfgti1Z6rnI0Tofsadd+7RedchJwc83N7hgyjuXg7NzoNgNgT6yJu9qDbAPRtkKs2POAP7EYh9cz3050Lh5jWYp1ykxr3Bw7KErEFjHB+xUDISL49MjM65f6Ctx8rXHS8vcj+PB/dvPO750plg4gT3aHQWVnuJwvI011dA32JvqFLvB4QSN7I/FMRSB/UrRR5GGOdmYwX0uAEac6qB0l8DLpyHhNDx/zT0yQU+j812K+1pYHj2/nlq8Cvde0s2Fzql2fjjY3+nChSmb31bGB7jBmsSDds7JOmjzxplte0r3j91qxPOQjmQpEFW/m4z7EZouzClMlZzac2LYYoiiRhuf3WsA8MLd+vGfOLKUaPS34V5Z4AkeHgn9MIm9WekKaN8onJbwtHtVqxDxcZe+zaPUgJmgIU3BzJfRGc0qRcU5EEdgDCoX8qLgbdwBO/GWRfw7PLIQ1JJfqvoJ6Y9C7ThnuvYxg2frsl0xk2ydhTDlvihxvSg/8uLJ3HPe2oOWIqvRCKTT2ahvwNr1E2pZ8Jv/UyapamKO9jj+mzds92jc97nrK67k7BSZ4FzviIFbELEaFBhzkIy11P2iBjCYwxkecucq/AG2Lbo24CwIGGhjkQJoDiflowI5GVFtt5UrLBnNt0vq4jSyqTlouKKkpflUAfMf2Hs+86gRKO07P/hzVYuF+YDhODt0wvGMKjXpmB26Jr0UtKjM6EoCdeC1DtSwNhvW+gDbwdiU43Z2V2Q+8FHb1yIumbQSNMQ/POm2QpB/e153RqfNbpej19GoCCEKW8gg4uF5JLH9qYMuXo7py5iRxul4iOhsqYS7O5qKihIvO6QI2VGbTAHm8cK7LugA4tmWUK25CDk3PQVzPKlNdE5HD7VuuLwZfksx+nhu+9ruNZF2gSsmF4s42O97kN9+G/3mwoSKRrZWkNsJ86DRcuiLjUtiBbAs1PAvu7K6ldD2pI50OndYQHV/R0lCkrR+HRW6lQloraVCYKOd4YTFjfremxLu9yRrkspRlUCVGiqrv8Qt5PxVk26Y4w3NP5yV2L0VCp21wmt9PkmKe/5TKH7tc+Wzv0Lxni0IXu7DYPOUfzhxFCqKYfS0O5OcLNFmnpss+lunWhfUG4YpLoALUA/Gw6g2YxPmpgilOL+eFpqyfFUU4Q5QcAQ+jDwr30+FDXXOWVQqk0WMY/p0ozjJ8rzan4d79VMZ9A1zSa1z3Z05TFQBhJ71JdEIBDsuZM5ZwcNeoHQmNRbFxuStHzCLwYoOr2IAnDoxVXiXIqrYZKZZ41h6jo/Au/7rFemwQyQdsn0+4oAjumpGraKsN9PfmWCNKMJXg+5r8n5vSk3VdTzZdV0yK4tJzZH/VprsGXZdE9IH9cfwBjhyVnZ5G3FHRefoMlo876OkL1CCE3+pXG7t2ZEKr55F1Iz4iYv//Gjx6ozV93Uwxaaj4jX5Zgm/0llN8PK377c6LX9hFPyIJPCPgjZIFIsaFNnMp/OjulxbFfun/cC+BM3wqXIUtf+oTj/sjso38ooick242kyA0QAiZfYb/vqmWczMRm7nL+Y8hpleqLbuSc9va/Y6zgJj+Y3Z1ITJlVse+e6nW6iozEL2j81V19OEPBzw3an7NJurjnNxUWZ5WsxFoYYNEdDBpZaD/2EsxejZA5hiGbDgq7f1xJEWgbH9CBO35q1mr933D9/RZTNvDVOXwvuiQdO92ZVcBkwwoEgmqrQtQJBoMao9CsX4bpx2zD2UtZtbDJTk7E5OM/gH/Ntg85CvSAiVxI4x4o94kWnh+v6aGpOOp/BG2V3GUz42uNeHXpQQ+tKnwJR0v88sbzFvU9YBQnnWacX/TDJLne2u0/l28Yy734nScfc83kc2M955zqlWg32DpVCGrx91SuYFgfoK45Hh4h7qikYtTgFGC++2tRwz2Uaf+k2UoCuDvBDepcC+eKbJTdvwGmDjgNeWt/i5ItNdrK9G576p0ktS0kzII7uGl4OVwVJNtTokvM5YVtP42/TqX+6rMSyAi65kATkrrhkJYXZUKDla0aF8JhWX13xYnb9OhdRqEX0n58HvCqRRQG7JscyiKf98mLtWabktWnJmigo27VAEc92EC482GGKsDgLkRju0rLzs3unVhUNxdn2LVxLqZZsYh+A2XTSnPnRQgVANo+XYl+6GF0Jg3AKmahEGa8gd01xaSmnwIfbe8DNtebKP35J96I2JX9qLVJi8nJYQqwoZvkSmsFJ+qoVGd8nU0NVsQNmgrXbwDd5uV0ZTqfJqEzwQ5hbLSpmtTTltGS1T3uWs4r87s+8ulodz5IUBi7wr+BqO0qArsXNX7LC6Cs7+AMWZ8bsoIkHHwFD/F+GR8iat2N/oSjP/FF47npwcTckWcnQN4+01RJcstsE6eyqWbljQyR2wJ1fKfnpjKU5Xj7oxP7+tRR/QcBDpfnevLy9bBWX5543HntyTUaBGBplKexTk7C6GMS8heRobA6LE49oFWKdy5d9ee5dFOxR9vZ7evyP15ueixtkmtso5lEnnfgBtsiyfzWW48HhBQ3wy4j9tQfxvLl1tSdSILmXm4uCDv6M37zX75rul0cMT0dtV4WJNjQ6bpeKm1BT5J4sz0sa5JsG18SUMccJglAGqoKI+9fq61F8JYAhJXJEE3JwA4ldQoAyJDBNj8wAdqOcrBrYBHjPPsq1+qqtkK8eh4dYGDIYRgJKdAU/7zTlU0Y6QnVgXLWZFImORRJE1Srj5DfsgNYBgD5WPbd0rzCyx7rS37ctW93PMlj3Lvn21Lsf2nq/17Ayii/N2VzCzhRBav2lOxjJAxDDJfR0YyKdejCXhemEto5oIWIplUZ2G++1M12+ChoWxRf9ulAfYyld1BZrci7UVlj+RPBz6lk1y49HO9g93Thq+D14pt/aEqkG/nFGgL3Ndxs0DRrsK/k5tpaGidT8rw2Bujx9LCtn9GTOSoSLEie6dB+wUUizRH5bGkVPNFiiKHBwc2O7OENWQzQhpxNUNdsdtOWJ7uGk2vQ9F8DWCIv+OIZFZJ8AW/KTiwLDbtsUlzNxDoJAZn+mqTC/Xnlkvp9LVLQP+WUKLVP1OAhQyV9LRhzl2ev2ZEqiw/25oNpC+zAiz0WN8MZsbjC5CxwtZjpAoUvez2A6oEz/5DNHGKHKSFb2ukt5oPUtnp1zIJfggl5hcK+QUGNURGqE51GHvXybRaed1QcquM1ZfuZsd1S826iF1VZF8tqnJQCsQAOu1nYhdqGi5czYpkEOeXHYfx+u3EsL85Q35/N8P7dcH+wR1nMG/zgys8C2ujW2JcA0QFzaVlSqJl/gt5Cz9PvJEFZXDoEmN/Qi1drIqfEGSCeqQgRELzHJmMjDqchiznluGGtPUb8fS3X2+n0kjW3PRNd+pSDigf6+J2kBFr/ob9trCLWPBFGuG1uompCwHs64b8F3V/uLtdPh6oacMRgdqDQdA8RHfIrF+mVgmjJZz+10ruuN0P9Ux3wEIbp4i//fnbc0sY2E8lFaV4dB/XtLJLTeW8p1h4hS2TSvXtRCKbYcrIH1UMQO4j9FBxLeJCrMnbxm8LuLfFFbCs/MIHPshP+0RzzF/ZzS/swqLgI7g21ZoBJrj1bMnkqumw8oFDEW378MwgKVg0HBUS7RvZ/4ODmaxfL1cc0D5QHLho7KeMc3PbyvbgV2wyrr9QZkmGxdb8PjOHqZSJz7s69ykfLlokwFmkNMI3fIJO2bQhjDYSmt3K8bL5HgEMPH2zK1SQj0RlzqA1A252EoIZq5m1WCJRQDRm7aKetKu6zB6CG3XTDeldGyXVSpsSXz5wUB6KkXhHhjZqVRChNhwXqoWTwgZ1V3iF58aOxyE5LmTce5Un4+fIcFwfenIXv2qboSstOKi+cayOC5LAKWTqTxLxk9Ojgx/DB21ydMr0YarpLRgA7yVLFq9rCKEyIHoGlZY8flUfn2KS62CwTO/MYHO+80OX6swYMVmJTGG+sYtD6ybgqwxsF2YosL92kqBsEHZF8Eq2iRKGs/I1a2Ws7WELzlbT7IWKSRC0dP3mIN+6Jl2siz+kEYsJnKILe3bo0DvsVKgz09JtQ7EMsCnxOS67tOEqq2N5sG+kkZupEgkHzRW4KvJuntepHPFDmDugbinwqioKar2FxhNeoxGp67bu3Jm4iRBMY911QO2mJ+ormTPaAn+82WoeFP+HjFsIaG6UBU9RnE9f6/nqE9x9LkFtO59uzaTDop7d6TdjvB//iIH3dOjEUSmIFQMNy5wqmn0Vj0IrvmWxZiVYN10AwrZaoaMwUYbcaM1sdm3zzpzMMYHg4/XmLGZVrTsYyJlOIsgQ0FF44RWe6GkTZe2NQ7a3gXI1A6nAGoYrZ2YrRmVi0bR9DCeKDXJLe7g0pmlNvRKu0giY+pEOcaocmxiqXiD2rGxESx5xE1otA5MtEq5ZbEF/PdJhGXJPWSy+B6oYB6NgnwZHoA1h0mkB16nRHRPK0ebKgfIZMUIJtPm5S4ujzZscQK/WRFLcKWcx73I9HddYxhmqmdpEZDsvQzQsf0A40lZzmuH+tRviH42kZY9Pb/RKVY+w6IUAx/q31a8WgjYCnS9xAU55J9/paQ6aFhwtPR2m8Gx6ym2Wry/tB6KG+7pI7Eq0pSVjpH/Tnite8kbGFEgQWWMJH/sc//Po4qogNGSiEDwBwE5OKuPt1/jsPBT+6mOA46OlMqUvfB1vXDStCXn+HAUNyZpXLpvvXi6qufrsDLCZcVniQtiB4T7co6td/IZANpTYZ3L0QO3Lm6fEpV2rraaOPjQsGOY+MlXTGK4jCnvNo2F29a8jUnTEk1Vz5FSmnv/3mD12WFQSZPfgbY/gdeMVPHKFEVT7EF4FGsI0DECxsFxZCumnUzl7DGHUbtdoqvjDcZrO6i310FqGuPUswjOadZfWXL5MxxnzEiONF380iVJ2RXULzV+IlRc0rEB5/Pef9BXiAzusEbwj1DmWdlmHZ8+V0GvdFHmQlOoM39yLxuWz0/okaFFfmahLAuqjdhhlh7hc7zZbhvryFN7PE7yXR7ggayj9VQYDAIiYqAY44kM16d68wrd0WaIltK7kYzNApVsLOzEwlPxGl+nSroF1wNJ3sNkTzoVXshMKU+HWPXbZgPdSdvb4TU/Bsz2RTJUoxcFy8lBGtIP5ex0KGcO2Kd//tuc4nElnyFx6+yF6VvWmD8xlQJkm7uFc9q0lAJXJdT6+AFwtu367qe0O0XABAMc3LSj7toOlHM9rmmDq1QdlfIyMvqwEoml+ua1O7KMCNqPYZBWka43aPBluCbodMg56NUvqyeFVCZYFQyNKKfWScTsrMvjSXT+03VZmCdVN37ee9D9uP2seXX4+f6mGpfSBCuMbHkUs9MDCWha6MXfzOYSdCyoUPQ0rE8K+JVkhZqzhE0WsVba545Z5W6xEr5QjKWSE2TjjIzMvVpOUj3K4a7DdkmZJTfw1JhgJVGqT+81x32/2sX+MWkk7X5tx5YFMkQooPwYsnkaiDzf1E5WoxUvI8nIl1dsU3e4XlrEpWRz39mbrW1owzO6cFucUYDuP8gF8SJdcKDAjvTB2UdinYfdlD1bEGlB76YaTNNDvWlLJDJ9PiSy5rNMkh+zJq4xzB782q4rehst4IoZVmmHGIZ+2xHALHde3TCu01BqfbLJqpEOMEQ7LlzMnUGonlMWn6R1C4qlhkBTI0cs8wSD+k0UWTWTuRYAKvCQ8JvvV8=
`pragma protect end_data_block
`pragma protect digest_block
5b4b4ff9884c39f5594711df108db43edf3e52a9216ac80ce3d47a3dbdff7e32
`pragma protect end_digest_block
`pragma protect end_protected
