`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
obGPGpXxiVBHaDjLZKlo1LY46r/VWIhaXveP5+lZHSACWzYeFGCNfkSvuwjJ1WcmE6mYpce4mlunUKCw9A4ZluY+Fb9yFzkIvfjTVqhqhWz0dK8Yhq8iXmTLvk/SdRdt7Q7myS2PRzqqCN4r67ose8h90MJi87NwNr1CKQgsafGtKvOoQtW93n+lqHi0WL9+tZhZUIq1KP+Mb8svA7RA0tRRmYoS4rWFR898OyiLJj6xqRWCUpzTvOzQJTIkebNwbJgN2dqCUNE4Db6PZdMsVvqgFIUo0/2QM2qyIM/AO88139lfqAhBBJIEqm6UEQTsKinTRFe/+FsYuUqEW6SvtQ6GHTF2Vlws4erE3cDRKOPEM1Gu68LPAg1Ir1MaQmcdWP0vb/cbSsyy+zHO7cCZLttkjP1GsDMl4pgj8IXSDd5S/SYxdf/6kyBqiquptlxQjlyfSYsys06jKe5SrrxSrM1EAe7fXDyVP93qAxaj6O4AMtKrjbZ+EtFtyKCHJKQwr7sjBszYJV5g9EDr7nhKqXATAab/Y1DmLFWHBXINnfWgHWy25KW/PFSuuEfAFw1oRoqBzF6Xe6lB/Jdfu6nCFoXlO/mtw2GXUFU2+rMQE2UCz2iRfV2nHA/Tt/NmkN8eJ3bJIfPkB5dOtsh0klIQA2xAonCthl0B3y4tBZK8KxR9nrW7f9NoLdmJo41cBh1fAO57dzOmWgcDJ7pwYMSJI+peQMR//l9NfM1jt62m+YdEJRNl+FXzmGdR24rJzTy6DlDywkZ6Z7Jslx4t9REZGXWkRwVlEV/RZZKzrnLjzP3daOvb96qKzOvpi4YysKoqqZ4ZraphIdI16bITcDwKxf2VFae+3P9ji5aGA1a/RcmzJ3n3Zpzg1AI8GBOErBcRAY/91ujYshvguEnXlsP6ZF+btbZIlsoWlNyIV4LT5uU892hsqPoZA+tuGurdo0W5gn7mTBnfWgCm4jDX6F5KtL2LjPaBAMIYzN0Af254heskWIH7ln1dF4qG7tLPDOZJSE3J52N35sS/zCVmvgBF32jILbpd0/Bdn/ilwynoUV6aZenbyNjmcedENnaNpQdaTf8LeU33Btmvvsltagd738DTyMeOef2F0DZ7z7MBeX7UpXRgvHqygOvR3KMN7JCCH3KlvaevdUFXG5gMr8jBuzLBwJZ5j/h5j1A/0AVVrZEHldE5DLTAWQOvHg4UtV/RePADqUqnYZJhbaLjN+LnTZlCwSP2O4s9z+WEdmusymOgt2V22oBBUp4I88XOB1kN7/LDtRvhM9MJzXHdbd056k6O0YVOOkXOnKuIzhLIg/eiW8rlyyJoCLJtxB9AiqKkkGx1Fr/gijF4cgVNn3rNf2AU2BIpYA93EcTswDOGvCGf6JXZPK67WV/szrWBumki2GcSHkaHBp474sd/1/RAsaxIwL++BveyBJslIlPYtuWnUjeFVLxnbtWDukg99xGnXbCl2nQk9pzObnvzqhnazpapR/erDFo+rcN4BVQzecGXCMzMjGShLvqp+zh9rKQ9pez746t7IO3o6xKEx+5gTbwdsNZ8GKIV9uQ9OKblSnJgXmVgEdIdOCXa9rIcg37F4r29zTMa461x3Uj0UXMNQcejbekV4JDX4qh5UBYt4fOdlPzs/Wnt4uYdPhpH62VoDr1wmKx0wVGozvBTquBI3nxYGT3JvTzwHnaC58jJmoB3xdiNcihJ6MDgLQD+Wufachy+Pg1i5g5aMvKk8qMQWwZB/GzdBLoyW1aIhT8yHXAaOMwqNDt7DE1423B6cBiPHJJtSWMnTCJzujV1+sUwau8uXCYqIjgkyfCR8/U8io0M9MMgancEGXwHAlYEGKzyHLvvCdCcb4gB8x9xMAWwt4lGdIusJv8RRFAuy6pb8k6ua0VYbTwtsFBeUgscUyw/vBmDf6BNGEF4As1XhOXnGYVxHfbqn7jGvBOnq13MEBZdRWSnHXB8EbPGn12LfCisxvLFh8J2K9DzKq0OOyHqgkg6//SBmTz8p2EkYv2dTszlnuB5pi088RB2D3DZHg6qyK782m8XOgAb3LBvut/4Yntvz2Qu5pPCCxz9/EDV4NljI38gyFM75GrNNEk9Wgmm64Sk5JaolTGoYRqRCJYI27Mg4N4grewO8kB44impStpm7Dx0eB7tulg933VnBp4A/FQrrr8nhnVFWPvCdGxDTZ/A0YOL3qQxJhFOBge8zloiS2H62euZxpWQKi2EnZOs8MKtbkPyWYlv28Q+S+RCb88Rfabn/9O+yGfYWOET5r39mCDDNsn9QLB+TAjtp8/wpvKQR+qgb7ask/81GQyLa26ywz/nZeAkyNs/liSCL7xgxubCcrxFXUnorjJySJyB7zps8rUgrWKt7uA/5ynuk+H6z7e1AdIdN2G/6kTkuUFh0sqs8WXpqsid2J4wrtZ6RcBvo17/6XpnFMl91qoV09+eV/15go3hUy5CrK26G4BOZ/07RuthouCFYUbZCR0HJmVyZCDT7AiWZtTZtl+7XMNKoEsYLfPNaribArf/a/PFOx0C6uYvI/RhLjW2aYNXusKxCkibHV2sXCTOHPc+tklsjtZEgEAfAUZRWuGrnFBQg13MBj5ysTTEVA6SodOO/e9x9UuPssu61qARaVlVyy5fl6mtyFx5IX38OyA2FiAbdTKOlCbkDufp/le7hyeZW4H8rzjISTDvniMycFXnFK73thXyHoq1Y8yi5eQ4BfI1SO0L5hC2x5JeKXhOhp2aQ6sDeK93CG4kaM4CQrStt6TsYhtog+0fT8emRwKecCKTIOXjCbo45t3xx61wZQrQMaR+5/OFWkdH7Hn9ShPoY19Ko+AYtkLi2xVYlXz4i8St5idipPmivHljISj3XtnG9aRuwY9/m0h/4Aisbe8L5+VHhF7Y09n7Uy81E7d+H8Hma3PXhnX6RcMUkDyyv6F0/AwJhcRYlw6DP+Dfpz/JRfqUp8zZ0lGoVR1e7jVHZcGozsCQfITpQeAtkOS24RwQq7KICmIaQiLKRAl4ksVSsJIcOJGoIqkp2CJXxIB+Gnj3Y8fE4yyi9poJxnMD15N4mX86tOkf3sPzpKld8nzdvl1prM6oCDME7p/SDNJpMkPFOzZ5XXc6wxx7qdi8VL8N5FOya89SMvu0ovF/erVv5FZ2BgxqYzmMpwJj9vDs+r6srkb8sZ4BUXL1KM6rGODHpsVRrrNkq0ShPTkOFaj9dKYxzHf8jO/seKIhxSIyOFSr+2V5hKEJXNUbM058UU3Mny5lwA15rV4S2I9RrWDgYTkVxQN2VGa+xzzaXGK5viF8UbVnSiuL+PujH97geiHFx0kJIJTXn978vcAizYRQKYiMkST54C/1IRfp43FKPS9+au2WdLhxAMmpj0C6IQryAqhKaY8/mZYhzBe+8stcyYn80zi7Xgyaek1/bdNOcdBNYEDyW1kPRagWV1mWjlCZeLUUh6qXUhregfnImapWqW68YsoDjsKYI8O7N7dHCOh1v2jQ7c+57p/bib3CLDKAYubvYRchlQM3ZJHufikMvs6pdtGEn+cOYDhcATmQfaSZ2OPnkkoIJNBu6iIVOPVvgacaFq5w3QY4YGmGFr1N62Z9u3ZOAptRyi5wFArsF+SnQBHROLccUVfMlDLidPOCrfPAqutiyUDdj+9MWwFEfogYG3argw8+oAs+pWB6D8YnlaOnTNUNagnjXGB2mKnbykjDk9b/FSweHONSLcjDR6S7A1jNhZjG36IqhS9bEfopCZmHsIIsV1fSVHZjeiA4iHXOwDDB94Tj3HWb8sBv9LNRcgzNKB/muYDQM9VJLb5N58wtN3QwYT/07bdmQFDNOF9w93CMzxYycvfQAgOYg15OBZP1vXopHd9Vnp4rMfEdEuiqw70QQOhrc2gYIzFG0k8oZTtfI9dz1jOqs90YlV1Br9uw3R0mFpGm2RcNmyjLayx03dNRyjV7RsR8AWE5UUYJvFLzkhwwrxMqsbjJR7h4y7367a2rkJw/KBkko+im9gFh6M/k9r2VHw13E1sPd8i5MCaf7vuLTEPekLWdrhu5NbaifAi4oecNVlZEmekHdYygEAYhdUDyyHcYRfaC7i7r5Zud8UAJ8px/ZEb3dRrApz0gmrJm1C18HPHzQtgx3Vym98QvpQmrLr2+JllW+7M1eeRSpo7nmF/O/8uaD7Y2yIZRxuD/kkgjt/NUFP+X4ZkGzuYjqTu+esLS7BA7nQTs+gCEB7NpIxks6QTeAsfa5TU96cgC4OrbuTP9bQvc1UdFsmAXYJvki4wiGCQ8hDj20qftCUzGovQtim/LlGXCxuvfMi47V39BeoNaQkytE3yE5xzbt0tnMIkaprryhbu0UbVPmFr9wKIQo7QSR7um3TOoOes9H1kQzLSkN371Tv4/V8+rN8Mlk7b0sXOzeKX7B4BUEch/mbwRkd91/4bfkZc/y0D0D1t+SwPuByUSEWbC6ECyOrsZE3PHAeHL1MgyWCcCMJ9mLOMlSSa4gi09Oy6BNEACJruOu8UcaTrrEVDv/N9tmAtCKim4i2fGhD992keKC4WOcwchm/lC6sXwI8Dph/lUajtEtWAiEcdFVLqDp5piUxxUmgsLZMomJ8q1LUHVBqPdAiy2u5QEvn/JCG7W2Q+y6RlsHuiBA+NK0wLfoCxF3NZN+zXBASwapAUSxiyqYArgfFegIRNBSzBpG9rYzxr0H8DttY56XXsfOBZTjrm24+a2j3xR8cjzaGsl0UV0B2fAaRpakiVEDNgPAxdQZjG7MRpbFWCdvsMgDl0dJa6AaCTrLYZtlrMMsn5Ez5M/Rpg3W9vCQilSszip2o+LZPXlT524SG/a6a4bSC8feZXnz9AOcpBctuUIFD5KkrqmxkPDodznV2mQCbGryKEnOdC4O6+eRzf/zWUEj6r06DFX1iKwoD4bDr4qGbGHLe2L5m97deCnRboFjsoOdf5DQ9H5zBVxLFi3iJ28po8SXdvpqLbLBFXnG3ZNECN+V+ZcYiQD0lSe9L8NHkodQlgUy1WuYH9PVlU+U5FLznKYwFepU5aeLjLfdFIVpU0uemEMvV0nfzKRUo6r+VnW9quKR02KA0Afl1esPjF0CgslQ+jT9A0+pVjX4XZLKm8QLMxe2dc67lxWoFJBwT9eUThcP16nUktjja+OfcBC0aqvp5S8Qj1NjtGJSalEMOT37H4eVfT3Vxv090wYelk2215ppo+OADar7UfHx82uWfFBFkOKyqLYXKi+4LHefZv68zFU1hwVom9jeMBTTYjAztFmdbRGM1jwVo6CGwJqplob51bQNOMF40bUKFl8qkyL1Dw/epYixo+4GPxWFF6aSM33IX+IAM0zaZ0c0wKZUBvr21ZbqckYrfxnzoU2dsKOBjE4mK4BlMCszoYgLdabctTJgolJjujLNQLlqIxICD/EQrnvOZrsHhAUpzTajcEv2qMTNeYsHSjdVVeQ6h3kdBVvIiLQI4gEECdvv7i/AFs15LI9ei+86/kO8F8R4fPZizM8txy7eiLckAEn9+Su7PDpQ+7NLL4p/ZnWOwT6eiKa3DrfFUkpVztYPIUGcLngV7y80anoS42wEXb4jMS2aPZfxmZuG9Q+mYiNQdaJLx0z9eHJyaLsbkYS8VZL5O1E1CbYHJjE7dwvEtK9M7PRKOLgvZdVKT5VLbXX4135Vsrp61suwqocsldLJ8ryxTSPlnl96BDvq/kfw127mlX46nm1mAkrEF+Bi7zgZpBJyCys82zRmiEoDU2R5hMpHVwApunAeXHkdzCheEX2O0GjsDeRd5M/KN+vontUB+3qalTM+oIlOtC5lAOsYY9/yK8xhPvaSCgf2nIPLq733l0a2Itp4fO8ADJwUceWGiJV6rdH/4x1EK+c+MrrP5rpBgBNa1WosxDpMmZdHhyf6VFW04WVJyxEgsizaBkYdBx3LxsWeboTNU/eKNdsFMFxI4R8/VNZu6gPkZxX9SF31hgGvgS27nfSRik/5HCLxlZlxOTryqpFH3MKmAgQi4VVRdE42V+fTO85ons8lVTe6qhoiQWjduj6fP5fxeN2TfTMBh78dArXK/i3M8QtryTP+wfShL1f6309BkCihGWxMZ2bX9FyroY0zwQ+wJo40C8HAM47va3+uSUF8PX+098gwK2BHbDkShjRqEZlHUC5Z9qC0mfkXFq4hrABnae4gI0A5yLxeaS58b74BPvETN7jfZvuuhdRiScBEf6XSFMZ2GUjgmt+CNy8JQHBia9BecMaMeq2rA1flYrsc3cfEuUVXlhNMcq+vBzIq30T5qbWdj5t/TZtXiCjUZB2yErdauB0SbhyBJSPYHRWCqYmqUFoO935JVTc5Lp/VVgpAef3IvwlOs+khr3+1sAXYpAYSLwkKKa1zOF9fvyrWHfSjcnQ7qbIy4kDKrGocD/AHUv3k7AXh1pDXOciuSYoTRQhZTC8qnqFGjysxCmrf50x8nf3t5N/2g3JMUTLkrhz61su9bgeXULjhcZBfS59LWTzuU/6RuS0dnqRJ80lLGIpo6oYkhZO+CtMkb1BKfV2KKgq/k6GOhpiG/kE6uwcgQAOkrnZhEhfeqHnMVPCJbt89hMUVavAxSVmRNBGrpbrZQ5BZoaD/+8W0FZ6widUga8ClUynIVFH3JEJEnFwl23Cp+e5Dw1sE8+G4qdwrPe6z/SiOk6lMFJodTWHPMgzOeSg1IF5QveYfPxJEeDZVa/jHE9PkpH8GxruP/6lrqri5GTWfMuT4Tx/obzry5WE9hmXZcpsXKuK2BjgcSLEnRNxbDBGheLphuLMy/mrNbvKn6Bc/+/V+QPnLnfXH9nTZt3YO0T6tyj+NYLnDXLCgPM7u8lznWhgRdWHnzhdjy6i6zZXwklwTNPcMIEcjkCKSAdajFAJw03o5tVtLTRlJlUVAnsr42prAw5aQpjU/a2vzvimHqf484LcTjN4wYRh6ONE7uWcDW/7UsQGTZmlNRLEM3j2xg6Yqy5ld/SfC3DgPtgsBiSwLVhGM4KYsrN6olN/5O7ysv3Qqvd8sNT+ir2UMGsbEHDHPCdVs1E3X3R5Ay/EuGtANrr5T2iv8OkhlQ4DepNXL3plEBEg6hGgD/irmRe/husfDJ3imFfYFPRt9noapahezgwfbSWlJSvHezP+UEYkScSUr/l3EaMghTywiFAOXKkwSChot2lHDLSOQ907kVkjCwf/o5rxPU1kToCM9n+m0T1AnU3heXJkllrlCFYSthPEgj+4KJWTxz+q3PvOObxcu9epwy1NJfPJI8z0Bpef9ym2SQSomILblajX0XFLjLS+CUguoaFdE2El/s8O+9EIkCk2m6MIZIqZxLtYUwBW8Xw593l4xRXjMcpp4dIdSAK5aANf2p2lPx5BuxWmo3h99BcUUMyxaONZLIIUKZ23eXtWJC+PHIbJ40Ka50xouICZ1ThQphAj3TnrGlUM8CIgEU8A1SnYrwWdi09JxUZuK1jG6QrIFZ9xx8QndJ1SsJlZwFRtMaQZAdf78YAyBJV0qv8fpYNmBV8klIv1ZBkWFnNUDBz4DIuE1ucvphW4MfwcM7yefp2pCzOwjtjj7bhDla1UxsqqL+p9i4cFZE0RsiC9F6pbIW1xr0SIWLuPAKSwBXKFKspIzm+L800NbVUnejYQSn1QgaCnIVE2xJJvz47HR9GgcCy8n8rJptBHwMkBKbKw+4dweERZjWo8S+ZQ0EiIE5RPEDdGAu2w7YOr96NRcEeMS3MUbABIpVDX8MJe5mPfWqskoxV3xlHxM8XH2Q8mMmYM56ld2xPXg/jYJrCCjC1wsDmZzhQm95XY3Va5IHs/mTf/WdCf1s15wKDCxR8t8JMWnMDo4f4/QjDpnlH5iiOvNKbb3nasRBY08zcINyhSPFt3YYXrAti1BWZLDR8JdOkzAqvTGwr+dyC34VK8J5SF2So0D7huEN+2/iC3mlIMg8CYeqsVsXgSejAmhXlRAp1YXC4KbXSFB5E3CcYVBuAoWSaON5xXEmU/U0xajY9QK3beEopATsxcJASh6K38KVBHaMjCnkLGMdX3Gh3vAG2sOtNmT0HWvDLRMQmyEfkX2/YPXIRf4dcTDppuvKU6Z6YyPvZsdgRlC+ifXjE2Yt6Is84BjoDWbilI1nepR4DJst0UW9x716p8eDfS/1utg1om3yWbBG5/CS3NCez0+KrRFxa7tjsJq2aRwZGAUcKvbsHYpVu9JF6EcclGWRZen3ShdfmBBH2n1Vvb87yjDXuDYAkmBmj80ci8YzPdgARI4D/3VCtbjsqHVDIW/oHgQZW6cvWnFBMHgHKVSY+dyMMwGBHKgRG2S7ZO4hrWuCey0J6lEtn+WZhtNyUC/vhcv10oM+Bi0tM3r0DWW8Z/a7VLjtCyaIeKDIOliP3APTED8jc4Baoym+dWGPPmzfkzzkBljUFFI1YEawZNCWk4Y7PQeUbuAuWZt8tlKILUv6VDxP4odXGy7nylro0SqcRQXmDJtght5rB32c4VC9EWnZz6Id6Ne2mdY/8hvoYgDyg2shj/oCMM4r1pCuNEKOtlA/qShFSzoBKc/fI+ArwCOe8F8KKvUwrwpF3O3nigQGr46u3Ym4rZilFJ2OeVJHpjlr+lcHOmQZHRtQdAB1fvYTHdkoalve8DSVETMs+3z3bC8Owcpekbllpecgh9R3mpV86/GShTBr7RpTYOikopJzVDYgHYxJzGAVo62cYpTuvJOcbYRY5PmBG0IZI6UrRLzk46BkIfCZ15HAdm/cfq/r8mwhXbEWz/gLPUxqJNA5ZJmnY52JxRm56SRepJsMbDRiV14/zknhuYTp/GXxPq6SpqLwCVQH4A/TAEl3NLVIXbRoQcnRI4jSp06UqNS7wt7bud8EvLP5v5svK3Q/gfY6fBq4P2yDr8k4BwbsD8MeNlFRDiMIFuDA7PwVhWPIQLG4ksadGoBzn96jmWaZNF3k7lUuizXpqK5j7JdUp902tt/2LRIiKPsZygz8dTOXQOwCjixQ1fLiNWHZIPDWYKWcIpVPebZTALtBbf3d2MDrFE80fPDjxP98U8eM1XeDWkY0tiOYfL/HueoEP10FZbIXPRhjzDyPO6jWXsFg6jnRMWziHOE8grRTonylmqh5qp+f4VcWq7qYQqWu/E0XbhMBH5TEUYQ7sK/MyKxDcoVCvzQO8utCHJCgs1KQBR+hW2P2/BBIiWu74fKCJpN/Jykt6xKHpVjRFVLHSvwTS/p5e5dXNSr6wnBZCZmEbVUxrTkFTfOKjQQHlFgTRGBT3nWleIotVvBoS9qyqEYixR94qzqp7/ZFrht143ZE7cdGo6P7yyJj2DGn0zpMqQetJsGwRC2g92RtIrG8L9fhwLraGdVnmfmoSZrlWT2unhHSu33fq0JILMcgMUGWjveAK4FWrr+c34aaIaxPr9x5AR8hoA1Cp0yjNUD85vSCsS/xbBUhbnSYX21tG5S1N9e4tqdFpARoaRPCw5FQI+6odM2bTqCAy3hp2nUUiESp0SUZq5A5Ik1jXAqHh7ZSXCsPECv5leV3mqRifXaZo8CoSymU/1vzYGCmzQoqIzUmZ/Gr1haXxM4/GKtHVGj2U6B3dU9iBeTdSK1KfIHY6dIJhXp+SfCO9jMS93yCK+7CsbBZ5fof9BR4jclyR3uFeg+9OvI66nZzYaEA8hT57A/Bt73obA60upyiJy7j8Wxwa+luhjkbXaL/MZ88tvVJ6/Y9xS1inbsetyS7woKy7PAIZAlAtYhvwPYchnbvZgG6nwyFtDKWocQinPMWg3vzqaa5j66Wn5RszETdFJDbfbuzTIxQ3j17Tg3DuVJdFHNrX0LgpzP58WcE6sToJ1b3Hzqw+TKsFS/UxHBnNIerkBVV2vicFqX2BOomAw5kWzFMbWc7wWsIpg3lUiQw6dwkkCet3pXf7GXbTxA6VYXMq7DjD4nFu8T2M3QyGFwvhKldh88S5MiAbRtlnsDuVxaLFbBciMa4pxR3FGVq6n2qHJeOx29Qp7xg+2f3jLUWb077SG7dzj7IIp+QvUgXoWyaNBc1U503ENw0aZI/oG3Eg0y3zeKGG7J8kX5hKFTzI6ue4z8kM5XeYfsAS/u0SOk776dxqYGT2TJrQuwtFBhfv/83iZhznLePGTN3ugyZy0W/QmgzUJ7HCMixh8XU41euLAELTivzGZWG9ftbHqmamOV2f5FQLgIVSMlJ6zftWuRb99sZFtLLKVddL3bcsAtl9QPQ149MMjpZnF0/wGbv8kCr+nLSmNpD4ThCxA+vUAXcIXjc5rnlqGUAGpKBDZ2TjkqzB3oQ3VL/TY9WwcUCOUEygrq4f6G8t+KHO1w6yxF4BJF6EfO3BVqT36WjniWLMjiR4hNUhfl5yaL4JrDzYKQG9gw1VJuypXvGduPNmtlZxnr8wjXWTKUoxjzDDhL73+Dm5oNq5fETemz1j1ET67fkHku1KpQ1g1byw4ITeoNYN00GnC4pjKLdv5mW+KzQfGb/Ts6n4dK/ushu0CYRbusj3owBekeZZry7R2XzanLIuZxAu3eGCaZXeb1MQigeeq6eq9HUx5/hRi26pY2nMZ3PgaIXZNehEYqrm304/WxfEyqvOJyO1hD4b38E3m6zoEdwVu93Z9ZNfrixF60rsF+KmYz1N0XAfd2qPQ/Gj1zOqst3TY4MhLG+n5JexdZ0iG4DdRsc/Vf82d0gTMuZKRUWcs/wbHJgIGp/h1rfxY5b44E35wXVD75zE2fw5FhJ9kAZ8F+Ma3Eq+hMwyY6FwYPg/NXt0tSdBFPT8Lq+5miZ3yZbQqkSmkQK5mF49BHHYzU0yZ1EWTQbgk9bzQbPNPyvLDUGqVCMkghY5op2HuRhXJ/RsBYTsHQe+GP8FWDk9ZxM06SQWi4x6KboHwcnqG4uBYeHjAKZ7r+x9zpKZ94cjhNC6MwzylWzs4oGF4NM83J0u8OhaGrm8r8Z0m5EJJejF0KS4TrhUWmpz6FdcETyVF/5XVtSFXp072z2tSbR10o7NaSNUsIqk5gqTHNfMZKBtU/SlX8xn4g+XjaRxH00hSbIiI7ejSZ86Y57ZigrUZuMtG7EPeErh65yaC8Y7nAzir2d+WsB4VtQSNrXGEt+LcVIcnM3h8JwFAfsRZuUdUS7u9DcvTzEiOp4qxuVk1cosH7edfDG9lsmjjEhVvzDTUQH4XtPwbFQauJXu4StvfoieKHFiWIleukVEX/ROFAssFtNWj4D8bklTsTmVo56s9bKSWkuiE0NJzrVX7nLBcokX132mjOWfcLBzMGLalUAywxowduTg0x3hFfLdhh3u4e1ujhv/CrkG42zUDTnSSml8vpgOJRdVSwwdrnV1EFS3xIBwObuci+ZJakqcsJvJYAYllgF5sK6NzGcGWotwfiVeHjlQqlJxP74DqzFYKaDmEi+DCKZ4qe2o1QfgepLa3ueZLnwuqJA08ULWdDdkC892UPa5kj+BfgjImQeRAgGgxp9ACyHBHApJJDt63dLXOp35TN89X5CIQ91Mz/41aMRlY7hpQikPEGq5GJA1rMcAV4ZJ/qFwOYOCwGNWz3J5VEED+sAmDEVoyIyi28qaCe9/JvJzUda29ZG7QJJTAT8h2CUMZB0QAhJDk/PCjqZTpAQOyIBlKbTCNo49USQOyR1AYxwqAfn6hYSBJmu7ZySt7DuSeGNQILRlNy0jatU/N1jmUBID2Eyc2fcXbb5xow9HzK64d9wywS9cTn4VQFHdP4dPVmpDXNJironoP/v32B6kBa2etLs2Rph+t3nyhpzi51tl6dFxhLV/I1ufiM2jeOi9z82oRxPlVgGub9Q2KT9xEBpemfWd6bxmH2K2EFycPT/nXPLuwTrhPMzkv2dKaTRNHEXsAdDuxq+Id+EwK/6QYLFenN5VPe2oRRID02K9YuoklgA4eNa+bptsZHtmRnwWLy3+YRAmzFVNvEro6aFsYj3oqCxHqa+lD/0I/TBRlQniXweA1N3G4q8lq/RMA7x2BtbZ84XwmFEOwSMUPtfw0MyPmf7VNihN0AhZy+hNVS52RE7vAgi+GYSlG+HMHK9lFOPLk+N95by+5dCLw6hXdL1cz9hxtYYhDXqK5WYIcX5SSwM7CpBAr+IiIdHCsK50Z94nGUvIzBr+WQRCmtiOkPNEFUDPMOH+89sNkHvdQPMJ2v49kqrJ2sATj4EHqgrOpm568lYno0jpeFxO/ez84EdvWnW1rUQp5DXY1rZYA/Ir1cSytr18Op6pjOieQF7qkqHgT5JdH3CHKN6E5v2pMeFTtc7Wj9H4DLbJya8HSVfsP6Fzpp3y5AIGo9jkfbDtXaY62v4isQt5yT0FYgV0hcGMcM+9Pgw9V9vgcxaMxgutQewYeACHqp8Quog5V1a4tNg/XObAOdHZKMAEnK3HRVMAPF5PNa7b8auqB5YRGNm7qb7AYRx3srobdg6G14CLfi6piBkhtvSW3ZAl/YQIXAnyh7DfcAxPUS93FQ5pPf4CowZifjoCLjPYJmM2+erVLeJo15otwx56SbdTX10EZvoWGsm9jbVedXzl13tNNS0SMsoIweKfr9Azxc6W2YaKOvIjDHspqBtJEI9Z7fbh7BXgiK4fV6Zh01Y8QUesm2LtPyx+uY76jMjh47nmJj0Po5CGXTDe/dpMnw/Q0WdJoIRsf80ax2FVX0wMbyEz2eg7tZ6UjhUxZ4sOFQ3MpnjYq7fJKllJClxZFnq3c/pgWRAZvChjFpDuAI0ddkkc2M1yb4fQ/IBp05rV6k1ruT+LjYDkipsNP3AOyTl2skRi6BYxea9hGhhWszCViShy0Bpagd+xC1+VTjFC5n12I55ss+AmsUJQT2KBcXELquZxXf0Q2k8R8jnkYTgODk9cqHajujFb6MiUFKBbMolaiJbmlzk2STfuoF8GmnwKmCp3KMmon6sCmflfQIu1B0Azk0VRTH3HPUt6VFEtP93VqFIprPm0TIMaJBCsyuvdz3wvgGM5qb5qxnIikYp73IO10UIQvE6Qjtqi+ZNxeWFU/DLg3+++6VCP5muDuX1gD9gUOpip6LLS8leAl2XfGXuoCVBG6WDXG5q6NG7KMJ2U759oNdk+UHUUyE7EHA5ObumY4gVTHmfi04d+7mKLU1pDnG5N3+S/SHHRekcAmUxFdTu8YdXo+doZlUMUtnsZSJSU3VfhzAIll3qM6GVl357ZlwaWEjAtAs1ibAq7wXV82zSSALfVftOe+2/v5PZWSTMwK5MT1UqKmiemYHDrHyxOCL/DxEQJzSMxt15fmt+moxrE7P2jpNd3tkbzWcVvl9wRFtnwHzZAArrE7T378wX7Wg+UiKat0qyaH03XrA/vUVa1g9wbFLWiCqA9gQJhd9eMmbzBp8/xw6SV0oflbwHsmSzIiPsbYRDPvs35wPDLWco5KIC2EKZ9/vTAIok/UwHOhgxpzuEHbQZewwfw0sijoy9VLNQHf3Qu+TnHp3aH9K7GC0wOBJARyGgtM99n/WKalIwYHD/+wiQNxMTivYg3RXz5LlI9jr9uMRD+YtYXHPgvfqrUb19RnaIgaAfht/Pk19hRO9TXYpPV3buYh7JVRkskR7+rKUDa4CJPD/dqnqYowxLl2Y7YVmXU2402/wXk9svCW0f7QVuvI1Dezv2qAC7avl9rFJ+2PlEdUrNAvnJzihgIUvxPeXUwA1ZndJn93wKyFq8d4gIpJofmGHSPlHawRY3ExwQf5nZfQ49bIET3byUQyWv0a33PWTwSjFf5V0khaWqbln2/HOLEs8s7TT5zGQBAw+t0wl2E/Uk1yIlYWTcZHrSPzmpHY9W/Ni7t7RC47SiYb0msTDurIISBHYWFtdEB5x9nK2xBNbBU9fFNdlkebPKJGiDijHCRfkmn8NKz4Z78edLBzuL2TS/1/XyHyOSy2CX9sHmsvrYeflMJzJ/W+62uhIs9kF6IuXZZ17hYwJn0Ep4s1ToYCXHzTt+fLQfY2/JXcL0pdiSDNW50CboYKl44bpwsGx2RBRgAwDMHciX3xHcv8770Pj6sy+9PETepgwWVzWprtE/zkw5nehfKG0GzEFHvH9O6L1+L8dBsuTq/cTogQFNdGihr14mYqs3guYl/8VlVnrnKqpTi4DJyI4XDh2f8YyRP+pH7rv0m23IpMEGyO4NMwcp4daPE4b+9vCxECpkiasFzYfCc/pFBjpOfmQuaFaV2lE/h4djgsPX+3JXi9zuUEzxFYgu+xpZO06x2j0XsC4xqlUOER2wVFbrcNHx2uSELQjs7TNeSyXF5v/n6H4XXSQOhHt6LKP8O+1+7Du3vN+S64HBOq9XSZI/dZYicKP1Pn463AC5VPsK6UduOxp5ZjcruGwubwavG6fV+WOzfzAGXpuDPJc58ZQOp5Dfnl3EzESr+w4+l5m7I+127cwJ0+V42P6IIUX3lnUE/Qy7g1FIqfxjXg8Q67HL8d07M/PrreVgqAVRvZLQO8H97Y1gsolmdf1osXQI+akfyxqBekiEfDg+27wfBC8oKhC4ihxdx4BITEoxWrUw9u9uMaR5WL/URyqzqyg8oDWEM9Q7hQh2YXivMOgRiHToH3v8zzdI71zUmhUj8HE005PHhLe6UE1noPbys8GDa2ArjXCPJLj/6v9jGpQJEb46LoqjvwbpgoD7t0I/bDG3dtdJYG8wbTWm/JaS386uZ83lA2R3xpvZm34kFyImin2P3bmluiw6M6mXq78TBOIekTFiu1cRzybLDy6CutclNmmNpApPxo6GnDSM+mDr7BZuOzVSOiammKZdbfEX5xJ7J69lrwl/B/48ovj7OIrZr6/RK3mf7st8hlfN1nUATFB2hNkIZYmhpfl84Rj3VQb/04t94Mns8F9MnWCrnb5Qq2bMQQjwKewAQZtTZwV/LE2QX6koPw7LYqSodWwzTY223n7zhfUalxWGnn9zAIEH1/k3PsizsIyKxXm+/RoS2YDc/p2XpgFHtOcPh/Br+PTXmpw+hlyqirW9F2P6rs7qPal81L6TVqgHzzdyfmfLTxnBoB8ag8FgS6J8rExX5IMOFUmabhXzoYH/DaA0C4WoQ1IJ6uPnNI7fn1HX6omnp1cMXt2R6LDmHphR2vEwvkzGnFSmYATgLb3fnHyNM+tu+MQjkil3X2Nyt06gVFvw/aOawGdAoj33D2MTbZyPLWWxCqPGrfgGLvpJFbrJAmlOYGWvqs8vgaRVKTqWbjzNGT1F00/t91fXkiA8ZHaTAptmHy4CgTPHlT4+6dfdNE82+I4MDRdEUgaOz3INrsWT6mOnCcIG6wyO31/6Ng3fYA13GRIcygEtVNmU5Hg5CWx4tVg5UC8Mck
`pragma protect end_data_block
`pragma protect digest_block
b1229c9d49b0f10c698aecb3f446f7dd6cf47b38f19dae1c6546ed9792cd969d
`pragma protect end_digest_block
`pragma protect end_protected
