`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
Q+2Rs+6MXoG7NIFsKJ1BvTu2POWpyCZk0f38Ww3C046VK2M8FyygspvK9YBYhEC81nlKkdC35hILUwLJnCs9xkoYxyJZAnJvynaEbSHXXwMyw+npSsn7HktDjmq6uiF+AX19iIBfgA1e5BhaWvW+dL36IT5qFIwugJn7EhSw0WCNjj3f2is2aB2g3Na/2OVVrbuZiy54kEIlnPyRf+7Hy+h6S88gFZLKrRd7un2bTEfspVtGjtO/lcHsyiZUrI9O2Vi+vvwv9FWZc+6ODd2heV5l5fmaxOGmpAUHvFSmdyAw29fp7Gec+FDkHWCh5Zc2GVuI4+csKnUewSEZkuPc20jlPkYLwxw3kEyS9KWzs/UI7mXEHgnGzb/tFlRhHZCOh3bsa6LmbKVQnIO9HMzzrHGvnoF7khJxcdm2vMwpE5zaH78kkoPOTo0qer7VkKXA9uozQ4ZqY7k/9WsFiuAX4buPYeZUtdbe820jlbtONfs24/03n/iQ92gnOthJQqtob6Hv7IFfSZs+7T7boUU/AolvaFbJi+Q898EOmPdWpkLv8YP6DbZnARU/AKjFKUzLvSDOZqVasteY2+uPoWRX5Iq5cLUd3cGtVA4EFRoRopiw0hDpU0Z9Nlu+8/rbbirqTEy2ceO9aPPo5UDI8yebGYhikDYcG3ltJePPzHBBIK0yMQm9Iec+Z4TqbImhCjzTFYpOc+sbnzOo5ggw6HVpLfjGxzQ6eu4UYOaKiPKZ4A4Uht70RmJJ9GYvkAsBnca/AnqszZWPdS15Cz5Q4HvSlT+/oOC19nkhyDZUrOUx6o7JxANJ5UC93HpRKkbGx1hoi+qabV6+JGqmvYBtObz5ZTBAhqXdvvqY6EkzD79z5dqXvVE8QaB4/O5trj5aQyzQp06T7gwZ9VLtSzgqIKdRXXtvnv4hBcyKrAvMm2/trY8LronKN7wLYtCs8Kixb0K3SwS1NY7tRK0UySTRx7mPGJXKSZIKyq8pz+z/KMXIG7SZw8KsLCQbee4uRun9jowbZ9KY361ZNjooJpwtBOIFNjP/Umxs/xpHl6bLnEmy5i/GmNmZle5yJ4hfdNYYTZ0ZKEBHWMU+yKI5DAhYkTRPh9GEZ5XSfuOCB21y6JGk63UtQdEeV+gBVF2+EQ9STPr+wxXS2siBN3PX5UbjYvzKQ38hnxQ5oiLgwbijuPPCihxzTkkmQdvwSCOJQss1pOVDVdv8K3XNKTWrt26mPrWUEjeugEjytoN/PEsZBcVxKR8/669jxILokg4BYCHFWokZSnTcQtGosLjpN1UZLZ/V1kbB/CILpE/Xwvti01AqWMkLq3jZS02xSpd1XiR7bI6P7i5O2Iy8/CaizAYRcMZPbeR8Aa+l5PYZH3sQKPgmLTAoGyeNMhHva6UjpDjU+ngOodm1oRiwFWbZ1nwoYAKqpjfWDIXETwtPduMxk/zhHyVx7195nYC35ewUk16IVALnolxSoMQaUYhTUCFDkm0uj7SS0UDXsSH1eD7kXJbjJ3om1GWNyJzeNZIibHHSPkBVc/0zFIIauZRxB8G0zX6QH/gRbLUuP4aiu20bE9K4KbsQ7xmbRNE5Ymy5h8mSYD5ocNXBIWfX2vc/IEnvUuOd+PlxXklAIrj73mCnjFSDrrCbo3X9HIL44s+/KbuyiUobpJOVLS9TNgKwD8B5UsfOnVIUq6gHSJ0MHHyV2xciPoy738i6+I9Hre7F+cCdv9JAyPmnbFYe1BBEHWoaIMG0VwLF7prw0tHicHHPVDqGl3X/xTlBPbmlkeTfnJPAEXGcFBea8nqZRRPkldlhDx78y7gfM5p/VnJMkDk+sXz7IpycDXvFGtxER2pMjXT55iNFrnqBMcdT7pY/ZKRWQGeA3jCfjKb7ygoGrJz5JQJ1pvG3grtveqDDAYoTKQNhSYQm5iKgYpWTxw5gfQtQ33YtjDPcKmsWGqfp1wr9yAV6/3C2h2ZR1QqDGloaBx6NaFXDkLgWr7E03NrmdiJrdxkUGbUy1iqorEaO+SzxdipOvck0kGSfxPB2jfb7tU6P4yuBh9YPwJNhROEjoXKIzG6QYKxqa911fVoKlq7RyIf4k/4DmFBxFjxeiSQlVLLTOJThAUAjSzaklB0zp6J9eEqbWtyjIGxsv8QP8Z3F22xtVtYbDGk08WnOupYzrV7SL5SrIMzO2S6l5Z1kOKr8K9EBE+WVxbyiPJOl83s02RhofzqKPX3NVLXjFXCS9qMR77AV5ug63a0P8gTs92gQaa4mzpgqvkTHrwP3k+73XqIvwiW2TqFv8PlC0mC2vbktHCqJeaQ33XSnaJ1IwVTQ0kOmF489M+1bjGJaA4Xordcdtvur2Vx6w2LZ6Sn8uHtO8vIA60R310YP/2Phg0qVW1w/RVjyvB3St6YDYm/iO+VaGTzUHJqJfqug/6rb6rWGNB2c3Vgjijx7u/mNWdx1mxjL01fTj7zYU17y+K2avhnZu/BagNVTXpL7jo7IjGPZfUKI438+oHFZiSJvBQwmsFLiJKsVpDZzAkyFuUD/wZZSSQQ0X233pavgsQsTsssf1YWVCMC7Bs8BSXguKwgROheSzplnSpFNBZEz6p8hsNkWkZYX0KJHhqyPIJg+Pu9glNN1ZN5xZaFrbRHxMZ7NtvNv8XYprbZsCsm5mKo7UyQFOS5j7JzAD4My+96mw4FE2j5wsCbeqsAxYKIz1rkfLLhFTLN7t4bwk5Q+anAk7jgXu0qQwBnGTNObxfGHX6peqJyuyFy1keO2mfVZbidLTgpOTMgGEpo4oboLkZbtb2EblUIpTwVuQuUNVN2Ic8Bfz6hDthBi9dEvi/roJWoKAQv1Tu5V0Cfpop7edwANAAH0pLPfDaOdhqCR8pbsf7FRjxJ2y0/ysp5dfwpRmPCMmRcJp/MmKoUcG3gWJR6criJj34OK+5w0MgR+5Qw06mBVge0J/1+GpWP9T0pJe+LAlVVK9ObdBf86+L+UpjmAeYCRpLQaSP3/0xW97oD9W1PrTatRXXh5HHnqvI5/pw2uZIlbhZenWC3JeTzG5wjNgTQDQyvwxGd1sPOz1ENrK4sP9dmbGvWiMzQd0GMPBvVN5AYZ10bn5h2te2C4PNOHEuFeze2LkeLdq6OsURkrA5v9xyylTtYcNbm7CBWmcX5+3wx/AePcsf3MW7f/TBiKtwj5CcP1OYKtAgDwCgrnWGL/dmuD1oDV6rw4wsI2z86TLsHfEyJKlext9pUBbwufj76Zvo4hp6Ic9BIqQxDDP318WAe5yOdQFOHXDgIv02SR4pvBAUrvaR0F/rLnofEDVZhR8tDHOfQjTITovg5uLBf/WwMMGsVZ8dQcUuEaZRGgtGv/qmiG6FBxm65XZDMx74N6ZcZ+IHtjok0iHYVyE8bco3C1ClTIURW80EZrs8Z6lhfh6fziM1xy30awZaLWUVtkrXuy61DjwGhaj82aHXmjXK4KVyw37VB1/qI5tGoTbS5jQAgcj7i3lmhvJh7vNro9hQlMdE6sqcSt5FFOZ98LDblb9Rhu41WeRDsNMQ0URyctUP1ecOxZiBWMOVOKgmiFaRQxKygQGjcqopL2Q+k9sYjep6Bvbrw0v2qQEC40QMyRbebSz+o6Ass7j3L5LJ0NBsyK7DEyDhmBKJDFdgIv7k82O8Pniiax4jcLaLs1X+WhsifDfB85Rlp1ZyBVoPjuChcm60kKLk+34PHqY257zel1QenpRG9toeZbfFkz3i/Qzp1lXbFpplc3faTOKXxlRP2Rt6ehjaDV/jM+1+HDk4pKaC9EN3qIP7E4wW3uzEgHjBC3TolXrA7AtqwyhbN5q33C5nuv7bCv1hrWXh6yTTKeXbgFXVgmD9SrJ/Rj8lQHTA3zT53bPfUS2JWbDKxV6DotrywGuDIsnKS4o1co2qe6Q3zLBkf6VnU7Z/Aiza/ia/JAl06ENa9ezZnEycc7Vd18RIsGC8Pxgps0hD9+VLtbQrp6GZ6fzTIMEaFHNaRAuxmVlcUg3xplrbgzCRw1I9KaT71LpwkNKF1F0O9tbpFwHfxsx67hrXLuU9lhjQxHZSu6suXinWZebh5kNJrYmKtnRr0rY6Cqz68fIsUZHOZM8j5FU7N/uFIfcxPnwgmpp+fdmXi3wOyp1k+ZZ+uIDVAr+mhpLV/JiqxZAA3pvnjZByWJg6HXVYn8VrSkn1qXZf+oeS0j6UMUlZidFsDyt78c/0LpsKr3QPI7y6uXlGHn45Ho6j2w8Yk8Vb+9tYH22mseDN8NNwKxhPYyg/lpPivinUlcQjYeV6Nf0vQW3QOGU9T2q0glw3BECv4bMdK3PSbgOc4Fl2aAk4EiFyx08f5PT1gxbL4yeDogYKujCIRjT/bNxl8gkFiZPowIBI07T4RHyS2a1R5opmQurTgx8JigQPuO1KGfAiNzHhjqjr9kgodx5nMMmbhNlGNbgJ0tEtmAC6Ha3e14/QInrKGvwVlUZJ/2tWVymv3RV1G9iDIgBKIu0fG2I6BXO0EP+gS0CWJM6kN4jNM5CbvMEmtGOzSQhv0AHgxu7MjkOSdmjLP8X5xPnZbZCwoeniESVtdTPHbP2vQUloLIdGaoM8PKzjrVKI0jbKaMrrOfcDixR/foL1G+IlqvOtsk6MDpskducNql1uvxAlmiWswS2QIDpUW4C0Ifg72t5jD3oTF6C72F3DKHqCjj1w2v7zTSUr9EY1VicYJM6MIuK7lAhHElML1W6x2U+tPsXEQLSIpyy7Gph+EmjDHEC2OYxxWmz8e2DiwhM3gAQAOJosqMZakgRypvWnr3yp0zk2c7na+j2XhZzB2JvxoGDzur3vrb74ZX2Yd7DudHaSYpcUPyRrD73VTDSFkJ28tFuBkBwEMTMLQPou5a95VYHAWzolEOGnrKxYrBpkrCiXHda4dIUOW92wMC6DHQP7WLQCDAvKOwoR9zgle59C0Bdo+ml5BFO1ZZHl1AHr4RNkdSyO+RT3C63g9MwxjsF5tM0NX6V9E9jpsahRSyCoyxVjog0z86TkcRN5HnEQofrTe1ZgdHnkeonWMPBJ6n4KRW5ethrlubsjMFf1kSq0Uw2XDbUukc7x3L4wllYxeoTxPL0oLIOYydredpHr5UtFd9JHEKgjMPXlFEnBcb3zG6Nt79ytZSjsmeTcfh9oWRSw80ruhvyAvsd5Ap4k/vRBi/5aErk0wIq2B6i6m7B5L7sIZwR8qfVV50xv/M9+AStYskWyPAEYMPNKpZNrsXeQiki08qStOsSaRe12Ggr7gosdJRWdsBXScAMYj8CeRCQmB7Xg6QkFRfBTMYVZKtjEfiOzkKtB9ZAsNAHwfIOdQMpbFRVkh7nUzDMgHsCMOh7BW5GNxsKSxejW4huZNzXvRYbBRG9lZ+fRUIvoTUfLUtDJHO9dZdd1VW3x9pDKNT+KpChihtnoCxRvp53KgFuLdAQf/6u9KxIGso0NIYru4JwoYDwjQjzBYiodMicptSs81+pYSVhAkD+g/k7VhKs9XtqH+qUxgPHpyGrybuet7PXr4Cev8nmQ+bnY/Ff5tZxNbV3oUbgV18YgTfTPiaLGXrg2hmV/4xxpmLpopXT8Fj5BF225OkYtslZE7BND+IxbJCyMwNO2qdpNWm3V21CrJCWuEx1RoTfbo3V10IK/WdSN2PXZDIS4qpXT8F3sGCbREJgzXUtyk3rsv7GHsXU9F0wq/velGRdXXupqcBiukxmKlAk4653PxMhKvc8k6AYWpXwkoOwsSYFrWPhYcWqHiW43AS9auve7MSBXmKzrSXjO6U6F5EIsJfoZfvla2I9O1tHtHdOkA00JUKaHloNziDtjmDEFq3upfc/45LsBSS1AaSzLDxnfWwYXP9tkpV3DxivcFXdFk6sMSjOVaZEcEgij6WD1sdtpvBXc22e+o0NAI1vpW1j9Rw0NTMAfsGOu6oNsYY0Bp3WWwUEtJs6z6kTTMmSI94jOCc5CAC/67k8Vb+MgbxLBX+p0oiu7xV0YsM6hNqCyMCtkxusQDqPn5JH9mzCCkbQ6EZVOyvRk0OFBXINHvrUPE5cgXqu/W5kjODqAwbz96YlBZtfZaq7XuPj76UmtZve3n1gYQzRl3YiXlG0MKkRH/KH8gD1YWdTiDkj5PXt7DoE2Dnlxu0GAmfVJg4Wv/DJmpsJnqgmPlxmXEYOapiyf+JSxOyo/vbnLcUm1rbAZM7xbj+U5Oo94vp56kYXXxQVOwjHzXPyQ5mj72rDtQUK9f2474QmBRlGDrbcvbSconVMvqE+HRFi9OWGPjgwKmyj7YRYd6BJT1dPWSdrIEjamTvm97biMSBB/GU1xG6kO/1E5XFZOekeX0B3jYt9ra9pDyFz/IxU/5LQSID+AF6OntULPOb9ER0Tljug5cugeZbg0awcWqTtQ1sgVStVdBd75EgbIYSmcsFCMXZYysv7sX583ZI6YZrwhAIxBb2VGCuW9XC/jiyN4+4o3hnRukUI8K+6oSQ52f86AOYRCPmluTAQrOatxvm0xvAEszFiOG86vcBUKRvQbgu2Vpzp489lPMY7dBN8vlVGXPlz1KCJSDp8mrYxd/lYNG9Uw511kmTnFOn+LrcW4xMu/VvaKlhBtOr6wr0D4AuyIBgPakPdBeCi5vE65zRudieULXJkgrainIxtcF/8JdK9G6EAMy1BVvhzbj67n7K5ppbpKM5WwrR+NMbskzyPHQed2pp69VanBtoPirgT+xAquynCOxIke24JL8jUZljD3LZFkdmM214adA3iChOwfoCOUxGmTmQM2LTZMmS//vFbXQaaopZaH9tdeHJRxzTnGTUDHbqxZPJTy+zJ/aBT5sXlE8kAvXadk7sjeG4U4u0hPwmB2MCg/KW4VRbFhjlwqh4C8noWnELEflC+MHDdtxV/KNQygy4zSHllXD0VKLTcrdW2W4xhf8Z8F5qiJFFrSlJ18aAr9oCEl1geGl7ws3B8PGRCq6nl1esS5lNs1mkHbtN+EXtRNYtQSN80099AYjE634pDkR074kSwb9gUYsYTdCAhjQLLCSLGWgqRGyZOPSpTLMYh7OR8ffdlIYRCimuSk8HBsMFS7XhmVH3OQR2fMaNkx9k5ZFKFYGVep/nIkPDJLRzw+jAcF6ryeyZVa2eD73JimpMdEiexHNo6CtLiEo2OnyxM74SWpbbGs+i15JB2kUrX2Yl+cltZSdcL3aYXtHMQZj3T9MiDAPcuf1uNWmbaiiv7kDBR1qdnRP/QDkFTRxrSHiVVsy3mQYhh37jUhAiTBsLq06+t76iH9brIojPJinttIalnsbeSEEHoJJgyUJQv0GXVYlCaCGFmCBxzmZxI+buz9YJcwGdte0kDA/3OTRIXljScH9Abe5Y4m0ajdDxYwqsTRUsBXCPq3dRBeG1BfK0sHMzv7fX8Dwf1JGkRZ6fBDAFDtRFxKPpfbmV/c36nE/W6IeBbQie+qz62W/ai+bw+rNEf9n1QHcNPm5iRtB0KzsyPuoyA3l1VeM+lz1vUSIhWSzzM5wLpYMoaurBPYjD4ro1oJYVd7lGtDOnIvcCJ9pnok/o/e0x05R+4wvQ+mGWItW0aWoQ0EBmYw166st/1Tt0354Ksc7/IVDiEA4ouIkg7gn2WCcqwXX0g0qjjiLr632NSx9T5ErJX4ulIf9BqUKBQU/rBqB/3TUzZCMtG3VqtGWs7mokMvkU/SR9yRxPWxHY7qEFKOZ8GGmYm1vRKAJt5Mz5WSph8oXWf5btcbdJTjjmUu9wc3kH5iK9jHZYhe/MSxHaXWEU7g7zAczGB+CO4bdPdYL+ocZUzmrfg3YJS2h4kMypamzTGdFZLuWzb8dtxJ4czkN98hGDd4Bj3TbF58vFxPV9c4lqDOcSx+qk+srqVHY5Czh+bgSRf8uTk/ivAsV69vBeO3EIYNVeoKa16cPkLAfwya+Y2jyhvwxBBp1g1Fi16iGfpv4TDVsobxs3Lt3Qjtjd51jIkvL1+ugkfMO3eWFmH8/WP52LTgIRY93ekpeZz9INighxImw/umsMbBABJo6ScGdERD2w2MPVBKiWKtKK2vNyK6lF8b7cLMD46qnbS+r3d6NYbiT7K5c8NHqNN662qYcDrprBdFV8MPNWu7DGlGgCqZvhZOinqWBnYFDVIcyfMMvAb0K9V2bZyZIR6IbrbfoybVtajoo8PcH0tbizJRQgsxDDqiKFQ08zu5lA05dRaLu0PTUHhO4JFXde75WwRotuW26VAF7hCdF4eQa8mtBg4HbHzH4RqMgxYkokvvBC/YIO8xCdesb2BQ1tT/WSPjGuzaP0zOQMP0E5ugREExlfy51Ry1euf/E4idF6kYDNBsq1b3rD4bXqHhrJHsUzIywBwPM+xaeqAQoDReuJKdSSM7/q8HbfkvNnA+WDystWPXXu4rgPyzLjObr4P5dt6ahcA56vUDhr6HCyqDckt6teTh5RmVABcQKowW7wPmNGf0RyXBwVC7FRC5LH1+RaONyA1f4Ygo2IgdKz3mE9hhzzI1wARPXmuXWfuQdnZklPtq+LSkOnvgFWRqtjS3u9sP5YY6ea7DKVSVugswk16dIJC5NEyONQu09x45pk318kQ1VhEcIAvlgFXkKlKlTNPRgRK459ggKYqPin0buWLdjrnQK8uW241YZZPV882sAq6OdIHzZehetAtMNUmJQuzOhGtxXWjpqxFnmICw/USyIMwVYNOGEvhFJ0Q0Gkjo73C5q8O/2x04RHTIVgX63my3PrHI/eUlQzrWzCveCTwKIW6d2od4VZ0szSeY5Tomi9LvhkizKWgzvzNk0QEbeQ2ewalytSkqGMZE9/Qs2sjwts2SSCL8MMtsEn9TGqPrcGAZ4zeFXO3JDoQTSYdGW2lHgYBDeXesWzMe4RcrvL213QCLgw21P8uL0Z+nRgF19+g1GDsFWuvJ5v8riHEhwEUnDAgUmUT+42a80grgIfQhPkkP8+b0WoUn1qYzxgHozkLQn4knrSD+JgeXtM8YspMMUM+Dc5b33lI/kJmpOCLabpoeUq1rNJaWyAJmXMl3j+Tw+YxdtBzIJKKs81s+hscuVc8A1jCesz41I2JLXhOQjXidWQrkhNrqqhd7umjVurBnmglNkMXBgDorpeIBe2cR7nv+DLKb+j55lUepcpndnPAO/OyAlb5e53fWPLgeBBj8iAZa1rt4t1EHw0SXYZHnHUh4crC4M/Cy9o3kz3Ff7ZaMtjTGYGwrTCZsJN77kzL9XL9qG8CTx+OceKlxe9Goe5dpWeAKZd1q95W+W5ryufxo7q3tVGWDNdKHbdjaKNw1UYmHKGRMzgOroB8d94cVH/8T5xsz68yWgshiBm8WXykRqEBQgXet8zYQ3odmNQLfUzhVLGhjIbYy/qsXHCSrwcHxmKOOzGcRyejbogOE+eE+wbHAPIKXhaj4wdpYttgx2HtPOA1331Hy2L+sbNm+Bu0Pn0UrbEuOeo/rHjHBK7lCNRpkKMXL7BcLS4U1sAGC9reomth3YLPNGqwP+OpQVrzDoz2phljBIUhJVPwrbX6Da7hxhVGben1U1NF2rucdC2OD+i0xLrXJOs/GAbcUkAKo/xxqKumWcIumpDtfypmGfgYCWy5OAmbXE32JhBHwtGRnxGkl5emrAJK1GoVEx6Sjd5MYB9cQ4fyF9mLB9Qf6qp7yzFLwN5AiOtcSGzswL/6nOg7eN4rSHnaJnkqXonjUOv2V+efFESpH5fECE2u4NXU5aE1/AtGg6jaGXNEZ0KuStOtZA2B5iv9Rivfx9gOIWwYEIJM3TZOcLfKsB+j60NFGn4id4BpIH50FszlZfpUVSJ1MamIsF5iQQ5gfgSRsSYk0w6y3uIz55q/g+MceVR9oy/2X+oQstnjc0XsoFzqbXpwP5cpg8moVZBm7Wpdto5tM3/j5S/Xu9W+ytRkt9ylp7HQdl30GJJIa5FksG1Nq5wJqwMHalAdHG2z4o3TFEIX13SO63VjUK2yrHOAdFsjGcaYyiiim70Gja9j2Fnd3f9ihAlpfhx+2wV75eeHXTWYCyReB2gEdvGLSbTAMK0rCALWDQwVYNJ3UfTXwPvXkaFRDyQIu2yi0Hm9uqeZlbsJKQhrNJlw5sqjAfGqzXFmIkAzZwjk+HA+g5n+IExgGnw41SvlhiLRRlQDurH41bKoLQG0XR2ujizdngnmQauUfObpwElkfDwnjTD7Vh086cV9zkNkr4VVk6AmBIuJvupcY9BQfJ/tK940S6mQerjsf2yV6eCCZRTqI730juaeUA1nFnYc1s2J68crlEwqO9Vjim/XYrCQgcaKHnEwA4c8z1vPXsytkS9s+5KSYr9dgR6OjFrew+sJ7Lh2k5jTupXJ/AHkeEC+yAdEuMSzSpiL+qXtxUCA7v+o9g5S04ECVDC/u2YXvjVvIzcDJJCGuXB1lSg+0nYH5d9/TSsmP8FJ69x/i5ToDoDzGd3qJbUSKmV2sOVgq6cO8m8dkZ2tQo/R3yEzXxt9uROpramMaFRyIW45SKe0Bvow44jAI1LetgkbtTs5WSwIHscPxwD7bRRcLDsLwistQXWenetUysxyumzG1Nj5V50rNTdlPEQ+Vb9ovyGB3lVAAWd5uGSFbrHB1CZgU673iO3PgyEivEdG6bHz2hKDOIGaW7yzjnGlneTsDZP1SAf+q2gP7Lw6wMg9NAePb44E+98zZroQGPAw7FqfczmQHoit4OGP3a02PwuAEC0pmsJWOJXocD1txA1Wtw9RFuzYDHztXPc1+Yixl1n4tm3+372/h7JRBGQMoQpnSKmxUdte0oTQVJbhKEXbQyjfyhXeh6H/AerG13nU9G+wyOHCVNak6ians9bGKoWMFZMLZ4PJHSugLrhFUyhcOGf2X0Ku1teEwr9ZqsgipLn1wQx6t/H3jEpKPcUdmwF6ncLkuQQzqGTmE+Wh4UXgaQ5hdHzdbK+IPuPeF8Ls8B2HwWvcRiusimLoME5LePVUSwJE8kI5qhPx3sShV0+kc9zQC/ri3fJN1SOVM4azG8DJh4hFJvH+A9V5szmrDiuTye9BLwVxEsXlljUH9cBVy2QBmlaW+AiP0D6/0/LNY4QKXpw7uk/PgxNRWwrEs1L85khn2GgBE/29ZxT1MYVOj3lKSlBK47PnZ5ppmHwf0THJjTKuPkMcFmxry1yXC+x/375qnkHrMzW9HP9TeDXA3xbLV6MGcsPLqbD9gjMQoICwCGW4U52/nWBQ57ags9syJYK/yE7sA119nXETq43zP1WK/46+BdvtMIyRkg0AoascqKJVVq+D2kL5VgGJwxFkqdHWaaJhL7OoWmyP4jPX5YOctM2YkLq7Dzr3kbJ2qMMW5VquF+UUJeuTgz1FARpVpxZBaVruHMIHtQ+y7blMOeSfOH2Dct9syotmOdXAv4FqfAVriVoO4f17vJwMWhFbOYwm76dHxn9t9dpCn9nOiA6eaialAG8Cehltt2YcvxF+c60kXUGHPI+ODF9udB4MbCWnZwC8AOSOtBS6IejDpX/q0ffTqb4InYlwZDHtX820aH372qpzRXTITfZJIgAox4tQfZvFwEpbSsDNDAAlJOOy6HlHwSY3CmATOwS4gp6sGvaOh+1L8M1CM667MG4WeMJ2a7fQbp3juns5kTTvRihBBqJ6chbrCE11Q9j4Xk82hpjM2dayoShpDeFeOo6jsKqI2tgTtEuXRktdXhmo9mu2M/Gh29/iI/0BfJoEsogSIyXp+jx/xRYb0IKOiaCLLphiDViWczZ0mYiWgCB1vCm/aKzYq52ot/gXIPwkaQe2cJO4xAlgowetg6UG5npkVvtMCJ0BrFDmSujceLwnnK2tmSOO1FBadqKyA28P6ovgrLBgjiUAQQepNY4pBxwxMMj73ot1YSz9vHax9IAZxTx2JgQNTZFRmeUmzXZLLfqco8UPuXp5CiZpLAwX9O6ebXRgknK50Mkbtob654VcPS1uHujmcZqUsC1OyXmUYSUA50Ae1g29gLqAOvRqfiXG6x2sunz/ejy3aCLTsqRHY22VJS13ng602m5dPoO0as3BOGe1Nr1LNPxuw7siG67zl2K9PsUH/r8a+5sEru0p4b0WkmChZK1twUNJsm2I0PrmYr+WpCCMdK/lH73VzCMe1KsvJo7grywOyhHQg1ti/86A4j2407BA4vop8L0lq9VlIDc69Yi5Oe3jLZJ+8XevkPm0QpkB8P8o+yRyt22nDLFfN94Zx3u8TcW43kpriWvcU8gR397lBc8M5XDOxhORIy/3UYXlGIx8kyEl/6FOQKlB2BHvxyGQSSihj6XDYXR9u/y59f8FWHEcvjcut+/jA0b7W5yf47tcS4rtAhUkSNfQ8tHeIHU0JszSvFqMmjl3eIJzP6C6446yaNpX7SGdn6XBlohIVGPnbig0TOcTVe/s9qxoYn4ZkbLY+lhFoGnene6h9RFV1f1rDYul8M8jpDwidwCYrZtM+bs+q0n4MCaZ+3XDGyhI+kM7WywMhhN6T62WZNf70aBzNLZ34SFy6rGCejKmlTEN3NOY5L35NJ+N+3rQVBkYeF8/DcCLup1E0zsBooQ0xjtPF8pkZIfYX+GgVDmXuy4qDAEuwEGSZZQ0sD6gYGLk3zXgLpP/71VjkFZ870HAYtfJIb5R6dcX28g/ap6B43mD0+v4ypppCY7Q2D9rEyVQcw6+0Io4HDeMR2MrY++1AFpEdZATGiMjOh9uRJGQM5PC78KfgkFqrDAiYVfppQ2SkzkF2cOx0hpkf8a2kx13NymLWgM5QYWqdMhKT38yW2VtoYoX7nOgCyNbohQEKPZ0oB2ivsSR0myHiVEywbrSk4acTOwPNPg+/cU6xtOaGyztmU1umgFpQIPLOMWS+dtoem4+a+AkFY19nYrEp2PPlTputwEcTsupuwVdfjP+Y8NRd5q9cHvmBIgBKPkNBc1eVVUPxM3kGFEez5Qk3UW/idGwwfFNrNHheBqSHc4kFBVp2+MHM7c3TF4jwjcnVTLca+FCDNFkXuQkWxZGExsUBTa18qRzYuGTNB5pPjktAIQsCxIJK3h4vjnRkyGRN/sMz7qifcgUo+J0wt+gnoNeNeumXUWEyKFTzibEntvbc5Nny8WgsGKQUkkIqM/zeS4RjnMO9jW3wJnFx4gehempTkoL1U0k6PYAN3JX6wbx3J4GClSBX2r+oVMAMt4+ESUJFl2q1Vk6CucI5XxbFy+hU9NIHCGhpHZz4bdlcOS/fGZq9EwaYaiF8gpC7hAipc0kT1aTfAVoJWBLObfq3Pm4S/q8JNpa48wKQhYIQnOnJWoxmF1Uci8qBMhQQkRaR8pTKVENFsyiw/bhJDpukNNIa4hhKvQqxpfhY1BdTw6kj51OlW4L5CMvraR+sDv2dM2P/jhw5NJPEp15Ock64XlnJP5D4Dv4VIXg/x7qeEOKIRs3aoChyT03/RYrAjpU6EYtzpljMxt2ebL0B2LXuGeL4RRHPil7SWSRJVC83kc1rM2BG0O6BB3nFwIe9SbNeRS+OG0mhmyjUVF8ZVEEWKh89ZoeINL98iOYhyV0lYAXv4V1l0fQOdMNiQsjnLLbGA/j37B3/qluEddzyesmcXtyv4SO/f27m5z+VRYAqhRP/pdOGHUfY2X4o2f0ul5Nys5l3l7mFDBuypQ6w2F4F0+L1AGaKLPGInKf3ObNtVHkJo/mikJaqw+YbFjs6mctUsy0d/naHa1yl3G+UfrhC1L75Dv8Y8lHL0zWkQpVRDgQH56ECbqA13At6lpO518geBYQQvSBoNVfPVChcuxI6S22T+X7FWlxw4Xvje33SlUEpaDxDPJgdVM9Gjxwmf4l9jRi8o7XcTTd/Sc8dKu1kR1U0yCbrtIckqpDHb7wvqKK9XsFkdcGoGsTuI3oQr4cs9nzuZ9jUh4R65EbowF8+gZkfcapOW9Nb5rD8w6CTMJILVv5D4STkVdDU0w5Yk5OtSgNQU2hMRDZcsUTCjwXgt/FH9sNezEUGHJtzHw3h3RYYjl4QykHS9YlCpLYmDmxnkl/Fm5LqlOSe39q2ca8SbJy6NYadkyEzA3CTMsu5TJx94V0Y13A0pUYoygAKTZndrYhRh2Un9Y4CDa7A4aZ8xM/AFvYy2TCmRGPyk3GvHzFIb6N5Ep4lrHEjX/aVl1pv6Sn+EBrJMm4YjkeEJCDfF0Uks7UmHASXU2t3pIXsT74T5/TwmUpRXqZrERtkl1R0XOBmTLAcpjbx9YCE2cVVLwmO5kREfmtArpHBGjxbsTaBmU1Jt0iJKh9lRKCaqnQ+5tvIgsxHwFOiYNVaB0ytT+csF3AWyknlEWvOsbkn5DyYpFhqzSlwYjGLGRd2YVhUC+cMH5mK6tIfYNBZoy0nwd6exFXVvRYGFt6IutdAHGMSdGZV/9nUnerSSAv5P1PU3lAD9Phf4vbK820rO7lr3bkMQDX91tn9kWg3dywjASedhN3crNYFcFsZrRjhIgLPc4nkvDktdByyRp1rYK7kvZsek0o8ytj2zq2x3SZnNrULnBFh6QXXqEMzhRxJYgyo3g6P+/6MMq9vlu6PRHka4fmqmNGMjW6r0/MT0lpwIRR9WydbiKqiQLBVKj7stwWhSMMCoYpo9nXpeakeG6eZcxufEfLIt+cP1ZubBogGDr/J39kOerlboTkx7oj4D/3apkj7gBqk2rEI8MnAPD8RJILZYB+6deeW0fY+DtMnXmY1AXPAQGvdUw7+hKNJuP85lTfJfj0+ewRnUaSUhQL8M3X052oQDg87uoNH8eLDUrcw22R33c/ZphjycQLM10+o8iNwVv8GJLPyVlJvnIR00PYL2G0nBYDDoggnJIYwOOGUA1PR9IpH+Bjn5lEJ8pZ1I/rhlhuGIvEYJ3130ShuEx9QzmRao8UqZdgoUFRVMLaZAUOiMCdFrx6JR4U6nI/af/o8rBrtrqHnIE6cNbY6yoZqS2uRIVpjVqG3+RvDcLoC1XOJGz8du4MbZOj5DIEmLuyWV95KKDudnhoixz7btvIZzWo4tYJXAuQ35Yo6XceaVb2H9I6RvoOVfNhR2yZFU7hJMtjIh9LqzAUN17C2NZEs1DjMJnJHg3ALNuFRnTfGRqEodi9z2+zfceQ//kwSMCDpXbBa+fl10Vvwb36Z5WBNJeChrzrb/gwxG7eSPNZbeLGNCrPAhMV6hlE+p3Q/Zp7uYQsgMdreUaMFMg4XPTmwCk0roKtePrA94k4UNxF1N7dPb81CNlOpZhDEBSJgrMlINZ7y8BkKxVb4RboTqdP2Wy7PsJvAYdBFUzWwLRPYy2WiuPmTV/m64EF/8SFwN9j8SY5lpGYx9XgloOCbiwIjm0bPC3O2M7Kuvwg/2ReEpVMZPlHODAez3pCD0MZC73NgEbqGbeVfAldeITg2AHIyKdAp0/xaefugHmmCOtcuJZ2G6IN3JYZ1/BFC9VnfZKJ4mNiU5h9tWPAcxk6lXfHrhhwLwt0xaywRluEGIfFELXDFJXlBwHspG+ADEBdBWDFP46qfzVlQ0OLOW3hj6mNQJ/fvlDDoy9tuP62h/O538u08ArfnMfIgMrctbC0CKcVxGwyyDMAQ/JkunHQnR5fTqNbih0o6CycyDbOnfGZjRHxpi1WSXaZwpKuXhq6daKURodnvSV79zVBfG2PzIQRVzuDJcyKljE7yM60Q2n83kA6Pn+HSqqBg+vkOENS4ZCl+k2ooGdhLfHqkPnWKnQvUUeEsImnIf2RH9kY6Z1kgha18g7psrkyt2E03E4WRsYtJ6iDJJMBGBHBwlqDJkRkFJrCbpj6ydV/XbFZvnIOhbzIuD1Y9qzmccugO2tfXYMPmMMkIbcwoeS2IFXbvjgioEiStSOZVSlPiqWzUcGaPlzFdSsI4bt2PxEdZKC59gUZFhPFleZudKnaQBIxMitt1GI4Y2m62M8zD5wHqkyptwUJ9S7xkrCgqRrk5CinBCGqh+v6zo2YiiBGgWGDoCpLjyjH91zfuon05KcrLNEUtsmRtZu64CsYDYYlZgA+16GcT2rxJ8sTonUksVYH4vBY4yqEoDjBhQsLB19Ma1Yqhm3EiClj8maJud26hI5QU8T5CYZkUHTz3mtYnTXCGMGFbBRYqPobuD9JB7bV03bcCrUWdpDLGG1rQL08zBAR/IrM6985W+mXtDtqCBOygCftbPBL0jNCFw9dpYisHPvkD+hrdiJaz/AJue5W6N1bfUzTxwH7bDbos9TaV8lbBj8qEqU+UEU17Q5w5JECyzmIfkiEbDJnxvwjsxtwx1bOM/Tz3/eyN/bA+HhoY0hUHajHcTqtn/z7lLRVsuixNwJZAruaoi0M6YPoaxo8eu6Rsvw77nUOjP5kdcXoQd30DEWp4dFLbafWv8c+Dl0AnFprKpvCrIpJV0SXxHgPN3rqbz9U6OcNGV0cjyLEUcTZ5M2NkJffX0UMMdzitzwhVvIWURV7cM7HQVL4xkmsdLw4d5k1qOCEgAZ8loT2YPn785eTuvClIkvxImqTCIWX1TxIkA8wyQCUQanTLoxGxVDfPwgBggEVidPx2QixYy+BkFMpUN684mOnC80ZKq/2Kwa9mHe/wzFNo/VL5ZRa4tCakr+7y5ELWLr14z1LxAGEe7pyvg6QjKwpPxg4HlRKF5TG1y4q9D4+LUIR9ojyFSUK9TAnj7U9YZWmi+TEkUDXCQDs0Mu/iWfA9m/Z8SpNzqGqbhfBw0+goLoc3cZRdDZ9r+Ac3GcgIKEAF5okKm8pQquVKunwaD/bqEBLP5AwqrJ8h1E7G6MQIsk/HTbhUyEJG+9DbbWYYHTVYxdqMwW9K9BXj/OGjkN6MwRMgDRwoGCNtE0AiJz1AVEpyJNMxhn9vVqdRTabaaGxBNXfT3LF71Qe4HO7w5zOsKP6mfDXYkjPfJOPFKltjIxusSOIBZDdcYZ5kY58iMWog3oGvMPyx3VQb+rD+D5Ib2gbvxFaNf9Hwsdfp6kFHFEkyTOVWSIyTrb1Y3qOrGsdWYWerN+Mrw677RD2W61i9cM1rIa6SYklV27fhxx+LpWdoGl2Axyy1zG/DYsgJrWtd7daTJcl4gJKR3nNenT85G201Io/YufcLaUOgGt2t3086zksb+zO66tCrzSZ2yXcCJwUGEC7AuBUAEZN9DvgxQBuq46i7OIZBopBG0q+wbGDPcXST9h4SQN1OcUsNcSGcYhD32svVhG1pm6gEZ73hbs/MHfGptyRea6M8kGVkUbSbmy4m4u5AjkZDpZlSrHtl5kzjQdF66H9e5YvMwr81EFdyVOUT2y20DKSGEf3CbF7b/fULjsgrUGrzJ/MK/JzGEMlNj+zddGHMZz7XY7Jaa8+AhPc4satghgBTHNK4wF8kzmzU0DCHik0U1/a6mxXw1E2WwuUMmvKbYMGHM64EbYCq0+LAplvOD7cruw/B78G3jyWTuIYAnR0+7uXgxLV3R3v1q4BSgKeedqJVRqfKfinL4wU4hwu926s8JxBqmeEyzBErs1LOvificVRfJSXwobljyBESpm0wgUO9OD0+HaOI3xC1dGI9tqZD9DY9UVruRKK76HmCBiyx7FgKfpb3g0fzOzw15SwJ+cSe3UR1JI4q7wuFzBESELfBNbxQ2SVjLO5APY6OimCODMAyBPWtpBp718iMWr7FMvzb+s4J2h40PitPWBTUI5F68Z+7GhyLoSGZk3F4Gk6N2Uweo7ZZ7q3r8+vACqZynXpIeqcqin+PQ/WjLV0TUtGJfoQx+qlVja5Ud82NDF7toq1FHanG0LhYnA7VTYBwyTobL6eKPwHO8EJQdCNfUof+RZX/nL0CRpnf4o46UcIWgUEp8eaZrCIY2vL2NVxvTRYEgXV4Ska1mOGsYPXKXDOSv8Hhoo6rt2CxdY16HsAUi483E1UPLxjUXTbZx6fvbTIK5OgF0mecanGV64iLcseWKS3WCB09v86cocpUk2NkqhcbclizKzkGSPGW/WbXjlLhzFP9bHPud3hKHpJY7wq4901emaafB/S8k/aT8l9FiwszYwQmvLZQ0WiNE2qVYup4CiZ/f8PCh2xp/YqeiX7th8NxrDGyeKdmgj5Udt6ibDsj7F5rE0gbzq2AOaMz1pbIXkx1aXqUU3GwyZlFW8lRh3Ne/MCZQbjvHR0QKAdeHcisVzScaOsKH8BtSYCXWOt1zsvHUeijUn3XuMcAY5zNGDBd6eyxwz0QUXV9DLGX8npY3h3D1t2LGwHs1qcE+kDNsLjgo9a/aJMa+Y54PB7NMWeQxK3CQxc+Um2MjVSp+h7PAv9VPzsj3OUtWpGGaaS4n+xNrynlY4HmD6NZX3UiHP8IB9gleOpSp8gZk5WZqlQZwN8nUEI5liz/nc2uz77l8WAqcSg+Etp5m5/mPnDqcZzznL6s4yka3XPt5nHpUFoSSAcb94IoBjJm3ERyZZLzUWhzegWOJlvmC9H2XtyVhIK7wr2pCOFzDHaPWgDrR1vlj/rwIB+pzhf9f25PmkEMSuAR/ZDtjbQzH5xQsWBmKGI25HChfonyaR5DxTcLnrMoTod6tmIV9r8/C3vIcH4LmD08tEzdaeQrJGehGQMAE7reFiSuwLPrdXRoqm5UvFUK+VIGz68jWm45BdJC+Ab6Pe8A1Ld8c6wizDen89ZeSuDmUymS46xJIzGZxT7V73PwwdPHRs0drJOkLo14ek1YKJnYVT6E+0pF3F4DLR0lhVzE+KglXszxJ8WPKCFhhdnpc7JUyPJAZsMdxOo4jzl4xm9J4Iv1heZx8fFjQywvRCmH85YYuwF/ztQIgd3yAyMIAoGPF6cZV1QUA7sKmQzmLpeJsLhRNc4amgjeuQuHHFiUyzlqU/HGGanx0IyWh5UPkWAg4cTyhg3QpJ1UfiPgPBnDuxFlIDsnDMtqPAEfF7niRuaDNec6jMjWVlOvS6D/53qkrchkcG6Z9i45zSGUX3nFK30eZ9rZMJ0HIOLQZ94mQugBk6GDEIKhf5V2Y/3fBtUpR8L7chttEemZ6jcNiU/lh8S1MMlaIQNSo3+Gd5fQg4lNKScJRdh05NyUSnl9WX7j4EIsR7cpCu8putAiz4kIL+SDHAaAUDHL9C7P7oyruOMDK94b7nC54XxSZucNtqIbtjIzuXEkvtK65SjB6zGKHYhYHgawUOO8sjgqD7Bpudq21PXn+g3k5uKA8NWefw03ZPVFCluXHv3yIHi4JjbxF59CAV0uWZyUYuRBFYaRrNM5gxfO1/Mvm6cV1d38GrGPnHDcIqsaSYv19xhABfR/luUicRCWby4Bz2/qIh2p56n49D5iDz4kbP0cZGHo8uiruZ3kBiCT7h61tTjTVFxUiEyLB/GVONciFF3MizcHXxO2PMg0G+AkjzUuk/LzjvRB4iWcBPfVLthw3nnRkuKOXZiWcl29e/YE5tgVVFAqhHpVQmL0yBHyDptRs4tI6FowcIE/+j5UX5YhRW0PJnmiEdT2DEZUeaK8rYNIbIaO6jrHhFx8wW2mB6sq39sqU8PyMv32VODvpBCfF+JgOCShQE78wXdTfr14buhyGxitxPdTg45johodHjLHfPTnfRInA4S46tS7BP4UWDgDM+GwnTNOzVAHHbNiyqGjKeCUSXMduMqZAjriEyZwT/iCS9Br+35QHIBtRXFuuKxYeTV9aKFPp//drNW3E8HEJxVW5XnZvV9mMlxby5n2lZC41OL3YY1edMGnCFR0HAhYtyusO0KBhVPHAdJALMfpyWGf92kt2IY7aDgkz4ICODaYpUaLilWEozaUUFfi2i4APTfGabOb3jpsi0ieQfIlTSKxD4Xu5BLrJ8seVgHaAMSrtsmSnitGviB6V+dN5pTfFNeEXyK1pIBIuJYmGE5bTs69egtalsCuqeWxDt7r/1rU2sLAyh76dWeVLZa/oCkKbn5MRoHXtuTRCyikWTgDehq7PHTXMhWifbs0HnP8prOEhgGb/V1nRNqxyK3cc0N7YauRO3b79WRtF8rlsgpSEufxR4JbYfSaJGd5GY4YoqcY3HVPMA+E+1Jw5vMpMQqqNcjwiEWtEgPy1iLqm/Xz+YtGSD13sxbC3o68wSXFllQQy/SOKDwDtAq9rYK5e/5jGrHBeb7uTwXaOcOWIuFtLLmbefbZMN7/Iqw6wDgH18QWE8Z6Ch0w0R9T9SeqrB+tV3aWOESZZg1tTWEa/qgzS9EHgfFjTeLwdd6onQiyoOridAalGVwreXcJdQTSk1gaV3iaA5hB0UteebiMe8tCSlWmhogsEWxfnTD+KozdU+sNyqAzB9w2WNeOFrL/JLpgvM8J9VASBeLCpWzfqOdYWSEBTA+lPJk0bCtHNQwaMiuP3RSknIlVyi+R9OyvLuWqq+1sH6XQBEjWlw+Zhqk98vKH1PBaEnyIuHcgAC94kNgAodvJYHaRLh/5GO9iG836JEXN9/2ZtVl8FyM7Pf695dM2D45w+M/YbcS7XTbTzn7/tApG62Q/6ctI55iAGbRfgDRSeG/yE77MRqs/Obs0qqrQqhkJPqTSv1XHrpQus9N4lz50dkFQy2mbcIsG4v9pOvr9ga7hu+qqqqAok0y/PJc/YNw87KCecZGeo7ZsfjPD/vESpgk/OffDhl/+1qMDTSiFQJkG2xDyBXXQU7px+1RoeMkRtfLZlaRk0GZ42P2augb8kQZj8SCpncPGwB8sx10yxx1V2Jk2qVYvPLilEXBdD3noBWK2AoeID3VKW5oPut5Sq0OmbI8CaNeXGKe9L9LSqfpDUMRDqfYhYpmY4e7yzjQz9jpmuSG1CCOsspM0fASrrHn+L0nvFkoKTjLTYVasEjzrOQe84RfvSAeRnfdaozpRYwC0QhXvoAfmYH+EhijH193bMADW84MJAfim3D2989RxWjZnJ3BiLQ4c0YtIiIawERk++fRGtCU4WNCRg7ghvJISYCrcCeCwmkZDOyLqNwxzeYP9FFesHrG1mgXTqKQf+BSqHiIFR38zU2tIpNIwhoUgEQjDYoR7ro3GRBTN4SFXRwm5A8QVNbQ4qPhALv+Jthoel/6VyPV0sGYKKrNsp1djjWiBjYA7UsMtTYigL2T3i/SqjeUcE/N8Xho1vzq0SyVSRIWvD/lqhLeIOckQ4cvUrTJ3mRimL2f3ACk8tejINdZ+7VD8kD4yJL88blg4JyXDc4dKePIirKCrKFPClXsVUOcdSgYP50nlpg76iclKA/ORM4XKGFE+GrllaaY46EFSNd/vY0LiDzTWFhYcpztnw9WreV7qNlCEPY44FmcQ2XwOtFdh378TUe9ORyabqrhMD9Djax09pEER8t01qqhGaKFFImTo+1jC5bSHZb6AD0eIif9yKxCo6eb4QTT72nERM3WfKTlU1Qe7DflQlV4XOFS04ahvBPIuoPQTIX/AiTu8G/0TbBWQWImG0ZJhFVenzhlHojVCiFE+Glf/ZB+sqhoKxLGHQHnTr5J1xAI3UsLWKApZCCxLd5gWyzb8aMyNMRpnsMYp1AUYSzQLVtqMO8stzVztcI7QppePbEQpxga0qfNbDSdtxBwAe7PX2meOnwdu+/z0Oq6TpQty3ps75i+qW1iZZ4TLAe531xUlFtTjqkUJPnWyn+JD9vib2sNVo8PjsDor2KyP8bVgTFOqaXyMsGIKrADukq8vENzauknBc+Y8n5BWya4XWyAC+iGpKrJ55XjY+2Cwh9XWSmDVPDn4pnWVgnPW6+cW4NBW78wXZVu7RJCOh/wm1a3TTPY2OkLb0k0f7bAdiMlnbjRBsrBDzNqQ8U1KEitHq99vwvxZPpB+BK9wJUtipX4JS4UWk5fCWhNNkDDo9/JWb1+6BhNpcCpXE8HxY2ryAn4Y1xKJIyJLPHLCAUsFS35FNgW77yDdlNkJdAS+0SXq7zjYKuQVrQJPuw9EE4AMxTfpeSIhGbKZcFvlP4uUD+r6s4vt+uWE+xrixFikef4bhimYByFjyLG5ZBI9NsX0Y1B1EoX2izAD+fUasZvb5EOOhI65TY7PVLPIDRyiMSxqi+uUryyIhzT5hsowEO0MNp0n1YcWa4y1i5iXx6UmAJMNTdiSPc81kVXVTbixIeLXby3bfYnH18L3pMfuDlsDuSmP0bmQ48OBOqr3whwTA4N0f+Daz/y6Wgp8VfHAw9wKb+ZYoPB8UVoo8Qz0+qVex7XyJYY3DjRlaSibPMHv7Amg798NuRruGKo+5DuOP8n1zNjHp5t9eYVFHuFFN8JcmaHBcapW6aVLpeKC2w6jYQ9KPSfnSyGEk2lKAs5xowwGT2/ItHvNoEHw8+7n14RpN7AwcAj2NMlfevQeGku4QypO53KiXcof/D7GqDuJ1/UMvciloXB8PkuROtWy8GwbQ1aHCGtWtt+60P+lTnrtWOYNvvI23LOHULGpusaNxTLMvA2AIvEaIr0rbPirwY9gODhcD6FKOsu3EPSIIWsZ5U9T+pp/zrZrWlPsnip3yxscncTECMmzvonw43+B8Bddlwo0Lq5Vr+B0ocpuMTGHqGX+NrieSuDFiA3LqT+ai0aNosB9FvToYD7bTkiQhjyIAthM+z0bNdbF/m6yqBSO1K6bWGq62adK8JHHfJm+0BnQ0f+uLwhQMUz35O/JqWOV3sMqyrYpLgYmq/pixdVm7cVxAgBDLik7UHjpTxO6nJRKnzX73XIruzFwLvRt21RXFltCjOnmFUqOTGWF/K6repbcsF8zexobagPshxjphr1PWkV/jBpNW9qN65XAG4rwG6wwDgfdAYb4zNnJuQzzcYg30FHQ1S/wZjRuNVfQhgQDTAWWUI9unvg2UiDbmSVhIV9+uhAYorIMVG2FIVApjDtVjXxSHoybpp7zDcTt2uLutWfrc1INAczkrFf9YkOL/AhcJ9NKBusiXtqnyPXNG42ImWKqdmJUGgpV600dtiTbhRu1i9HFtn9qtFqF4qgQCMvVCvw/iNPdG31QAwbyE6k5kHM2JV2HIzsiPhTuvUUKbORi7lO5jJOGV6RG5ZwQIxNUBQQ3QaJ+NuHdeHAmRWgB3weBSA+jT0MraaqD0WtE6GNPsKtvkkkqXqvFnvZVVPbJJCzOhBpKdlUdCoOTUKUXpFyrlva1aHQufQyYTSDA5gezwYKARVrVovKFzC/4FoYbFpL9eE7pZ8whpGZnzQwzkTF0n/5moYBcZHcTnrD9aUmSjcMskBgK0K1jEtqeCRWp5ddjVulnmXI77QGpi5ObJJQhfxVO4oj787Hxq8N5WbVV7kiUStph++njdLbfrf8bZLBRsFxJpTkXe/T1sDcMTsENpQ2xtvCCHrjSMlEjI6Uh8fduzkD9MnrWt9j7cq+Nu6+B4LgKA2U0KHzYWIjn+Nz9Y63HjJGXhfOEoc4M/YEWji0MZW5vu4A8ycJ84wBqFKGNxLD3q6a7cuS8b//8Tq44oB9p4zqnE89JcOxUwzWFpcEYvY0B22bOH4YjIyeYhoErJ265RA4kvH4bj0oZdKhz4MR2+lsDBe9/mMqp2PCGiFQU69TcJwSXhSlv075lDU7FhZCKIa5omHAZAKyHQ5TKq0o3ekDcS2h4G6Pt9eyTS+jm/QczT4v1+bfUC0zUGaJRPAKddir0sO1sVU4kZEiFKQa2JAfuaIZaIGzRE/21fVwEr8ivAFJgPICOxpKvxTLx6ttGL0ZEGtm376MnXjxd0dcNpUiDIEb3BWxSvRtMrTdY/3pqCOf0YGTsQ68VtgE69hIbtkPecYLL62mJwshXt+8CmUqnulA7W4ha4wg+PFdNMjFyOuwit+qxgM9w5jIjeXjmN4X8YKNaWM1At1MjyF7KT3+w6oc02YeHkyARjg0N/P28+ewPhfOozQwUM9sakKo8u/BSivpu10LLGijjcKRbo95GIAHXdT6ED79EOBIJ6GHhR0U2vG23tkuVZPJ7gKpGBglE+X6cJCtpKTmNfzyWmpuXAK6S9XwDMz1ZT22CguFrWKJPs5ApHgm741dAIGksfTlu5XJDNQkLYyYjJxLnLXvH7iaufedEU4fQJ6K48lLtrl619NE2uElx/mXfiQFKSnGOUmHPnvDaopQPNQ+UU3c6i6g4iBWcXcPoEhEFX8tFDIZhBQCYViBXfZDLGjm8OCk1ZZxmoRMY1n+dqGph1bwVRIv5A3LSlwnQth//+n08NczGkHooDPOSSdOnvWAJh0z0J2iHoAFmhMe0yfanAomO2SAnDOB4o0IefXDJKCWJODQHwnyfq1JNodFerFl3sxmMYQnf9bJf/3CGfzk8F6EsccTaJ1VqJlA53PY+vDn1oVthqq9KJoF2kZ/wIzHbGDoPm0W28oLEUuyuhC1E3nMTjJW4Sb9U1lbi1927lOs/Clhb23lZHYdWdvYrpmaa2+upOLsoJXtTR8+t0uK+TjuyorgD2x+/DfI7m2MjxAJ93TMT3u5doI/O5iTB+WCSVbmRuymel1205um0zWJlFHbZQgGaf0RKhOdYrj4hTMtr0kY0h+fTVlH7Q12gP/MblF06OYDPy2Pl2412/6MxBf6imGURIa8i1o2GxBBWlRr3PV/+wkn5e3FWG/zTCbqLkul+AohAsd7+233jCYaQiRdNeIIDl7rYyBCp4jV8aB9MH0724/0/GgtHpNYfETFdP6z6F4bdpOj5fLiouNAjSXC+byJ4Ln4ora1panGSY1X5jit0ON9AYUuS9P6im2R6CJfgkfce8rqAltrfpbCVS8zIxZsu/h+8BiVwWiQ/W2t1pjW50M9Sxl/sZ92rUUGH0rjXzIbjwK0ueJXLrmYFcID06R5yytz2bnyUpVJFn/MMMwlK2RbTFVbUuG76Szc42L1Aa1InkUyZq60XqmH/nHHHzmgn0ajK3qvZU4EXdW/FgB1p2UJLKzgsYapAeVSjcbXjYtkbnNTC/NkOYb3BtpgwaCzvtveaMBs9QFtwkUqsN7YEiS1s8rBNTO5R88aC/BndVdQgDVn+hdRXPktnmRCV7jdS4LQ4qdipBKHb3ANtFCfeOPB9xXa+kJZiFujGhueTfBOsn/RKu9Nl6vnKUPrmFdjnXMzgC0TKojEuDjTMFDwm4xCMxf/3OjawkUyPmH9xc8174CQ0Ix6/KIUDeYnvdTEdrJzMdJqaGhazDdF/Gp8/pGLYtoeQddGqfG1BSrmBohfCoiQs/lp3DgBRMtENYS9qqLi95l6FV3azoX96YuUcpKr67628ZCmls2L78BDuakFH8j7Z96VsLz/TGzTiEpOS52BTfKBOIPWZtMFTHxpmMXk8ZyZJ2bITCJxj5lZ6yu3MaUUvDN5JAUcqr3C/D8HA7g4fT/Z2c6Iqa6dc5maVlzroPc75dhvCo39xiaL87PkI+ZVc1oQfOEzKBr6a4lld+FM3a/n/l+9l3glpBmPxZb8CEquJZNaL6K8zF0WEgIqS82v736XAPC1zaqScE5Qi3lLKHWc5OxpWvxW+5l9KPRXqxViDXjICSDhMLStznH+ZqnvVqvLHCQGaSnEoc1trh+oF/34c4XXUgikS5eVzyDrBsBY8qEjc6C1d1fLqoTf2f67I9oLhBkclfpLK/PG3JEk/TzSzCBUD3T3fchzbxNjY/cpggNyJJYe+hZLXHEq+gkSnoMVIBnWOdn6Gpt57IUiPH4uT9vSzB2shqk/k6XxaV8vKYUW3rHo1jrkAy8B95h1GDLQAKlZu+7RWNM+d0zFfyhh4xI2N8sU4moJiR1fXyjis3aNKWJgRd5/Wa7gadSuBU37avyH8CcHJlH0sEL34xxlMvxLA30VhAtAUfLzxizJm8GlPwxyEM67purF09/MevzYXTE2CE+WKpnmNUDguWUerRYD2OnZuR82dYqN6nj1pc3gO440eQQaWlUnUrj82bhDQ/4H1bCkcyPWZ2MBsCROPeGtLWSqEZqme7vjenNC/s/ZC4UKYsG5xlXhEgRuBYyCpHGr61s9zOIL7pHm4MlzM/lduFxoEq5Y/QQr6uBqPTOVZrWtun/B2gt4OcmKimmo3GajL+df9jCOGiIDpp1Ba1nlYMV32QV0q7RgjRkVDQtYegTfAdAJZAUM3dQmzcf04XbafQbzzm6bQ9d+DBFBKVIpVK1CvB2xjEEF4864wDHIKVgLXtCmwmpIjQKpb/STM+uPcaaiavWxaOcat9wsfcnWAykgqMn6LaGfioHBUOjY+2v9Tf2ijhmOKC9Ck0o/lMDPZ9IBUhvGai2XVxrNSkFD4gJ+TxTP40OdhhWFJjrTCLpA55w5pF7/CmVmfW43DPQVqmpM9nCWHRARkGAldY/2oqhtu6PPWwQx7FrRMXQxf+AUIpcywJSXHJle7BuJVQ1nStHy7aN0dfRXyLjX/H9r38mrcdeytafALxz5yqTfn/CbCSy7FTwfqF7eGASHbY+WCo7PUPCdJtS8D2oSQq1DIQv7daLWxR2pEBgUmA2wktPfudQ0V3q/DJuLGGcMW1ElufmoLZ9ZrgiFP1K3NCYK9UcznVksZEA01JpKaQ1R4VTaGMMEF6UjbpwrQcJB9DckLWoqE5PEvvSu5404fJuj4cZk3a86uHKBB2P6/f1LtWqAtix61IwpNWVVLEreML9MfCLwgxA5PdN2BtOi6CqRIp+/roVljndyVH/hLzzeONpvvYlYTZDSRbtDCpKTaEIpjEE/QLtIoAHNkMQKJd6sx1TrRiV6cJaM75XyuP90bGzum521KcwTD8tBrgPxCuxLibblF0vYzhx+9fA8C+qKsZLntjsKEYom4GqSk90HkTb2TbkryNp8hCpRDheuLo71gAIjV0eDFWNMZzI5sJB4AbCVccxnnbrbtk5ZX8FBkKENgGdAOd6MTmVgOoNtR+8OeVtIDD2pfDcnbkLvrjUkEBgu8xSIPt3SFFn1dnQitsQH/Trw7JtSyXGrV5mRDMtJOPeVWN2jk85hs3SuCJ9sX7kJjMfjy+5AOv+iXFw4OYj814aYLGg9bPsWhabiR4TfMKfO+CuSKPG+EHWFywPPiNEWYWBA53tMKZ8qXv0GlFpVA+VbuEONJQ16C0TUlRQ9hNrExm+a4bZTUOGdE3IXBjd3x807kwobnmjLuAJrTpB9NeZxsBC23iok6IbNSKtMpp05dB8vGtAIjP9dgnSCGn0xustuK8kQHuo8r7y8NRZ5aLxrqjf8StrR9j41zuyl8dQfHt87qCY5dUtUnvMOrz5QSxpE/WA0yxQoNX7nm9PQ6mydK7XZ2OAsl0R0yhoEv4PfhsySZMdiWdIKDhjwescfbaVI0HOyC1SFlOqr4mVriuzMOmkAICIh9GoJ20Bh7vDIuIw1GdWMc9SUPfUiSHuVbPlzoriCnF/1OvsmiXApmy+8etzTj98PVSfY7NpY/n993r8U96sDplu6t/bCT7oMkeE84Bx5Vk5sy/itE8A4yHUFJA7nF3v6UT450Vlh/Npfe4OHHaasGzJoYh9TykL3u7tZK27W60FWVfdwpExbsrVQYcvIK6ZeKelfXbe+gQSp3HW/R9PnRSBSwCyDilFIZLE1ZZ628U8HYtdzBqw2IWWacKB+NSgAy3lt/mimlppidjUKSL3ag/zxeqE4CQ8X/S0ByB8IuTUl/y6uZvtup742QJdDsBagb+T3h4aStuw3qx9SXEJkySOuw2Vxewlniw1XgLUuMqs6hsJWqIKrd4bk889JGf3LxTaJjteMdVtVDMN2sbhXzIvjInWMTCdmOQWtobpdGnLQ3VY0WQ4OiVsbBuAUQYweucU7CyrbRxkFM4ofOm01Ufzu+5YzuhT9+e/T0XYMNosPjXseTAG7BjFUtt5U7Y3uDZZnndJPG8DDEj0r9/uS8HWDMkEx2Kylg/qIEa4GHtocENuzP5PgUbqaPWZpKbT0zc4vJLvM9TV8zHfb5p0CJrUBatQDncbx4Cxn4y5rKpp8c9tG7pX+w0w3zONfhBSrp42D28wJHBqaFHDIvEMouJPShNiyanitPohl0CZa/2OokPIf4hw3uPRXnLxM6jrlcGeaXYDXaNkX9AvoZOCgUHsg/JZ/c8nbjzY3AedlJ2fr5pZmm/IO1TLPLW8Ecq0mTEheyR858IX+bK1Kw7z5ZPyO1j/T7doe0LXv4ryubziPWh6ZZGYf/MWHcpsUKJVrPyjWsj/JFf9qK75g2t7WpgU/JTUQHV8XMxrzpxdYwTAzvOihZzBqaC+IraUhtvIGYbgedo4xqnwMK5jSvC+HIlkzJ38zvQlf4StGrtWLGBNwfiXPk46prGbuiA2jSGT3ZQEmW9Eug6Wa9yA1/6L64yoP1PAKIWRXYWglNA3/yxnIzWn6BLe2p7pmLpl3XcFtxxUR0+DNB7sNA/3iPrJOL7QztsF9Br6iHWAdk748XdLYmi2xz+i6CSJ3/cBLuhhI/gJVbTcsyijPRSCjSqOuIjyQgZIkNuinbeFByyESbv71vOgT66uAmLltEnjZ03FUXDP+JM/wVygVpsQnW+buJ2gk8nMVqDGaP9xf3CEZ82JNHSCi8ME88PmErKEqY25Pxnjiqb3deldotMkmXD88cgyUsOvNVJVixb/wKKhWYXcCVVIoD6zMvdG/rmQ/PpQxN473PahvkPEnZG8YOLZoWhF0p7haYi20x6H4zhA6B/xFCp4Qzf1Z5mxEA+N9Om3NPpiBohdt1IriIZsc24e370aqvya16Txd55GbDijRIoN6Gbo7aRyZi4Qfxx8bOoHNfwuTSkmVAiIn2IvuGVAebme1dMGsQiy/hE/L9lse1FYKS1lJSBVHf6UC8VFIBPBSGmkNRoG7OQGJn6MRkD1hV9i+tgVaovc7WM5W5Zp7Z+nezUSPK5kMGPqEMKpJfKGCbnFsHRJOS4DyfpMXXterXAZwQ1qw0NT3msPyn/4bI7NZ6AGKIpwxOp5cPgHYkcKvQmlczDS+XcfUsXFfZSyd4RB2sPRtVjMsgHYHBtxPWV0aTHRMR6szjL5Vjv3pqyOfgzUDpEZ5NTyz/gpUfNg5ptqqbgZuGAfu79jlGFtIl4nWmmnudWbk/RI8BVUYqeUGq5ZN/BYnERB8dWyXhd7o1Rm3XPfGZ1h5bixUTFzXkDY7EkBKuDc4DmH+sF2Npez0j9Vcu7B5uCgSaFZDvjhBBjoe1gRuxjWieEGboDaty2HTkWcTOe0O5ytd5PbBVBxyvV2wry7IFhoB9cPjX8gWLOwPnQ0AaDwv4+UVz/bngr8W9PGgFT0aZqmn7vkunbeb5q4+6rsfMpO6c7qQ3AKmiwG1U/pNqRpHmu1h6SV43/rL+PueqDNemTkq2WqKADIcIc2CQIWJqTb57sFwaBtQEYdB5vRt4GsRFeVl4DckjIZpCJIJvEbGwjh3Wq8hs3CmTZvaxMCQFPa8doOVzgN+yEOB0qErveC29z1xWv8RH3E8ZqEhAFFztjRrt6PZcB10uMTQQCSoGbO7PB0xvZpYly3V6whHZwjKrcsnOclaPj8O6hlf5r6OQFfMCqk+udw5bBTwlOC6EwRQUf2Y3vzdATd83gXG81HVlhX9aCaN28ap+UuBEa1fXZt7c2zirp1Q5105OOXFqEhyjiK/R1kEcUDeWXkvBjPFyNF0BYnN7eCfFU3cv84iBA0NWBa3PLF5sJHRkFYZn8K0d5G5i48lPEkvr83CB/8FET0N4t44L7f9VobDrO1ZyLlquNlv22yhoq+8e2ywEsIrzOuAeiiLsrci25SRCz6Y5a4NYCz4u7nJ+480pvQTMO5VFNNm9wPE/lWYaeGA5MJ0Eo53DP5Trs20K3u05kKBJTVGDm8Mupj8pJHaQv5S4m6jArpZPFbnArIT5E3Wwrn9KJHz8Y16CqMaVlthp7Muf0jkRphSTYJPzGVrNswcxxNBup35c4W0YZkEgw7cyww5AvnDgRYT6t10Ljjj6Yl2tFdL4pA+edCwXyQcPghh7vzT43GpCkiTzileE9e0r2uBFqqLZrd7qmgxDNCbzUpyoFyW248xTUF3caOlTpSkccsDKLwJpbD4ndt/e560p9UG4rDAvOwIhn9cL2k+yD4zb69RdUtA2P6mJKj6fCkvu7dB1oZdSZWp04LgjfoyqKZCOEg0A5basqWmAUQKJy/w9Hyj1nRnEwR4pWACz/J/8wNLN6OjHlXWTpTGf2j4wfISrnwUJQ0WpcDLnTFj7fI300UEeY9pf4LK+E/n89PYGPs5ReP5bmCDgqjejmAZ4cmzWDc19gzEawQp21Yw1JIuYvkpLbQGz/eOXO5crHKxocC+GA88u1ibLqCMxKpVLQGehg+srlSQ8RPy3vBB3ZYDzPV0zJXHOFc8j19NpUpYVlbsIrfoHtGgYsu+hvRDiNAZz+vfaD7p7IsHmP6D9EbHVJCK5b8FauIG44YTZOUjH3qgJ4P9u9vimwU8ng5PF1DITJOe7DgU6t0KTOTcGmfZ8zDdemxWYDf8VWUNdsIRA0tTzcBe/UkQxEDjqnh+pYfUR+Gg1jUXXzLAf3uUyPj0iA+uTcEVIQoWhjLRV+tLfoIo8RX8roC57ME4yi4abf4wPXwQiCc9gifka6J9desqgdRYIMdVJu3HG+icSYL8X2x6FYyq70g1EgeBnC04kS9vqwy5PuskkfKj1geu14yXrl0BohEGxFD3U/1aYRSnXJusWYf6BPvTn0S6f5yQod07CBPHSHPrHT+LzFunSTjo51FGXL3hoXw1HZZ8JiRWztIjt+I0TFFyTvtYQdMVAReiu+qw9DsD24mMncbiOHvfkPcd2TBlDPB2vXbBAAZbP0iantLbSHKFWYH+6V6zMA/9Nb/16kLElV6dTbcXOHxUVCKwXwQBsP0n+Q1RWQ4MUuqshuWt/S/p4cE8DAjyOJyv4QOLyK4pDZIhTpJfuT4PYGWNl7wsBc/fwZWyJsX5I2JLj+7KxKYRwPmfC9yy3QR+Y00uAcCwycgUAXfL74vvwynw6tqagPS/Nj4UWZr+f3r0AYcbjxxMoB+TPCu1BPqMCHXIG0pCm/wB5cNTlWDVmyqr2XZLxrPkO7HDNw2Ho8k9dDy/zXECQBG/5dItrBFNrR28D2ut647OjifCzE0y8A7s3lMG77W8WDZAsA5bTLtQtMUHq4GCygblJRXSfJYhuix2LRRHSSp+fEmO5QNR16aJJX6XkSLJ9BAEaSP3TRe78YQxdq1SNTWSvwqr1fg4/tsWpGgbxm0OBNCeQ5fWpB3ui4vIYccolS4Xj9qHoobkFyjNco9644fzlafL2NvtT2Y7tgpNyOThosK6QHt4h9ioEGHJdSEaiufFKtW/RHJHXTergkOHUnArWg7Fzs0DgFqRw6iwrzJUtpPd4EntiZk3Pv55y2KnrbwgSaKcSeQBPJeMHVmmw3kP5E7YogjMescQu/ddRUto4PRSNOOoX9SNhuhn8nW1OibgsKa3RLHXeaSxU1wp1CfOTq2H3LmTnKI8xX2Tl+bzUSqaFLg2svw7AxK6/RtiY5l2IRMZzj/iu1HR2l48SyVDy+d8I44tT5a/I8jnYTv9TUKWQqClb42k2pYBi+uzG+u7AUGWQdDO7S9Cx9S/lCZHA2e0SUd0b+4VQ6dwe2hB2fw4puJtQPhA0A6DAqIdoV7wy+i70RKIZWMuRSGV+WBamabaGc1tEpVGWVeo6CDOu/yH+ofxnUXLIe2eacfunskbtJtXUSsFc/GAFrueUGFOxuccYK1fbGPT7RS7cEuDhdglPQ7nR7Z7dopvc4gbFY60OOHTZjGt2OH6LAnhVnj/4Z+P3x35BX0x9NtOl56lCdILlQ1a5oLt8jzKgTVp/lYqtpBrkBY2tGN6HeL12uqEVLXvMBq/NYB3/Q7MKLwIXLgqGrBGhBw9NHLx9ZOYrMk5dYqc/CsOJ0naWYwt3xOhvyhBFF7LQNjNmdJOfrThKYJpfe/pRGg7LuSS5ALAzDGZndLJpWrsyh3WXC9AmHXCooR0JnzOBPHiLpJb5u0TNyjtJkjdoLL9mhcdaaGjxlhD6B++K81IKSV22NDoEphUVNt6uDrnY4jMZ/bGQCaXohZgkjtuhEQUAsqXVNzRL9495XpfF1bNBK1YpHau1uG4lyEdX8yCLBVt/TJ7nBAPBJ4SbKIDvhXmNHjaggvwMb11OoIuOJC9MwMFIozJP7DXaAKhev/8gq9ya4hQnp8SxXQs/kG52XFHluqYlaMDu0vcWWJo+9+Aaqsewhb8TTPYwvhle9d41E8TIJTReyEeBVjs/icIOnZ8r4C9EXORN2eoBboZtVWxUkAQSC8FWACjdRU1eUI4xFbmFVaKcpaFWvACPdx/H0Ltj5nN/CdFuyApONsRROVoTawT6iKNWa6vGLJDdsRSpZ40U60sCV6TgI4p/AvzDIsOMrWGqe7PwRuZWDy34lE7DArib4reCTK5YZILToiRTJmhcYHeQ8kMYcI4EN+N84+g+CfG9vE8V5NrnPYeS7xPNtxtHI1Pfop+aLnKPTZX6tgx717IU4z79WhvakF/bmYL8YG0otMpsyquchYdeGCoFmNOFmJ7eMTORDodyNPWLk8RJO4+S5U0nGhIxTwDYixAGN3DNskC0zKVLX/SvVru3ixj8QoJLQ6ZI2vIhMH69wUsNGh8Ed8UJMep+kF5dDdCvxJlyyNkpVIsDaUOWaLHccH3mALnSOwlzo6BlVmAsD8aOmyM/kKnqHvTnsnDnCDz+xL5OXNh4RlP+nH1HZkcLiIAf5cYeCJQfqnEE75u6nXrmjJ+gw/3P1ugIX1wil2E8xPWkkHhbF5VYP9oospSU3CLnPeOWlHKmEG267Z5wewX2vSxTPsfcP03ly0yPzLwT0Kq28gtRi18fYyp7dwy+o94cr5sbPTl5H64sabtpyLYyyaHFIE4EasnSRVEaZsjOKMdaf6SGlJliGHN4dFnOXqCkl7Ld9vAm2G4lWK9mn/nava0Yj+Vi7v4ys41WbSyQSPXEd9rJHlsDrwwasQuYSpM2lp/8k7X6PGF6MAdAAsRixngbgUpWSkY10l70xPCOSNpwc/Ijhqvsr4/OubspoF8oQegmOPzyskL3fZRUL31ObDxVwTna326G1uPORcrVLzlIbyUpKqc0Kv1D07hc4JJy7vYZMSYIcNKfsEQTuFrOIIXHP/Uw6CnE53QATvA8572dLiTzDaKWEatil1IvPtskL/BmDzz8jYn7ZVyqqGwAod0lhZ362aN9/sfST/xbGw1lPQnfLuDNi671TA4qRPp4PPFMr8aO4g33+sZmU2IGH44z+3XYvBpkIq+zURKiTjvT2cmopwkLw2RfAPcAMM9/UYZl/htdC9/8U0458OOfSyTwtYMBUDCN3sL37EWFtI7I8k653In3OnnlsBMmIpuYqZnL5Z7//A0ybMbWMU6DByeA6KZyLlFpAVvz5g5hc0G0cJJnZKfg025n55SnvccYk72OCDCQvHVzWVLOgmipKmWmWmaFUf4oqjUN88On2Mu7+nJwWNswL33TXM+kkxnbZx5Cx7h2ZxVngtBpJuZl93m+yjVSmnbY/OfXkmjKv1s0UGfh6ECvGrMzi4Xmd7LH8x5xNNjz2U/wYlThjaTBvBsiq2m5ZjpF3K3Iu65+OmOG6zHoIpIBiV5hioQ9f1G98dohi0boRdlPS4M1kNdmui7sZWAbqhXpyJ+xYSNuhk/jcxwLYd+NfR1T8+reIWR5dwM0VBYWM0B+3V3dkMXv9GgAsE9q59b05W4SH/aOt46Sctf0dlCViwQftcjT1Q3BJTsB6Alsg+3E+RIROJDufXt1iNuGyeKKj0jLQz6WO/kYRESxNpV7ulzrUwChBqLZ+m3dtbeHbwsMKkNHWSw1crFo9nVENIyjSk/jI29r/apFjJ0NeDBsZ3OPQC2fRkFHADqfGJo0HB5IOPeK1gJX+9nL7ErZhLaXx+J2uN6OQ4fcdD5uciHQdY09/gL/amosNgBEi5Mkmv2KoPLPeZTvEoZ5S+zHsN8LnC3BkGExTWQnZ4CYUEBQXsK5pzSgXxFDV8vwabsNK0OQtky7NstLFzAL+e7SF0K1qIglUEPPFdAysTjeK56n39JUGUqVF6bHaJpMiS/7aGDTrOmQuwwt06fKQJ0HkteGF2yPZKMareYw3QluY7M75VrRurJfuyAmotCsmj2sDhJWfH57r7tWY2d8awTTClnzY2HRJgbb3QkX6rxAxR8suX9fm5HyXwNrxnXF4iY+AWjmKoqoRdtgychcpZ7OMoJVv4vIObZfxV1jb0+NorIm4Y8lVNwMX3CwobUgje1A+UkNqq2UHoKEPR7DPb6N7SQ/Yz517krJ8Ty0EsYDO4PFK0wKYUIw9dNiy9ZzCpW8tAHtah7FPo+TgXKUgDeyh9EPR/5xgoAovDmMKh3QYMhWuIVcdoNgx9qB7E273UihEEtoy1QZBjUFyZemHGQvCK07sBpPOfR/3qmZLW/rte+jOh3yOom/GdOQ+IA5DlhsL6dlec/r1P3YITP8R/DDvnyeS3J0ppDSdCDS11PcRUDmZ4Q52A1JKQhxRKhNo4Y6mE7zDnttj3QvxJi0ymfQz4GPqGUVhF/5UjtO40WefynodQtda/joK3txnpFHeKwtlbkmvJ1oLa6V/VSgZ43F7D1HrmQCPAPTly7Vxd9v4ehucVybxDiJgqailSVeRfaMlTT5gT9pV2Wor5FbrWjJIhSvdcVSqiDccAWOLCzggCoN2xMVv+Ar4/bnfmJzgM09FinhSegMlHgq5yQR1u1GZjzPfn29SIqNt55Y8fiUFERf46zqTmFVSeGPwocfO70UvJY/krG5S89Z30BPH5ncT6BkISkQp1muucz3/cNooo8VtWi/wkh7Zl8Ejt3o4LKQhY6cy5ChIfhZEdd51VWrSV0T07c7aL4NqORxVuQF8USQmdLZzVerv94HZjXmvSzQYfmwxffSfNzzBPeCwFwKoiRoWu9IlXcLfss7e/nIe4ke0g0fiCZaySJL/zGFCaz547Vq+p2iKjKbPan7TnzZ0U7Td0pBLl7nX3ebkZTW+aFJoUFEtX5Xmqa0oDiAl2R7cBrbHlZlpP2AkGiawtV/wVCmrJAWmBViBdH1gmJv0nmBpU0nNG9J5ZetLciIuptugBR+S7JRherujfxsVogLvlByl4UDSf5x3iN/gu53ksC+HutkdqeVbBFelsG7ohoHsqkMKnI/p4riGDw004AB0/E9jf+cTKPRbR/mF0l91KWMJJ6LZKadIu/iXflNFTYoQo97h0Itv5g3k1fxOhoCxkDFKZ7Nt84keN1sNthveGvW36eT61LavsMUR28EAZRqFqqlvcbpIts+b3cFoUc6eOs5bMTHFy17nFAYQisppOU89j4qmjFjFUvoEAhg54dTcU2/11iNiOS7Wu+Zlb+hPtD3E3YEF+ChfCrJa3VqNZhq95ZT9XE0CJs3ZNFN8f2ArEZyJYL14I46SvZoekEqp0+qrUogGj81xCLiDLu5+HZGQLc71CzzSIimV907ni1E3lTNzemCOUhqSFHhBvk8gWKefFyzTcCQ0ovKLHoVo2A8zGi8qbb9JTk/a68fl5Mt/cGzU9YgWxJ2dTy5tWy1oz9W4PwWX0cAn5o4XTi39izgUIjzd7zEqpBTJ+TMANqPdwAPMtmWTcyKJd0v2spZyQYypFuItqn3rRCjspvlizpSGXrahQpzIDX60IvEfNue1NToQgt1DW8WMD45cNAHennPD6LdzrN0z4eaPG+ju/E5i8hYfn25vsSFwlKppfTJwJ2igKRb5SA2p+O0RfJLBFCCFpd+UBNesmIQhYsJSA8sdp3NEiLW+L1RPZT+IsPpJnQW/ino0kdiqlpkJr2Hs188GXSIBdoQaRGbw7WMY8dgNL7I/hfH7i+93k6cILERfOcKE3a8WSUSdHbIb4KN75g702nKoMvI7yWjhU3n1gNuIppXizcfJ17YewPzl7pTzvmR/msFmN2ddz1IEyTRpiE/A68UT0IaDkbH+UIOSzfKe96UXF3m/7Rmcryit6Qe/T8TIsnhLiB0I9b1i91fsngcviHkHTdc0jtnmfrzIK8c/LimCcOSSBZMMvxZn42uQo1c114ntKr7rUr+HI3OkaReIMUCisnb9GaE+k48KzW8E0hf2lUU3yDSz68sCi8rxV2MZ8aqwDMUED3xsO1S54SBHPTrJpVWd8y3B85B8jlqaAqy7+x5K3g0At1xGty5gyg0T2D54ygh9fbnZVH67I7YMRPDyu04XxrNHwN2rRe4dYDBogAyFWaPsQe4XeNLiHJ7RnRsn1dncZ2NTKslW7ZzgtP23PCrpY1vZHL3zHSeUgUrMpdGU5LBnm3BKHQiixhGNIZaP9DYNeECqYmX86aXaS4e6VDps1byyHsugNYpHRZ73UzsH91161tLAg93Cu3lR7h2Wi5BQn0/XDo1NWzChg7hgJ4/K9cwPPHWV+5ybtbFq8XJvbtP01xlhtzTPlZBCcb52P32AvSFNI7RJZOTbVA6yeNtUVAk5W094adzbf7L6hE69mEQvBzHnZ3fOXhvao+P8wY7jrv88gPazcnkTM7Y8VlpF/LJ+BVRVD1tym2L8Jjz4YUmtLusYBHXbcg6bxqix2B//32PCR2lA98wsOUgKeU0Jigr6ULWyKvJxzae0VSTNRxYhFasGGQH0kDpyOot8Iq4mVpv7iuknF91zngS1n38HDXeq3rRfGqgRnrB/NDJo73jFPttmEJVNaBMMYx+qk2ReO8eqWHTDy14js2GHdBnxnFz0OsApVB1WD//Bu29hSSQwmHxwcnK4Btp4c33SC8bVSCHh9el/PbJFX4l4wtjIUeyix/yGlqY7Uy+hwzU/kLNuqqJn1i+esrcwGT5ZUD2esxMJWTAc7IIK337b1PEdZ3oTpEslBue7C+4llF24yd313mUF7RJfqvazgfYXTCt6w4eno1SqXvtm8SW2KiqJWAWqBrnEuu55Q+Hzy0CvTUaNA3/H4ioJvj3NM2bRntk1lmD6S7JIZzxHOMU7/IeJg2mdEgUU4p6yMtvSLni9hzYkR+O6b1hcw9ivNrSO4kmp1+Mz8rUkPJGMHtrJ/fPUBdIeTpurc55N/VujjTv6cMAZTUh3Cd4bcK148MF166qKD9Vr2FIEcNTeNf+4sYgYOgPZo8/1bKJikehPNbk/SZdZ+voqUHQmtE2PpevzvWuF5coVeNs5DjY5mIuukXdlNDQgyDjRNoP0bTgZQr9qaIGH05cqEPFZfuDoWiz+JEdIr6F9BjEV7eerEhLIvVGtO2A0+JVQuMJaeqG1K4leeaC6AXtyKqFMi5hLMkXyOh6/aFrH08jmU1IIjJjbHxVnqQaTDXB6FbGF+bzzchTGjvhVrb/kdqXhBLRklAIaYodpqL5h16zK4VTH80A8DtXIGw8E0kaIa7UDlVEr08UXPKAIONgY0paniaSsrbE7ZMzmxq5fanWnvtJzyIJbKcK4QEFMM3Goi/IlWbsaOWQ6Q6Sk1/iL/+PxF3rrpt3V9jZcrBuIQ6tdFxJOb4ktXECIiIEupUDcLl5modrrmyVqSmDqWiAF7xYcquCg7ZZ1HJJh9ofwAIA27JdJf46HEu3ZLrDg6398Bur2erKG4TxczNUNJZdHAPE5SaYD4jY/QuWyUBKEobMouAWNPvzDjtlsfSobiYBmcddZfdfjoic66xh0YwW+iL5ubCvq93lkr0vHjKfgD5oRROeaAQO7Rw0AaleoDGCr4Nv7j9Y6lrOamkVvKrCvhsq0mtLl5UmP+LdoCC0+wdY2a/JKogdPsVF+Wygani5ufugp6ke9r5BUV2yh3idURvwmOEc+3Uf5ov/K0SA6pZyZxiD8eK5HABsRRiINcUjXiBeIK4wP6WLOvopOnqS6NLisa6EQMYt4y/znwGUW5OiYwXEJ4gY1vq5pLqkTARmSeCqvzeYKQe5Q1J+rA+JYLRF3X9YasdYp2QKBbmURYiRXztM6Ol02VcMq07Zvi4WkNeNXLtecvyH4oK/8zzCG4HTHsyN8aAhmuZU7Z9BknWJCmURCTD8lyq/UhM+KCdL0YiySpMTm1OpvMvhY5d0hw7vrFyutx70e9kW4bx2Q631t3MGCSimZ5xz64lukuB44T1SkZmrhjwvN6OlzGTYKQWKlNoa9STJ+E3ajuW5oMCpXz2U6MijTO4ko+4BL8NyGkTs2U21VzIoS80nS3DacjxkgK9YFx3TEIWFfnHKhPd393sxtSggJombSLpXlYw6fNWnq68Y2jUe0MnTnVBuRCPBxT8CLebbFFSENF002riebOPZXo2LCCuakJc2wcEziQdkJJF/dDZeJPBOWGp7pY4Ria6rrMrAGmCHWx+RLpd4mkQT8HhkYbRY23ECXZHo6lreF2epqtBTY+2E4/QDfsHY7ftzhlhxDyXzASvF2Wq1iYbelOrTZ7ITk0XDxs6XL2d45eKr01Q7q6TfwE+5xnc17ePBP2JM1krXMq3RSZnx6rh8F8No/R/HAhs4tJ2GqAzs7M4iPO+/154gA5/l3CbySD4dG1bypkNG1GQW/qcwFOKyyhqH2kChlr8LAWS7pyzWeTxBX2HQ0p9qQqiexJPhpGtVg4p2qmiFbWcU2RWcyy88bCv6i+uPNMfwyTwnWpNKFLGthasv5i+aWdgT0FcM8dfNQCwgXkiguaCImR0pby6LvDOOyP8GtSjzcmec14gN9mZYYNnEjkPtpH1XR5FGoBtmyFFQTTiLX7cjeY1SwunMHJRDNNGCHOMUE3Nf1ho0fux7OOdwd4hhyJ7oZ9pgB+TMZqdf1xPySi4SbAIeUx/KShK3yCc1mPINAt2DvYQyt+agiuWDb3cNClJFJRIRM4fZzjcTti2u2wpYTvGApKm5nLF1aZV+OkY4CS+aKIzI07BUJkHVt8lNFY8U6/6apTYUKb6dJP2FQiYW5Acs5GGZVQqVoB7oA8iFrFFwpahe52ig4EQYWp1kY2OZyVgw0Fp3sVYCD+jYzKQU1ucKPOM6KKDfgpj4stnGcBEEszgEYSTxW/ZgEzIDzQ855gTKxMl+Ufjga0kFYF71rYJhfvuypKdDBYVWMzbzG1Ag6Df+pEG5GeTUHoKEZtMIoXRZ+B1zSVUU0DDyFn/9+pkOlpGCgXXRf7p3T/B8idb3wnjxrz8WO2L2vH2N0cZ8uW9aCbuTqW3yk2r3tl/jU0mmK8VA1UbLBqaAyUxiHgIK5NsU+tTSJ9MR1JlnqPPoKs5LvBhLVseHTAQD/fiCrV90VO6ZBD/AcmDXDLalQkKrlxu3wS0HHKA6L6wGCXv6UeXr4cP/PxPGp1a3FAV3WeKH/+pgUdZC03uprudZ6D1qtn3KpDlHAEYP7lN4+lZlEuXowTj90UAzs1eCJECKPZIK0KfcQRbQcuyGgQ2b/RH+UVBsSidhZ3Hewv2/yEl4sEi1MbRJZPupmjaTyYUrbxe/uH2AqvKyG8mV+x4uBXHGGjS53mDKFZ2o25a3EeQhYmFSPsAFoYn3LttTWSeAS48LvAFUgruTDU38OwRjmemN7h5HAYeYK84cv4Tx2dmn/dPjMf7t9SlEE+CKJr6yykpgB7ns+AenTFqxZnyDI40Fip0AVW73mw7lmJ54lJ2qa0PP2OUYdR8LZ9Sg643l9mflVT8btpCou/W9sZvVPFrOU0qN0gkS0EqMWrt+Ck8CdyU5CS2rZs6JxtrMzb5+oegPQWDAXaDoN5tzNCgHAQIMd5zqM9pWgM/SH3x66/09NZIH2Bgjbe1JGNmu2a0jrxhndc4BiIACBKJOKEUlAF+OY2qo7whk5Z//97Sdd4lAk5qSukukUooifbfBTnWgG7dnqpiKzkIETut41AgkRcQkrHuq8S6PCtlQLIeRhnuHIemOBv36eyepRF/dOKfZzvADRbAyaSMjR0wDpu2AsuRGLCH0Up79BLDXoMqxqwOHnb7WOu9yCZb2I7wT72hnsMaHyscW7lq0lUPzXYuARivYAnVCiTXHhOhVBNHJhyk+Hygl71iY/YzozqsxdHVkPiWDE+Ljvxsy/3U+4d1hP7FyyzdB1rzqO1I/Ls4TvkbqY5t2HXc4qRAHHjRDA0m/KN3Ulp9k4rKPpXUXtASEuop09PNSWwrilaPqWSfNStfqC8q0TbP7KsX6hd3CdG3zTuhea55c3R3044u3BNQryXbkViKU5rFYJ61ztcDzMCQVaE5bv2jlyZi2h5SbT3YbLmj7zHgbr+07kJrqgbwCUqwOyaplsaOVCEDSk14yconPs4ITLsfT8452NipWhNNtKJf4ssip72JaoRW23zYqR1tG1w/UmsWEs2eChGMUOIKWiDKTlMuB1S315yYAF9B1gM5NbRN62Y61iDdEX/XCPtM7eYw/2Ngs1MC5gPCOq7/31DbOxCgWmAtsRE+wENZcwXrX608KSFJzrrRFN4uZm6spzc64lgu2LSTaDAMNxLcHlGG9M6bAa9nuN13c0dHZE2mxvfM4YXcKSCtLoaeLYvOsphtSzfipHYgvpBl2u+0cYTOjFYTNuKpjMcRD3WbauF5eXV3msXqo6ERhJoSnk5cTJIaCk1zRCFNrpqacDMt7q3ys4aky99mTF1U4MF7fmSzG+qp+0UK8A57aHv75WxwgmaagDyJTEVQ3iy5GuEhQu0IXFJWBDDehu2ddHem7WhJbJNASa4XyQyorjsCg1yevirXsqvrbLRmyMUnj7mJqeJ2JavZLIVFAyseW9Oe0e75A0OV8olV3ssh59oCQ6/CjrqDuqPSAWabH2Mi7HS5CGLvzBZ3oCx4sRf0WiYZ6Di6K/BTq1aNzCuoKJw/Mpl3tz+jMSutMzZKaLhGPQ3ZxDJzwOmQkUKYnqa/F48oMRfdO8NLaWn3DZhJB7SBpS6PEm7f3wDj6FZlyf3IuefM+mxQQtIis9H4YSPXqa2qT4=
`pragma protect end_data_block
`pragma protect digest_block
544094429e424b4f6173dfd8892ce194291b5f958391a4df37bef47a60da75a5
`pragma protect end_digest_block
`pragma protect end_protected
