`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11925)
`pragma protect data_block
Uww+6JqSCcJB5RJkZ2srrVrtdXWGHaLbgVV9RtjwPElSRhsxftF2FOCTjWGPMNtKGYiq8yNFQs8PtHhYa1OGVI/FJTZZ6YD3KgRAnZonZ4Y//4PseYU6wp1BTOrZ+JlvK0otuCo8y1Fiaa5QhDq6sUhtnuVaIKtXd+eElJE7QeuFXJZ+uqTcEj7aO+Q/T3hUkty0b34OMv3FDNrOl5UQWhdQeD48b4iY86XGA8bS46moM8//x8YyYgDPUVWapuC5Vvfbg70qB/4WhvCjPbD9MuiAVJCrVAeolF9bRsJSsoE3MZQWVjxzbiILmjwqWuTj5Blw5ATf8fsvo1Tju4FGGq59z39A4Z4qiZdOVQ5pMqdqqQJWF9JfHd7pJH92zCgVKHQC778lkTBahO+4trESwqLsXXK8Ahb3woEP5AWbOqc2nSKMvPDhqnWNnaAl8LmEN/4U38Vh5jKAO0bvuthAc/yugWbMuKhQ73h/cY54rGH8mjERyN/MkBw0gAFIQp/FqDodJLnukQFuR2mYPQuhBhEOGmomAWR4wVOPgfNQ2n4ZQs/8P46ssajS8akqEF/Fz36aIB9wkWCoZAAnGUOWK6HOaI9+fXC3n03VUJqkswSEfCIFSx6hA4rmQzq5E0SYDXacoLbPyiKtyCAp8WRG+6FtmWovhD3cCTwXCBEbUcJJHJnaqgBWR6UQ4E3PeDSAlvurTbjB7SrMrOEwESqZSk9XrT8hAjT1a7bAewMvYrwCgIyYOItMzKBoE3l6Wj7XHPxP6ujKpf/f2f6o/l78SwtuPwgQAjMfv/seuEWe4VAOX0pJZ883omaJ3fLJlBs2cSlrX9NIXZnhQMqFk+982mUgEdk26YAMmfOveY11XSS3KAYjDHJSW4uWFpMKTOhLvznyeE1cR1HoNn5PQVqs2I029EvJeLcLFYg28cj/NqN63l7EUW80hpyWcsdCv7WkypGOE3cJ7QbYRgJpkw06x8O/QL9XnoZlmXEwTC699QqTixIuZJMfc2bY6Mtib5hmoy3AIoiaq24nr8BBM6FJ3njOrsxxaRV3eM3b3QNj+UBnaqp3ewURVNQTuFPWt3IJrwne9wiSYVbVTcP45JmKAHNh0zExBRAFiOFKbCkhPyPsfElHzoJ3eYkEA+udSJpWyIuxtahotuBBY9AbvZRam8zghlMczAkwTckz7rK+Vt7IIZS3kizJ5DIL2ayAl28fMiKQdmdDEa2A08yLKvqMDqWuZF93GrArqkU/LGGTITNjsvSiMIV+3kf7iDjoFekOXTbOgb89XRZlamueCxZH8A9wCqRjfgFmd8rYQxag/7Ay+6vU7TxxA+WTF0uneL/ozwAOiC8pkvZ5XvMwir74ASglNnmQQErCjmTSSxiD9UwL/9CBns/gZe39ac5nZAeee4RraE7i+Oi+1ho8RJ4GwfvUUKMbpSUF8osQfsdB5jM3J62sizJW3oUj1+KelNpZkmnnffmFS3h8l9dxBTKnwYKiElV/w2lkMKvC+ei4j7YxPYUtU03fGupOqi7IWG0xu/RZRlQqVkvwOXO6MA+Y0bA6cl2BJQcXGlOiZjp4cTcxjC05slKqU6JtaaVr9o2gEJkcpkfbEiWwdQwD9xjNLzFmKi7MJFLjxs7ywpmUzrdl9TwOrqZwQhXuOeBpnWZKTUfjGRa4cNd/71l+3iFniRlBI3DpKcQDQuqAwLtD9Y2TqwWK8bTM2EJ4kEC+8UaQfY0/98Yw7pEXgnDFMh1t1HjzDqiKGBbr5J0ebdap+7D15vE+qkEAqJoY7d/nY3Mk3C2yBNJfz+O/a0/tSuxaYrTKsyekEifxJSMNhPIwyo7D1mwtRL08Na7iQOIQLX012Tzx6mnCoAhnPSG0bcLkhqli3DMMVr1i+El6AEDWQAJQO+ozZOEciuEBXqg4RjFNPzAOKO8b7QT25vZtjqNfCojRd+VPG6ern8rYjrDGv9eQcFZljR53MLejBJyoTGJFZwE/c9LlgU5GJ5rHm1q1MvdaOKENAcsp47Wc6ZFnz0O1oObwp07mO++yTIk7GMhqr3PXPG3UbOnmr+FTjkyCgtlJDL6AeEArid+WDGR1LBCHz75dfHbQfqK8rWgIe2k/i9SoXhuUFS+5rxbj8d2bw3XvinoHRNd+LroHfwI8/59Hcc2hgCZkGQkU6ljbtnwA6Cud2dKsG4wTMab/gQpBkjhjwKvv1tmeLvgeX8TBirmCvlNNRaITIw4swVX4LnxLGdzjzFlvRHrwmn5lhbO4XBWP3vtXf9mKB4s8BI9MKmdjDBhbve5O7YPyZlvx5hsPVxnXzI5hcsiEe+8XGgWX3DDOeWOVRpYzpdTueAwoCqb/kuil9LnC1Ov5WhTHncs909eCyDJCr4RxFbLprDUsyArfmx5iAdvTMThqStk/s+6eCXDIDeMPMrTB+UZW82vSkCsCutJYsXVWxd1k1jKBXSxGoNMvFZsNMJ6coub2/ELwO9Vbu+Jhmg1Ug9tmypG33DYeBDO0j4UCf/A7FFyRmZfSgWv9q4c9M0HN1SjpdVSPFJchz9atkcDzbHGRqNe8p6raNhF9B8sNvURG5lR/jxBG1fwK0/URsv4VJxJsTowHExyiPp8GhabQCnmZsh+wCyj3EaoYYJkC/rVhTOYKmQCT0I04vGs674TslEq5EZjc34cU10Oxe/9roBzyjafGoIOUTxBIWkz7XXj7sgPSA6DR1PTERr+ND90PyBjzoOnCMrgee7WZjzqaOstNy4zeyLW7K0kndBwugKGasXt8BdKJ7NXUAeOVuO20f3I6tjbqzB7vKfWLzYEMOOioU4e8/gr90UA42dxDU8lfS4VdLU2d1MnS9v1x+WU75BFPjYqd+ZZFPilc+Y3Rn8atlhynBaOkDiWztc7lF68n99k2IzWsnlXwC2rjmfk7RnGnPd1Tzhd2AxUNJJqJCm3a0XItA5xGzuAo71KRr+dB1eHeRWBGbvjiI2CQSty0nAaPNNPUouvaM6Nki7m5v7Q4F0qV8/g7ecfNe0yfUiJ82D71/bD0E1VC3EWme8wejvTQSNgiHCxuheNNET1wDQdsiMcB5ZF1FT4H0oV2sz1M6a62ahzwKA+JP3K14NK4I75ZGfmxwSdYUmgegU4DB8YgQpAUuR7Pf/dSf1ror8gbQSmkCD6jaDYL2ftAKWjYr1prgbUB9W5A4n4R7d2aa+K0m+nfbEWE2ffoOaq0g9TdY5pd5StGVevhF21kOxvffCUMAEmOrEnLqaLo6aRzDrzd6CjiIKjGNaDpdp3aH1h5WRkCA0Zz1lHDLPLdJFmRPvzGNz+2fh6Onpo80irQUEvesyYhhWdNtBh0NK6phbT2QRsBCRGWbrfxF23cmGDwGnu8Shd4q767/dhfQ4JZ4Yq7Waaw1XocWgVB2npoTrRlctj/snxtji0Uz202R3n8Ec+afIsPmmBNM+ViOoRT4dX2JmsB/h1rkaegs4O8x00Rx0Wk0G3pwbvq8CFH/N4zf7FDd0QPKUya4sSEL+SvUr3TofBaO1qA7PcUfeARbwFo9ye7U6hH2F27G0PLntIVwX1Qm5pzI4eZV/raC5sbDCXlvG/J8J+8mmKxzRzzb0KGl/8yo8rne5qzThHnMljPMN2JMXxFtxnnqY3Eff9Tg88ZMxvtfxC4oAoaGn21w1hskM+P8GhyXa/5BSS2LcUuXWERtmz/8UUksvV7cA46XPq4DEjvMUV5wv7ug0FAKWGD8EdasPb4mReslHKDbIqHBf0+J5d5appIx9GtwPWl/dmBUtKT4hCpMnTBmnnDPPgCcnUuWk8ajBy86yT1zvB33TX+l5aec+wRFlQdKVN3lK0e/Sruk1tx4XPUCVg3a3qqEgsNLF6fdE7krl4KjwddorFUF+Dlr18eoNpdhEBa5U6k8Ad5oX25ApPZ/b0qN0s7XSrueKnatyM1u1IJud3sdaDDudvFCCM34oczRWrDyWWtaie1km6ptIYwBxDz8VZe2X7BBT9Wylc4J5LoFQ7i4KojZsfBNyi/VWQRrcNhn0330PPXT/HB+9sDDyXCHV4mI/vm/aNGb35buHD9FbGreLXiMdFLBqeub8Xf2yzdAmtb8gsLIvwripGA/ee2VxplXdQl7duuEgz611RfkiOqtmKKycTbMwMzpFIC7mPUoevr+g9BWZ45yzOLBUuhA9uueNG8Ln05ODAgQSVd8gsFJ//jeliU9PU06vHGnPaDYnIP+3mlxkrWtW5S8pUqmAu96K+Q1PKDtmiAmtAn+yL3P2WVK6qr6HWeZpEduq7QpxYoGGPbgjjyE8JFUTJLCoqILrSEYXm0/YQil4Ygzytjfx8y1dVF2hicA8BzWdrwkYPePWv+wtvaqcj1tQGn4IhGIYebAb1rilUE5Qjdmuq7db+aJ9IqGmmUglbfDMRGtqM0pJYLA3mxmAGKSgTnoN5ZGW9jVTnBHHFCEz7V/dAOzBmjU0O57KijgwPmNiqdy59CqMsaXEnwSI0boL/lOlosls5EbreXIAx6RLKEJsNd8uoZXMmFd3+Z2PHemDQQSJbLqviV/97x1O46u0snljEWifL9beNDHjs+LxStXIUh4x9e96ICcbGnbl+ycmQALfGLJ6CPSW7K+mWI5IKIXnknWdhFDo6hQ/6WylpMcWPhyYmIfO/iKUJQPIEN6vHEJ8Un/dsML77NadFS6urm265hwzDs4pKKaGw8UdKkJ3dgw1e9I7UWdPbHM2ll+Qxe8u/NSrwm5a8d0YLVbtVlq8kSXvLJr7gJ81lNJa8I+PBmiW+gX4HpqxqK2ejvUu9lhkSqWCbKIbQcYB7n1eXKqGefUCq6yfCzFivfc2fiq3NUaXq1oMV6QwxT1GfFiQWREoh75tRnEY6jhwpPrltaKqetunQ+l7UukzLULOpLzJmIAiRuiJpjdxQ6YyR/2bF+gkDcTwfEoa69You9NQaExTnq2m4/ZwbkrQR3C/F82Rk2uCfyBlYk73b8yE6r7Fj4ngnuDyZ1IAopdI/BBPw9ASRKnXibI3x6lFjAmUlYNldDTHfspJ9lPniFigOd2+/cC/LADYS6mc97oPSWViNsF621CCSbxoKQ/IMku8fPEhuEEIwID1qHocakqcL/Q9uorqoKZD/dPSRoYmREDZp1t4qJHdAWz5BWTj6FP6LCcr+m/OaVeq8VZrnJnKh5YYrWnwcII7dZkja6RTfXA9l4y9r77mw/atu7SKXT46AmrnyFRdMT0Tjy5bZ7VTBNlozF3Enyek3xtESy1U/4sEOgT6GFqdMQRMzCcONNklAPI5shxrxSE88BbQhLbwepV8lb5pdYld+zvgaUDgfaaGjxPpW2JE6QAM5oGQMJCzUeyJAHyZykGXJnr4UDg24SPH/1+OVBsLrFNfyoIq7uJlGSSquO6C6hCYdSfeb95Ii6VIpeHzhrmyh6ucMynSVwNKLnMcdQapA2PHl2a4bm0SFQA3+cYZ38Jl7oNQF8NosPkpQ8NQv8hisHNCAPY4zIEejD31vzTCUgevs5eh6yhtjhtTJrZPvfQcJJr9PkMSMlWM+v5NcmCo5+tQCeK97krLdI3Y7HVfn++ogX2P1Lj39FpjleuaeGSLRzfxqA+R0e0nU8NJc87xtGO/ylx1jHqE2r7562htBZqMc3xHpcYFmXpNRkWygzQVgloUUxbBwMA2arX8ziYz+sxwjliOVgZRnuOFJjdT0oNNrrL9hZXNce0SaOSIUHdKKCu/Iw2jua+Dtm2pNfovzbP6lueUsaUBuWw5ILV910QSAzpl2VcU/KLSvhmYSH8BRZ4sW3SNUm30FPk1PK2CtuoEFcEx0+9Wqlafe1Kp/CbzcG8ImbW0noPpnrDmFkkTz+9wpDp10xr5UxZ+ffZLvuY3amEzF1umLZxvvrzySK7H4Ci207hBDrY48PUB2xWRWW8H6mpYBHMzblvVHRnPZWKfohbnlWvInzpoWb4h+lggzKLljM/HrXAIAfcLCzNUsgUpYDHWAh2yyhlGY/YLFWlUhZpSN53RpvzmG38+gfYWa8aZ4Z5+wXU2/k/uGzt+7r3MpdLR4njf5DkRHkBY328ZwwDfatz0qIfPLGSS0x7czMXyJphhFIg6aSGqiRIcOuPfR2vIduHPNjcy/mVlWZXoGC4HUmRNVN48WCeacgfsmssbUYApPGiGAZeg6sLP3kARUYvq5nRDgmTcRN6ZNQQwqWUIfieyGKp7F8gbnFvUs1ypKadBSMYo22q2t5YV6J6FYQOGGVc5FBBVZ6HF3TcPZ4nqiqahQGyS7DqSg9cFlzXydkOLfEaLA+ZRSXWu7RAa3oNELPnqXw0u2Idt5dhe2FDDdRplIjmJAfoH0CA5f5zf1sXMf4VfQWIgKiYqKMrIScao47ZOPjU/UHWdaJy9BLi1alECjpf3XLC3VpUb87e0BATflatprI2Jdb2ehi27Tn++Q0W5DI7nal+hBcfmG3/OCEIvkaNWQeMKhmjL67xXOZ5quaDUIrO2CBo9G9VNvwY+fETtELCm4nd7Iy1VOQgvDxpbQQoqOo2UJ+Icr8blDh61CeNpmYsUezion4ajafUepebuBsb1c6pv6+mDTw0XfFlIdtiHu6FGqsRtbqloVJxNyavWdBxqKsYnUNYF0gaTOXTaerAlW7YRI7+5u/nbbARBqLXM0zzX99WhpAF8KKRc/o81+U9ODxuwsF94O+vvAY2siXvAKnOqBslMJyWMh5q8S3wjhovdegG6riC8nOa4VngWnAvijAG7zoWqAOzLeYY15AsWKmvFMI4oWPdJROBEwld0nfHjVMaN3zZ+kUddpsRqavhvclQsin+F2YmloMjYEQtXiPBJYRDXNzq4jOgsZfQRlQgvB8HEg6jUeLexgaMiim4v/GxnkPZtnClkN2ONsWw/mYsoPdZe77gS/XOG5zZ/qLoxUWyCO2MSOcmFoETK0o2FI4ZBQ5FsTikvwmgDnsSJD65XEcGlVgFHgkxQEglYoqEPiZdtRbWvnmhxTl6e1ENonWiMVgoiBdJ1K0VD1rDLLqrCewYBpTWguTwTMnkL4g5JOhR6geEHvL7eKf40kMGOqUPFPu+YbT9XhripAvSmPLewTnmaGS00oR/vi8At5y9eFJHVGowcBucEgbdHL6DdOnK5A2kQ/edZzRlWv/KAiGgoBJUveGbcup6ufuUDImovvos4STOI68zG2GYckMh719x9+Z53SwYfrvsCfAFk1brdTzKX8c5THJB58qQMCfD7QfiuU8x4Sqkdk5GMBU38hDwLzvs800hNkh5q0HEkMyuZHnRLFyDU5Jr/v6+im2cfxNebzgz/oPiHREKJHOW90NtoaO0UO1D3hyhBfeFUEGrNtfWKBvZl5rLXEB2tBdSzmhK70S4ZHGUEirMvDh7tXtyvnT3/c6k0rQZwjA+5U+LG3Vl9IS8vRTEkpyI68wMVKZC1dNLcBn/2vT/hFxW5hSWuVDVXJ4nRelWYShozALZx5I/Q7UgP7vy/YZSEOR4yyB72Glu/bXUXC9MDIhwG6yhCQ729NQ82X1HpNCQl5hZ+UTPWmCf+303MQvL0j1/L4PT8TsLF3VK/SxdphmNSHZqsxWFzEeek5wEni5+KuvC05fy3TUMh+Psne9V8iEMMpV+akmZXF6SrGI7Qyn0sKkgl0kUP4p/URDGbmPIHjcm6/1mJYdRDVJm+45toyaQCnrlgKwcAAwp0/bJP7QImJDaKfu58rrC5KeQ1fAjI3pXlABFbTCymNcxPG0m8HWNFhbD09iBYz8AXQ5rIcR54sKkNC3BfP+/9sz1bwOG2PRtH2FScUSEtRb4Dr2e+7HyrBPyVj57v1ncV+fmMW8b2fsbTk5kOH6yzjClgMe+SWeDzxIjiTF2rdHZZ754BtUu3gMnMDxUKxg4DbdL1ZouRzIeuxElqSrkWu4B/LBF2OfnbeaeIReWSxx73EVhFv2MZSCBxf/+6SZJuAMjGTJ70ZmELUN9Kxb+JqX7zy7KEux97G7Pkg7d3hXeDwrIz03bbeENws/YoNPsF0IXVZgjUyvEgs5kEDqPo9Mz6svK8lj1KYVS2/waimOF/Zow7BX95Y1UN0OlJsF6wE+km19D3BzrGrmTmPmByHK4B8Dq6JeOOlHbuBVgd/MG0riggm444ZLRpOJ03KVde1PDexyUOZUUd8aE0YclqrTQe0hy//99QpWtj/eMDdPHI0E5Ku5x+p8XBmd3YeiLlsc7etk7ilS4mpEdvYxMsL8g04zh0lRMSJNB/m+L+LKZ2uJQMZblXGNqslXjQ1dLVrFIbbb7ZTWTk8uB8W2XVlHRdZS2Mn+kPT4igINsXhKO1gANkmiunPy+Ik+wlVGHRwvLC6o6Q5zqtMHky84LzIzt3QtkC1nAMXryURnctPPzYw7UbLzn0gcyou7FGc6R3qukNfpNJ3yuAzU3QY/rFSbtSmwzacdjYI3dW8u1pyOGJzhwHY1MKMMCHrsr4Ou0fCpPpgCUyMyzAZ8RFmb43kpZ0x9fbYoh7LvLohAUPJE+He6MPz3WrkkrwCwIM0A1i11XLGCqxyU5801bpbf0tMesMJiOxwHxzmR73baPNSsv8N3Ik1FB65bHe7a7RfHprfNwUR89GZfFfDH1o+pNEHD6/U9oJ36Q+RVrPRXJnmku/1vE1J9xBy/djv6fFjn3TZA85H0e6vIu0xnzWkJGTa369maDsIJBS0320I0Sek6EkIAZ3QVC0k9nsJHDyR3Lg4guH5IMcZDaBUYiiXuL/5aaVWpjD40OPEn2e4B2h9L5lnfF7a64XEmXIuIeehfoBN68L7iR/XM/8GNj8rB78f64a/T7w6wsCsB/4MWjJvLqnDUHaXWr/NARD4NrgOjYip7ybgng2tjifrREHiAY1g1AdUFmqsJt9WPEuPbKVaEJrhoOmoJZnorc/QU1IxRI8Xp7JJm2LxvgF5sfG9Ev/IxjBSia4ZLNATJdDboMssUwoafCTwaMqgnqiU3ZT9HkVnXGwXcF/5FcgLvixLMg4fo5snlkv6HB4wmIViRkTMP5lf/4OxTsE9GNUktLZpSPs+ZzdXCoylZ+wudb+6zCQ4WT79CXiWhsaYoLaC2hvqmuvLT0KSFt3IWrpN/votZGf9mdo1mbFZk27Y4VErqwV2Hz8ebE3BNLOpBQkGDP0Whvtg+1oGB+OaJxZPWFhScpDoZJYlWYSvesvImCUWGn7TsvKx+GyLfiDWVFyttsJ7eFIoHIU/+6KkKCk/5Maej13PYx45Y0o5UvGln3kJYr6U0lATbl/jsyAe/YB6NF5N4BrRDiPnm6TanG30UiaQAtw+kUFGh/C6dJ5sd50kZxHiezLGF3N32Wdwv/jKumAvzkuSwnqgNfhboPG6wlrV/2BxcIE7ybA8fBI0ugP5IeIM/KkjF/9M12K4ti+Z39XoRXawTVWNknqGaAn2VAZTLI3DPgNYRyK5dMqWSWy/b/vfWhDELpw4TOLfZZbgE4h15GmV9N8fREhRvvGrpP1reOAEzlR7v+Zj5XAxEnspHXgNG/ZC7+DOKOAkxAuSWo/Jhn16/kiOr11gUQY59P0mQHSJHlZ4SoyjO2YgRGu7HxI9pFBjM+z61pE/iGtl7lhV43EYrzFviP1UG+UwOOZUWTJAGwjlftJeYEGUeff13gMdZX4IiH4M54QyDW9lft9hl8JUgo02SzIuU4QjZmV/C5iYJ2ZHW3fB1d9IVOHN+wbFC+QN8OGXw/q2Y3ftxMnqv6d/TP6wIRHObcdLUTCxFnfLBHyMc+laoHbvSdC/LLDAPs0pU1z0mQNDYwKOnLn68Is6hWsGv7b1ywOqWu/1ppKtiU/rzD4TJgrIw8GBOw80KLsjWs/1ZSV0ekLvFQ2j6XdETiKE39m6ODfs9D7xYva503+X7WdZDb+9zVd1YuwWzfl0RQEv1iMMeTQfbwejomJqBzBDrTXDN7bkpqiom1WpQMNv0w+tNBnZU8zWUZd9jWmtEcRfB3gJmKa8hYTkaciDlIQeZzxLTCEDURefUAwC1fz6+Cn0uOCB4qILQK7vcLVJUqTcjNOVp1VYqRPnJlQEbT1nFkt6Ns8Ll9fb6I/bKhPnTcL2glbX/okU1TcNuMNDjaTxyREsJfaMps0rmuAVu9uK+DJX09Qdo9yKfmana6rV+R4YgWQ/6yPqAxRCa0JRjem28enUw3SX0ZDq1WhBo3WBke+u8EVnUFZJvMkD1GzxoM8qMSuyzrSJnyCHhho5xWtnDodH3p+vZiP9OVrgdfbHU86eO3Z3HswXFXSFKRDGgmI6HlFrrZdQstt7+izBLNkBipL5ua2nD8QPZotlabIOsqyXpEtRapnJq7MQluXiZBQ+sgqqZVqyHN4kPAn/rAaRjK1jgLCP04xIX6ehi7Y1wbBkmzklokktnyL1ZsRgV6lBRc/MHCyxB37JDKUAff++QhlaZ6nbP1l8snPDcR8HgtCqlMRiplK1fo5kjyXN+LCC4CVmClhySqaGCVNDyH1XHU/YbPOZDnSLBXNWNTX7l858+m/SWcbXc+BQcKz/zph2QbZetOoxQclM2W8N+WuAHjb6md09/dcQwbugQuHuFB3gIdKTXR7+0c9b8W4Y0yGJeGk4lS9qakJm5qBdqTZ6PjtF5gOVb32fhLK/+p5tvBJEIxtUwkeIx/okNKek8nBHNiePO6cYcGr+yUXsGGqKhVB6sfYI2bojD6ldZbB67mqrcc3Y9c7Dea29Fo2CGpcvOYUDZYUJ1bm45uf+KzO0DApI8QWhIhWspYiNKhJsCsZ0dbnC2tkZwhGUTnweStNyA6Ae271xePJPorkGTNSEa+Yy/4RY4I7C/uv1lthVzH4yu+x8pBtQfhPRvAPxB58LUD4ysuab2jSvSy+o5cIbXfOGbuj5UraH0IDFiZISq37+FkRiISrEzVXX87EDvpJ+XB3CD53JXucS4NQWR6/pwId5Olo1ZO3hJq9F7O0pTjH+keIoFrZDkjzplmSYymJniFWMinP5OBK12gRHAcWKzHkIn1TO8HtS2B9zPXtHWbEACFZ3fihJj2SvRKoX9DF5cb0nR5scrAlNO4t7KbWSSXRSENNS7ndq6H7yTaQo8/T9KZkiwl5OKM98LNPPJ1IW1/YxfDO31lrt5nVkym8NzDF/9FLMHc7S0C5eTvXhfKWpDINcLPl6X+5UjV1UpDfBVC0zpFGucZYL3guidRdMlxe1j0I9MSxwP6oPMg1newz7ld2lm8MtVungdIYOpr923e5AegKG7lmVGMlhCNPdps+ftN2NOsID4nUAwsOnVwwuHZve+yJwHRQEbck40uK165k7IZPsiDwdloBehjZuegO6Sqvhl2gAu7Kn2hcCCun1JV9OM6l/HvJwWHNL0CqDKOk8dt61cXxkjacHesXd7majsis1P6NwpjjqgMmMRSLRiTfPC/xMKtga6kS2gjyH8MvR8ezwh5P7k+M6fSv2BjOKaKMtKvhZ1bENBoj/ZKDdfMa8tyenGwJ7l9lIxj+8lKYdcFb5IcwQoUNCdjkHFp/FKqlqrqMGgHiogxKxrKCZcLqrpkvRQzZScgpQoFiMRatnpV/f1/2DCqw4jL6f2ouIq3iz1ZXYds0Fbs+NYd9h5YuQdTIecPRLvY+ZDmdfsoX4xr5nBclWjzhAaJqMHaMkl9ZzXETu10oj93SaNGgIkLBATNlBgWIZP3QSJdNJ9et2JztfhPYEgYI3PVjnZwYC+2NEJHoXDDDTYlW/4C/rjrhsB0B8T/avz8NL3Pyx+hn+jhgPU2eTxlYGR/oTvXJqAFOTYp0wTETA3uuf6dh/BIuvp0s87ZfHxS45ONGymaVIGWBKjxxGdtbJrGXVlT6QOtG8EoqYgNo8eNFeekVYS3g+oAPWXLcUoFS1FLrIzyzYBVXDuPORKyB5U/qLcBFRnq/4FJ33LBKAVlSxdJ0zlmAWIey92q6s9dz7U9O9A9ZmWNuRyRwGE0h0KPY+ogNjXQaXNT+ueY37efHOBODjZIw7joViSuoh/1Q98PJ8E09O6ISiHxnW6Qd8hOlsIuN9U7V8dFza9Axk0Y8L9VVCajm+qwPE1si/v5/U04T8SIAvQjNdyCkWNzML5fYGfuTBJsZjFFH9AKAay0iKglRXrb/X3QGK5qgnC6QgGzsGhAuLgj0gMmEIsi46RGqsgvaCkI+KyXQ18067N5RLO3auID2HQRRhWC2KOkDWojBY9V133RlzCE9gEUaCGSZLIuaOedw8y7PItfomJ7iJAMQgnKsCi8Hh5dsyqpyA4gZk+WzYG2ly6tfz+lz+f+3MXo58PhbqwFWaahCdUZBgEksrHMRiWRMT66Ars0DQax6T4CADjS6Ty3hcVHk77th8K+6GaYyE/8Gd3nrsq0oVuu/L3Pc/1XUZnTwL3EhZq1VSR1N2zQKcBTE1QSKYCol59IQdDPfwQlqLn2+oylrgBb0TYBfyvxYQekVzF+YZsdztfvy2POu5OL14vBaSG6unVDoWGipndpsoTm5jsi3w5BaVboF/s7G7n/sM9/raelVL837L5ShI1AyyIPd8aFbERbGGLgDo0+uHh5iQ3oTlfmwZVuliWSKgfQMPnZNWvNFC3IsLEfWzYN2SKO+SvXy/h2xxGCXHTDGcUAVDR9YG2ZsZ68dXlkznd8Uj60TSy86dsi40W/RJFM79ctq1tAfu3QMgM482uNaheVObGM5IigFxvh+v+17zjc5p3jEFKFxmkHGszLeTvuAk/mLgE7RuEYZW3NPJOI86o3iw1fFCJyRy9TduScX5KvG393fPtPRy7BALV8or0/2Ssr8dB+Ni2465liwY4QQ2ACYYKuev8DryXcMrqTG+3NIm8sQKVp2z+CStC0vKeibrbbnE6G4ncFl3xSZ2apQHba5Kvyzgp6wD9Pe3e5ofHKZyS9s6v1cNPOjx3U9YaJiv5ri47znfjHABl29JFRR441ee0lvnDT6dilWxnYdiTguQollQYtiag7+kGIon/7vNfQ9NdHYset1LRTf+Kw6FV+6CBDwKxlyUADew06yqCqZpsAk8k+Y9JdnvBW99++PBnNU8xSKDf/yYfywmOG4bZuY8o5BnHpclwP4rA//lS194MX/WPwDE3HBpQ1tfzDtBM+XkxNQrowXBst7MmC6aXI9HPtguOcArIvDDiOlPdGMceTx6FVBTW6S0NdJFJck393iu3qhr8H9tA56ipWTxEsssLz7QD79lPnKfFJq8SOJ9rEnLRVLdK0rPjSKv6VRxGlCSrRRIvJtFnsWVZL3drt1qiBc/3IfFZwYTcHtRgyJrN40t/6uuJAd82/+sS8mveNH/DhPEBiVDMpCigJMGiu2maQVHggeO5ycbowHegD1hWVdC+l1uNAHIpWM5Wokq4fGvRV8ttgKbVunCUVvOL7MMcRdaadgJ1biYINomlhq3TLNn2rVl/0SJEFl1th25iiFIL4Yw2WHBbVTbIUYf4j8YD85/oZkbgFxSatp9zmiczj7SO1BalZcsqBIOBt6f+d7fJe+EwvCmzwQFiKQGdliLUOb7s9SCHEZNu2dNAqdPk+S31LwlvxCR+Vi6LqRTs3xn6B4OoG5XIHKX6BRv+wkovJUZZYeFKnu2UEdxaOhNu3oc9DKzc4g8qZcVhPrqmovOh+aNAUGJCsqKC7wyU4QGXgZoOgGsKkAuNDYfNHA1UK9mAHLyOAGMDiTnTeaLMPoMF+Dxpq6H1kjuKvRgKydJoGUaYSOParBSZbPFV9jWDxKY51RmUD/YI9dWlSVQby3bi7Pnfdu97DaEZJTiEBGHEIlKgVxfslNMKvNdnOKR5ULUMTDbNZH3O9ussAASBTipk9XwesckmKlhiZ1qfnHZYUkXQzfh5/hMDgJz6+jv2ip97Y2lJA8tfFfDKTDZr4LxohLT4yRpdxOXcmr5bqrXhqzkk7xdfcyFHOdlDSdxE63NYYEReRnd41h3ohjxZ/n0oW1qByidW9MwWGrzPM959EMRKXRzbU2sMlCv8xXZaINgBbz9exwRhX/oN8pvt9S13U+nEHnBQTepG2jy+oZjtFE57hT/M2P4UZhby5BWTokdIllS+7ekyNsQxC9ao0BU1yvoLr+E6skjyaAq5E9aF/nXat1YvfTRifdd3l9B0Kartir9YKQB43Fu2djCsA0puYadqXpbQcs+Sq5Z2ymlA+wNO2/4UKVhe3RCimbVthMhjodsTNbPLpSZFcMRK1Ym9miJurI28sulRGW+gEm7i5GIqf8Lid55F6J+BbHHL08coFWPR9lJSksWyYRyDgXgRV7fvLvAGMOPW6CANq8WUgD6QTLjxfLBpzqiaxpWVCxLYwJwQNhzio/bxkBaUKhuVRcJ4GahQTUVIJyi20BUoyERdSF39V2JMDV37sIl7guwWnvJVUbV7Y3bwdH1NG5dIlKfD7Ugpz80cia5iQed4bdcn7DOO8zRmQMB+rYKO9rWRZu/gCfWjWGN/QkNfNY+1U/46oY3qeFnS6wqXr2vrfLrq4EosAQW4+X0wG2rQLcO9o8hqb1sg7TmokRxxDhMLp6hs8mccI0XpsqntwEs7G9L7m2lQjpu6ck5Ciutfz0vgop2wP3qaNlSmVFBGtnliT2lcIk2XBB79aikhQTGv6z/ZRd/95z08CVtc7X9aZxVuLP86aqaIAXoJ/XOHxwT00pamVuf7eMdd1TF+wURI1fkETkXJYj+OXeQBYZQ99rikcGZAPZ2SvN7TFAdDi3G7K5OdasQpDSlnP1UQOXFZCgdf/XSsbpkTMgNpgrg/b53mEovSFj+x9mZRXnWMNUuHt8iqPxPjcRFX5ZDxWDrHF3avZ8xikAMoY1eN471ObgWr7ziFAZmgyL0H1aAC+TeTF5kT0x3Ysepdsnlf/q/MZTetf7uDwLE2I7G2+AjXxxtVTdCIe/qtp6A9uIjEpWyxszTwQUhUmw3i25eP887jW6i28/cv2phZaI5j4CusfXarirelMFKHyzCDwdTAZcOYNt5QmGyZxLC1SIOT0DiSh5jz/FEDeW4b282aXfzLHvKf5s1j4nYIyn2nhcNElOLu4+lgKC1s6bOzpepitS0g4eD/I2Quwv7pLg8NVvUf82bJlAlXR19HmxN0pH6vEsgWy/HWUwIsEmjkFAwzpgqS5pSBqlVDWa5splialylRf3+9lmXMpcZz22f/oAOIn6Ljtt6v3PuAfo2cfhT+75hJ2IMRCx6oibJaZp3NNVeCsxVm03JMx3nCShqW30OXOBd0I1jR7r0Zm5+hdBbMsy0fdanuoml0dL1yxWT6Z0JL+pePJPT2bH8fMUs5L5/cVUsaicIV1xLEs++dhuZDVrn9338QK1xOKn910fbtsmo3HjLQtIef9qbyAkNBShUzIdxBT0mQqZhDXYRNxGuVUWyxikeFTr5onnT6700POlSlPwP8nk2NvVvowf6fq1COjcu38x2MkFw6eGIOFFJtjjcCDu1JqEXW1aEhQmZl8JU0bhs+acxnHZrpzCpeor16tczMXC2DYlSSytAw+4klwUm/JONb8MvSx4xQwUgHhgsY0sz+vTxm0jot9LVI91GX3HRMIRd5JtJnu8rHBAuCUDeqzLNjtJ0wMnWcAWOx1/YjvJv4lPzXDRuSPGcsVWWA79un2lBQDn4rGiK5OV5MzmFGzHwyGPOtlgKFurf0QLyY4h8mlZmEM9lZUMm9812QuBbAy7EXGf93bM4fkEjJzYRTpY9aR6GOJkToR9plE/9B7ZugXO790zKHLSUpOievH7akrcum0XsZWwCHX7eZY7NiatLScB2m2x8M0sxZkRZzQEaL90qjc4C5tFNKlXoD/AJRec8Gz3nIXKKP7EGHH/aAtjRLjj9sokS45cBTafLnn7mtsqpCi0/6pDpNFAD0GvNKmYJ5HGnJ1F+fcB4q0n6/mq+1jV5yN8ARkwPRJUvG4igEbx44U9A06C+J3E5x0dEcIgcdpxs=
`pragma protect end_data_block
`pragma protect digest_block
81a3b943f749992a7c30f60d9a0e005b84166cd464876090e03a0048be9a48f5
`pragma protect end_digest_block
`pragma protect end_protected
