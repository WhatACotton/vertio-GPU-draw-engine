`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
tl6ioTsTYufyzmZGRw4NjKUw9muPszUmuhmHR5Na6VS+hsZkbmWn5cm32vHfX+pv4rQKao14RWDqHLufjKrK4dbqpI3uABAjQgE/I4wXP0ooUYTWF4f8Ys4nvKP/jWo17kZ25VWzk8/hD0elu2fvO0jJerClDGmKOgR+MLM2568eicNDPlF30E2LLZcX4cNKzaQonfNmI/D7ZUf0WxDF0hKWPIo3zKjomcj4hOgYvTA5LvYZhrQHCs+QFj+eJp6SKAuFKqw5DwZddjHHsWfcEBSiz0koHss1Oskpb0eyGFHc2J4YgOWTARXLxdc9FiO4VrEYC62mlNmmBezfj1s8XwkR8swhQPbW1ChKD+p33e7lqmJfYate8NyO59UR3EVr9uIFbOeyZNvgrUcZan0EvokSgVB6dJUZCSRth7C/wGQdkIprRix0ktgS1mEIUU0LtQmi4Sh75FItpTU1crB98UYSsHmqbroNu1cD/BwHK/OPCLKLRS/SYjMQ/GJ0AZDi+mynJZWrsXAn2OaU8pWS/TrXgqGibIrQ1JzqnO8c8GBnM0iySQhlOryPOjLCdiynO2GjMs7BxTal6RKe7zWfQ5c1miFdIsBl4tDMxonK6JVpUQukVnLu7Yho57s8PUMV12us3uHf3Q7FNdPx9UkhV5c6KSaTjjpKxFR9ND1E1vx+Xe12NralAUsbwlg/08Kze48LCXc5VN5OD/we3WfdyZ7/fmZyxVSo9We9umsiygtKJQbrLsmDRFPz1kXnlX/ctHn3r5zhF4Fi3R+nmPFaWFXJbPhECpEjAF4TZVgSl4uLNHcvT5Pdi1qsgFEaK3FbjSaQHD5LLHu1FZoW98AQBS4SLkExuq2jXK8cWAHKvNRyVuThOA/0qdcB7wcO0CcTcpM1lYVu1HHMn7S8U3AlenrnUusNpSGd3csCR74Bs4g7lA0MebTdcWghG4eEuDXmFtBDl3axqMTJhJRsBZYyIoy5JYqqpmgo7X3FiYr65PdwBHG4pSULRtpwkrdoiyLVLd+3B5keln1VRhQM3oMGTecSPdbjFyewIZbxsfRhbc+kCRUlCrHXxFcVeXbiSOAMsQl0j9MLyycoSzKS+0wQBIspjM7JJun/5NQrMyyiBl9alcW1x99b8/ECy1chPCG7NRi24zP6kAGx4+d6wXedlzH0BqKb1vcH10U2hY8kYZmSCputekJqGJ7pnylvns4LmCoYYCniyS8MXTrlylJM5TLzYrC5OSFQr/s4gfix83Ngff1XFatxI4uUFNzzUUtzEqO9tRXPG4MccuyoKVc+qcZXTPeNE0TC05+BE/mDE+TWYfIV7nFbanuCKoyV9luqlTL9JDifdXzlUIItl98VohB8+E/XlOMo2qJFd0AqD85sexOUvNTREXAD+XJ8SvNfsXcLfTJ0dtcbmtWVxv5qkzJkAbgYhAKUZP/QtXmoK7iZYgmJm3UsuR7oJkgFW0jrmf2hSFtoKAtXdy/7FRich1A6deqcbqJQ614w0QfO55mKQ3kcOJwADzMKl5yEWDQ5LA2SiW4GgunHtgFXj0CNaxY5jxMCCX5MXiXkyuHYAgysKcPTIx3T5n6aCX8imDJg8mq82fzP9FE4bWrx3980N21NcEnIbX74Z8lkpEIpLxkm3ohyDkpLAqNLQsRoFsbudXSr4x6Bw/zfsFud7MzjxsPfqxv4ALGyaAU5Y5qj7JR1gtVFuchyPa/fE7BsXHxNyoavK4hxP0LMRG7z55WAElnHQbrayD3NnM3REghouieznTUHgMNc63prUOaZKgYLsQ2v82brZLALu//ekF7EGvPdtTMqaoLoS0P7hbIsMXyDw0Oj8or56Vp5v8ODIwDix4wQq+SvzELpSwKaqruJlbmjBFX2psIQ3gD3GMdOiGtwqYpqcXvv1cfCrM861/FwwH19HlFl7X8jLFe6cqAViN0PGEj5qdpUTSoFl3bOCbE9CndcZHAeC9AVxk/xA6p1MJxiJJL9WygzT3u9LYeVa2RTEQoxT+bqJUbVGha/+/bEdqUchwe8FUpNaeWvp1MW2mfrr6K2x5kCpqWj/M5oUdXOfsz8Gb7TJ3w82UT47BKJCnP6MNHVKtyaBdCe0S7jjL1bGU14rKRttVkhaNrg24KnNVYiySBOpihvK/Cb6YUMRfmpvBlNe/HL5UdbQ8nAHI2XBex8qXU9i9EgjjUWLtnUExMlaDA0Gy5Pcoz9QBh8L19luGcGMWoA//lqgdYEFeJQTmZ2Mv06lKIwkROj34ePe0BaiVD+ax9FCpRYXBzLzI4yhGp/Arm+FPWKoNBmftDr8M+q8F+sotOJz+ymxvTJFpk+1vNul2N4LRXL7/MS4uaqWl2OR9mj+FAD+kATpYOdI5vcXYijE2AoFVldHN5iZt2v2hvDhURnd/d2fwYQyYFVsL5J74igH4fyNIPeJiFP+wPj1ZUL2mGEJYk3e8RwFG5/P8KtM13wZAy11Y8Qe9SE3d21+kCcIoXZ4LTfrhFj2VQzVZ9NiUPgEeE1EHyPVGU+9w7Ao5yd1th3Rfb3j5uWYARUjW5RBLeMZGhaqdM6dsVHa0qX0r4lxy7b0uXEcJA+R9WknDttQBxWB2rFMWtAGz0hP6cgloQlpXZusTtXQtCY92lmFGc3VaDT5qQidhWZkftQIdcUpebyUppK9V+MW9pxossnd5Nxl4S4zgjMhUQ65xHGKa3jk81k3K7IeL7j8WbVkU6J9DIBkKzrmjDBIX+Z/d31hPBA0HsoDWuaYIYBe4VTCNOu1hQiR/YwThimO0U5HUiJXDwWNzL8SCfyuLSB8mlUaysPvcOIzeGSuU9uHGJRIv/MlEHVMjZtH9vwlaslHvnZT4ZB3nlA0I1PKy0uXiWqcTLdqOLRXsaRNjjZBYEHMBeOE+qcFschPt/CrttrGCIqYx0VL6ziEhhFBIKcd4jHA/hP+2+lXHKGfVBf6xsqjwu2LHryCuVNpcMTCPgthC0yzkcDqW8QQlYeTjvgwLVAxk2vTDbdYxq+XfIceUmXDJjhRa0HTczNLxwlKrfpOKo4vLvn+LY/lWMp1z12vMAwPS22WiLETsZldsdFFy1/y+YdwU84U04GRIia9wzj6HQg1Rbj9dMfviR6daG/7TTGw1jGqyPFPUfW5Y5R6XBTb3mBJn2ZWPKlK2N0Bo6lbWjxecRjYnD32Al+oJa8mU3QV3le5qe2Gvh57nq6SZlGg6gFVp6xflhY2GNJVdNkE6vww2CVlEMoLXzrfJAEJmLpxmZeKStr6YWAPNnrCc+ujGtJw6PgBUzSZzA47x/moG0+ZFAWyDVxT17Uc9SdsLJ+E064xRypeiI1iK8oqGblFfFoRR6szAu4ChFbxnzlFTqKY8G82MYPe3jskeI7kd8/zFm8mlQTzxlxjGonNarmWHKA+dsS1VnqziTBV754H3oFLgIuza/ar0mjsVTLo2Re4dKy9UrlaVgz+8H8cWGBu45it2ep6m7FDroaT5ZuylVGwF/IltzSg8ojxxqp92G+XwD/z+1KnSZL7PKeQaUuSWvih3a+8b1RkyGupOKOFOrA/K/LyIU5uyCfhQmTVDxZUbHr2vFRqne6SuY3aKZjKSkZhkVT4qGhuoXrcxQamAHLB7MSLgWbsRWgeefR5HjVztXjTMT3XJpvXdw966BXBwfpvhob1ejCvJGnpIbWftVR87rRJfSlD3tvBnQEFzV9Qz9C5HZUeMemxpUKWG5ht31tM3w6trgszwe4nZLO9owLfRosagzzMvnJfEKFng4VO+4tt9L/P/7mvGQzzFnZ/fLCEBESytWPFgh4e2OvHq/HaY/aDivYyyVgFONHZbk22VkMaTtQoBkDEz2GW8Bee2l3KNO5H2umT2prtcfcHt8zZNogP2+VH3XHXm0nDO9eCcVsCFlDk5KbrTtI9vl3z+2SHWIqHeoYpiSGs5Jxo/RNBNUVf7ihCAF0EhRD7CuapyZnITkKRtTH669n6vK92Jgm5kLo40dfuRUdJjPZyUafZVRQM69VPGoImGFDCvr55A9XtslK6e+o9+UI5mvxbW1W8mW2wHb2g5pW0/zccZAaZotvEp076o2XXbZ3lfJHdNAyLANLUs1R99+kW1BpPLMl1p1DPA+PHUfADdX22GNpuz+1FIuDL2gWPe6F+quWD7VrAtYjWNeaKD8WOtYw08hJXs0Z/H6LcdgGRLgdTHMVKb2tHZO195RPd1rzE0ZjoQrDoKqIjBozjatKwcE3L5CzrbeifF1hHONCdOyVYd4ZpO6NMFKy2YpCASUee36T5NCSHvkq+rL0bCpEAF/WRgmwFZ9hdHjdXFoeU7XGL9wIRkJ3VisVaoP/PgRkXnFhETs2Hf7HWiA2UhhtTSgbEt7Ib7p6dC0H/9sXIhI9ErtM3MUIg1ZfOkwNGfkquUMyVo0KD0hJ9x20QELxyUTiz+iGqGpS9Wd6LNSXz0U6ZrK3vBx/ES+A0jRdccmHr+6rRDVfqTdYTU8rfcWJ0JYQqbqu/qdYS+Hqgj9kofWCWJ+mA2aiZJttUvhqFCC7ym1CRjeaCk3uYmeRXrzrQIuZREDF2ePEieDJr77rL34gshTltMK2Q7NgLY1E9uI07B+QDY7EKBTkC6+lL/ccFLfnm4KYk+woBualhcgYN4mmx4sCYWpUiQwxtXo0ktNLu6/Mp2EyDWGBVKiPnxSOMwWYDmBLw3lOUMSheq0qIg4he+F4t7Pd8zH671DMnKY/dj5bLsjFMOFsHMZa0En0vYYbfALvxT2rBmKNPXJZ2523KoIQLfe7WWaNZ0rxRa/xMMT6TabN763xha1+JD/+gy+g6Zr10M7aaqpI59Mmb1bn6mlpbmPKWZEMNSfNS9tCjNPPlsEKUzWaer9AKpjX+vQMAMvfTqDTFceA632zGisvNXsbDRywNa3Umw4FTn1MbAeNdzi1YM11csfHH4ZxFH6jwhFXaUBxIUSRu+XNOYxdvbDtgsBL8z6twOj2IkbbqgRf5EDrk7UABowAzQrS6Oy+krSz3dGVUhZKlKaaVuFFpI/f7jMyGEwNGxyq7ayF1DKppYEIRwmp4MSTxtXY0HkxWXmriHV+IHHgfXGC6k9+B8NZ8fOcacaJc7Ym1ymcbe2mEJUQ9k8MCPoUWrpXfKj10MK06o8kHcF8drjfovD50ENVvNPUstnocu47dKRMbuwPT518yMVC4q+pSjnA/0rtuq5U2HDZ/+o0f2yfKp23/3XBaGyUue+RTJYa/UjSyvEFJeE70amz4eVOZ7QieLQoqAJOemhFyWxfwz0YxDUSDm0AGHKTPx504w24Eq03OnbF2gca7tDnh4OK67mYB+r2b8ZmRaXu/qkSjA39rymyVw7yHNqokN0l+nnoVwUC8xzj9Atv1FyyuzWOWRDTmXL2WSfZWrbMLoVDSdoxEC730RYT7vf6QQVgiH9JrKMa5PLIvrkPWmLyWMspPSb75Z06TRImMkEuMvoC6q13sS+N1BSRiQ8IPwaGkZVx0iXLRvk1Guus6G1cU3hKr/DtO+3DWXFV96Y7/h/mEMMc8lvWg5avOfiRVdu7HvUwCKfCccH0duQSkteQW20snZJ5xRoc/ehOVElOH9VFKlEQnG+WKcqqfclELuD1pb5eDKz5YucS1w75CX5Jc+rVnsU7a3/9xqUCS0s0GkAdp7g2H6gg+eHd0J2gVl6EtH6z+kfrVLDVhJd1DSO+GWBQesnOHZkZE5a50bdoRepmIymaKi/7N2LBwqbXmnu364Uzi8HRYe5+eXsc+5xvLEjJRwnHjdJa9vpAKgrQGmuvHYW7vzBPVXev4ErMyInnjp1aJe6LZJ4DfciwG4gxzEI7KfUSjMkJ7DSDFupsNjXxZGVWX5luc4j27zLYnruGAqFORlLj5eedT3TmL2yU7YqOIa2YBiWAH2l9SEI+IQbPHpCWq2K0/dlLOZRERDHe0l3gRmZjZE+1rrF6B7rQ9Wzd2kmzdCOLN4mN4mi3CvWTE4Tq5+O2vdYn1p4OTjMiWdes5L/F3ryy6YOTth7LaMAigHbTjXTKrLeTDVcPlPRxmXqKbYiwMksTF4h7e3N7HEa/tUDtUYgrfrXPc1Ns3kfn+jthr7z5aKMHzhdsw/jT+tGu/KHhvB1EB1KMZAEuJOkXj5W/E2Jeh6G9XorVqtgOgJo9pBv0stpHb4M+9JcFyr6C0abXLwix7snP5iD6dC6/gxFpO8EuEDIQKFJ7T1eFWTxMgu3yJr9YzHsVeGlidnr1xNNfbWe8NuHMWIYPo0xbMT5npYCrkgTW8D4oW2N4C195rR3Jo1uzGVOx+6U+fuaGhoMBoo+geEdnGwgs6b4rW+Xn2CYgjlXFQsAwYRsKWVaC8vgrLr/oI9PnZIa1mSgqdPrLPR91xWsx/XWgxJQjp2o2oPGJGLLnRxgan6GBxsPg3+XLa1G3oWqYDTM2vdHHpC0a9NtYrJknyV6J+BWQL12Ta1mnRmorrwZ8n69IZTfYbySyOaDmv7eOqbiPM4v7yufwHydv/2s3BbXZCFShHtpFIy1axm54xOrd65R3yv2oU/wyE1DkueIZqcSMybmNtA1TbJnV1wzbVyaIPh5QV17V88zCVH5qVWwjt7vDp0qO3Uw98vYPOt7MTMfVvIYA0vvNU5T68P6gASvof7Le39cdbVakzTaBEOcWIi2xseDSl+iV1LOBKFMUMpLTwee7ATwAgvfoDORIC2msxRDmOOhyjRO5HYEKc7JKUrYp8YM0K68jl6rIIQuiMC5G5Q0H852t6xwdaDteNktnZuWkV4P/ji8strC+1PZijwuSZA6eyLSPowSfhwAmtMNQWZC1GASSWKMmqm3t7X4VAqTpYRiHf5YeAUbR7duY2/8bRGdctYJEvAyPmo6vXZnAEm6uIdNaiSZ288P/eP/3/OBbBAJozxBMLuEj4yvaqgr3Rm66u61Bcxu202OZ3WV2btPAXEBqzReXZbB+VcuC02YtIwLNNurKMlevEedUdk1yejmEleXXMGFu1cLAqI+6WS/Yf51Q6nx5UOIvgo6huZiJnh05rj0hlv0cldAMVLltSs6W229X8Rgx7y1Q2HwY0KUOlNyqD9XIALc/fHxD3EEw+xx4zzPJhQzc/OmVHvng2nTXu7mJxx4J9kSfR5kTcbmY9HZylfB9QojFrSsn3+uFASPfPdyDuZIK3eu68iZjjLc/+SKgL7vE5hkQXc2lNuon/K75mXgSAONcVzD5UcKbhqtm/gUclz9euwCbcTqsT/yfgthLh/ms6NMHKx2Lvj9E9Y788BrvPttUbYCLY/99lbUEjAcExq1UCtYy0zs7lQKlXXHJkE5KIwD0dFjiHrB70zF9KS9qBH7BYmsEYbngJCKm49HtYkK0+hv9oHA+qrVs+bxs5VsA0rZo65+LCi0GRtgtN3bEhMkmJGjvuKI7ptGC7sun1ZrvnDZj9uxBLokA/T6deFyacO5krgVgkA4T0RHiuRiwYztBQRW7CyuOgwgwnGoWj1lvJkCzbjSEguaYdFnQSVQFy2ZxYPzh+aNdn19l1Nje2rXK0QxhXR17XEJKIkT2n9U9tvDe7Fe4OOjlhN00VcrHfa+mLdrEqEI1sMovBE5y/qGb/XrvBBb5FYcqQ5nPRaQEgNUJTH7b1w+a4Lyy+rIoeBohFLvirrjy+5EYNeXagC48HdQDgdgfyVhQ7MNHtJRLWivH9IKBc177dqbvExfZc60GanzIPs4BTVvDaueCwt3BUAhqXIYEEGUjz99Yrp2Y4Iky/CZKT70d7bZrcWAZVFSnw7WRs4oWizzSP+Tr5r9GhmSQfqDzfyzQ1a2QWDWyUN42azwvUxdvga/aIYxlxeD67CwOEBuy/gwYElO9csRmyqUyC3Kw6i8/KzQQ90jafVqmT+CHOQdu2mCsvKtKopvJvaqKXEInqmmpb1fZd6VNoEbik271Rt917F8+HDpq/VWWt4lVZNjC6AFkiGcoRI1jVdzVGxcXmAg8CIk6m/66d7SoLXQuG9ABdKmk3wXEswMWxKz1ewn3qjW+7W6E7/aViIq6PmWW7IAYv1yLkZeo5OZ6gU/mLmCv1k0iSEMBR8Q7uFp2BbEOt+Q+KNY+ORDDJ6V+SZ5htSvXxoszkryC5BYNyPIIj+jpjNDPP/8XwkBM8qt4mj24d8xzv7faAez8DEUW4wtJRvV96gTiDSp6yQQChfUe37bxFSrHyjqOLWbkSeYO2mnHNJIIjOaCmEetuHYXniiR7ga43EdJ2X0rJElU6G7h5dfQl+gEAGCMMJ1G2spFMS2Qb3msORK3MzegnjJn8vv+m02U827J0xokmt7ZxPfOM+DP1SAQv0chNp5gqwhHfZtPbI67xipYJpn4v91bnkmNU55DTGCQ1XfFXqdLPj22az1Sku8IkWDmlOF/C3KQzG97qKWNqPU91dCD7ioOoO9E7aKiFpx3NkaKgCPItboT5EESpenm0nHQRdTNzc/4k2jfuF1+vhg92ArlR7HGGdehBGd+bnjsbTgFuqlc4Chh0BOkS0ptKhCGpYO+XMucvyww+UC+3kyJnB/nUHTB06G3RxHwM1qQ20x7BQQg5diEx3UJcK3B2KRtb51ZYOoFGwvr9QrCvVcjcmXXTpvBwwc3lFNrEtbGgUegbAOfmTrmmgV9G6GsQ+mZKj8CGJZbhhCyED3pG3Q0rV7gQnf71IIo0GJ0SvEnwI8y5SaYZ68/BuFXraKBQeafsTrj8yEVEn3jiM3KuaQVNMy/5vvdn9jiH2sq6cDasMhtK7yghkW0WGnyYGEUe4OG/+OSvWIn6gXu0eNwMxVH2/IgKhBaXBadvdpH3Qw3cUCOuBi8uNDZAl5oS44sM9/lw/cWTL9oOkq09tUSwE0NaX1awxF/qMr4bTM12xluWp7fu3gP8HhDSnjei9IS8KjaWt4WmB5f0GCd1A1pwxHXbyzQtAHdFhhwVYYatBStnWxsetfpSQ/aegn/lAUqhmrUu6wZWmrB7NkVxGU3kQTWH7XGAz2pmuRadx7YXG6YbRE9wKi+BNssTu74RaZ5U4tpOfrfUPDuCPghTyR3Adt+1I+W+MIKGLo7I4Xli3RL1UmMf6Dvn6HIp7RKkQieEt1h3MNwolfMXZL6puJ9hmkwZ6XHpNV+4htUVd89UsI11/6uobwdLVqrfg+dvrB7XuGSbZ6b4xsxjnujoSkgwTVHzb6EG2EeD8WTrNsyIk7Pxr8wta5sUV7qVU33sH8BGxCLeG2pZsSvlSSYKAD18BUHlxwRv/B5j49FO96vPwx+B1oTfkDamULmummVMx0ZDg7PJld0SkJar+2lXFXP4J/qYUSV8o39yRQKXuZ1PktypM7eVM6E3z0LK2DOiXahZsgvhltiTBt/PbK+nAQUiQmHRdOkIMfNuWl6UXWO+eN6YLUNGk0L67p8LVyX1LEnDLa1BnEU0R++hfarLqcSLnQtLzdPMJ6g4bzWadO207ak7JFB4WgKlgMG6m+W4hZPHiqO3CtXUPpIXgsKpPWO5XXK01uJtvVSEqsPXnnCradHjWXcFGerJvqNn2w+XVTZmneFYu1l+14PykWw3UOwwiWCXl0yuziAzUKYtr0taEGu40+09dan6TN7mqMlmd70K+1rMwmLHpAwNNj3XmwhaViOTNm+zfkPPoNSmQDhtSWCe16NGLAPyJVfYCEsRhMggrhsbbojZKOL/vbTygv+1Dp2z3Q9e7ELNozsGTJQU1d1zEVjibdD3f7K3/8sW1Xvl7pslxvfyQzpqN9+7hwHp4u05Mbzfzy9s1rfZqAw/Q8U/UH/4IdWurCjvL3KVaUJaQYJ61qM2lnR5OMSTv1O0y82ydAXDl68xJVnfKIXpaz596lkZvI+nIStLDk2kNwcflPawfLh6Pv0FrYmYmh/m1LMEVxQWfHclR5nWVzJdl37lXpsMaWRINu33u6JtW3er34PETjTx0795my1ZVIPH6yBvTo0y24JEHn3dgIYbZCtelGsHV40H8CAe/cvzVTfaQIpAp8Qq/KXaJhA6EPd8JSXxU7FkQIVDVXpJ08Qxb4Nc96haO7TGliDFhY3G9r9MidDigHvjrWv2CPUc4racfMUmYod/ujUFx0xpovnFTTJRknftBWLgynzinTK+oeBsGnt+2UE2JgEflxT8Sdq017rQcNCOj3Ix/VpDu5G8xG0vcjM+/g0O7tZfddxX976B+D7UzHpQfZHsrkBH2l2dgGakklKIOqRtJR/6PmuPJ8jSEDOeL4DmB31/7d1GJK76wOWu85MlmuXCVoYvn8Zs0cKPxdA06pw//riQaa2g7jkfMTU3CkbREb7PdcolPBfQ6xLZoEME6STQcfM0RJWnDYjG/HsVcpv/1cWzP+S2KgoFZz80UOLjpKaDt2MLibjqZncloD3WA/kxCqXpUSO+cbJBOazAO8CsZda3x4MBvC9RxHdD+jrX/tUyfJBvhwtTUVX7ZmvkkEsr52RrTM2+W5k3ZDYX8x3JcpSSr8Pil0gEpaQxiMQX21BJAooDvfeO9ASvlxx8QWMzAPNsTUELwBYbbydP5YeEysdXVHLOAH7Gl7JcitC1GjNJLncAFgxyRXlWupyfJxIBCxCDdCUS1r1IHrF09BZZ3TSDyLlO5phmtbshBgG54lJoGxL2lrGcyBW/hbrwg11dJlUM1vDN3XVr/l95WpufD0umoUTx6/2mwgbl48Kl+V05y6V4Yy8VH8IN3+v0PG/Pe62QsLnvKOCgZvDP9E8+0ZZ9xH3Uqus2K0HTzeVo6x1uGk+/yubQU7Sprp0yolR0OuVLgk6a4E3/s/90ctedDMf9rWwiEH4yxhGRuxKH7sWKNezCtoHTbCa8Zl3kIY1G2ExqwSXQ5JQbMcq3QlRAgxwaHacXX/bUUOVWygh3QLkTmwkGFzm+DJgS4DRUtOpnRs9oPFUNRh6/7lVBePeRYz8chAVU1lH4POnnXKCVtYXnyuW+V9Jfb91Hs/M1hEFthvKQujWHU7f87SH5diTFki/z3r7FCXTYBwVrC0d5+NXbllyjL1I0W9SRiEoI91gxAmXlyKa+cFdEGcHKR/M7vzC4ZsUuvp96TNPSpN7tW6UZT+LV+pxERX36lUPy74L2he3ACK+dnkO+4EVNkcZhb5+kmp/xcgX08S6HphSpMY8mpfHExG7Ougpv56+rvBzuF7cYgV4VdOAWhstcdSpUljmbTAaWu6tpLn/uNbvaWjMJMwT1kkJ0qnNmF/py1vuvS3fGx1ufK6QtNH4VMyQfuWSvcD1fHmim4U3tpTMn8LGiafK+5Wex4uymtWG+CPcfPTU+WL/R35r9qvVTFLx5hOyEKSqaqmw4lGHOIWK2AHWn88g8zKWQyrfoPctR+fuR2EGlPUdH4kcc457KHdqnV2fqriO9K6ZUiOHNS5nCZ3afxUPnlUDyGHpfycTRfYVBw0+9L3CLL7BfdMrUQG0R60+sZwdWA97N7aQvKvCm4wFU7/Lr5Ual4vPX3I8vArJ3vfApR9hGMfXZptdD8Q7Avyr7MZ0bftQ+Qv9RUhGwFFsjN1yePk6Y848QhaAWxLKQf/ok5C3ng0/ygGZ5vwyRbYQ2gtoyJyKUY05I0jf09K0UBtDpumIesyXpg7hi8H18QUvZjYB77kliIp/7oBf5YructXf7/bMN56jaTKDVL9jcNCj0gJbdVBsvmrmT46ELR8e2F7ZGSzxlH4KjqsGIn2R66uSlSA84r6RSKU8J2Bou/vCx5xjx/C2lB0dWdwDFw9oIQns35waUMZ1hUwVrD7f6rlHL393Vobr+7V9WfUd5lXWw9GaYC3L1qUglV1pfqy/sacDYegHoKb1MY/8JGG44xGHNCqVEwsxgj4kB/PoqyHJNYbEXPDkn2ODRxPi8RlIP77w+6iOCXZoM30ytOHyD5tyJk+2zF+0jGhIcBg7UnUz2Hz2hNZSr67BVINZ+KqCx2wiTtY2oGE27OLbnXiZ+68E7btnS6d0fUTtm+pQn1xY6q6wdN7JDG4O8LKDXGonfaGp6WQdwtTmh5tlYhGKL2EH4KWI3AIxmxxBdaG9oOikMuxgBesBdSwXM5c9LpHRDhhEC7wd/18LtHLFe4PIzAGnKrcWnvaabN60fJTpDgjG7iP1tkf9CBZN9LFo6hR8Ge6x5AQjXQx5fb1/CqkOTgVOJdDCwaGliZ4Onyyo5BattSh4aDrFUtmwhACZACRsfyIpj4pio4hhW1XQZxYgdk9ofF547EK4ik/x/Jbj/w1j4bBrTqeWySIxowzLXx7viBYl4qzEs/Rsx4nO5aU1EJYE4ntS/UPYekjoQl1tkbY0FElk8WzNSUOIqq+pEAaboEmLk1rvyenqhHu9RoLT7jnCxhAXJ2DO14Y/yHt1rGyC6sXVi6zPOz8o8XZ1LQfaKH1ljvVLlDKuLeGlYZB6dp4uIhUBfbnrkLDHi7K2O4IUlRkdtFUD82Xum0y8E0hkNv1OjWBUcBy8wpoImqOvYMuxRBGKmVpTNYrx/Xe71JHjkYzHFp1q+nLbMDyexUjc14vX/AhnbS+wkCxACUfOKblrDPW/rTJQalXbvsm79mX3wme4jhyPC4wi8gBX4GsyJLvd2ZdcmB0REbMA6jOZwXULADV3QPDAOPf0phA862csZs5AFdACltLuxBNwq5T9KfXv34QGJ0PYG5MpvNFdmbSAP9RkGQ2Cxs3aZ4Qc9/VZYVNtftWOGoTdwENmMzxLpvCd/z5I9U3t1T59XnaXpnJLAN4AhT3W1D1HvA7gMcGbXgLDAnkiGwcsegXmnuGzmv8jqS/A+NNS40cQG3LxzqShOXujFbuaKbkEw4AsUuxt4MctBertj/iAu+ILyYCf/I0mKl0zyrZrDidu09y3MgUWifUyelEL/19+1+7VAXBHS3IqJ9IL6WGKFca6qGWNFuR/iiGVbgrZULFUyzY0y8lImPVrBC475KGELwdUJgnHBpwcq5X6VR6xC9UPZ6/eQOC5x6kyabyp2ogkG714yE6vN4sJllbW0391ygpDpwKcsbIgMjwscRUC56TXxGO0V63S/bHfF5yI6JeALABpWkTKVFFQcnBjmZTEE2d8aB724JpOf/HBqGdnjBA5ViTOnAspI/Jj41r4htdqNqFaOKM4LYeZm2PRfmov+k8G0djUiZLPqfjch/jmCMJp25JlW/bj2HznjZSlLFlAhsd4/6Qy6pLUKiuIBnUAFYFptQSgFIYvllt/qqbMgJuxtkws4Z3CLdzp9iVFMjN07ZgP0dlnC6m0fGGAvaz+hqk0K8iECFOnNyMbo1zp/NBsZWxlGHIBLt4VW6YM5MgNFkp+g37g5SQDaKEObvhLZAk6Xt24eyh7S+9e8EtVxEoBGTyK7FklEkXLTIb03nn4+IS3UOAx6sV8oM1j2YpKfcYC72lmRqYfgadAHl/lxil6XSzO7UUJ1AAWkQw71LkMjVmqA0lofL057YVIn8PONgW6a6A5DUnv67wz++iCMRXnO42jQNhBdmyDCSHErJMM1VOoSCW9s7EhhvOAVOOtzyGFb3rmq7sBUQ8d2wBuXURRHwI/GihJeaUtRl+33LxbslD2WdkMAwzdyKzv2yvwLupQcfCcw/hoisjaYZues7c6mdqIzZfOhPoMQ3S5SIOJ02nkJxDFz9+f75wkEBsM/hVk3oVnGxOgWqE+HDIBLUbUketnJGp5V1+hohZjp+a9v5ScpnN/D8sCL6kGquschMsKPh3XOeZZl6YpKPT3YJC3q9GOYN31rwP3gxvcoEzQq4fggg+E3VjNG/uQFIOUk72Q3kDurOCpmff6jIxCCGVd1ymz4UyK06yexyiJ+efc5Yz3+u6+xEazeS1zgVbd5MOBL019wy9pMda8L0oh9gHWD+PvXyB6mcStbHGUvHrpeBxupmwekJU94Px17fqLW0cmVk9bg1TfiVudNRBwoNDPb5dDVpJR8Dpfa1Lzpfdwb7bAFWXWoxMKGmIw9qFTOlp51vZphLfLuIxYXk0UKlAKPer+KtQJK/52FbsGMShPBu6BpIMfkNhHOl+3CKpHyqi22v7l+sZJSowJAf1wWnIaz2EY8qlt+X48GapLkCxZweyjLBhBOf443vXTwzW6jtFUfCblu05RrqHjsKbzCAueP/12Ss0otHE90VoX9KEkbx1P2WuvbrtITuA/tU8kUL7m8ODtgR4xOASOSZfiPlfv/K4E3/Yp5vh1nDD0T33dYquaJKTIsON674zBB2nsIJhQyDGf1pMnSvxaRIIRxVstWOcuOQLfW7cL9pBs5I8r7pOylTzzqEU9uv6RMh1HxmJ6KoiPaHhMW7yfp6IbK5CENQki14N5SviQhs/mVksx6q6Ak3/JkGIfz4UAN4Nr13C3ZGodyr4ww3WNcfBBiD+gtFtVXrtDyZqADF58W1jmqNjMs50KRUkR8yoRgHNxjLpi77BTwc8WTzozfPA+9I0vzxY2Sa7lz2s35rWCvvKW5mttiJhBvVumJLRBnXtij2FYGaVDmFA8VjH4Q18vWwxsD8wT9/p3LE0u325/E7c0JfmYKPIB42VdjXlbMKiKLFPJjktu7V407PaQVyifb04j6qlypgLk5uwzvUkVKpb6bXIMzmUwPs9OJFAVRDLjDj+SUgcQTaa9I7r+EvKNtuS7miNKU+/tNrdr49EpxdC+5d+OVHMwdwi3PcsV1acjpx2nglWnarOWNmZKUjqDR2fUMgC5Zb0GjAD/GxxqMLrtGntHC35uP5qS0jVeI2ugWvJd33Tuoy4ldKE1XZ6ngqa3MwNnkftB0k+xGNwsZFFKSI/JK9lOe1YMmQvHbqiK+WLduCjoNyWOgPC91R0bEYvcm5VUnMmec9C/eq9Gx85flj8fqKzoo/N7c+fcctIt7gpjLHwb9jyWsECHuqu3C7cR+YMOFggRB2KDFjerSICdza09l2mLL2K4khdNrPKkc9LE3ieqpbuDxJP8CRJgYtN/75I8MrtNg2VdJNyntTOrz2k5Sh3Nxs61JNkKylxa0x38b4hCmunLsgngr+2lpmJu3elzW3tvc9CCsC8BKgFoQz1vqs/HSRZ/pJiPK9MgIFWnGPIP3yWcRkNMulnlPm4gxWm0vL32VJ0ZPFCH+SeYHLBS2ZDGd6eL16KZIa008W55fArcssRfJcoFHBIvCfIUisUCFPpUHw1Ksux1QRx45r8ExaVdXKdCwQyen524NvhlAY8hAPaqMJUjNMPtk+Cu1pcRBo/ZQrKp82U3SmPkQLPVVaD5xSFBfIXsyEQzhEtGAaWU92MO/cijNBK8HbuQ6B4Gv8YuSrFwoP6Ht8poSpPj1KU4hrFNhnT6S86kJL7rG16GV9UJajQc5FrXaPtMvuZVsNVmdoGLRYjUnex+hJSudDVMwxfO7o8XegQAl1XKDzp/oS40gbKvl10QDlCKMoGgQeQa43N0ICkOhEOCMMMGdu52bfs103CrdyDnt3x2R6EqIdgBmV3/nLnXNBMulUaW1xqsZ/TSdYsheG/vmq+yjw0jjbZzdIYAdmjDomLooULQWViKf3H4gVPAiJphu6hoDL1TnUYnedYc8NeNSst1AK7/HHzNwIKxNtgo8PgQj2MpFculbZj27dym+8PuxpajotI2VVD2L10KqT9/3onPqhnz/YqzPTpsb9MZFrWZ4O0aNideyyAwTn8qtTBqe9Omde7mCjOzhCBkOCZprpYnve9nIdn+0bOEUmvjn63GBG9zPPHrndvrsfh5Xlel8Tn0mKWdwMJ4qmOtUwa0fLTK3opZfWTPQI65ife63KsifMqY1hE92SGg5OWs8JjtIk8xJVcx8cvEGVqV365VKdX4TKCPqOs65kEKyUGjbD9I5EjycXavTBKUAoVJwa7BAD6tJGvs1toj9YfRLWs/mgdhL8RgcmAn0oDagkn5XBKHDSqbiJ7FfCwbaXFOfqkd71fooG21B4gdLgq1GwYIFXNmJzGFcJQbxnrAUCRHQvrZQjf/Q7zgVo9Ut3J/eKT45J2Nrr6LerhJudj87946f3A+AaLtNj5aCPCFAG4RQ/KA58ZPcZaQmvBxLBMrcVgaDNQgT7ncPdmzQsJBItoRa595JR8+yt7Xcd77AQGQ3plcgKJeGTTIqXPHEAcZu4UhbXQ8YlIe9yBodRRm2/aP3vILdlzv7f2UXD3c61N5/CMmsTrNqlTIxTCbKHRqh8jSSWsjw3nEHb5Cyld8OjLWV1HZuwYVDyfPqtOZhRUnhlwAnF0mn7aWgBHGPIi5fdrhH737YjIQnrYxpGdvaOL44g4F6AW9nlnwSuw8V9lNNPBrZGIbNaXzQDaf0uDR2XaGvJ/2EMHscb5lstihMhhC7/baD7C6oc7LPtxUD1mzFX+NFvW8P8HHfNwvDBhscMZga595Qht0v+ifY3uygr69XK0El2HrmYdisGBhidhmLd4mv69T2V+PKBc2AxG1T3EteCbC7GgQr+5yoiiZkU3K2ftjfD1NqFSne+WsPw89gykIxVHL9z+IljoSZ00LJ4Ilb/jjp7Mkwe7KLEAMFnNvxVBa1L64aQqbqRn/COxHVY9YC0Xv8c3quW0wkp4H3ccpAzIZVt/jZeUdE/MJrQjYMWWh6GzWzFKfKJjchcdbKHx2MwUmNLZLaI5m5ZZmRbZPgFL/m3cHpCMQe7tZMeS55GgSkJavXl0VspwKOZiofoj3pEr1vktsEbQu+3QVb5if9MepDlscuUqz/L5TsIWX44W3w7ATrzZ9h+Q7x70Nf35y9uU/5Qz1Fvx4jk4menGoDV41hY+fW8s4vAS0JgSNoi7ZRnw/Ke42fBYPp0g0ykTePWbM3AbC4uHQSeGfWKuoVNFtOYW/5TEW2id19BR5ZIkdmKPc5qw4TiLsGNJXoBLf1D/HT8bakZhkkkQVoX/6zs+t2VrQRCg1R04f21INmyW4usNLgVK7a1e2JjO6mg9oZo+AuPL5xhnG8wJ/TS3HY+5GXRrv1xrs7JGZjMJVeOn0KgVPpHoWCqmnREdr8+dGwzJDg1iFLC7/Z2wNwr8V4qOJs0pKTuj3XtlmqOdExvyzvr0JWQ5eBTGsbLRfNtuD0uMUERW8d/4N2TDC2QqfNLXcE5J6WgXAj6pz/kQW27Y4ax1sunKuHpvtAMaDUN5a5MA4vwJbGshqJQClq9M3f6JAHvxe1H8gYL1m1hOSHynD4hJMP11LIkIfoEAxJ4LvLV8KB2bfBdkw1BTSVE5NfOd6zxyn6WBjq49okhQUmCctaQWJcINLMauHH3wZX4bX5UmQyldK9Usv13vNIWwMmASDRf8RHpWAba8mqJfJtjCGGx6sv6j6QEBNL1h4CxgKdPyU3CFTdUgs5cbP2jBiSBh3n4y26e2cEt26LpzlODJNwxmanHixJT8L6oCBW8K5Ce8NTZG9dqhIJfcrd/vXwxxr/dn7hbHzK29PlJbuwwy6jYzy+GAdYRzSZL3QPwxOGzJaojtG+iLA+hW4agUNrcAaamq2EjEOxRmj3a9m6fs3NqSaFgg2mFTdLaC1WlpFddqNcPDbfmWKTAX3ysUtTXbOuUgfPBlgroASO6QA8oIdzSIYOSRqySPlPqJEbkLw9bxMYeg9+UsZ0c9D/zNGbS6AaMxBOLroc/nrtLqmhGQUiKdjav2lXOSF+qGbu7B9Ng7PD0nqKhC8nQ2+qcB4wl5e2X5huJVWeFGrg4MzE1xYPY+r/g8H0DwhA39k7L0hWrLBAvKYH8QQgDYU5guxN3OGvl1bb2sMymGp0HdmmMgFjaxXJUNjj3kwlxRnaLebviEeZZJ5z/kCpCiprly7UgT6anYqBpOPSZgaTt6TU+uzeP73NJFRI+jvKlbLEKrGjV1Yqnl8bFWwcl5u6+e6lHM7nu+eyfCrGgYdKSWpQCpm4kOLJbnNGRw5TYEqjIZoz8lbAeJVhsMMGt647JnpF+Crbp+S+JMXs+xkJZkv7unx9mzUlR9HHbIV4IJ40blcTamm4/+FuAyx1kU57NmNVkLNo07kOSg2GdFyni5kk44QW8hsem4fc/hIdGp5Q2jByummsMh+c5Tv2dPQYuyA34lm0IXkzfauUhsN8XGCROxExKd+lQC34/4xL6kJ5Em4COdPAbH7a1Y4LqnFWW0NW3fdIjUvMKhZpGD1VejFNhld0VKoeksnyGg4StbvaNIE3PpFmorN6M2m7P80qgYZRsVzEB7L23a9D+0KbsqIX67yn7X7NzH6PhbrfpyVdnnUtdCLS1AFtQHSijrcXw7Oh/YPLR5c0/H69JpZzOKDV/yMBTNAu1IXmDGUz4uNKsr8sqI0q0D1plTWhOMwPfM15KmVfMiw3LeAkYDi6rsqpfWq57eROk6bETOygf5nS7PKYFfcAF25gt23zElJ1oxLIAMo88MmtE0yfL8T1mmK8PNUSvaWmMF6QlAt63ID/tf95eF+srwtNFRSVKbgwFle6eh6vvxAs/Kn9kWfGX3mw9IFgi3W6W6K/3NyGPS2FURTUvWyo3X1VCPKCqzPZVgvZsNkftcFhK6PoSy4TkJbgTwkTp+XhtDYXu4lSC219+7FS4HpEAcQkvf5diG2fCZzRbrnFHjUp5UxKmzDeWXDbpW03rPvBLAE/6Ab3l6sfhgzTBX9KVvUzxp0qoPkL0I7UV9FtyXeWkBL/Ng7LXTHzixeBnqmgE3JFtqN3iegE5hzy60pp8g5TcMZrCgn/RxbBQRIot9tsEu9wv2d9qC23DOkrypfAkNqCq4TXK+igiv3NyNQa8FE1mIyVlN6FmNlqkBKIOlb9N02enfQ0mvMLsfFeLpWgHOcd/O1Dyv/fF0Nz2aoJYqLLvd9j6r24CsDNQtlWJfo+7cSjmbub3sqMm6Q5tl/VM0f/aoBGAqSsP72meeVyXg/fGFTXvrQotlBF83hFOTEBUdepmzp31q1WcfKCZn+ZEuqGTx+cyL0LR8rw1Jpq93CDotiFTfZx4/ESoGkut8XVXevUM+s8Ir5TDN54T33JpIEfHFg3YRG3TaBmy8fow3CMyBNzKMkaU89I0ToZnzS/gAQVZmePSmEA0580wbZbqjKgYN7J7Q7WTpKwI1eGSowE2sO+ZtF5EFTRA7e4D2gXLjgIwbzoNWcxFsbo21+IaMgCgmjiYCCcyCqU2JjIRjoT8z5g3Uvgg0qQe2ylwyu8jBXjhiiPPLjiy7S0mwQ9RkC3zoWYnnL6poelPc2pdMnhrYVjh8b/Cg+vIK/2KBybf5TLNJxManj45+TuL+bKTKbl6Zo/MJv6w0oGxcYSMI7y655VDdarQiJ521DPFCRNX2OicSRDFmpR8+hXeLODC50fJk0pl811Sd1gCmaY3q6ltIp4e/PLEJat6i7HGp6DzhcUGKCaFB9ne5Y3A2vdorSfLIGbM999xnkKEq2y2Pp1Xr4jLZfhvJXyNIgWZSmkqhLKQVuGwoBC0ToeLakYzhMpck2M5Fuo/0gCzDxmZyP8FVN7wWcEFY7bB1lc0hV0z8jcEkPW6hKV698u9VrhSzOUS+ES9Zeii5CGIQJUFFRYSrbdML6Y7HjrbjEo7jZwCbSwuz+XdxUKDlPhWKqxI6kpxM3Sx4fav19dk+IhHOtRCwCUBGJcklS/FHxr57PYR0XCSH/hsy6HYOtbK4BVu1//YGMJKVkw0kzpO0nW/Zgi27wdFZefk090uU704DykjgRQI27lSPPwK7XefQmqHy7U+IM2mCzlu/CuXfL74ctShnoGq134UO6Z8EDlWZmKFEJloGNUNNJtbTy106FWL/sUY73GGDQrCcw0FLRFInprWRQ5FKMfdzqkLBrzXSwnIykoy3+PEHGrqxnVUNLDcktoSyotZpz8duY/WhsoeWAmgBGbySBi6eXlqJINUV+Brv8z0V0bz+LbtRMNOI6W0K1VgamAtA81aRfXnAFXvmDPSLxfuS5J5F1krQgDA8n7AeFVkEnUXy5IE3U3yQ07pqbdhfXbmt3qa41sUjrjz0euaedBKGMQRU0TuBBthR4MLottj1//uNy9Tj642+dhgxE3XmZ3DuPvZ5k3/LkjuFQDTHuEi5ew/RrkcHreC5KITaDWpZjUPhF7oRf3DqFq/fPqpZAkZg=
`pragma protect end_data_block
`pragma protect digest_block
61df3b47686faa6485fac1d93bb8986f21e16ecf554deada27673ab002835ce6
`pragma protect end_digest_block
`pragma protect end_protected
