`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 1079)
`pragma protect data_block
y3MhpOk+ZjPU9VxEwjenB/6gu5e8fSxQ0zos97V0bX1YMK4M4xDyTUzxgd32MGrWb6d/tbuX1v2rtyka5xdqp43s+04bWtidcrixZ2l9DoER9rq74tO6mjRUNxCces+jI6ZZXDK9CO4b13+EgHjNdo40RZoltvDsu4eJxkF4tQhQLLo38QbtFiX+hZE5xO2AYCEwzEJfgG25sy2Rh4kBtC/Qxcu2dkXK2gqVNcVbdI44pYOnJLC5HJW/qxR24qtrv3+sTJOgH3NhK4IkhdkEHw7YXmHq4twxuTM4piwz91mXABUyRMxSw3eQY4koIb3A6+he60AGp7PYoSJeXig1L9Pwnr7FuOUuJIfJtWpi0ZfsSWUObA2AXFiGP9kuXXPFu/fBgC7c777Pm6AGz8Er2kGoAxo37K1pFEikKokoX123Vq3nyWEIqQaqKJTTrWCQ1fdl2PulB6Moj2X5Ve4aQX60mFP7uUUVQbF5CGcE8miHMmR4HaFxW+KHBNIyj91brjQODSJkbxgCSpHoafvSIyFzalC6fyrKzC7BgFPLFSN4rm8RJeJTtCrie0iLGrx/IHauU0DYuoi7h41Ph9oJ8aIzm2RLkJsGZ9DPGa59c5ZRue3LNVxx97RWjYOEO/IE3EJAigJuXZR3fs3WH32WwPl4tehnikeyYfBorB/A9NtbqVOhn3t2qWOUoZpdtjTo9QOgRz0POiivlbLa5Kmavadm4gAeCJYzvJVo5npQQcSHNaSy0ffucoshDUJbipFtWjRIeWN98iyBsbxF7NtLxrt/5u+JNgfgiNCmXpsVqWw72S5KGW8A/FjGd/2Vxkk6hpUvhjQoMYFni5z2MDXrt3pXd1dVgdDToOGkUqiAA8JBHlKAtiJIZJaSV+EZINcF4skFIQn2SCjBVcUTgE+WqIRcm1rbZoX0kmHvvrtesyMXqVrFOxaMHouFBjASOiUY+IjJ++jHaGn4LqunXYinaZn2Vw6Aman0U0KfN/TsgIRNKF/GVw6S/Ux0viAZrwL/47LtXgFTCu3cUc4Cph33CfwVj0DqBAo8VDC+QtGJZhx6Hfi6QIxfvRfS6i24a70Ea8DZhYmcO71PxKQwExr5uQLq9FtmoezH4zyuNlK+WB0t35aLTD9AT0f53KA+gbXlfMK5LkuMthEd9fg/mBWWIfMwSM8ghx7yxlIGhx/yYJSYd2DincSXpSDK3i+pnyiCsHyly/Hgv5H9axd9xYjgGjPYhnmir4Tfl5h5U4nqIwPBNwx7+TlraELmKdqSF3BAXMRkOnEV5zfdij1yexsDXbViNYI8qy1W0NlSrgUz7NpHj37Dv2eLkLd1JMoWp1giF8i4IRl4qI2MSosXoOLyJ3nL0TNCQGUA692fhnnsSlsEn2idBflLRt2njJjdhHzSWkXwtDy7yq8uzI6bBdk0X1H/JMfUq3A4yBQTKGT+N/o=
`pragma protect end_data_block
`pragma protect digest_block
57035225f7caf6faa0682678da00f63b0f128b58a601c41eb30ab3b038551273
`pragma protect end_digest_block
`pragma protect end_protected
