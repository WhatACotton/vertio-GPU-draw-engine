`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
KPRxUnZqT8ll/yhEwu4wtKJfisjGzcJV843JN8HokmfkUdTuv6FhwtG6KA6o8bu3/hIApLfxELCnNe3TnScr/1GK1Wd6I0/LqGzm60y8l7UApJKXMOtoHrY40c/CtjoAxSzvMQ8AmS1JENkSSDc873kkhFDG9afSpioILqINyBWB6Vej265yWuurNnykSROx3j2K7B4kyAQeve0YaaySM5/q4M3f0MjgM4R2AIj/0CLBKgOL3w1yOaaNkPKN06VkIALUh5wBVsAkRvYTqBAGsaABbZgyxKg9Fum3Wryo58zcA1BxyjDRCX5Thk0vkIoGh9MOOmoNcBpAOTtAPKC6zfuVuIar9Xd7jjDzHohGVPjKkOFP9MJgfA0GGvfJ/kFYWmXpmnHn6Y5lvh0Dc65hImYtDtHwZagt7SvUsyf5J13WLlr49GiGJel6eS0SFdkOdBzYe9KIr2HtzQj7s6cowcLdOoB0Oz2pazAriXtAjHkSkHwn4hbBVHH9nUhO/qvh85IX+YHkqB0GhCVPpltRXVyZ1lNelCsvT+wgDRjQs9Z7/nS7cI+ycUjZmp6z4EglUe5LDnvTVyQjBjdIV1dSQFPknrgtZiOUJruBQSu7rAsb0seJ02bMWqnmNwS1/cLdY/4Pw/OgtyscoWDy91QkEcHlwbuqTxObZubOPSh+7CTkL9T48UD/+ja1ujPQ/ToieD067Z2HHghkax4ofYQWtjlQM21pZHaYNUSkEK/zzt6PMqgMvpi5tlBHu5N2UeZW0MkdTICj4L3bNy3Nt2j3B0RqqJVshnGcIk1mjn9gaHcygiZPTRGk7x/AE1EjRZSBlblJPldhAHa0jLBnsXpYtQBA2uaB+MbGblZxpx9z/bQMAHXAyfXtVZZ3vUeqWpWJy5WuAMJdszyfYzDySYx4OGhmCmrgxBhY2QZavwf5WtNMzLEhicPc9rpBdsIcXQi5aMyfUTM9pWh87mj7niVvz0MZ1KCBqCMGCE7AwhE5wbdfrtafW/Y9LSttdt10SdooAFE5AT85ol8mS3tSNeJBXw0a2rVuC4FpKdlhMNOvVRPTO/7k2OUM9shY58mc3N0peoJ32zzl8RE6nz3g2PXooVwhhALX/BFfyfaFGi7p0bkCzywyggsENuUzztZx9mFNGkgcxr3R7QHIkBpPp1N+Yam3Jd0BAB4UG9wyeBnMuwZjVmfoYSYPjtRMGaxNGwAsdv14C0BeVXDrlkH2RNGGqNxCCIxfrH16ArtCH5UfwqrJ7c6WAALc2qTAtqEnX1y/aEqWY/YHSi/wE+DyvaQHzZtBEBCz/T/TqJEh5SI36EOwvrTK2V8XZo6SigTTCf++wABEmYW122RKW+tJeLwUGqNgsYfmMI7phnxoK3dyyO91hCT17DdGhFyqiBEv3fvNpFsNSQ/aI7Sek6AWMae9XAxgD4O5/lPT4nyO5HQmhbBfDKF9A6mwdnXF8EzjaAEzNBSuUY01xZ0D48OyVIr6FLcuQ5QpdG5Vr9KKpw05y6bdLZXZtftQfCW6o4KBNzIi/j6/lS5xqrTWgPqbLgLJPfLZygtQkh/k0F/UwhDKnfY26nqUckTtvdSmvcxnCrbi0OtIG9wwJPFE+2o6LcUQSFy3u1RHMsr8l9kQE4f6PLd3qUNIIsEcBukppUx7Obb6LMgm4eYqqgnBMGa2zCh6Dof+orT8RpiIYQpoztgRvLHZn8dqkwFKVOBnWS/V0uZIEoY/uREQF6D7PKnAOsJKGRUmnLn0Pl02rGFrjnObnrerBVfWMeWJp3VHbnmizDXNCyZKgtm/4EdbWpX18Cwr64IAKboNF+4ZW70w8g5GFAQl3Ym4DvTnuNcwBsDgx5D0o4e1BGAecQmzZb0UYfI0U3R3Qcs/YQtJNBWL5uhUG8pyNL0ARD+aAbmw7Krwx9gFzl0s8J5vei3n4Jxad1owbArfEEODp075taRaKKEjegw7D3f+PN4MJxZ9nWjFvli2R//WelcKFrf/tmA9NdsOj65EhgJX2QBKYXxzXLFqpjRMgI+RSj3Y95dsm0tyHA5fCafyM9fiCBM6KLLasUKouo6EP0p1hH0rWAo1c5TNx0e/ly19glOCxdiV0Lnrf+sSjTAJoSxCzpJmhPX/9EbD6Egr28HZKQx0rRzp8d61UWqgkzzggeQB2xcIjrMuRF3lsxnY/ERgewjIsFPE4ofvQ/iDqg0uxbkL3zCsQQCQEUOOqN7Sb6udzocuI3V7HLrvD9tVuq7IOJwnIL/LCc2Ubho3WFpmmO0ARpPJ8c15mkgZOkL9wwnsPSX34FX4nj3+Ds+f3qDKiwAkQhwzx6OaeQi+saOuOXwUWlt+n2gt/npEObH25GdpDrM+MO7ALFvriJjGsoZ/wIZzXFsdvpOQiTMfpc2eU6Og1kuye5uILR/Y+8qBwA/iqBVvCn3X31qTgdgHYw89f4YrVxcNhjRJrHZ7jQApTiUP1e0/vgDbgeYpgv5/9Hlz/H4skM07FvOlr4MFV46fBvoZAqOpx0c+5/1y8JPm83VcCxYeYVuyTHOzYctsbc8PCGRIq0ubWRxDnMnEV5gXmyUfPzUWMVGiZdWiK7o+aC4vp9zsy8L383L2b6950FD0lM02ZQip32rmWNPeddyMVYQz0MEBe+fWIbnKQWta+4VHbjMCnGZrmyx2QtnAjv7fMvEd8+G6p7E+WbyaVC9sgoc9hh/1cuIF5PTj5mDIxcdKTOpQ2049/gkSMyI2bY4xYEkzIbabsuuPzfy3R6owTeOZOdQFIEW13k0TnapKujEtmm3Qr1QK2hAgfQEf5AN9Yl9OQ08WUbc6n8KOfldGENnq5b4Ppyx7q9gTGt7wtGMeSSWwv2pic6jWavTnk9p8r5jXXpJZgG7YXVfoKNKb8yYIXFG6ID5RO/c4Jp6aBELDADXL1j1nLJMvOb4pvBthQq83/FRsZZr7JHKp6hjyVxW881KI0M8Dgylt2tinjckyiyJj2hgOPL54LgDezNfep2eiwPjCThQXdLpszuydiedt4INLoqXhdB07gXKpm4tmvJ4n2oKhFuTEtEPE9QyWUp3XLMjMnEppRgqn3DQ6BylWo3tN4/eMEKLEwcGms/67ipwpsqWKchVD3KHstUpB5dItpew1DhaMY2D63uRkuKcSZbKVt/8zfSve9pkH3af4W8iyAaBuubYdqnMVg7pZ27t6hmrWGDUQdfNoW3zDx5/F3W9R1LcWFwCgdGVoifqQ9gjgvqTQCoYFU03anBVh9HDJFeoblucGNcCn5mO81Kj+gcUXgr6hzvTsp0DsazRihBVhXMsUJV0BLzTeXL8LuR8u4J2aWvl4vgLcwNAOuabKh/D4hJHxeOW2A1Ov0aNJOO2vg3Ggbb+h/DztGsLEodzhFyCm2/tXgJryU7BwqxZNcCnMifvyJVk6tW/V4LojYU0wYUVFGFSBnoQ2XbMawc6NnLgBHeaVeMOQknzewPTznRlWD7iibTvOlRvfe+43HJIZ7Js9NX8PsDakOramkd/6JNQb5L0gWEmVsx7bWrjf3x3gjS3roS+Uu1imbEUmeIn94Q0PAfnKTHjM5XNJfAitMBF5QcpyguPO0nNxq10XPKwzVcPF0t+iwXGVpB786U6ad+pMqu6mEYUKs9fyUh5yhbufrFUFOS1YeiP1ZsdVLNdcRptXi5w69wD24LrHzxDZkBAcYFIjdE2bMuxEDFnlciCLc0sibZ7XdnXFQ9y+HyMV42BfzVH4us+cqXbqYQlKLh1D5TOVxVvRjV1bVSnMTXKjvu11KCkN6MrVgnUwprQM5MTWiyrX4ilmXz3Zu5/cYkXRgLDS5tw0dZySkZRTlMT1+lEAqtQ5qjdFt/lsWZuEcMcb/SOM39gJKKuNmz6etRBxg/qHhvuSUz3KAnCzhOpJ8SXiDYzal6d0mAXf/t34OFyogSO4PMSuR/3h5oQPcC/oY1WKNFmH8cDTZSbvCketmsPXXTbIOWvrzHj8az6OQdiAcEV5qvE8V675Rmmb/IknD9oMZI1mwguTZ8ex6tS4+y9QyCjH8l8vKLmAB4Fld4sMNdrQ3VRtqsBQxF//O+JdyNJ2lKQo5xXcEcTUwv0L2VrNkAO/Laxyka/4O8u6vw/lLHMgcCVjg9HOfX/0dGNU1MiwLDNh78GS94G4LeYTjpHV9cF6B2CNbInrLqQpFvmIXgpP5drHJrIKygzKxdx5YfAsFmrMEA7hCeubIMhXvJDiKoez/fLMyETjbWaTzzt1APlF+f2bou5vidgXtu7GkUNqym1rLYyePaSn7Cqeq3dLdzLxjjvlDMtVjMDoxhIJqPSte/WIOVCGudYq4VeUCMLR9+a6VcF4GJg0HmUGWzdhtOoLJZeZl2XRzKpcNP0RBTcOMpEz7kPLFRPLB49FzYu0uS2J+zqcDPvp9LG1Va3npHYfNtK45SPovGfNjNaAap+ioJdRD1w2M/yHvHydQHZNyLYfJz07/z7oWFBgsAHNQJBbdK9RE61AXfSzUg/rUqeoMDnODMNlE9aHiS/SQjnhpLN0q0Row2tVA2K6fZq+oRKovejfY8csgkI6+eugdRoLq5gWWA4NX8NUCjfmJW19AmNGFEGYryLjI6NRQnKm0fEa5pZvpAmAY5YGlQcWbwbttqegLrGutP5trOa6Gng3qSamOmSTj7egoHhnqf7kiHXfpq4YzeaarRi6blUTAcyDhkVu/eH1ZrTfC2S5iyJyL5clbBLqZ7b84AGqdJKrSO4s+DLdzjwwQLZn2xYpk1oD5jKmAXKOtntNPiUrBvXo9d4Se2Kl87DGe3T3aZUlbb1g4Ht408Q1m1aasY1BpNS/S9pUG5BhVbXMSYbKVpgLOwaoe+Dz8BZT0yvgEM1uy39B9xGZpB2husJsUr/QLlAVzH1pdmdp2Ml5E8m1CrmIC41fBgkEQ4yYiHUl7Ijb4EwXIDK6ThQQuP+IH/a5D8/LR4IBRPdQUwBjPBiSP1Kftf8wnoMHsnXqXBQUUsxm5RK7QHxGoD95vP5yd097ehQN8Fq8mbHRb/hGyROyYKB2hwPuXvo7qZIZOHuAPLzfDmXMmBtfmtF5zriYFBl//a1ctGXOW9g8I7CZQOw4xL4ZE1wXkImgz62d04EzA2357Jh0KkZ7hyuZURhsPvxqHiaBGTF+41NFZc2VeZNCwzUhHja1jYhYBgVkEmhbqXjaQDxcCPNcdDaSoZu8+z8ksy2HGeB3C8SdDhkjBlkhkPqslvHIVDseKMLiMxbtrskJVGohb+3ujNuortY05ApJWX6G6WV95chANHQANU4hE9mweXVQgat7KvE7o7Y4En3Cl0+rk+oCM/tBxANFWuDXBGI6DqNL07iRMNBUHok7L73VPUtr/A6+YO2VTM4M1Gc+a4dMLS3fE18m3gcNjbp9VuWuKuF6O7648k7CPlACDDZc2zUd0dLu2irJsrlR6E88R7iMUwd1Ni6+40Rco8QPHWf+7rB9vwhth4ZgmCVJxE3Te/OltNF2J59iznTLAaGun4jBl82bSggIbxcCfYMTuFh02kGVMbhNLMDnHaJ7uowsMMcNMO0J21c7K5WOqoQJhj8QgZVxYTfY19OS9jtnH2zwI3m5GDHrZxgCctldCn7NkEldS1lEFExuO30dP6Qwkm+jdqyfnX9hj0fApLdR3mSAPiansF3NvnkaCcF+vtYMSiI4cDdrQRt/4HTu9SSwH8csvBZ46j7YjPI/4ZdvFm2iUu65cNn2ljZhtw2Opaqzz0q+zdRlx1hYnzSemqgokQgJloWQPW3CyYZH085GID1xu1XYPn9gCoFUsBQeEdhFzdAo5n0H0CwBFist57ybB0MAYqSJS4Ig6TER+wR6yjj9jifGjV0CvV4b0aw0arEx0VAUBHjm83wLBlTZ7or7sQ3kk3RfOEEjXjQZ356Oxaqoo1iGBrb+dNVKoIKUAz7cvGFyIfGHPz2oQcOF7cobFtd7LK+5huGq6cgsLbG9grG1Y/Zj9bM+9g9b/EyMaM9D/zwm9C1m3gBJ0BFIo1kxb5ZbFj5yUYgJMSKBTawRoGqPZzZtOFv/V2P0pASWKNaERca0j1kpKpkG5KbpLj3niy+W4s43RGuhvxuGjxStJ8uVgJeZedhTTUHS+c4WnFIvE6StctCl/KFeL0RLDp7iPaQssDHX51e/dJwA+vjdl5yuabhsdqJP3z9LjVM9sK+zG5RH42hXeAEE8RaSvQtDW2KcUUd3lyZAyC/45jjrxiocm0NPWtGk80xc2aMo/JXynaz7wzZISjvdCYM2nl0qMNx8FtuonJOXKJqDXdaWfglF7YgMCqiHnFuoPhYfhOjnIFpv22+bVigaEO5xvpfymXlBtaG0Ch/x0LF+sipNN8NKMtZTX3b5nUmd4ImOxQUsk7SpyKsLxSfrCrRlmwr9q5D5vhN/zixT4FKpa6O7WQf8FeCni/fHvjOzddbgpzLlrD+kn8iqXiHP9djDCubCeGh70wJVgPfeA2oKFXp/BwpxM6vk9WhOaxYXgZlNsl1vgGGjbuO1egvUACkXY2AFhSm/SFzpYFtzM2sI0uUFBz/XYZNLSPLpTNjk8KI3m9b0vhOK6r6B4W3Sxat34geQjoeJj4hiGVzc6JT0fTcUyKCS/wgnucKotaq3a6z8SleK4sHsND1YTp6X5RMXsEm3X+yVPESgYGqrGz8W6BDDK4lP/u5QRS1c8+ZFZ1VOeM5RpNBdE2Mwj1MZ57WTKt30VJTir49/j+DIjiOzLo7urlIPwsD3ObfnbAV9Hp5sntU6RMd16U/ACUpAPzWG8N1QplHD4MMmGSh0rsoofbtP+Q3PXWWW/6bWx3Y50l5qnhOqQMOKwwb6pC5GY9Opdiu3eZKKVKVw3BQa+RNZ7m8887iji+VBRH9wUDytyQThD3vRWMjF96hanSuS4WLmmosj5IhjxOQxLO1FL5gcveYvzU2NXr+2Z3vrk0zInsvVdevQwzLnQ0xUI99moJDrd4vm3dEXLrXQiVjzmZ7rvOOS4umxti9fgnaXNSJf0HgWEeSHdbZbeAEI3g5dzvkP0dFoXAQDhT7U84KlxNNd6Fe4r4ZDbsAaUyikgyIy8AoXBVQtS31Jw2BzUhcYLcb4YZpyjbGGBSpJGfc0yP6gvy7LLeebi044zh+umxC3P9xzV4qevYpd5F9Ddxjv6TXDnhcZF0GKGDqWSn28CujDXK/gP7RqqdCkRlhd5bTh00v7GAn5+FwBBbhuDcZ2zK4Dxx5/zkZl5zkPU3+kr2SOBAI6se+kDMzc0+anhs49nz9Myvz6gaiA+4hrTmfzimJpocbU9/37hXHlVRacNN83iZbJaQkZsjLa+TbERE8pWqeKcRdCGwXN65l9XcY17M3rpoanMdDIsavWFH4KgmPn76RO3rRsSBd0cAiSbFcy2LV1WHI2Lr0DB+kwklvy9KyAFYRD+yPI/sfN+BoVVFOCsn5LoBmithHQ9fQKEsZ8nj6m12DGCROiuGewT/gPr16p2hnVX+3oB+EJucQLOcnKrTS6lTBR1q4ECR4Kvzgu/+Z7pn/SnL7R1MO3c0Lk/xm6ipFXlapgg1/1lOk83IilDmUCPMuOwJ08XDd6LIVkCZcFT8nY8omtqxHc50OO2upP9d1+ExD2gvLifdORsKtqlE8T0sABaoNfqaSkpxjPYc/Cw503mz1HWMuSsGrXUzsgvUd3JyIUb75haAixaxSsWE7FBph7B/BrPwS+KAk10U3zfQSIxXzBABmCEV60Ta6dpanldzkltpATP779joXOAYDSJtNZ4kCCtybYjgouCLREjxIcES4drUbT27BdZeh7O+Y5hZoDKKLTicnPnXhUPwg7JoW8FtysrKj9rmfK1S4hEgZAQqVZQBNFCxTkO2ydbPb52dIFk/yi29ya95YHLO8rvdsrYz1BXpvneExfc6qct4QzXT41AsQClsa5Xk1m11mvcvTTvRf8ZtPOGev/YJBc3xzhHi8cw2fWcOXYD07zO3yXXXlFCZR+BjTSkRsSv4+1T5gZ/tLRVbjkT19KWS7ORfA/+unth2ctqhYAvJCGWMB5Df9EOBxzrCgo3rncyYkrrUnWj+ardW1NJrTuiNVSIK0QKyjYjMqJwhP+NlMhtTae3bHROeAy2qH1yBRvDMM3VQHjfwqT2K/0Oz2SxX7XVXW7IYBXN7PJ+lYPTQ3YxPjs5uYITBq4zyQ/btx76H5xLJTXGwDzS5B0dV6rk7TqyJEF7/dqhNURdHydu+o0Ny40ViNvNSiOVTzhdOFqhgnuLWJnlJIsLx34oAIqGNyrjJabktSkH/6jhwgJSfKOtR3Hq5Yiv+dm6T3QnXY38OmkUNGZXh5UXDqvUxL2CMBaWMpWl9pVWNFz7F8gKBYYXFK6L6JnePt35JBVUkhIfTjANTYLCsh1t2xQ/UeHMEX1LqOsYIgLOxu2efjvOiqZ78FUnnYDYbsq2wCyFmvUmWsunq1K3jj1G2AEVqFXOXrHmH2E1Tmw2pU4Kg2M5xmB7JWoV0n1rnUvbAM/40hAfmIp/aEhobZHuj+tDBAZjbZllosF1zk3Rj1nu2FQ14KXe0Z3cPiiGK/bgh34KYWTye1OKafUGtYY083YE0SqKs8IrPhiDXH/WBs43oO7tAc8DfDsOHedfPEhdEQ+vuXnBMmFrGjC/uC0xr8XtbkoGxB3A5dWa1o5RHr/iUivAyKybjOau2QBiyMQ45ugg6B7ezITiYEpDrsu0pIzE/OzwID5lCh2a4W2j/mcL9XuXbENc+1eZ85LOM6I9hZD8MZRysQkmIpl/Y67NQe9zd6sF7hG0MYjZBqHGfN8ZYX2UVIP+ZVQBrf++GfCzMZCvEdyntQfAGaiJhjWqmJCxMEOanHIm2D/ZwOUn4Rb5H0V96cKvS1d2NuYHH0kVaEfCdMXCdMwaosVYk0oto3Lb2uBgF8wABAc3e1LcvqcxykC+rwD9hCwm0vqIosBTCJxvBa01uBKCxpz/lnkNklfpi2CYHKYUWx+f1dSk/uCUsa9mqO46tbfjrZiSmbyn7dcBv61VMK0wXWGqlT2gkf3dL9aDbeJKGL3RK7dQ1L6mv55T6ykuBNqyM71L31qw9aq3TaSRIVWzroW/uccI6rLJ6kCS8nUC77v8TOQCBw+RHdyAI6AApGyZU/ysIW/ZboCt5njyzXeBsp/OqHjo505yZahteW7FHeAk77Yg7aJk0xbhkFgBfjr9DlfPnZAsyhg317kuNMCD5yhWd5/7FtXd+FYp4x+HNnVz4mKsq9ANvQOfK2gza3HT/awdd8PdQBAWwADTrQwaZVNcC06TYI3vrVeF3iwkWFzBHHmN8LgPjmpBRLflBJhRWtcjzSozN2uui7D4EC+K9UUMRsVoAupZiUUKrFK4SXcwIA3S11BN/IXghw54X70zgjDpW9O/Mqjxa7nRlpUpIif33d2HAg5w4uCuqvDlpbMGNPx0gEJwZQbG9Yjg2Zc+I3iwtZnN76VU8kOC8VvTp9798X+pME1se0qxAbluC6PBSvF4HRt3fBxpXYgoARJC2u+DoyZTppO4vuDWtep7Nta/t1C3/heHlIZvuZ09iDssP98mxdQn9f3iUoiM/442y/42eUwvfx0iNyxlA7+QJTvNICLVUr6IfFrbC20dZUMxR5uWJhh7jSYaDDL0e/enz4RDWfiYS9Xm0LYHoVQqlKGx+5X2SYIXjeuG6ie6ib9qqAx2Vi7Tz7iv3TDcOLeJaHGOGe1DcPVOv5ZxAirywMNncEW15Fz6Lqn6T77Irrzp2Ncw83qWOsF4wESjuXbd5pTuMLeibArxvPqdmzzSTuMdC5bM9Cn0aAAjluj5/9nJwFboJlJtMg+jTECS8Ma8wLxwu5/itRZ1ShsD7GPMRBlBzhwHNtU6HEATE+H1Pgj/E36O5gbz61kILldVlNSvmDAncjiEDIj3zB0d7+Kh2FXamLTTstdEn6dozgsFWB4K1RWNrcTALrM0nSzFhtl2eXn+LQsr9LSd92B4r+UD/Zh1N9RxPkAHUeidUONhtAo1yzTH2FPZVc/xRGOJ/vF9y7EMAyaghUgY0W7gPGdDZR5O+DoUsQAXxZAcsSy5vfnmeoJSvDXsEUw4vG7C8pyZPGxJXBVMlS2Pndbm1lezdW4QRTM3vhiwavUCRjn1Nmx4XUJTw+dRguywC40XL4yallIeO1XPn0EkXxvAqyhFSGmvQisOMxEmCa0wxJvOLCOX7VBxlr8XcuTmbz0n4M2fkfByvyvvgb58lTdX20ZKcBsmQHsrNms520DNP9XvkPCAFEh5h5YjfIMIKMprh3uEjG4oQqZahtFuePF+e3Wh/NgZkZBcPWknlBgTN40n1tEimB5xOMgx3e1Cyws3JwUhmStHbNYGtUkLsSAIMZA19CaroF4SriSo/IhBx2Bdm5ntnydnwFUliUZR9o7uoJhhbYzaiqsoxt/dHRU+s7IvC0ljScLBU34B7a1S4rcMbG7pENu943qB7vW9vtKsCvVIGUKhwCTfwzTIZKbg/vI6uqkoyg2N7Rkz/UicU+ppEW3zYauLqMTnrqZnLoKQSKFSV7POSivM3eBpsSCxvXcxUFw6LbGgOPfAxysKyZl407l4wqH8ZWknoa/CXv9n0uEpYMuokvmBxYIAFSsR13XoTegit5Ra1BNouioGf/DjhHBkAYmlI15ogtD0MdKK0f03lnvLuyemDIlpNOezAZkXm3SMT3aamcrYxQyIC8N1kREx0HIrQ/pvk4LCIbWlO2GDGgvtNtNtWwF0TEBKK4cKcaM1MlRu6BU1VWF5NSk8tuBBItIb9ZZiYz4DukddqTfUhNKesvFGpPbAiSgIUPGLznh/xKgoQ69QWTlXP4lkfPAFCciYKRPqM83n86Zqt2BHC5g9vse9dcKH0ebxd0BnIyEQyLYI9t3nlraXXwmK5snF/EARTK0sVjXr5x2K7fouDa5bdqXsN7f76DU6muhxOi3AOza/bhguC1mzWL5DXhc9zcpeGoWy+3/6oyo+gAP0j74R6G3jAjA06LZGWl79y+Wn3fnJg1RO7Pb+iuxenMDptC0F6DkA/SKhxoJ7OYictA1ewKF755nKRzQEnEbxZbLBHfT90abZ4U1El7idP+EB3WucHLMohhhwg/peco9ks5kbPmbbZab4qmuWIY+43+znQGmuR18/Rrgta5oNWT2i8TVclZY7LspjTiu1df3/DmruMUa9BGAR1C+Xr3WDX4R4fF4MzaLs1ysmdIHLlBWtuejZrStlt/miUewf9GuXAwSQZxFo0zfMRduCG3ABN5Lb0PMIPC/WdkROU1eTuXVfX61jrz4d4OG4mibpUJrxMl0E5C5MRx5CExrmnlO1kgSje0iELeh+ae+k/od5qT9cBaLPS2+lLbAlIC5AsjsgiVaDe8phNFZjVu+/L/W3fKYNd0xKwYWHKFXP7G+tX0738Pf3XIZvfMlE9UHlg6uDELRzmH0d8BqBkEWzUBUI69g2JYfGMdJMb9f3JDVyvMCvu8oOJ2Z4cND0nokTVDLh273mMvr+mlenT2uYlpmG6IJu/Qjs/SZysBw2yjcfxK6E35tdOGM6gM2g0MNLZVBi41jOdNjvPS/dWo0PUa0x4KcQxBiYmClrq+uo8pIvfl/F782P6gwM9q3JTTl/PTXx/2Mmu9HY++0gjoEdFk5kbJi3VPTEFnETF78pyXkbmcPwq+8JV0/sNy9hZcZUpYnllABYhhwgj+GzUFAPtn+3V5I1t63uZMTylSo+qLJ60QaSS0Xa0e962iqtdob0Zgc2QlZiA+NUyPsGVr+WmeYpZQDJ/No845Rh8jqBTR/QPgyBUK6RSC2OyU7yr+gXgLQKOoc/6D+7qAIAhfwZip904OMPskLG6dl9e3OLorZNj/Dky/U5zx9LGXp1yz3QrT8JZ/v/KY4J7Fnxa0rPOmbCjtOqhxNbDM6Lvd25l5pZSjKnN2O5X5Y9peBaOuyF7prwW5h7FZCGk9dqMGd8mvyTuf9RmHETZFtgGvBQbdeZPT7ua1zHJjTAq8x1KoeNp/MgQwZHad7mZzABEYdvQ5JtsuxfTn0+BEJmE4/Z1bDZImzecRoVfmURNLx0/cWwMmuoi/t89nvlyhA9+7Wye6+VmsvubCGavdvmdbRdAe7JH+KUIm0paKVInmZiZRvpDq+0IIKIp9v1BRrRgcpIOhxIcDQ4D9+rpDkoqlDLF1AnWldcr1FDE/uZhjVQ3XYYYFFORGs2z7kPLTqhxvkQaxprYP2gmRkvIaCB/usNgQn6PkLHPSj9GvMPZmC/GbD2wGaZXF9Ip1+MpiwqSgkQjr03IQPdPneEiraqJD70NpP0yIsEkjgc2rXyvnJyUZtekDQ8fjsp2j5cUpVWFPcChbHlzWqOaHOryCMBt+f4GX9EUWriAZFI0+HkYEUDsTwHK4odSDPTxLYVx/m57qNcNczluF1xasj+LCv36WX6QLHJzvypH/7iRpm3IBal2OaNaWMFi7t2nw26xOSPiJ0HIEiTQ6zTnTXvrlkNfeuJr8THRCRVAilja2nluAzmQ9Tlikx00vvkugAXPDkDbDFubhtg/2MjpTHdxiJrrv4rKX8v/LnmqY2tjYNuqCu33DZp9EvKJ25Ow0SoXozTzvTG2ggEuQNc8LsjuFUEEvjmF8P5ZUawu6TRourOV/Iq+f/jXtsL0l46rw/3SQ2zQKOzJpr4RHGBtiPTeHMQht0VrjC7EN0FaBk2cn1ucGl39TnWzSdfr18Z8qAKhacvQqC63ZjapD6I2vUYisCYfw/nv0qJJHepU1TqXyucLPmXBZ+6ZaT/fuUvQsI/QOIPHbUWtC6VYvbprCCw4yeTsfKOJhurE3Hl3oAzH6r7vLlLz0Cps3Vvha3l0UO5OckokJc/rBfFkska8ZzwU11xOTwjbSQjjo5t+absVX+zOqp4d32sWSO5HGU6MeZ96zJSov872KxGhXY14hwdTjHBlJYdeg77wOuZKdKYvFqWi9+XT1xWFi2wqevMmaIzxDrkV2wqD0TA/FdUhky4VUGpri1yhiuxfyXErOfNaDB6rnXtnmqUsVFGnqITGeJnNwAHcB8slt7t2mfjesy90t2VZAlP4VxVULT+0GhFP/8APgaeEOCydAhbRRtGJYmlbQWnou9tYL6njm6IObgJzE5ZGkzmX6s0C3kopuf+VOCTfAqeOr6jkX8Z76s5W9BMZZNdJac8tZPgbBi1qG0xQezTXe9Y7Z0gR18SMlvULMTqo+4lEZyhIYHmwWEd81Hqdbh1XH9n3lyggGvYjUyv6BlY034T8Aj+CdRYTcDijP2bg3RHYuLM2bXUvUUlSmqnWs1T9C5nr01StSrEDCAhTk4ii8ZJdXlhPDRqlyzrcSLwfKGuQn8HHKzEIF+Zh/sA+GJmk+3jdaY4LB3u6mJxiKO+DsiVom284OK5Sq3Xg27dTOP0r6Cc3ChDyI5WP7cXC+B4x7xLXYPyx1SH3Pc69q5CXpbnWxyDUi/LtijpWMOE+DcuF6W4qrpimsXHo8jTDqFVNPCJLuDzGfYZNDeeSwQFdWX3c4ajTghA39JambfjjEsRszXFxdpwag7rSFZjfdbjHqiD1j4XsMIBnitgQuBhEa6X1ZOg5jPHJfXEA3lz+PNfRpn7IKKPExS17N7M22PdOmYaYXE3ALvIwkcMbUVCZ79yk9Y2YHkldslNwm7FU8TusO21W8/YMVnUmTnghSsBF+sYoJjopso2SBoaCQjtOZ0mgdraRHUEFLmG/6AzEQEY+XoYFCLUl2seB5O1Ko4NpLrJPhzFKh7aS0uzanCv4Ws55/se8vs3l34f4tQg1z/xXnGBVa0FhRLIBLDqyaTasMD95l3KJe+ZtAoXtYRo+zicXL56UjDtAUjoh+jvHdo+MUsNPz4H8CGuIWmqR0XG/JZI5rt7Ag3kwV5w0VyRqLZS8siBnx1Sud56jCdNHhiYHkXhVPnTdSC4cBMhb4N6UjSTn/UT1P97Hzjc93ix/XFwweeG5VqifhfgSXgJcrkV9fVtb58PKjmlCR08NM1fuXn6RUQsbCI3Hs8MV1VaHnSpijQ3IKzFkiKfdNLTf2MOKe0qgk5kvrO+57DgSXxWxkf6MEg2l1sHic+/lqJyr36Woj3U/n+aeNwhvB5ZETKc6GJVneHRw5edz+9wPwuoFlr8xJthoVCfeYh6xAZiTddcBOSYdbWRo98YlLEw3QYqlXXwLo=
`pragma protect end_data_block
`pragma protect digest_block
ad67e738fcb307e097cab72bb72fc8e7536cab7a6fae2cc52f72263fe40539ab
`pragma protect end_digest_block
`pragma protect end_protected
