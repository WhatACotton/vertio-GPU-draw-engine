`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
CLx6Upi+SAZGuIPS/V3LRyprbHOywa/CW4ogvkmTgb8XyITttH2aq1fsd+iQV2I4BziiRSeI7V9mUTxDUtRwz7G3HPxihAoD4dPJgoHbvmHeRCS+UEB2DreBmjFOWZ8Jifhx2AuXxXZHjbIQVItElrZOWynubEy+pSrBuYwCwTl5e5AuFlPgpYRU9dTx7p2LTq0KJLR39kY6mBpjb0/2MC+3RI6HxsUCBk5x9bvRdPFTJQurbbH42dtnTRcu6Ql7xxh5Wz0zB7lyEsV1k5mPpO36H1MbmJKxghDIUtRffjFEOjsKYNPNeB583xvu5UwCxsMOf75WiscwmePMtPcnR6i8Drz5wUMHlUiDG5ZQ+tdh8min1iTvScm2FFJHxO+nvPHdwUB2365+uUouThwSxVyat4pM1U4rH8bZ9GmxjI5oYtV/4eIJWMqS0IVvRbIo79OMJfNx7jGbEIbovAfUulxULBhsjN4MydOL8mP17FV6hOnDmEhqdhd48HO9x8M/txuIQaFb3pYipggMCGcvPpyZxTs3k0ypzDpBk/tnl+QZJajK0nsphaOO+ciYuzPYgsUMb31pfSCZxgZQzeUaKmYkE/20YmX9bG0t8Ln1TgPGFNrM3fX2AgdzWOKs9A0Gu1b7Cj1VhPhqtCjhnufSOjBdgjB9CfgPIZ5km/ngyc1Avl24MXmywyytaebEU6nJuGpVZbhAYVeX5veCIzK+uIbQs/NADMW3qy/iy0P1OW44DlNJswIjCcRb6DdpbQG30O8iewOv8wEua+XFdDQoDy3buALtgkyuP+T1l3LtO+m5b2aJrL696eD3icxd2mBpaen1+RI/uHCbDq0K9wHRVDUORPY33ozsz0kuU55ETQNGrprV4Q6iV3RxEmlpnKD+aaGzR0peKGnetpJIgHx6bNdnLx8Qp9W9GZ95ZwuqvauN2m8IITg2zEYH7HLFZV1HUCusURIaeyDdWcaF694hB7FTGZAe4EvECEmbFUeAAmS+9G7E9JyVCSYuPaoQfusrS7fvPbRpMVa6Mx68UuuObx41wl3V2/s4yBWNc2yZpwvpEOweB/1sQ7H7JmEDwvYAp9pjsNRbmdiPLrqlVY+3utWToaW3oqg3XjiAnKPeDszQcV4fThSZAwgUgq+ZT2ycOi7ZHvFz87ELV0CysVj0FlGFw41pwwIKx5tVE9Oqmj+OUQKEDNOQ7YMlHmQKZ8Crj2ReEFPb8gkxuez2OfRgbRJBmq8pXMC1hpKRKY/EuO8SbnUEIu7wlHpdX+7yxtfC6itUFB8VKvL7SM3hXqvbv4u6nWfQZxDcbB4R2VdYRRqTmmNWWv5KI0bEmDSjvt1BvWpwBTB3i8RZxNiFUvMTPU5lz9Dbes0p+X1sUHRjiHcn1hEBwHdZWUYV34MC4YKUpZViFul5HXaO82W+yt46eagMG8sJEWtoTICOb5d90VfW6ja3WOah+UqSoYzThm1a104tTrk8GX7OBU2IM5hLZQnFnn8lNcnD3Qs27Z24ymMH33jfLDlY8ovSLr3X13s3NF2gq6yalQ0kK16mva5Wc/YLyghlMP8xwcKFYv2Tz/le85D200ACUNnXDfjLTlvz0e9EqQDVkt1pKaFvsZejQT9uCFhwMujuC83Pa8lE1ydYLaHsLwhZ6Yrv/ClUpN9dH1gil9GhsmTtBfkNrYHuxW8gbkXroLRpIZvNuKkD2Qh5Xu4cAd+MkDe4qMBl9mn3YpYjS9xAL2MHxxxZjpTlwFxVsdPCcR6udDqLRBcNOQepJrSLE65YD5/bCsR2MG0FBVs2EVfVVpJ7Dy58zDKuxrZWp7psKXfKsSZjkER+ytwwMlfrvqoMKmMI2MtRvV7pizc0JFVGeYp+tAxgtZPBO0vPJfrmlZGZfddCH3bJSqMU/g+UnGMLwrPEvCO5J7tJv9/0RdGl/Yfno19Xl+G+ZTv8RdvpHLdPidykVEHCFEXRu0aNye/qKMYP9FK0i6kHw6de8chnWmtD6Y9t+7ZD4dYhkkqSJe7qZUNkwMFq+Oyd0EQl0/jbp3ILy9arqU4kzrhlxg3Y8MNQyTqol7xzaDg0VUzFBMcCwSf5+pYzlvWt3sOLOfgNcMdWq6NKxACaq8YFQWDMv2g05CCOqo/P5yR9dxXgj+CNd08wkYXqY6jtbNc8O543PVimpHlzKQqEnH/xY7UWFpls0PcqPzj2zK3+mmEnlPZ1BA9C88p8hTbw9VwKrvT3Ygl5UbDpO4X3gtr0jYCLvuva4jeEzlzbPCieR6iMB1YuyW8q0PQpzPs1CDjjmX13lnJC8KeMx2h75Wttwjqp+tpRa2PD0cMYYed89PpBoQ0A22XTPzq/ogbrv3H6A1gWxXi7P+3sLPqAm4L+pg8iCt6vSWQaWzbWPD5nW/bXdgxM86Pe0SEiygdtZgrmG5Rngke0DepoZzKZ+XnGFz/AUyaEBqIYnnbjOz0+YtiypP9hSXZOJTByn2/NyqURIMgsqFOYD/evdiNFSFe9ScyCgsN+RGf7inx0oUy67Hw0kePoT+xE6mSHUROKKLAP17qbW6lBtA8/1AJ/NLYA5W5BfxrZtYYr0tdWDJML3ddoy3BCbN3RKxMUMmHOs6JmSCYDDjh4BnbIgJxAZElb33LfA4h1wlVFci/0q88VEf14ffrxraR2y98JQ/qN+VThZ9ZgkadStrHR7Zcq6efAU0uAXEfe59x09cETEQcoP7oXS9mS/Y+7vzCCGJvIlVraQasV180bkTY23i8VQRLofNO2gXwzpwGhDm03HCt3JXw/DRpWahqs77oYAuHcWXW7zOjLj7kaLMBXlo/nrEL40zYsqeZJ0T4ysAo5tz1vhuYD09ASiN0cBgmI4I9Qs2rNQ4BvmqbCtL2euCEaiGjavfd9lzEvRGe/PR9r70Vh7W7KtdNvsI6cXqFQcTs7fZ/+SLg6Pi7oxQxhknr1GvvsUkfdEezpryOnMzwX9h9KFZOU/BigxWZnPE16GRqFwlDOS0tqn9kS+EnSZ/1TNtc4kE2sVoxZUYhxmNuNLWz89SCmjunCnGxVuhLYfa5DjjiAzl7ulA5vEpBnZlfcXoAQ9wRBO7qocJYYXXPojhPecfeOgYhFr7MDZzT4upY1od+IIk0VHBexxq4Pbx9EMEbbCUiYsci7E0jDIGZUnSFMJq+x4Qq0XpschY+BzzPTn3sgoqr0OPW4evtbOb/xYTPNyLvqt5OF1yO5jl3vaIFv3t0dmgLMTe6ssVTSwnWNuFPteLh/zlsXnxyQQota4OlJYddbZ1tudhr1KXSWpeo7bXT1kO7275G2SpV2ySNl+PelrvZAAOfIIaBLcSFGwnkwmwWoKAl+6we/iP6BG+R1KsdrKpHmDP8Dj1sD0AWuh4zr/MmsqBt23LW2iXGMYqmriRWlmSI8ejFyqR1dw6dh0byYsElIywMP2C7FCfGoqJtT2tcyC4qBvT63bGmEZOVdIRhmj909IDbocrcvMo6KuLP2hpH6Ls6deY71c7w=
`pragma protect end_data_block
`pragma protect digest_block
e6c8fad20f0805d611df125bf3c354666ffe425c8e31b07a4897bd9b94e55908
`pragma protect end_digest_block
`pragma protect end_protected
