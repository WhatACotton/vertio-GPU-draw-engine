`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "31a463cc4045fbb868cf41f5bbc62317"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 2615)
`pragma protect data_block
G9NOsmIkFw3ieNNwTAYWxjUx60hy2Aqn1Fp8/IHdfRU6A7mZCNVPHVehjgnXiRb3lXE/katl9LXGwu2WbB4grd0W5AY4dSoCy1tT0eCdQ8fqCrp19rpDovcJTsjtuL0LvHoP1VhOPpPvdUej3ylffUVAVA7CldbO3A7PlyLLysSJBoONC7sQPnZPvwxf2QPlLlqzQ48eA5KZSYLf0JtX3YohWfHJFZPJSEFgbPn+mAkxwwJ53AkKwFcZjl3VvJngBFy1FqnCGCwwYiI/hWOVnVafMSalTD1fVZwKI41znrC2GuDDLanVsaKiVzQ3/yRa/8JRZkGV5d2JJqLTCFWnCNqSxCNruaeTCPyB+yLdyiNtzdCzILCjs7isdRQ36OSfvyou7ev2l0Y+n7/68Ws7NbI0V5k3NCYxS9DOebFAVAYZUOPeeAkR58ObUSW3/oGMX7m0oIz8lWpueDhvUAnGjem97xUys+qptcX0GQjHy7jUjC41A8cB0OVAHFRT9woU3UdzrsrPffAdkOo+BUHLkmwpJA81immbxv/9rV5/MIk6ELUGHxSaHK54+fK2DCr9OkswXlH8krY6GRDIxYp5yuzqXR2hogF2TthHN++nlvLn1BXdrr5xHvWPUAHZ11klCCuqPQEaMeb8Whu3pbmt3u+78EsCGnjW+BRtO2cd4OT512sPKxodiE+3UJIdtOx+3WCJjEVWsgRb4Wq4sqrs9JMzq9Vox5Fr9YLcICoaIzobSRUD7jXRXkfzeMY8P9gwym3OMxm/wqjhCLrSeZntqDXBoKQs6hhqb57WbTSQA7uuuWQ0BILXX7GXz+Zf6qWI0UMTrO2IrcFqRTzQbguPRBmiXJlkmkdINh+YCsrxts0ivZeISAQEr4xB4U8ZuThjSV8QIhnzgtoVpu1eMt2y/kJvb3fi9Fj+vSXVnWEL10ecapH7wSXHG7VAlGxX8300QUATV3kOdNFTufxpUhpZPnhf8BynmlcMKyuf2n3gD63RQZsIvK2HElNSloFNM27Qn7dZ8ggV/dRDDILDlW9gvgZ+B6+bgT2vHuhuqh158enQI+3qNvEbZ8YwpKhs6o8/3KVoPir8SnIVQDWuzEbUKgi4gduIkmyniOrw+0tgATk92CYfKsB7NFPSe/8WbX72Jcq0CghzQVkhs4Dce0s7vN313P6OeHutFnl73NBAPrJdknlKTchQxATtdoTSuLhZBXbJ3IhR2sB/NUMQEiOyiJgjJRR43IlMrkt7vjhUoGGWmB2rbAIE/gXL7frLMoZhLLhFzj3XwsrIQlIOaetQfyyhLYIaBjTsa/wrYmRkREi1d5XsDtmVa/mjbERtxpnpzj2CWdo/lJjfB7ppdOfPC0KC/uOjcEzfVumeYgkzlj0oyOnyKLSI3MedsshKEBqs+zK4H1yUs7cw+EbuvsOArBGqM/ewMI0VHqolcl3XUPRjoAe79+BE1SSP/t6i4JXJHb42O79bqTV5c55ZDXrl4xNe2sWfuBmZhmZHMtDuDiZrAf7cPUtqdCCznIs3AosWE92xIP6gMmzRcFuCypFybkLe93TsLxxsyMWJ2hJ+VwWrWZiHthHuKIy8HO9SshnjxgFiK5kYfYwnoJLoM2/dRTv6S6Ew5iFhe9DfovzojUwMSl916X0z/3r1zYJGZZnbV3tCMCUVXW+ZVGym2UNIHJG4aWXDfnBS12eoSC5qvMlPmxgvJrlsvK+1XgZGg/qWpPcL356nSQlvqxVq4IisLjCNrlncLGA11RY8iHgeogynU5FGz7eZX/YwrlrEGwYuYCPIMFCIXeEwWUESzQ3mNwUQ42/xTT/AM9McIFy+EuNw1cnGEw1rcmGfmKdb5w0NyQ8eUxZXPxcnAq3bNVlJoZBtc5xxdgiAky4EeWyf2qTQI7M0UJpNkv1RxcE0rThKGAPjN4zBMfqs3h+gzv3xwX/HH0N4RCLFtnDDYF/2nuFRl8vaM/2W434SdOGe4HNytseamigLLjoRjB4bSIotX2XFYvH06AwIv8Luht7h2R59NJ+tzfAHfv0HlqvESKfS86NvY1TrLcAvyd1rvFJOzC3qG/PsuYujOSU5gdszuLvQXUKwjxniWn4Ksh6ytvCOKM34b9gQdwSIafnXnISYbXbDemJmqQKaY4DGbR9+JprsUFFcPWi19Lh8yj9VDxj9YJu9oXmwKDZkAmlBjIT71WxyoEWyBwJFkKryt/Hc5d5IqMww9HrL6gWDLlLONGuY+aXmHeQCkkLuFRz8BVp2L5aUFWZc5YL9r2x77gE2plsNM7lAjWIeUAjb+rEUkAP5im6Xw6dOeHS3N6NSzG0Mbs8+4As4/ebMXCUKyOcNc2b6N6NfT99FJbhQQ9eWYDWHgarJL8FkOo87RbtYtIiSN4TSWlUZ45YYgAMRusWMsJkFoqGIsqDJpX4qNxOAWrXdn+esrO3K9CosYlVMpGmvnh6qMoIMMl1Lr+wlVjEhQnRc2Yac4nQn217AtL2k6v8RMMpG36h71mdyFytgpOMRew0jgHUvje012KxkgtBzRYKfTqdVtyTouokNJHIUocq+SdmluZcHf2jSS8CVh9E+2v2K0Qq2s4oobvMGcHcw9bwLolp0Naca2JluMTsXx+XPju3HzUHy/V/KzKHDYT5CASURbE/YPg+47GFemwA9YNVLT7XiqY8+3DuwkDkNwpAW+uU3QOePpsTABhgKn2aS72ZC8/cbEqtao8rylqXe+BwDUyAFQu0x0CS3bTgchWNWc9G+Uo0DBFa/6ZccXbT5UEAuFftGHgC2ECZeFBT+HQl0OHLP2GHIYxpyec3PI0cO4/8tOQrjONJTeiA/Fn5+ITUj/XeSOD4W03HwaZSXhN+Q+tOp6eLo9ngzdFx+iGMncjjksHG7CQtpXauANG9eSBuYkCc52OwK0SeJd7lflZCRInd+kHFzeRmWnu6OSRryGh1ZmJWIxvSWsoKzsxbIqGctIamgkgjcsV+Do3nsrxZtZ1OsRTpMSIcucU52lcrdUB7LeqebJIL+9EvEuLBVgybm6VKwydT7VCkoMQN4R6R/gPKNcrucO4M/AQOsAtXcLE1HEQc0f/8/D/qe6HCFqM7QgcQ2/DsEsXZdj0urRnp1+hGthTuEomjl7H1thdNvfSb23H3o7/rOAmchxY3FT4NJwf0R5BZsdB7R5vT3tPasUrj3v1x5Cy67w0jH/CdapswQGRho26DBMKQiAds2GiYpX1aXQGpyz7Yhy1eqvob8iq3IdOpOYAYWY16C9bK85D7a3cCw2t/BJyOJFiJHmOQmoTeX1JzQiWSkkOmtnlaQBGPCWG3CLR9ChW94xuVGAsXlGnLCkP7VGebv6AJdDeJxh2v4WjzKz5REAnztOVUh5PnruK0wiyTGB1vq0rPPL6eVwRMY011BpnIKe4UqqRmvv9nQI30Ar4hl9CT0gLSkGVoqwVNbsc9ycdZJqzkBITTdb8VQrCdxithOkfFt6Ji43J/dWuHAwC3ekEUouD4=
`pragma protect end_data_block
`pragma protect digest_block
3b0702225cbd917439b8766acb78a6ac7f3fa3dbbcb9b467e27ed7811a64bf3a
`pragma protect end_digest_block
`pragma protect end_protected
