`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "baf0c89a2e089fed858ff0691bcbccb5"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 40673)
`pragma protect data_block
mRWrRPheSnqG9K7Ossko7qqR8k3zMHx/KiSvhfFMcmvcp6NBcm0QsHlzBzbFpsoQOrjoAwKevuZqc9KVhVZjsXTLyki7fqq1e3Z5qEyVsfbVyTLUBVOPP2tfx+UNvGtLFPUXj80BCoYCcuSKM+8qOQdvnAzxta0Ne+oLM5afI0txvhuoOSDOc03JnvxvI3vAvQ0ah9jD8PiyIByk3eZeEW4k/Pk9rrUAU0XXYjJMAqf+fvuGfd/xMoUTfmz5NPNTyWV/BI1iRroub2jb+ajattZC2mUemX2d2aNj1a0kh/SPfApr0j4FIOT73eujCvBK9gD6Vf/1jd0aJ1LNycR5N19v+Esjt+ICDdqesI+TUWPmf4Db8XimW6ngtyrN7uKf3YkIUaF0WYEPiNGHDa8aWua09ncJV1pVHkHzfA9Hzd5aR0iaY/CHJc82BSQ7nnSCCPC4cFiyXMDGr/Slsngt2vlRw47aGz7S/H2jrk4Qz8VqeseP8VIOinYWyg+bG7/e9BY4VDs5uw03z+u++1j3FcZ0HTRTXUhABfTiU0OEi7tFjHF4vsLZsrHwUR9UW40EHNGZP/j7X8XHljNQArwcD9MHDj2hA0EZ6J/e7hBRdBq8Oz1hFwVu304Iii3NNHMA3OwNkHrUWEW0+mWPLsqJgT1ewkAB3NgBeXC5hkx6tKuDtEEbLbil1LFFUyhDl0geLegkj4GGYY+IepPUtFBCMHuSVSLd3L83IBXGTZnYPC4x+G4AKDLFtiBdFhTEoKENElk7XlDOxTHtDXTGPQF3cKUG0lWX1DuK+6afIAisOMFNSu1kszbhFrDo6/RAYb3qs776VarVoW66uDmux1jJDIxr/TUD/IQZnpHBbpVZLf9O1UUhQaO4J5alwhtK3XP9A0qu0mLDk+Ya9xlPDed6/JorWoJ3KzHyAmhrJQqKAwOHPTb092WcrRfmqDN2NxYs0Gjf+0ZGfv+VVSfkWm9EH4uiBjfNpxmNExNGYbhB8EngEKX6czermUgFXA/NJijtWvKGBh5dB2H4Zx05nZngy9r7C1b7npTzaOqemEk2HOqXXoBGzcldtIn7Wi+0gnUM7xxshekPXkL/MH4mqwbgtWPaqIi89HdaQI8DQ1JQfvD/d7XzB5xWI8jPqoytCHbhv8iTsMQq/rAkSlSH8EjGGQtpkOCrOx0FGh8ywM2Ipihjra+kw9VpZVpzE5egatrwwwGq6HcXQrLQ00eB4hs+Ia4oebQdNZr3swnn83lPnMPD9QcREzVZ1EHbgzJ7T/Xn3/6pJfjbnm170I4Ig/F+2kyKOqzkKd90Ujulxd3xqKfPIzBEXWaloh44z32yhcKWL8XKE2GRW3WIRCBRqBj05swJzf3rTOwuAp4Lm6GS/TSIDtY8FQPXmLzoeDLZmzRKPrrfN3wZ/X7gJl7rQya7Dv1l+iFuxf52vwPd2SQmuLlod1ZMZVKkuWi6xLPvP2/EkLix/bD95Do3r/Tb99jpJ3LKeR84l+heXWM3IaP2IGViO8X37VnCeTdGLxzQP5Rs3MdkGFYH4IgAD5NX0UBGw0Ws/SyBnZCM6qye9EmJEye2TZ1B5Z2ZoSGmHiwl8rNf+iwSC0n+0EiuEdCYgLG8XUwOEcsU6y2Y4R8qVtlIwGK1+Qa15oYXY09RD4wi9Cn3AhzdwbRJlcc11NqtkmslbjRPU7ISkNOnJsMD1GIyC0LRgo2PKUoHme/G0DaiHzdHDTWlrHIYe1mSJj8QC8/9BCOtBstKNFtsjNrJvCq/yky2eRODV6LdQqvTBD6zyz5yLaVVo6QUVG0xzevmvaDt83nIhcDNYB1Sogd1xCxwYDoUuJ0NHc9Wj0dkgPLXHbCsMEITUXILLP/mSpX2Nwcsp3HJ2kEdPI6oa65GubPos50A9i82sycAItyGR+WhA3Cv5c9P4GiNA4Xqyza+G9u5PGwReNssdK3/MFTXLkhGtB6s48Vu+pFg3l+tIoC4q/gVyH8aYNmQhR4DPOoRpH3BzrgkC6TzTyQ6SltqNtafNs7BgLi6o8z97CbUZs01Mpaa0p1Sb82pFG7IioQdrmhnw2RyURB/x5A9CHpRVRlFZFc80Yc10WsbGb1u50ouVGWEoSh5PMkA905Ww2mN7smcwwAEqO/021hAGZ/crZRPScJ7bBWkOgvYfMgSqdLnJmEYQQWxeLfC0bTJn+hYXrDs7D+QwksuggBUMsGTyGm3npNSq+kV1nQsKcYBpIk37v6r1bDqborGPLSSWoZTUJJZsYGajTl5zBpcG5ACfhIqxuIl/cyWn9G40xRYlYuARdb487WW5RfmuRXBIzaXIgp7OM0wjmzdId04XtQsyxSbopxusLRFRjNzncpU2hABB42WEvIfeEoT5vd6cjG0+U+0jfWzMti6MMnekbvXjXVEGogVVkPDZQJI7LJtbtduDsPpvbHff2BAO7Oz9gutdDEwslgtyZb8L/0SaG6oiNaPQrJ4u13wTlIldip9bTIaCO8bjAYPTQNzA8OOg6Gd4LuMul+ES1oSQfPBoAVWqM9+yx2fxZEs8cF6fLmf7j6PTGa9qfYt/bt1KmdF5LPK6fEN+Kbyobl0AkxVIV0D6BzkNB2QhtFiUwjF05Wt4s8ZSEQzmYgTS3igmRazokUn+UNgObUPmD1a0pS6saSdRYDnXVRWrrjdVRJ8LlRPz0LOrM9WeFVFAZASwS+DLcjRME11LusNDhY/0U+0CAw8He+mjsn4uGiWY3zKZNWZPnNZpCyi2fUEh+euIp0aRp9NNQ4b8uKufPpDnFSHkaOjRNHxRfhd427woK25jA78siOJP1lzoJ8BmFOFWTW3PiHY9ErUeiKqVGDrFEGsg2SqzKV2VFFir8hW5GoVbnE6r9l5UXevuprh6X5QZdX3Bi2EsdJ3hBLQ87QSsRORX/TjCGVR6reoutPQo4b1BxB3hx3Pip31EBP4jvT7lTUKC/QdonWtx86F5KCAl1Gl0E+DfUEimBFgKWPcEletAenVLtz1ucr6xPzE9TD5bKTgh/yV79uooEvzXT8TsPVnn7Dmnt4l9DUSk9R13Pwij8jXN70AkqWqEJyfEFVJIhANFoo7CRHnc7alMl/AMDmRlQmtgzdP/F969qhYQSmQ7OUuspCd3VnpbvN7TbucvvqWp/RynddYjxxnz6+H+xdoWRCqn7rEwhnXjAhxLTBCBQfLS41GBHSCCdjcM6StUntcMeqZ5uctERm+nBRg7F+QtD3eoHo7ajEZSymS1Z62+qRW8qIK2wfjfathbrl8slo7OF3CWfNDAaL01+d8L2fNkK4iDYsVipTsBZnNMaDzn3QSF7OxfVixPij0bcyL2zyMgxNXPvQi1KbPVGMjlW/iTao9XHBnJseL0+QH16cyx41gu5UZBT8UAyZLU2Kv4sG9uX9j/XCL+TkWtxHvknc3TPevO9vuHANk56M2vP3Gobbr2SRgTux64WFdd0m9rrG2x8mr8mw2SCww9VvNiZr2ClmvmHc6rUoKgdTfRvF5o4sryLxzrOhr9Lhe+ibCXtcKbwEEG3zEKtUh1iVt8UeW+IckguisREPtgtuYl7/IVu6l+ynlbZV8ACUCQzepAHDQeROf7AA44aCvZA1SvTD8TINJUFWcdM7ro8Ic8fMLxjMq0iBUu1c27shXzdN1P+sEqyy6zTZZYAe+DGZdvBQQ9FSgpobr4ayHgp4IcEQumd9DkDHpY1xkYwhwE3r4p3nMu/5srR9rK1PFnPc0oAwwHYSu/0m0pwlqQuoN1HAPgepH8wiCr1TQF7zyFFNxxtsR34hTw/Xj5zxPQ1tjZwkGUYCeFXr4WGIES6FP7OcXgAG3fMghwLg1IVCpXIbPF3cS+RtEWX2UJXQjznxrba8bhG1XOK023uj6NoH0tK3O19W27BeUCd6tGbd84sKJFgE/trZ/jLts7Vq9hmw9IKakfFDY5wBgaJ2cOGMcIrt4Hjwio4dHc/Zk5PlUVxrAqFmQN+DythLhrLRK/QOOTlu2CAIknJCGUx5oWBFTHhTAICwcEjxqEU1IQLOhBWqXqsN6mfPm/WSXQJezmDZlLeobJr1AK5AZWTJC2d197CZINYdNQy56eR38sqiUy72NqkSrU0LuFLabT2TF8fIrf2kWDU0aEvlCxfEtGC/3ZGJYu1ISPUzZXZC2NdZecyEGyEvV8JDK2GjQd9PhqgtHBGvMVYzlfjHdUE3gCYPtbm2vldk9NfHb4NLTMoI+R7LTARWM0a9PhfGZxT25NIBAyH8mRoiLz/Lqyv8+zIE0UuRWHeghFLVb9AdFMcfpxMVdF4xrpXQU/1LKVsFrpJfpFMQC1w5RFopfvCrMbkubUlJRp1PEJ2QkGBprBCbhnSN7bb97VfNs5Awyl+7rX4q1dUtyYdQpEwdIDBa6RQZGoWTHuLamGdzI2tSqApfrbqX0EED2L7tSOZv8JlgSOVckmlWodwnEB6uGdOaM3598soDmFjC0ao1/CvjFdlzgdH81sKN2pP7Qoy+Apde79ndr1WMPqFi+Aa+6TgQZeMoysijzEL3WsLNrzSmHOgltW6mUiFhQeJKAqIkP5KGkGs/17+dAEWslTCHKvrzoKtBPI0iM9VvPQN3pQb//Z5oHzW3B9eskdOpOzagvzXqPJ3aBSvw1bR+pum9VzWAcqRjLZ/+j5xmIGXUE4YTy4Zaoa89byfaPXw/mQeU36Bv8B40/ukQ5wbNzSlXqf576jvlgHki0k0IDypSo+2fFgjFvgb/AEgDfDu1l6axJlOwnjwWoGVtxXd99DU/uAPgzzVKTlYj3WKwr/luTm99fDIN28WNgA2c0JJF4zinq85aUdEavZWc5swEoH/vzky0DUJpl8i+YMrYxJ9pYAM5FcPPZJyL+cndjugTg4fZNmBQ5BiONdoMw3lr7WlH63xojHHcCeKyS54m+CCuqRjYyj772rfMceGfT5FGMmkhdAfLO0DWjLQwYqncNVZ2uuctzBFwU1Q+sPghNBFhMpoBdb4fp6DikAgDkaxBcDPA7O8vd/BfnaepntKEjMPFpqqcvb2Ka9hoQY1RCZPF66cMmPDTMFHJbfZyVgmHzR7/YlKgYxb03X5cFhOAfZt8Ya7zghAfhvMErYcBYe6w8irGl5uyjBpolQe9tflSdQycWnGaM9LShv0iwNyHuSFAWA1A/GBYjIkJWQZma6NHb0e+hYpevkMOxfBle/izHlloA5utnzz4+Gg6LexT8ePL1r0ugZujuhR7rUZe/NkiBz+ZcB1mHwLI5m+9SvyJmbHaio2COOawAxYeIIvuGt69NvxRirjBhSI+J/Bl7AuLdyt57llIbv/X1TJZsKJBdVsSPPMCFm+vhMbBqPHqI40d6jkeGwKqb6iVL1k4kbcupySv57GtXSD3KVucaLP7G0cUVwvLcWVEzKSAPP1cuO1jpWLAC491Jnq2MzSLNj19iCBoAEl2fBx7WU2D1CGlDMQQlHgNHV96sjtwLWUrl73zDX4Pt62sVLYqfGsOxWZ/a5NoIMvd1bVpZdEbx3E4tZ3XrF/Ix0a2UMiAB1D6V3igfa87tlKCzrilMG+7BRsyGGPu9dSnb9He8Bh8MDmPUi2YhQ0F+R41ExYCdKwmmN/WNU4XDcGwShqaSaFKOKZZ9xiUyfIryeqgs2XZT9Xpr4nd0tdKRpMOhuWRYsGJ85d9TKq744q5nLPZCmeUbZPGHOAr3TRP33lr9OPU/qlmFl9uOCtdR3eTL2qkcAPDelRZdOXcfjOvCDwVUvPlD4iG95+sgvOc3IEcN8u9iHcTEgz+2QrdUWfMJlHIE7ERkpMeCciwSamssMbZ5syILSVODOHREv3d1XC7jVENxd31v88D4C7eWR8zk9F6IlZPtMoUhsAoj8oYb87N9dMbZfy0bs/+LctsowAfzCZGCTcj8TbSBdMP1O0kzuqCMc4JDWxvQlrbxlsLBHT7Zn5hlj6Z8QJ+7EMCVAlDbWW/+Dr4FSEjpQkD0b2SXXdKL185qbNPcwMnq7+xRk6MD4z+pyyqyCNzSwK6IpI3KhIde7CUa3K+NndCuRwUK5LVjMQeoe0hFOWZZNUreRGFoRGifEY8p7vDXKpEIaXxH5jnRWWzKzanEUtAQtzgk7TA/1Dc4zyBD284nl3k9Ak73vtUMDAvCQtw/MKAOk6anUi0xrOfMqKcHexw0xECNTQ2HpvB1W973m4TIV8yh6W7uJOe6O00AxRZTDxOLBB4GwHY8jCwH0GizDy0yjkXijVD/pIqMoJYFCgMCV+p749yXBw5tMfzsDfTjQpj8ThFrLxG3wm2ODscWPLkymOVizWaUeJa09xbWtx7oEYK7eVZj55akkpmzJbmQMRLSeo/z1X6pg4fQogIxuLW1uXwivhCsEBbfugFAYzhoozw/r1qSN1jW3Wb8WbULzFyPZjdRx3Q0qbFQg8Xr+ryl04oEKfy6clNKdgRIReabQkEhbkIYuakRBso00IJCu5gri73vKNeciIapOwV3nDUOfxNqZHeuvnJ0BD4sE5tMuSoJykmOvMvtm2QWq1X9XkqaFZXXd3c7xHaywuPlReq789Nw46e2uDW/a/1I4RNsr65GrBGWCZjE8qvqR8+nnXACOxGt6lyxR9RDmnjE3ntS/dj3uNpLlmf6OZsdjKTWQ8LI5TD64U9oXX504D4LBCoEjRAGGjoNS9N+BQHlBlBEBJH/5MCqDzyOjVOBl98JXReFRrBxTy7lvkFAVHbbW9VS40AcpougQmYHs2t2uMaO1MbKc+WC+TT/E79S0G2PuWhpryHVqT2TnYzZn1Ua2HiZXqZMrmZ0QjxnWWgbYRLGMpFXUVjkLhsFlstWTr+c0hWBkuINgIyT16YpG2a26f8IYfyKl92cjo6IkIGvsRZc+SCjqdxKioP02GXFbQpXMZ3Y6jiRFUcBhp3DENYPEZ5oMtuA76tTcwVX7mbaK3fsi0fSTMIeWXDZHUP9Fbp8KngQY3FAWmTY35zEQkTVqEIo2wiJhDuQcpVnsjAAaaML9se9Vo63Rxefc9VTXkdjin4s2+F5gDVNTVQW6Z/4j7HjR0ugWquWsiKUompBn4j5qDmWOwERZGc6o6pjvJRDhywnSXrAcu7/TJV1/NqGQAB6zVKgBZEqsLiPvilRSqZx93+1a0mL03COBrfyR0QtchzG0J3DPHaj5d4jW4sN2eC3IFrH9gtifH1vth+TIxaVWYVtF+SiO40aAXkv3JfxF+hXIFW3BA9N/gU/IyFPcw/0Vf+HBgFzunmvTs0Gs14TWMaO7IrQAvAp15prHY4OPsQKBnuWgapfX5+0tOlvh9+hMa8jHI6yytCE7zz8pLN/fl8bAotHR7VGWzaDGLvdq90sq4qyPpl+2NrlaNsdyxYcPFprbGixvUls/5qJe3KaDlIbzUT4/9b2AJ/UFzVMTi7WKFUIJC65zW0SF0dpoIU1gpUP+wn4Aeig6P55ua7WMJGkVJ7NTJ7H53pk7TX4Kr/NKAQxHuE77iqHn6blyfqP5CbFNEq1q+fDE0lQcWpZKAZGyYJ/j1BJN+lFUCxC4qj6UQ6MJgCZY/0+yajwWGKX63vA1KmuRVNv4ZauYKW+uia3CfX7RPmHErTvyv+jK0KEOWvJPTUpwnQSTegwO+uNMdcTzZTesq/gpcL6Uws+gp4Mj1rKO3P3XM6rR1GhcBNtf5M9xzY7SWPhJVS93n5jWoVoZ5C94+027NOnY3L3qxOq56HeYDGTCqzc6vqKWf27JJ9m0ep48wQEATzj6DLKmY+FKycda4DSaEjnG3u51aJPETHLxA0xXlEtHLymhg6UxNDGwori1K//JDoM48oobHfw0eEOKyKO1dV+STyirhdAqTilKzz+wkhAgUUE2rlR7Fho3r5J44e29kj6jTpUiFJkXJfE6o+//8gYDhgHM4IP5pgMQNC9YGNHRVsaza2jwbttDAmbtdi/tswrwDnAnS+YzJecnP0NwDYvvuJSSH5071eKmFXpyrumhMdUZRodzcIJ68z5OV7CtDH7mOAn2fxveYq0+nm/nMtMJ0mtpfNjQhe71uJrC9Or8xoPr6iX2Q9IDJ8Ac0DcmVmGGaU6wymu4ZEShsd7U9mpojD7zba6xnDAHIuh3EyCoKvmFe1yJ+DSesfY1bPLbzciFGsg9mGj4w6sC4XlFeY/spEuCqeVisETHdpvtFKSu9GadEc3K0K9XPQQ9q8StsbcWJ/GNNJEHMFl08XYPU2z/UuBfptP5obSeCf6YuSNnNWBWVyggUjwphnniucE3x61p1+/aasc/LnYCSFj/o2NSU0CGwVBO2lIeRgpHxSXSbNG0FuWcwjMr/YFCa3lvD3Y7roEtmbUzSpotLKEdFWdliYO0i+2eqtc7l/zZmbgfZS8zzNEGalBtb3Rc7AdPpivifLzIFYUrwDmnFXXL1oU26T4D5CJNf6VFExIqsuoWcOZmFOhtGBmUYef2bSPDI0u9v6mq4l5ciM5hHR+67ulyFecu+Jwd19N5fI3sYyoBEGCpxmfPchTFv70dDiNK69jsmNZCxKGvb825oLi1wXdyqq6rn1CmxgXH9PMaI7l9aJJzmpm77gvYuymSd8pvIgWWPaBlmA8o5OI0doo2J9f1P+d+9yLBuR337x6yWOxY8Uf3fJOR6YzDO1CEAU5aT0EWfFHLcxD8ghKhJgrPjOezwUkzX0d28+WMH5qLkhQ31wjz1mVv/D+pDO6I6HEqbJbYCjD9zMndPQSGHrq7z2VisKOxmOx6qNNPjwp3Ti0S1sB+1ODh8n2QYUsYQmsz8tYPQWHLtEOKGYUiUNwyphMH1R47QfEwpGLJKY5sHC4qzoo8NZs3tc5cpGg/tQEv/4VSYPKP9r1YPCUasZlx6X4G+GUCqbXe9A9SQK7Hh6OmI7uarUjOh5dMvoBdI5S2nCAHc45F3ICeL7bJdUX/ZoZQ2GySlJ0uAcNZFECD4IlBEcEjCnYR7ye/t5L4Wib31qQ6oj8Il0pQHPYV0ka9oKkMz+Hh+P+wSNjvYQPeZS2+hvAUIwYIXs54q+k5YLH/JvjIIHh9anhwR+LWq3Ww4ZIUcdqXxAlEk0AAXg8yftA+0sTxz4B5vZV89czlJX/GTyceIFw1UJNi1+Ij8Qw4S/4o8mOEmVzVKRjgy8GrCfMVP5zb8EqBIxNN55hgrwfwy6NznwicPvoCnhfyadrERV0fbrL4tLZx7nIPyJsYxb2nLkL6dIcmNodXa9Mx3h4oi0WheY43y/y1Ir+/evdXEs7iNOUlFKMNwSw5G5UUX6OJAAqYbwXGVAUvhzgKpUTzy9gbsxZ5md5g3O1NzxiOpzb0jEsI9uoqzuaiLqfUy/PJVebjdQwgw5bB8xQ4H6iTyBdi9SQSXANtmeecopnkFGn+gUs0EM+BXaOiq1RYyplOKFv7+ztpE5V9MSc1yn4PLtU0un+v6QtYaoHom6SG91kluE5gegNSBoKDbSUZKzhZakv/tYDT2VI/rxsG48BRGrt0QpvdvPI9IledlnhmnVw0kWVnrEfYwx4BLbRxgFmwNxoJabXB87kDukQwIEOe6TqS7nwYyGEO1hfBbdf69bAj2ybMrXoXhr7ENEjIxCGhB7/VPZEGJzAgWXhLwUx4CJoXTxPOHgwF1V2GBjdZtM+jgb0XkT1uNjL8Sb+1BGQawDZnLQZ1smGbTv1Mc+oRVTep6hA0mE/3U0vQ74FhFkSTPzH5JA6mPwKqWaExOZNVJH4udUsrQlukPx9tBpwP/zgGNWMdSf0rlAf2aPP+io7SFAedLL9toTXva6Xn+T9BMA1TbDAZ6iltLvl7ggAsSLL7m9HnvM7Ok+SFQsT0+BodNNvQv8Er8a7Sbwvp0JxoxRR7sgnknSf2c+o8T/aIPcA9dLEr3Lp4j3NgFB6XY5qWomea5Pe8B1sSMNNrY7A3Zi93GUIOhaE4cpLW3mMEJ5E7WVfmERoaSAOu+YgeGUbpvZoe8jM6VeYARmrG8zhSgoyA2bG/gufJYNFozscvRecEI8TrQsu0LjQnRHsSz8zMGFEhhJAR/rXzxANG60VdK9XKMUD1CAF4ZIqb6P/sf7ggntdWL89hfeCjfKvjF6F9QTWJ9JghTMVOsYkubdhbO+9mjPOc7bDG2ciBol4TdkkJGV70r8X+t9Z3dJCERhKZ4lYgFIi0q517OBL3CE/FQ/3Q2lc60ciTK3x+Ojnnfx1fieya/FYEMnXar0Smw4J0VPbsiYAwKyUfTxc6mt8CKq5DXqq/miYKB5/eW19JLRD7wJMsfYCXud6tdXxF+8wY7XoaoW8BEDY/bYbBCJTkqIJQTUjB/ELyAqsD38AoBWwJ63mIJCnEsWtkavLkwEYN2TVaHMRaVdos3MCczU+lmWKG+TCm8Sa4CubvNsTd5rNQ8sjGqOfuGl98gNTejsF8Tq6WyQ//VF7spgW1NitkXPPGh8BW/SizKpWXNbqMjfgx227d/edYvW02H2EjzcXDF456nEGOLbvAA1GVPpAAId2B6EXv9xHMvHxZQLSqBGPtKofUULa+BLNuElHmdEIqP/+EVkVsqALMXKm3P1iUJsS4lNTIUOk3zu1F1XpLeJUuDSgfVXh7ftk/rDrn5O76xqlHhJyqnsMZN+u1nBqTl5DLLlshh2uTrH1EsBi5aMDkaHe7IbxJYVgVw6NMBUni8OvO7o7wAcSf71rhjdk0Mldts53h9KEpifav+WqcAP6bQiscyeRK3XUXw1YmRPpNl/GfCFkjMLJlW6TykoJ0guTbFUBLLz0Cxs6AQ6L7zv6omwoMi+GJPnN4uu/M+ShfZyxpK0bWVCj22VdZZQouz4ysEHTog+DOfyaYX0aWvFGA22KGU6oXIFChIcP3KaCLX5jYhAUWyNcMCfFALcA9qA7LMN3iYzI9bZsQlMTVN2iVj3ETvFsubNnL+ZP+vORGo3VD0M+P8xRXemgjLzR+CxqL2V2kVC8F3VYW5TP8rhRor/cJ0vpkmGK6I0i52ggvWNP25dwrBcANTdP5uT2yyur7huW4D0JolszGYw9WhPr2VU+uKu6W5CUjyrtVcTQaL0bLgxvudvl+Rhmhmrqo9KgUsZc04mVZjqdNvnIZNyYaIq1MutHgpbC8KEhsYGRKGY+hF79LTnpPyp4CZjViK43RUQNkpGeS2XLY0Y/kk4oFJZZLuJfrshM+XEsVfn7zTf6xBRgs5WKs/8A+CBuTi/xapQuln+lmeoEulyK+Z6yce6p9EKUoJAs/FmXhU0uQxGNWOQi32aQkRfnOOi5Dy0ve3HCoYIZmEKucMTmsRT3/JgZJqjNlr5G701YTXT/S7ZXkCpX+QGY3a+EZbDniZG0XTyK86X/Cvsbe2qOcCwubVAoYrkm2dzvOgYVK2YeizzgBcttzfIroCXrFzAGwq4q+ldeYCHTClpFx2QX1mRJHw4LH+xgHFE4V+lUnm089VEivAjSJ4+i2zhEeIHSPzG6ed2KjmTMq5uPrB4oBlFL9jzV0zW2laDICL9ivIFjeTI+FLGdjHo3Pj5ff/4BiEfBJSWRAH4dTtLcD58DxQUp1LSI4HoRePUgJ+ipjggIbtwKXSGV1FtP/rc6YaSQCcPz8xvISYL6HoqVXJ689n6m5Os5ptJ/Wg3Ai0Jp4mNmX9IBx0LLjJPb+7577VqVzpDm4D5IKMmqY3dlhXiRH4+WMxe2eJpB+rZ/QQjfRfMz/b8u7Jtfk/8NrIn0RhQ8kCyCBmDTXWYpKe+FW791F5h1aFBSYqW9cuhzio386Gjy/sEaj6DYRHznYcMY/dxl0giFQ8BPh8evWPfQfcd0xe7XsStG2iQNm6lvnWF7IjQNSeH2fGAwXOjX4pvYuYrNLtf3J+1RRseGIrvEqTxGwqNNj9NFfCO/hWGc/mefp/NGBg86DuEb6/K0majuYw2VeTRLIq1ne5QMpGLaIGcVIWCGGMORLb7H2T69amUA3k5Vs2fCn6rxB2UVYHDZzpCfiYEDAjN6AUYybRaoSR7/ack5j9m5pQWJaxCmpf07KtIJdBkBpjN4UU7piiTReq3ecQQuKup72EYOiOtspRP3U5+i2xFIkZpIF3v6Xpg1cwqG0f6cgnGJHA2Lj1uIbdSpxPFlrVb5O2f3cf5NeuJehtb5fx9eflaLyzD2k/XLE+EWZh9s34uK42K2W/+Wo1ie8vwnF8iFlNJOvRGRnGvqb1Rlmxxjy1iEjj7ft3856RCyhW7g9YNC0ufi+JavY9NaRxx6e0tHV0vnn2cgwYwcPwLc2ISPPea9PhG5iHBrAQGYv50Tk2b4aHJqeyxkrzByAjgY/D7vU3RAKnIirBz7n2jtdggp9KCSJPAfO+vwl61x54FtCcVBw0N2HoqDxfU89A72hvpQde3vn5VgTmXNxradpKWdABUiIkjcInXFTYTCSYIPN1FiSVRhWqX9uQ4jhmtkY0tfzfOb+Z6JQGAe/6g8750QTbxikShtsXF68FE0keCcEzS63YdisM/upAtHgF0SCipkdrEF2ctmpbVPBi0LQvlIYIiMNUdzx0iDVjddrs3ddAs1yUPHLOVE5cO0yy6lDzuajltay1qz2fP7icjUrWDjDrdRanQ5nqJSoA3g4k1+JygtKPQeeegZnfgTiV9caFsR+hqpdnQDhoFHNa7mTksXMfu4fMVsbzgFLNBCyLuOaf536zpRHPCO8hxyLYVWcSGVxge/RojkGLl5Z/1Bsa9axi07nt/bmX/aViQY/pqQ16FATQIL+RsEVFPywSEq1MIsV4o5PWIQzlhENSdkMQED+mgtkYu8Lc+lLbylptfJ5kzTf/QrpxWgQsmazM46n5geOETKkpAdakBTMPeYp+z39oUcPWvY9cKdLD397FGsYJB1YVQsuSIfPid7ys1Nd2jHYss5i6zBlVim4ItT42NLrPTYfl0Y/dZl/dUAtv9wgTiqiH7ikBGojSXvm5J4i7BUtoWgRRL9ekxG161nkc05Ost5Qbk5e+Zn4GhT54yKFhJIItfreH5lgaAzmOjiu33kRic1LGr0evlxKCm1Z4h2921d0RUi/81JLRQiuDSHKJ5CVaGleoRQ4oVyPpFb9Ji9p/5ZpXJ0ysEjpLgmJ8pvXzEjuWuZv5q6+IQMHApbscLOZADNrYQg5WgXUVPNrvE9OhK/pFUfYGgzpzteiL9rW60wCya4HoMJlCCQWDxXOHIsfGsve+s49dLfEP8VA3/ct3FQ8eGgsoxpCVmoiDpr5oyolfTkPUhAPxd/L80/j+mRyKg6LXjmU6rWmRsovc9b6tHlJ6Bdw4MTdRXCgRCLCklb2vfryY4+RVQePxmRlXUWlwNT0yliN2S1j2s3spyY8/B9RXIdS1U3n2Lu7htE51f4YFB6ZJDraN7L/KsBF+po4+g8G6wZ8EWMpvek3q9tnpD5GfGpUD12gW0+JtrgR+SWWXUxpld1UOpOOyTk6axaNfi4SL5vRDS/mQj98Y3+AleAC53hSIClZ/JlCQiN6mKkh18wuTp48qFSc04V5xcD12RurWK8Gi7zzAL8jH3w2UmLMkkB0W0NNKBxtRq3aReFCFWIOW0it4C9dkUGxV97vWlX0tH2Q+f0qdwUb+nQQdl/ZtqzClvBJYSOEC9j79rNgpj3bT1IL+yuoKF/E57MXaa34JwOXgKpeuSq/ME2FrIvNONlM8AJ7eijALI12TxJNoLQ9k5uK/V6xpU0eeT4zSJhSVL+ssG/RIZImPOcCSxgZQIesPWb3OfHdynNA1RETM6mffhWdaHcN50M+dQ+Xqs9rJIczVJvvSsgiYryemCuPChdeshu5BhYZPm7TiHGEO6TkdG8fuVmox5ED+QxHpmhkoZvfP615fruC5akHl3DrVgPVaAR4XAQC8At/zvs1aSe1iaMtrfe7ycFtukyP0fU1oHj4U5kP5esRK273tlypJ0Pd4H9ThlULNdvQDwukGL5f5BJTTD6Ih7R5zo1K4rJtYdp01fS/yCedTffQiMIxpWqhBJTrvOSEh4aBe811LRuQWP+pQ+th31IpsIaOrl6Kft73vtJSYmU0nTaBP4GA4kQ6AsTKPgdAD6Y6BnbSIsyAi68JLmAcWrMJjRfL9dD3PB6ZEM6bncL+UsUpMHvna3kUY+2APQXO1BJLriX6plKOHCEbrJcQNwLDqtJihUYAo2hw4cMJJpe/+09GXt+mUq6K8qypUqjHnvOu+p2pPsB2dq07GIbd+7kjLNyNPhhCZaXbB6Sc1cv8hKDjQWuwOo42qePKtYgRBQ6cwR1+1BlTXFuErXTs9vaXw4M8rsfv1XznGVRuNF3ACNfBkaJ0Xs7iv1QtfUoE/IbF69AHAfC/5GgkdIIuOv2xlWrJl3K3+Dpc41PQFKR8VqXblGdE1ZK7WEwiu3ByCT9shUF3WW05xVz1fIg6IfLeTU41HTyEHh+fYoAB8YqFzmC5yx0AE7HQuSJuMlF7vu8TiSZxWSjthOJGyUkyfdrjxuqJMM6uFkO6hbdnxtLg8if6JkUhIUj9It5uvjt6BPQ6VSejl19SpATQMrBzahqB9WEU0xVqC8ZIjWL02Ux5crofmkiexD9685XlB5T6M7xiGaivTnQSfJLQkBqPsw9L75eWqD6qzaxS6i3RelWnSTmr7Gjyml6mvx8shkVLUDt7U2kZR493vODlElIn2dzmyWYZSKLEofZsypQwed90t8G7oNqi3RKZMPPF9NxWAIgQFJ454/IsG2vHmFpd0DR4uRoYXeqkyxq3bYym1QAnaCCNmbTvrFJ9L7YzSO40zee7UREgHAoXkgmRc7l4/xHH/5iJK1oseA+eel9x+6b4NuoKa8jaOa0OU+YP0NIAmFkskft58IWZd+uObuJzINnoM3kvkZLtKIYfp2rzCvcLiL+XWXG2FfoQiRseyB75a+mTMOYAfbp77SX6ROI1vc3IOoup1/GrDFBZwv/dC6MIPRlL/zarvRI0BReFM3jPyYtKpcpqF4jI9AWUWmfAB7FwrwEJ+weH+Se9NMu29bYP12F4GfnssslNw1qkCbFm82vPriSp8MGEggAIgPHXpaeoki6nHFQnqW75gMfV72T1hIfXWNsL0ddUiP/2lEJNSVMCleQbDdF0oozbE8NY5OxSAn8wQknmrbCnANUpo3eoIal1YjXbWQ6k39CLZ+yFYFXkUnFbTqZICJBrjI2quS6BTta1FjenTEs+OYbCmlY9Gy8I6xwGt6QyDHqLUHiEUF67v4Qi7pnM/cHyFALA7XvqwKA0wr8zRh0+9j4OrDq6NXColeKhbGV9lqLg9lOA6Mv6nV7xmn16nTEkLsvuE0Tlrt5AV7TMC9D5vbWl97EuQujvEZSKJyfRR2wZGJrwtkk8JI/3p4CyT3pyiEsU30vpPI5vlwbWBWG6PXC8UZUftAsiiVEkfErqqlTJFGqDpTLSwgkBrjDHbe0rOoPGAwAXYWVvCnAXrMM96lqhsbwqGNfncVq3BhqnCHxqU37JaZve2geMMF8I7HqhPFwdE0f3OXUTVSCENfXaoogOQA9AQBAQS8/Ix/z76t/yPq41VA5egvASatttmod5Uae055BUCdGmtiXeIIuqA9WDWZ0Pdi/5Y6nj0RQmQCBZEpzDWIJlBON/4RdlqmFzNMQDVohZ/NFfEju0ZjMlzMcuHBb2LjckhyVOLPyuI6W2T0aHeht7HHmSe6VdqAKnOQxPB838Z0eJC0i6b8f3HZe+z2d9dec8QZmV0ESDKtryOQO/XjZ5dgqO1OhyLSCD2iKq/UXuvKH41VeRLmo2EuRcRWps0CFmYESbDrdloDchOTzT+YdlzvU9jS4p0zxGrLYTzLt4KK3Fhb4AtXx6LZB4b1/OsO5t2x4/3gHlpd01jK5hPhQa2ln4odEGRZ4FDp1rB6t0hDXqsYRzSryeKAAeKwjD3iPH1lOTGDr4x4oSNN2GyY5cdo/aI91PmfnkRx2xkR6JL8uKvJcrBr+vFlN1eYMgMldZcbhKHpPDPQqOvM1MqjxZHoMtYRUUorxYG4G75QqHf5EMocqQ3wsITuZp4LL7vt7aS3CkqBGhOSW+oQmhHKu2Bd7Eg0JjNATvkBeujF/QOcZH5ZM54wIDYiQJcFQN4vuQnwOMRxK2F5rgOphWCHHSxkW8HpFikbB3gdie55txDtcOWKIypYWvglxEQlk9F6O1xNP5li7/yOEL23Hw1gU/gb1njHMcjW1Ok8zGnlFwnuZ1CSjFglN7ejKPMbTJL9dIB9+WpOIRFOC2eIakxH0Xq47iiuuzu8jiz/rqe/chB2gOKUOMGqffXnFB0ElWulLNhyOdz/wo8N9f2mgo2TxRAxsgx52X8LDTLfjioYhhuK6968acuHViR++5VlFVoj8DWLvZwl7lc8XrrFub+aCQruAj5ME+f+JNCwSja7wRA7JMqzARabGhkx37RvFZrK9O3/pzrqt/4d6wKdCvKe+GHtUnQmYiDKQXyMv5xAthHGJWfD9sCFCUbYFDHop1oR34x7lHwG/lxTwD1rnHgPJ1nGFiaSFO+s8X1/ET6B++fBIhxSKSuJI++rHcvKXuMlzSZ59XS1f9qHegDjoYg3v2JjfeQoNStcmf59qXSlrPp7CTBiWEa6M8efWzFPEY3zHLp2O8RSBwBnnc61Pm9pQDbLFHIt2VWXm67Pl1mfUI0uNQraWc1U08go0ielOyC1Njh1RE71NTfWZ/CHXhIC2P8We8iyBFv65F0B83en04A+sAZ/w/IGn244ejK+dtn/ZL/fo/PMdLathNvkGfXIAcKJiML0oSAlPamz95ZGy9BRgMv9Zyq3bZb8/IEsc4L9vmCZiYYC/e0VzaLetLSYFPU8n7YDOp3tywNs0+vjN85e8ayjZD3b+sfZ3xXE+eP9jk/YMzk7xal12UMg20PNn1nQ+tNaAQnDhhefJ2hBxtiHEQMh1NfVdwx5qpRB/Gd8DvHDcuI9iFFbvFZl4zkkFYsFZtz99jMsDZP9OYd5tZOT6AJFZiOPjqB9g6SEVXiFCz8sWGdwKhntWwUaNb+wCS3gTIDRlHnRFFV2tyKLhVfztLrMCOe0CtQNsnZ33t5omJlmJm9b+xZDSvdxecuP+gCiFnM0YYjuBV1DXvuEnmrFsGfBcjGSdA0gP6HFarqpRRiu48XQJHHF4LC/g7ZA4ScXJs8TNINFQlu9fnuH//qWaX2Hct88i0UtkycbYlodc/8H3mjGiCQDBs7/yfWpjo9Y1q7rXShWQgyv4HDy8umnl2lCqMpEsKzbogCjAHEomE++jcNVB2m4cl6+a0ThZ/AUZ+ml/r99PEcGxQw6y66/yIFFU2tY4sNlhSL5055zyexbsy6iyuH/0pYDMUNBVTbrIyKmC3ApAhBQ2Vab992rGRc3X8FC8GaD3a6lugrsdvAXoWxzSqGhWv90e8oGn+YuWlUBP9+pGfWDdDiNK1kMYvQ+jXVoDd1eeh4hyReS9GuemdkBc8K4XYfW8Sw6/clkzKRwEMcLcaohgJza2syt9iTEM6JMlthmnnRUf4xnAhdwYiXaM2WBOiE3CaqcZHmVnrp0UrmnKck9GA4juZvmXAiK2gf4ET5mJpgSqeuKWzkyYoo/XZMte1iAaQKaLSV7YHqAPkJWjoJ1ua/CoYM3iBi3ozvHPVyEiD1oUZrkJLSXOQq+63zq69BMjIEZBN52+kVD64pUaBY9HL+5pBMmOZfWHTn8hhszwkHfbecsUUPmpi+czDVNpgiKBRyCwlzgF9jur+31EQPx6NnU65SLTyMeQPx3liJWE3mWj3wpa67HfPWf7SIJyL7OxWELWKAp+y8v+qNnuLAJruL0AU8JQV8bGlq58ROuCbAynfCsjW/3E93PU8vvpclQlYiXg8dQvjsNQ+nsJC6eBvv78WSSYdwzYjrQqwsBmk4wwMwh8QqWyvJzYJ/HyZIH1DWXdQRnY/Jbw0VJo6fmFpX+IhUR0IcoIywdPXeIT6VZHJBeppuK+ndB+mvj/E/2yb1wpFMGTYBQDZSJbjkZaDG4gkCaQhQS+dcEtUxdfUhDHe9NOlcv6UDuN4Lc2qct1JU379tt/wMBPbi2Izd2m8uZ43rREThqjdRBv3Sf9tR3muBNcDUqLBmnnYmHDPKLuXKmZr+XAJ5BmcvEkH2yHpxXaoynXMcw5euanoOSfObIh0LrXIIA+8o5gP7rBDD74pYY6dTB1AOeXij7UBWYMnkTk263fWvlzlizw/hsXdGbtKcTFlvTzlcT6x1h4ClvKAxtbVz5Du5O9ZGowhHXh3nELvnnkX+0Z/9ycZJ8wX2l1vLce5HO3GcixsKqEEV8i6dkHEWI2YXWqkFa5px6BT98om+JN/E4pxzY4fztGMS1RoG2LPwYQfXt9D7bwb+vlE6sZQxMV/2bsJXe0vCNKj4/IllVqm83bTVzPKIQa5pw1R7z0pu4CjbXKHbizeKbUgmWORekI9x56A018jH4lhjymUhE4UyLeNKS0OHNX3dXSO7Ob1I9rCXMR4qDiEYmjCsKit9MiDZR6YLGRw0FFRT1X50jMGablyi9raGDEHEPCxliGsyjLkwNL6IpSzgxDs6KHPO2EletKUHtGFQcXhLsHVeNLE+3kevi9K55MUr9r7Ol9txIL3ZRfsCLx4hRULmvZ9WcmAsCreapa+Mh1NfKl3DQUMpovnc2o/kpFb6fRYgPvsOC4rN5EXjh4tlkufRaiL7fchXq1hNB3DrIREWJdvm3835EEGk7E+JS1yjnZuz0/0P6arD9IwVsnJ+f1E9p5y1k9mORzcVkZEVRF79ltqY6UACHBwtSpddzOpEQeczkQpg/F1dTM4H+HVQGSm3V3cULu6WoLeO2srtM2Zjxb5aXi4zuXGqia/wYiLCrqoxYldWzdE5kUfJydvhE5n8TG/bVD0xIVnEaoevp3eEI3phu7w3iy6LFz2WZFnRcmlyVIMQp2Clwg5HKslcTCcqpyZt44TD5bxMnlVN8tiJMQTGGZEveyKyac8nOldgIswr6jCtdakNsPk/Lurg642hsdekcw5B09rNKLmYjQlPBEB2eCa9EOCQb4UtPUfFDYF5bCid82ulWcJI14G12rKj02xiAwBVKot4wuONsxpIuGPXhLeBJwTCYaf45yNmuGUoRyvdSI0MZXaTnWf4A4HK51NXr/dWAN+MrsNcVy5gvYZb7XuP/x3cm7lfuGzXoCsx+TeRT0nG5M/ts6uvq5n6szHrhUoVEpFVXHwolBOUwlWgsr4oXyjWkJOFHBB9lJMMNyZfy327JmqDwGaLObOApide/bThZaAfjNdANEBMkVakN8ZUP9kOPbMdk/LI480wTsgwaBe06eKeVK6GLboNe0RbHaNGx5feljTcbYf0sMUie/glkAj/JnTSr1SiS+LGNfzGB8sokQ+TmgZS6H2hnxVaxWI6RmhCYVdJfNek45wgm0fkTbpDdPwq8tMtn13YHx5r8+4B3jZl+fKA6Mp6+cnO2VwCe0aReyTfWGLdx2nhwY6iuIg8XYCXnEQsq2GlHVFteRT4Gud7pyxnreVY9rQCpDH9oSRJntaSPisW0+0iKa4D7Ah5iX6e8jopc959YZUSvlzKgg6HSj6lANfaBTM26BrpthRNrtL/NsJWt7NNdSXvnkeSpRw26Q6tBdJtQ5ZR22EX9KoyMrsj978BYPdaR1SoaDG/XedMM9qEpwvRZoeTRIRARfPPTdyuT2N8b6iZfoc0Vokzh4cQd+CmGOZjOoT+6Hr9w53qKK5J3vchlmRnMQ+74kU6ZvXpeq6VdP41zKDaE1NZpc+r8o6zxOrwpfyhn1pkG/gUurXsAqT+rRwjoXuTmGW0v/tGdrazcr0DMewD+058n32rB39/DPU36jhWOjD74j4spTy6dddCDMnZuisLjREohDHq42LbCiZBWnZTTGsm5/T0KC18yKsxldIcoITxDZChaD0c2njO/+3SF18X9LqQtW8S2shaD0kC/SlPNfpa5C49CSOyJb0Pqf8UIrwBF4g99vDzs5lWtUvI+ZcPaq/sDnkMg5rEcCvVgtQdeZGUULmRw6m68jgWIdi01YsqoIDQgSU3EHjvesOQSb8gSVdTu+VxwQFbXpGFUto+W5qjPB6fU+xeji1QiTEwSgS7DNzgn5MXYgx3eJ2+JOjDGalrDOG7awUjerYCs6gxHrZYt8YtVp27LSRpTlxlCaySfARShk9VTxkFKTv9b+JHRejb2ELwvU5Xk2q584dWSjJdG0NEd0hUpV0IE0HjLxmT7Y4DJ3eOjEpEdhXqVmgEW1Wf0zDgXoVvipx/b06//5J0z262hwXACKlpnnnNVGL4/UG0L1Tg7Fx/RZ+VwzXuzRXrMMXYZoR1lZNcQk2UiKLgbH3bFPnOuI2E7peYf41fFckUoGfQ4fH+NJNkzOuyyN2E7BRbFQX8tXPJ6O3Z7ssyqXzkrEzmng3j4cr9GgtBQ8CksGahC4VEG2DdZdCsZ3xNnNdrIFyKBAstD4OGOPKx4q/NUe5+aJOHYBMST7+mtB7cE9jaW1FIF3tmDOl6tcX+4lpEE2HZy5uCfmJR2qQdoFD6X6ZynD7i+0BvWMvbvOaZaWN/9TC+tUTEPDfmHwXPKatV+DpS85Ki3j0fkz6GznrFxSXZm5JrfsjFfyIY7rYnFMnWuG0LBih/7LXTGw3uKopvFsZQIN8pQrDHf7+WkHoV5IQZqjltV6TJe+dA+y702kHzP63gxG+1ScCduQKHzYRI5cVqGdL4Y0oQd2CeC6IGU9yRy4ZUG7oz53z+BDM6mJSGtSljCfMHY6AFnTX1yiCZJLUsppkxg0RzFNDr5tyShN7Mx2HoOyZWxGJD9elC7EdLQCR8ecEhISc7IHZX3UH49nA1unYkvMCu/+LA5nvx5avzQAv+3T5CH/h7pW+2syQ8kMwvVtnzhNsxlI8hWh0kIqCpfeqX0Of5gph5UMcbQdIwWllP4vQRxOeN7iEhZHJ4iJu5qJ2CgcQw4zn3Wei3uthzo2BJc2rjVLiODod2kNOXfpcDHCNFLZYAON21PpTn3I2OCzbO5vXxNbtHrymNUoruiaUSnKxIRGZgz3tHkrvIQ405AcwyyN9Rb9Acy/meqlyK5jpUEMiI6NIgnc/dcih+h8JIGxg5rQ5NLbdo/M5DB5O1X1f8CxC4erN97vvXtvCzkyHclMDGYJA/WqmVUVaSXZq38iTzG2R+PDlhC3bR8OEwFyAAb3C0+sWRO9U/Lndr+USDIui06GWrlkog0pwZXjO4O1YAKPPPpvEGVr6DtniN7GPg4/KSIPohlH71yD84SK+Q/Co9YMytpB3KxoW57YvMicemCxKdiWDECvEeK8OTcfXznKVimnUeVmpB+idql8ELM16ENeXXYe1+LqbRFM+oUaimF7P/1J8AxsOCyGouENMAhiknUcrK+CNF3GDbhk6QS/GWN7PFuqKE8ELZ/5l+NUUIa5McCSX5oc3oC8yUVj5J70jlKYLdZUSNJ8rHE0MrO8M4cAbE9g5Jo4086XOc76GYN+1zc8ImJ9o5iH4MBON1mYvm3daa/+LZOiD7zCcbgx8w6sN0VulBoRXbu7M4NtRZsktINGusDSXOdcXvv8sqCj6bQVh0Fllv2CLYimq379EZiWLnwKAoN8E4e0uXqN2F2Tvp2/lMuSDxAyZFQRzj21MS4dkX8/OgAuNLw+q2o8K1o3YHDyERGdHg9jAbjjUBvmx8cjQ3lY+8WsZPStEhoPbmmZbeDkTkeotdH4x7iA+zPKP8QLPO25Tiz/wa+S3fHUtud17aPfH33VaYuSzV7DCR0jutY1IfO61MF86DXw2AjpzJjWmtH4KeklozS6wh4CZB3AFqRY6aT+u7SgqQCvGqsdOXtAkPYto3YEzX5ZN/P6YeZGqxXjMxyyfs71njU7YWEWv6YkjY6FnJXma+wlE3sVgW8w3Lq8OzbwSHH0oZLmJFZhK6LQOCRYLiEFExslcKnObVtzqVEhPNjqtToNnZAWAooIAbhXa55zcO17H+oSV6xdSZcTg1Np8KHRBTeHoY1axFQe1yp09gXp9jczH5vM3HL+gqgU6QX/qtdRzta9gIrCiPB+2pO5va9D/y1OnweJ1ieB07biCxpImYtZgM7/tcJjOO6Q+WO0GSZHz+DLLMbuc332YF/tHI654GumpQ5kSi32grq27/meyjxhmaI7sOJDZuYKXWqu7aCiQ5kX1GRTkaF9n6HsWmmIuI3+4OGErZk6JyXZjj0ZrRCDn3K3dCWC8hCu/SSNQwWUg7X4iDxTLZZxaZGN//1n9GKpYtyavVjWzYj4WtMDnF5hADmCCtIreE745ZKK/rRKVBFUrdZ4yrPHquRMp+7xqtDpNb3wmtj5uKLy7KoD3/B4L050mjph2GqECVwgTZsMP2botcnx0B6mVng85BI7qz3bYuhRPG8ipNHT4o6QE2HnOhl7HJvy/+3MkyVu2fijT9qNj0HwOKRQKml9A2dxj6xHaNF4Q3nkQuOxEbII0zmpZpvTka98ywFzeJ8SQRZvL4PXwq9aXWFuwFkQhCCTWl+COqbNa8WE09WUE5f6BYPinkFXivREJwEMhX6p8kjxMNLKZn1Q1pu/J7htZ86YKQ3YHqIcITJXVbCcrly9j9+XWcyP0cRl3rUhCZiN4eL3lT9cQCuipF4Xa39FAs1t83MWccSdNBzMGuv15MQPYDeamvb8xZtpnUl2KoYwLeJQ69FZ9bnl0O+kjNL2zxQIBPlDoR05nlpcV9T8dXGvijr63eCfluKqzihIePZrKSTmFd41Lu51aIn+wpPG0gHjSFqPlyXYbJJ2clsbRa50lIBthbsZauJcEbk1d4F3mk7un/kZPTOe0eObtHm3vi3BEFoqCxio3RgWwsjVXwi//D+hvKFVW6r+iCxiXsIzmqn3e/FGbYzt8YCntatZfBCXu9WvMYvDBxliD/5fQQLfUqbPR0iuY/XpsNhI/B54tKEyvJWsXThKvwfhjhrTBZQtwJcYkAVn4DCd3X0HHQOwju6cEUgHMxd3xFfKNQFyX4ZANhVYqGUQ5nwUA4JelRlw0LTJ4ZetgMg+XNaDXR5I6/nxNKLwqDOMDozhtT/7NxEZl1EJ9iVwRyQT+pIniLOhgm3jEsFM7kpF1ueI1U2eoONytne6AcMdHZBYBV08UKEwd3TJ3UPB15FMMTaGhJ81Mp38AYJSF9kDdrp/YR7mDJ+VCLkLVg03RSl6f8mYrhVQkMn5HHIaAUwrDls+6z5EK46XUwW0w5XQoWH/fSrIE8BeN/uX2KTrMiFlTi7D8H/6gqIHWQSo6dHOdkLCIx3cSaT4+WDToSGP5VKDuKCVgL7dTu8bSn0vjk6Vhqz2i2/8q2tITlJGkv3TWPqsf8lqOTe1E2SfIrjfBFQpHiXjSG2SHbUK8n8kzcg7xTBpYxofDegBu+F4mfrTJMdhWvVfDh90jUMttpXL36hcfV9R2anW9LSMobbhEsIQwMGOMPgB/y4Bqxfueujk76xMl+UOD8X5ttPdEXiGS4vat+xaJSt7VwBhA9X+3aO1Qvcp9tV1NrJzUfjxKYzy1ncDgrac94REfVyYEGhQ0HdbDpX8xQrZAlzulZjmm3y4RWlUK8x6UOtMRJOEh8XqXg7r9dZymjlXoftuDOuG4+BmBxtG4+brBm7GpGMvWThOINjhJuiF9p7j7ns6ujNM5mhiLH5FC3IGIb6Pps7FW6xsPDuYLOYeEwFiuE79NVih+x8vydONYuemTf68hAbvjrnwvSBW+tVXcNzYR82n8wdXj+a6yI9x6IBPcTJvdRks/24xZ9biQ+ivm/XN6N5BSByyej6EBowX2KJdwEdER/jl/hLPt5h6bVTt6lcJyoAymspuYsnH76NSDsvWIqjU8VGRIlYLYbQX7yfsvHNjJZ7L56jkNKD8yTRFWIynpCh/Y8U0iEDeWOQlGmGAxAZ0bKQUsHhqwX8mjAF1N1w4Fz58TJYoh6UNhR+z2vRTATJ9p7ueYZGh98MSJ1YPDTgLMGie3Kn+vfQC4lZGDUTdbwxhlDOv1AkFTa2Sba1dklsQYxdStRG+ARWk6rPkuqzO9lbn1N5QNi5JkhReaAik8eZdDOQePz1YOFjyBHO6XMp6KBuA5wOzQoivH/7HnV8e0V//Goy87ZCJGsykDUmBgOliFOlbqTxOmEeFDjRDyjWzLvUuFSvGpXpAv6mtRMIPyWTZsZWkoaNxgMGqpmRwbeaDAKPRE4g4+iYh/7GuF84Sgf+IZIDa2INl+pPXABGXSAadw8YPLCua4Z70CsRuxv8UpZL+IRcYswIf/AmGkRi71ewiSScP8+7Ne1if0tpjKjYIVnEd5qOC03KF1H4Xh0ZMS6zAlI/GzaGIqMekUAzlbV6aaTeMaKhFi4kfMrakDekGS54OHxwt5MYoU1tbPmbxK11U8XmQp+fuVbsYkNDL5wFCVAMxByatWnr+LdtqdVCczPGOcbd7j1ny7CZ/XMMxYRgE7vu9RNH7h1m+HTCBMwm5zP9d1GB0brFTHJKwV/8yODW0AqIWj1djSYAGhsyNUVNCIiQ8y8T4CqmCcfz1wbuTikaXFzGf3+QEDGsKLkrZjkGgM/p3jw5IwtpjDQdJ6RrsKWIfkt8FOOmvx7WL7GUTD4+KT+x2U4L2RL7ezxvevNd0iFhntA2gLVf7yx5Jy2qVAa5hXrRAIV1pwZ6WLcr6ZGZ7DTxyu89bj6N+Y0jF3e8DURP1Tj1cBUUOeDDRse++W/bWLSrrdK/YwWGB5q5D2edW4IX0id7aEWwKohbMV9SHI08gtNfo696OZvbWwEUTLZiRilZ4nrcNBiohw94+ZpXLlPig0eWfW1Uydfeu+lTAqhBH8YYtMM0iaTR62ullxuOIXWRogul+/ZlfRdlbY0fidcZLkX5bPAQcXjrnaGLlw2bsbmsMZcEZ8l0W52erUwnYHTVH87p1vntNVlyHXUHf07Bl/Oe2mgoe8GW68AW7houINHuPegLQFOmI/L/aZr1QP0j3f5tITjOuBY1AoT5sY51+FSeZ3NgPGEniVM03Mtz0d0YkYlGAFtjlC93Ra00EseHKvaaUyyKn3I82eEOGyq708LU+I4nG9fG2dh7AbCaVLR1HGWd4QMNb3JnvF5iVStNKL4eU8d3DSvKqSv66oLlYAfQVPI4Gxo9SlHf4TYNz1CuUxMFJZQPHnRu0oY6k/HVzu/Of2dtfT2gP5gB1/Iq01xyhth4VIOHf3tV1q7crotx8JyEepIKSyK+mRDhWUtD0iWeiAp2xn4qVuF2N6HMTkObKTs2OcKQ598n8hE83SRF17pKzSYwRcrvrYuUDCWuU3FMreW6FGW9G0Kr8tBPabm60qUuXvzTe42xRzhpKx77D3twQQ0CMBHVSsihE86mZqmY4QmU/f4JUzwfDorWNrqfDDeTV1nSS/qQy00D29lsGbOVEzHbIeKeM6bbVuERYbO9jRoKYhx52IZLBWXISLBB+NGzAcNaGzv4Kh24EMOwjI098UHerXA8WDIRZiBretxun3+n6eR5AnkRwPJF/6YEDun+D7Ij2vCjsBmMGhnxv/e1Wvu1ZpzhGWJjVstixY1gQM4DLQRWNcpEqG+D61VczMJxqkWgNEaRAedi/JdE9lVtqB4z2jbADBvucUk4J5Jk6xRPYz67Gxn1Sm2fcEo2nSLW+9tOkmM/KJ5M3TOpeB4EoehReQi4DXeaTFcHEajgMVoG7rPkqcx616lU4Lk3+Q6hPT3mX+aH32uL1yal9lM9VWvagvLBm/HOnmCkVa1Gd/g4wUR9sTXdrD9PAhXbNhZSK0oz/uR72MbvpHym4n4LRxJnYfjq0lZ28nwpv2tng7r+aSMTcFuSSr/8MOoApVs4xSG/S8SirOwj/ZncdoM0ntT7rGa9v6RUZ4VAYwOoj8dmg5IfieYHnzFEa7EiVyF3sAH207Uw0NProFkGpvA2tc7da3fKWUSBmtCMikpIJuVpOvddqgc3/NbhdOD5oio9fRyivMr2JBhuKBRjjoSbESR+R26XslUFtFGtOWwqBorsGKhLJqFxVwZ99JqR06xOOQKe63zkO96AspRdUeNJSai2I9j+Ub3l/EfJHoaJ7SZgP7fY3doeppqNHDalzgiuD0ogIkPk/ZxDvyTuKev9YWp/65QwA5Q+n1QWUd5hmX8ZjdjLq2oWhVUhTMxHLuOC9YN/oRdfl+Ise+lrbwa41NUXjpRGGKYk3QjRWLMHCKitaCiOHDdVUUjynhCyR155/rk+5BtHLb+RN+me3B56q82ppYeZL58iNjHc8rIPSXCsS3+ikDaxF3pEjdDVjp/3Z+H2LHuUEjrvpTMOkJsBe90eTODPRyIfPYlbpGgX45opsNXiV3BOh9tsFCtPMjOkXlKooOwjd63eEX/KPD1le4/7JnMOrOCwJOb1u3GDeO1ROlzTpQsG/71aB/i9vp3K6vkp6rOaFpCA7KjwbMBw9PsGtmo5WEPSHrWYginI144y6h8c1vgHsDEIYMdMu/OUZIITTM2OAoTioHQrqMtaSUeNddqwozi101NPzl/tfumLsCR9yX97EesJ3GKfdAbq2ODKA+6H/KvGq9H3DCjtMJ47FtbYF/XmcNVUo7w8J83rswu3igfHhGwpi5sTdkWqmWwlcleD5LWCTCHPcbtGD63x/KbrzypU6WnmymTMllYrBtDaik78GsAo7XtlELM7G8H+qnvQOpsbxrxiHtH1Jdm8DAFOKpqN302HmUu5iSOdSq+EygYTDtVa8UJ2ReKk2G1P+DMAz/Qu/8MSbffhi6Q9peycysUhzg3e5dMs1UIGWnwqP2qhHAMrphF47PvAWI4Cnr/zcsxkj63knTnc3vhP88c7bQbgI27mNd9LfF58A4r8EKAxevGUiZGPZ4d0Ci9IC/DqrD8K22zv7ZQBM5jImmQJdY+UR4CAUsQ9swUj2SlrZS8K28SDa2TB3b9XAyMh0TaPaW6vIYfk9ki3OwmEUp1aobN7Ju3PY1OoeSdyW1AOvZWvGnGxrHEZ7hcBotkWRypixByWAHQyMJXlGlBhd3e5W7/M0jP0glqkh7/m9IDRn4D8jtww2g6x2p9PvqjhQIdt8sky9Bwh33QQTE9XFOr7bUcUkEt2YEoPez7EbdC5TS6I6oTJdNVFexuVspyDAlyrLrMqPLknZMTXYnvxE8nUoYRqzZZytPt71YuXuGxX5NPFZcbglp46UrSOv5EW8pEXjTfd7hqfRMyInXlExyrQV6iNTEMQhjhpzcS2xgh70Vz4Zv16VwdIu+DIQ3yIHKG8/yw8xcMBp0YjSDoUzs9+PTKUNo3d1tHrFFjmu5pcNb5zXGk/BVigDtCy7ar8mo5YW36iBUXcEMsJhgvg3XlX8Z1OLGrfO/v6RMnALAaYvv58KaB9TVjESNr3vYMblPAW7rA9CY+2BhD4C2lfEAKqwEuPl4rxqZB5GHY4LKwlqLPuFZsa+BtMFTdbLdzEhlBejDyvaVvj39Xe84/d6nxTlusjN1udUM/puR3M5/zS1TDK6WqzaMSxDcRQEA9Al/rGhTm6D0yvtT8cUamgpZ7rd9nQDK5cEbPJUg502FO76cgvkTkNhE6WqlIChQz63akKR/WVTFHXw617g6t+pP0YHIQzhRNd06RC4aOLCT9Z3kB4z0/MmtounUCVfL0EUSHQawduYe+72e9OgGgOGU1renfDaxrB4KFB0/iJXXvH5XMXo64TcrhGgQpzaewGtp5ikmFEr1Iwnd5P+PZrSUU4qmaabrbf0MqjGItYHIzzYjxo+ii8XmOD+cYlCaxnn+T5t+tysXBN0jFMoE3YdbA6HlB56KsOjVUJFNaPPK1sT5S4tW3z+JvQSwndZcme5P7AsX+tlXNGoDfNGklbUgtfCWuDGfz1HYzNOJKYmjL+lGT0x6RZoeE7eWPggmYlUf0C8sBjkssTkLHon8ttBRmSWWtRJ8COtCUOkFub/vSIxoeZR8rW+QI7DnW1ReMsEe8qYFQTgQF2zqBIjmYE301am7SA6uTxTxS3Hw1zcKcMJ3+BijMIC++zUneWcsj7giM4QyH4ZLKXyD4R2HwqGVBqCmNZWDCBe3KWb2yudzeLnnucnMUFkjtJ/rBLco52PkJn8SQKu/ozQ1cdoaf2W3ynVNyG8rNUKt9XRMNcL4iBkVOPC7X7nnW1nk+VbOpewc2iYbvih1h57nzZQwp8CBtXYRoOEMPuE4SoMUagjjuRKTL2PK4Rb4b3hvfPzT33Qm06ZAeHbRWTHxxIkV8W5MLAGqg5jHWWIQvoucA2RHDpLccVjowcvWQ1LVjJ+aybr0mAqUOZLnQicl7bGFgRXkmHHKfgvRk/CKXwN9QKOHF/R49dL5ndUILQhS09Ns6E0c71CKgc9xmlwrfnlfuushp8igcaJ22bsYePj+27ZwMy3oCSSSIhF0gDKykWhwLflPcXx4+UuZuiX2vtOlDPgBnpLduKRO3e2d1FyGgj6gmkPJdceJJfoit74YQz94O0xxppH6GbV8bxZUtcFzYiqx2KYUcRA314UN8m3HqdL1mbarNHiitwODG2Mc35fr/CfNFbGcLPPQj0fWt0uxDFgttOo+Bg0/FBpopINBgGBc05iYBgxya73+QIaoX4dvsicI7pyP4Cc7Zi0qcb8MDJa1hPgwao+BNi0iQI3NYvVDeYzQs6u7+So5NJIu4MBr7DFUkmfI1++LPFqe9tK1IcqT+8ITCGNmn6jF23TjgP+TlNQZvyZsxjz9vyzANr+JRfKJbtRB49PK5R3CST/1YdrP133bZzRavoMzOfRdbMwK9WvKgtelMzrJoLyXFRHriWqjpEfPC3rlTN5oI3/zRuNpJS6jwM5af6N0/nrrlfo7IgXILZ7FWREqKpHYLJ0jfkOjK6Wbj8lfi3jsgQPcGsDEK6fnr+dsm0ZGSQFfrbOHO2JkIz5mJb3BEAnedU+XhaOP0s/rRaFHVHqmsNSpaocZf/gZBgSAemxJNedUNwvfoeV4IxkLXHlKu167ezSj1GC2iOn6hgXASlK8YbxEU+nBA9HSpJfcyqh21IX1lbubv8lBAqseiaN4iWdUvAO9DGdOHXUL7OkpPcjGeoAG4ZDhx1htvafb5AryJC/cUHvfKHkgqmLveUk+ZVW2K+NNhjf4sLd6e66Axw8PjI4DEAcqg1+m0oxBtiSELIMLBFi00w6eGkCXIAqUTaBv6IOqBVIy2eeHW6EVR+R4VXv4MyD6Jg75g9XPivfrh5PpmQV9Qm1fidCTqUwluLeqn01p5HHGk643Cj19B6fMIdtyUpvhWh7S45DGa2GwXQeVBXDUbIcHssd0IMlRQ8bsSlEJLhnpxkxoYW7J43AMlCvNX/RC2goK2pJeHkhkSnVWFM6Ta2abcY6VAMmBA2D2v6lGLnwmxORPQVLBlxyg0iZKv2hLxp+FXXoyiqWEaPZ24FapV6bJp5DC7PlfFG+L4kNqj09R6LdH7WbP0WwkYN1qPCricQn3xDu5nKweLZyV8h0taU9BRY4NTPp1+6+7A5BpznkKu7PtcD/X+2Vi5U1ftCCIwh3gFkoSs4eiPZMDpVWdNN6eqQtsa8NGpvP9HXozLFq+Jlha7hmMBto2FHpX+HwOfqIHcO3u3ITNArMu36SdRkgr2uE3RuYLH2Uhj1b4dIW4uuB14JHhrgE87USWOD8KSOuq/4lXen1FPFGFhZrhuF6Z5iSodFCLkTfMvTZGVHELrZmJcyzsX4iD7/o8rePwuZKD2hxeY92vytcqYpbwmgSUQ/emqM7szvESvOpz2zsPzD/mKgtdNX9aEYqUaCLQSktV152NgzwPcNYmWQWzLGJS/nonOeqET0V9SJhEZf5g/3UaAtQYQEpJbSHecMWuhLHK/QtJu03v0j96oziNF9ZGg7XbKYnFL3tGXyPCC2A6kW+Zutarf+mQDR5N6ISFa6fRvgAryQUHkv5G3sLE0CjTxOqe32C+U3rFtD3xumLNaKEpRqAdzqaDjr1tbN3EdBjTpGuCfmSuHVoFcw589weRR97bl6R3NkQdLMu98SmXiUaXMLnR6aP2sWP7FFrolO3hDBI5b/f3wnMiUXG6Y63nwwdaU6W6zpv+VRXBPqLhacVscT3YU0vvxwY4KwJQBba/4KR/1075M1o4QysgDCHkeWye5Er3p8YxJm+1v+LoMjpZfFx6VX81HAVwY+ZzFtdGte+pfonF/nY5B5kRWBjvw8kLwVKo0md8r4840qfYTw0H1FMsaeX5Ba9qFKcVG9Mss8yxBtL90g7wNzi4cVp3NS1g4FKc/augom8iT7cIxFa+24jOY9fEZeEdptrhxXLLVoAWjCEkePXhxtiSVETcJqBwFMyXojeqMBeWZw1sFCGUboGGM0Bh6XA4ugaUsP3SXcg9RyJml2gBdCcLJbD1zY8AZ8TLnP3dP0nfCMiRasEe50xkyP8cwQX7F0fnBu7zdGDjgUEmpanssl+8qyuqRCTUj2uzhO7lxhTPrH4GPmuAIHurDoLdXBiRFe6T6kSOWcATj7R1kC9MGMw3hFeVcGGRFWnaGEdRZpln5slGCEECGkZPCnBdqAn8H2dLeXkGQxiesWrnQm9M1+uF32mTJbvPL4gFkmPcOfd+IudHCeEUJmR9ASfaD3AlOjNFfRPOrxAK6EFLt3V1JXbi0c3+aBDpCU63j6bYILMBDX7DusHJboCS1XhSqU36awxMYA1WZsZE3kVQeoWBrVKfoVrZ7kbgm3QeiLwW7OPOCOQZ9ajJbdsTzdl6CpOmJsDFdt5ZRnlJTLNjvTzvazI5VqQgWImUe+SvIJH4LZ/9r8bPoky/P+lMnf4z9HrzuDlzUrro17cKetKGQ9ufbcWAAAS2FfbwkcG8BpxFXqI16uk4LwOXxwIgRi+Qhn6oE3PCnesj+WfsPepbq+VsGpcVZtLei5MbsYQc/0D7QbGwUCFTZscL9fv1yGNsZ/WkGRytqERvSSRK1hhLrFc7Ko57c3A/1q8z/rcPx3kIwHagIDlw+wpmUv+iLA0JTN68euiGnY0rJj5j7706zataQ9ZMoPw8WMNDknajk7eVRGXIYVp+lWEyOb+oDTOmLso9VU+shKXFwhEmgFZgy2QxKg9axgPk1onqz+SScgvZHyUdVUAvL9QiZuEIlg+LH2ARZ42eS2X+PHzAhfNz3kr8ZZ9jSR8D4p9UO1dPFDNFCK8el+lTU9ntOL0uh/9t8ve0512j6HO3/70wTjic1bc8gr+CFI+CndODOoWxMy6wneSspCyFJpVzc6BuBfxWB2TWI1RiN8wZCy99LbnkSxf2vgLRsCskegW+AH383HsZhDVIGoCjZBDfAq7P1WxzKf3oAuhckf20FJyoUTitHJIfRdAvnCF6zTWoJtdf/F789ntH+TzfGcDJQ5CjN1zHX2CP/kmSVwUy3qs6VM/eoKcinOUR+XKi7co5ZfqBW44S2+zapZzdv/xjDeJ0QUkJFbWFuriR0GpXdzwq/i291zZuE3SRMySkMqQg9Uo7n1TKgPZNe91dbfdCfuXXnJD35fnSgUU9VGkHz37Iw11Hqg5otQB4Isyc9QuGRMvpfB+a+Izxfy1oLNBEBEPFG7RLSGLFOWazMuTteiA9JdoN/Jpf0wqoUDbUm6SxYbqxQdwcsdS3YQRQOOnl7exq6WOCsALSRn5EhipdFfMNeMhYHBDxzDh7Sd50O68fi7OSBwcQHUdvcc+smxnbIDsFoTlc2uYSsKs4+biin5sF7FPvPjfpGywWJe3wwTZXfAIlk44Nh+cMvBGo+jBLIQ+Caw1eLsfPhamgyXOy72Yh7cKpFqpN0x5j4uRUEC1eUuT5uV7WSicoKMKbWLuI5z+xga+zCT+cSg4Hvvf1ukT4wTM3jFgV/c5gszIE6Tn5f5fS/O3hnDI3KygnOEEVWkCNDJNdAITro/4gafqlkBYfQUBRrSOHxFsKpF86y00hJpvctnBJZrnTVjBVC0OtA3e9cvgbfriMPPmtVxUIQL09UN03UXpPUtOofBNB/edWCiZa97GpqOLYDjAQgiSbjrs/VaQjl60zyH5VHKFekg37UOb8J2Lrj0/CSmLpc5mEeJq7CYMjNn9E5cVZfSzlkmYcYCk7pzQ/NOUW3zfkINzQgSj08PLGN96fjwbo8Te0I7ntAjBThcyIpeIUq1Swge5+1bPhinDjXa/+E6cJUFZoRXB8uo9JeqzgLg4bNaz2rZ/+j2uD+4ZZhrp1p6R+Vrmv9wySd+iU4QCZb7T0u03SEPMMIQUSJMoUf7e7MPKZqme4NV9EbTzFB7F0TrwKB+gMQDZMDd78x4SzeTPcgnNtDqoIvmG+56zlwIQ3srEqbznx6+HRtHj6w6tIXMX9V7MHHaHgM86Uu9DtuNaikZnX4xQPWD1dbWnmNc2gm0FSgzVbgR89ziU1bTWZppQghmhUuljC1JSB/+ZhWAkAEqtfwZRFQ3DNAGGBuu/iCXXVKYY23tJ/GL+wIvGvjDGwtqZYb3ai7SOIGfE+GGegeSBqnv3yexxuhhSfCuQtVxh6Fzvvg0Jr5mMlkHFRaLLoVQPb3R6CMHi38l5PPfXWKu/nUecEyZRoVqZ0NKO9skat6jSBikCTF6mySOInDAEa8LcJ8sNG1jF6J4ppCkA/XA4dozXOi5zYF6hSW7dE29LMOWFObhvVs+R/spfFexYrOAkBGNWPsq09PW3NB/6zqngBQupNN4UISqmUJHp4bHeLXsgc/nmEX3dGdxNcmEf0rgopNep+Lbygoy1BP0I0slDCB0fmtjy7MwecNaId+3GkyS8xC1r9h9VCrxOWqhLM65U0RB9+cH94SITdXSlRcwVjv5Ia03GWCRYYxDDAMF24q3L7LJfsABKDO7HmbkR1nbjBLHpOFp5z1qgsNavBjEiCzxPitWlfJiWvNsEU6/XmdOAR/M6cSBUbGlFOTPutR+oXd6Hb7ms+vCYRiW19JRtOz03wlJvp+TPvcy/sEHokQKSTa4TCkq9vchY+xcAKN4ptH6d3RZGA9CleoCMgDOR1AtEhbSAf4ZoI67TfxWRAxmDg4JO2J/P4FOElEtQt+B4Giw23Kpl1Z67fFagNNEMKljCnmrp51igeIkJSjlJY1R1nVROBmN+EzF9mlapuG5UdjGiQA8dzHBSUSIc2pKLX1g5xf7RY1QcgaMZv1IL9qQxwrHhlXLIk73p5hidiSD/P2yzV0q3NHW7fmY/z4jU/envA13qQwfKYs+8yHTAsoOx8tKmnOfmNuPIE3bmkgZyjUXHL89Rxpr+Telkj8WYSkNkNXaCaFyDXwinF/IgtfZO7Oh+nJV7SHzAJ4KfTAgKOf9Ybe/thmlWsfnAgprEp5ORwmZZO/u0gw3hlZYInnZVtyUtsCUqoFUDgxfAZiLdU73YLpJX9YPGOv3QkwvEn0BY50bETDgKXa5nO1bTvbDntyPVBF1FOAH2GPZxv0rf41ygqfCxY0KbCSzMFJTKY846ZI05vXyK1Z5Pt4aRntnsGyd8wQZEnUHZH/ZcRMnux+9OJQr8aZu4/vXkosHr1eO7efFOfPLufX+RKdj+TLnNMqnnMGT4HlUwAXzPuSzSDUuVZNBjNi4uB7zSK73cvfFcPahOi83wiKJLJgNOzTof2xK/Msp/bWQsa46XsOBygAmJea+18DGqcAPF3Xfw0zoHbPoGuezR+OKfSAcYlrem/c+GW+tCN9j6xPbqPGPWlGiNHh20rpk+ianNEwkSDtqAEPau//9a1bs9zGncMjSQ7lLY5lS/zIjyYzu/XqfFEuwSX9jQ0gbfyXQA8eQABSM1PjZqSTqWwIGBO8qSR1W07q72NhLLmULnQA0TK+Ry6hpUF57nkuUFC9NPccimUSibuWdq0TjaUvWnDUOvODCTEBalu09qvGYFE7RoTcJvA9DXSs57i7JwRhyQPa6QQv9BpptmhOcDZAOt0rl8waCUe5pmgyWmeraLy7hm/V83ad+n0X75g+GpTw4UoaoqvS+eiiyRYhbcIA/j9ftURfveD8dXDxD/oJMyoiM2ppouo85KaMLi56yHQbo3fyJiTindYIQPuHlB+zY5O0+lX0HEpKZpTsdMsHSQ7uOX2tWXFRXr5/nlRMRf6YCOdkDnT57jQ2P56mvKv5RvGfoT/WNnSQJM9hUb0DxZl0juVyqRY4brv4DYVom/BMtm23FU3neCtBKUmUeiCGASiDkqhRrc78os9bmH1xgs0e0JdM3JEhRxW13hy49X0b0oTeQlWEI7w1DasHvRU9dzq+/dssCPgLcA/I4AWcjbofKoky6QZdHo69MervE2L/SK3NM4i/qAGMqvFpp0AT/aIxseEtxSQm2DIjm4Ks65DRUS9vAMlMZsbqFj3GOmho3CTCS/y4ARGyIwxMVKGUzcND3c50uaedn7gCG087kPPtdQmk+QkNDYfnGDFZ+WOnHwAlYCjBk+gTIOIKp9ZiIX40eR3ZfWGeXn4jqT48PIHFtoaAmmeGTCe/4YaJ8VTEM1u+gnvRLuWuGhYMpE0947PAzBrB7TpHDWp0JoYwmwoD1efPtCDQJVPCy54KaPz0433Kbe7rgnIN4I0k7gjOXVw5lJkciS+aL/jSDdTeacy6ZHD3IL475Xb/9RCOUKZXalJdlrhiDTS64KPJr1JOrGbAIWxLIE+Qo+9eGVsSfjndgsqZwro8DJyvlWgVlEK4It87GivUBDsoL7xo7iWFte6vJr/Z6ycGLX4NBWafcxask3ul/dCQ/KKJ3FT3zx/6/xKNVCI1LyVsnXed00xn8Tab+M1ytxfORNveJdHf6SMlzPEAmRdIZHpuDfA8azJ6K2B4RGNz6o22K8jW1fLV3lyPlS5Eu9wAz3M7gu64wXJX7xhUGO5XLquG9J0sFhINwzKXYF7by4rFc0bEyYyJwXlb6t/OblTRvsgQE/jXRE88y4O4b54HbKBf3WOevYw5z6VVDaexueeh5W0B81N8bUoQircFak+sLSxj2gFIaP5IKVronT3wY/emBJofPhpWTw6KEX1l3oeG8SX4GsVoFXYPN1XchBQX75tUhC7CF1YeTjJ18xSJUGjS3/RU3plo9YCjp0Ci0kaEmlkrs4SZnpNVyEzIf9qagYEraHG4iwciujJFI6KPIMpXGeOyEv4tAFUvxpGNBngSIb6lFNwfaG+vpGmrJhBWFMx1sDtpThIAcLuAN/KzazpUYx8rG3ZWx0vyfX0BOoEq1rg9bb0LiydatzVsYSe+6SyuWj7xY8p62Gou8xrbwPhetHER1qeqUQwxsWIP78k6apZGEEPalTP6wl+GDyI6Ki5l2P4ZSrdYj5cBHm9PvFjowbERih7eyTjaHSViFLvRIKa5b7z4gXIxyyk5d2/iHoCWE+/dd8cfM8ut0reTQTih2Hq8xeS4BWUvjzRn14wsIAmn3ql5uyMxxHOMytW/webqplzHQQlu/tKLmg3A9UaISUkJX3q8inVgQ+hlu0Ke4rDmKITzzd0ocI+SzdozBbg4AmbwFKbCa208I07MCO4nffLByFrs+aDD4Icjwe22m88xbfcVQfd4JLxytsfjv2vEBVaXTFAlqnv2Wo5V8YFwnwjSkBEBXFROui3kj73wBoo13hiz/DnZaln3J7KPAjNPbQoDIw3cFnp305Uvs9GX5GxNtTGs19/1aF/PX24/ThSfwIfTlUa71dQ/8nshuObd1Dt1BHvfH9JcLrcZ9yE8S/7CAwcSyi5CYiryy1nA0K2FoSzNn2T5NZ13dM1F8bzwzBwOyJZjp2Uhyf5ntdxvhGTBD4Wz+B5yc1YbC9eW0VTRZomHvSYtOhcM8U+iVpzv1RQh5eMjqWvnRXSL52xsmAneLykJ0+sDel4a21+9grlDmMCWWKqm49ecxZWnm+HnPsZoxe3LGyYmo96zpPnkSW6V7Ot1KtgAKSInmRm0NX3jiMrTFyUXyQRLT4Qj1joSwY2zr7Xh/LtjtCwOn3BbpWzx4WzHsR7IIriHEcOuJR2q0Y8vMqGvF6qjThjHcgYqpu6Ek4bEGna6qRBBlrwZcSiY5L9i+R9NaZDT1soTYXjVm5BVchyaJWgK6oSt1CwsojanheXV2NIpTuZ5/O2k6B2mzFdaPfOko30amjboVxgVFq9+1H1ka6HLeNNq4j8BTCFf0mNEGy1hHKX6biNl1P6oRDVmYvv6YplbMhZS+PPFV789rHaZiKukDwVZT+rQjk0TG570hhO3PrOqm4IO8HMdiN6t3oZlbXAvfXVd5R74eAcIJnc6UPU6oLu5CmHP756+/iibcAKjqrL4UKAidRwn4tttpNPvZv3p25RjRC3oQY36UvP5J/tGqE/Pm3U1+TV5x/E/lezKcNjbZuM7vbFtIYT1gFi70lj0LOTl4BXFflsGNRzze1lZgSwSYiWXcoPGk2VGwqs0oaQJ4EzNW1BIvqoCyD/lO1jj0ppwT7fqjnon8LK6oISdrdKJnCwbFMEKHZt8iXWDp8dFtd92zIrj6D/MDvUTjdhrJQqKWupI2jPWH6n4TIuk2dqo2OVod+e3tswzOFFCExYPGbixalKf/esxRmU4Uus7mD8gr9UkLcXGhfHY1n5idTi8839rAOBa67tNhEnOUw4VGVfG3WA6IJbASQoL1H0EO05i0IN0BOSWNalrH0ZfI++E4IuHocriSHXd2xQsDtresgfWfrLuoD+7JRI3ojoOb8UdV4mgFi/oPzAVK1i4hunzh9T/4GxmaayiuGWyvGYdorv7VBPbZI5X/+Nvl6W2xAuO1TyStCgHAFfjKL/SL4RmblgK6VkEmEDzEHSBpiYoEvzu7+pMJrLiMioOB9K47rsGC/2JZWvvqsMngreW7VgVY4gMx1sUOIK87KveMLbjuiiDgP+m/NDucViM9f97CqzmhyRsCSFjKcSTdy7CCzlr1WN2P/e7ZoaAf2ZdqHoyXzaeXnUouzKA2Apd3kaCP8nQ6mBXcp0A4QhqAJT34vtKxl+ZUIZXZ332veY2DN9vxse5qxZ80bSRbEFd07sy/CDR0wiGazTUez/jneKZdSrWYFUW408eGlVYp4iFaK8Ec/yOyntfkFsfveN+j8F7KqNOwOsBue4iYiuBoORUAFv6zS1VFLsiXTohhFVEDSnMPuFQ0UeQKD38X9jiOlf0AKnzu0goBBrnBARdJ8TU+Ygk42ZwPJvbE4xfu/I/vEYCFPXkhAJHdM4ZzJpni8/5CVK+cEwgbPO0W/vfyXvvDVXsdXCSVuor9Esg8kNfrqN0CVp0SHb1nIHq4Cd7mp5421gNMWnZm1NdxD68Ue229EwIzb+LLL+Tt4HzAZUMiKRrM7ljhI39S0XLQkUmuZpJYx5D+hBB8Lx4lpjN7fp2sgoOull1rsj28bPu5QLMDJ1LiVxQiSeV+fN5UmXlsSlWzjVcLNIwJDOip8lgGL++F7x4oAgodlw4nCzn8fWI1y0jsbYkGbhd1nH/nwuLYQfIjZwwvndt2YcdnjjqQUPviykz4ic6XbxydIdNv2DTNAGKAGDPHmb5ioaTqODSGpECGSHBVXyUxrO3Cg6XTsEWBfYiPKfAru4hZC/PgOjks5TiYZaZTInBhfkhyfmKJdKxv1OYlHYUnwh66un8VZaD+FrGEnjjHDBz0KIG3mynPQuhArNH0PHf7X7CUtY0uyoaQGeH59JIAod/DHMtIbhvsnm0f9coOFwcP+yAfW0NxgVwPfF/ocYWV1UB6hXcc0KhqlCV037pAmpSoWgE8SnBMNH3oKzzHbzy+CLf83JpTNeB1Ek/a9gp5vRgW1eYJoSxuEqAOGhcsYwV7TT53CZb29B2GmG6q63W9R0LhSZfuUtJCkelO1nnocZuzrtTyH2oTMgJ673NWXWsOiCBbGJOunXnq7GTOwz6QGauY7M/HrxTouh3mUYp7weoF3cElzsuEsiQdbSUs9w3jmrV2FvPJxwGq+VqIZVRJiMBhvNda/CaUIT/2jEln7si4snDiRt3RUYM9U1zfu8BfVxuZsAPShDUqr0TlDQgP+pWgSfmH6Llrfl/ZIKvTqZVlnXfcdC0E2xvSEYyHnUwY37ZjtxmRVeLRsEF/tTZut4fxHat0K2DCTFYJx+LNA/mIvCO3Ysj33/DRC/tKcOxabGD5yLGnUK40cpK4iqlFGJx6zLZS37xXd5r4dYOZRQgFkZHoJdA8EhNu6OftHba9KKU5+by5/hrzfRRErtWOj0uz3BVEfUbZ8sfbF/wRHakAZ0bnbogsNNtovClqwiRSXKr7jiE0oCJaaH/tv2R/BeHuBUwmrzAQLqFkWohElBNbanU4g6HUsi0vgL0KoyV17trD312O+96db1wHDrDHAp2UE0WHozYSifXfGmLdDuyL1RslVBc2YkQY/VZTQS0QcdEIHdBeaBWG7w9RD74vPi6u5I/OOEg/GoSdGKLTkrJu/UOzb17Ieytdl7plxCGvbqZ7qe6tTy3NoU0BhBv5VbXOu9lWyDDj2KT0s77AJMzzs6TumjzNqiU2Xr2PoqpbUtS/n8elxh6dHVIpJXcTMQIvJyO73mhSKOsoTb8aJhJrDW1GOyOGQRiUpsg/cB8J5yWgTiERl3R3pUY/qKkaItqH7DxYiRCCoKiGN67irRVnr9jBXd87UvRw8c8Cxqi0nvHfi0rYtKChuwacCxOjaRVH+0W8LPF0VBrwjaUIzhYp3AMb9cZdj9wjlt6/ohiIg17fKT1PK8/K09MwgpOQ0ovHl4l25n/KUKaaD7kQkA6VZtsiEK37zzT/xo0NzopOkBFdZar49XnqPkHesMVbmmIWpQjo35rOkIIig1azk6+i792At9CKDPFFqnv8vnAEfKH1ytyIZlwgit5pTZTS1FjL3ak03Re0I5IuuFHrmhDbH6jWhyXAQPJJGwHsBuBkLg/T7a12MFTu+qZr5KmvcvMpC5YVm/sbk069d1y8h+osFLbYaJlyMcmQleRdy1sBOwSXljAJyMBON91Ji5JzwplpLCwkVoSzOjM0h1RX4tFbCgX3sKNHmHauOni7ucZfArRWLrHKz+Js5euRa37ktoVez/6iJLx4PDWq3EUNan1V23SxSibZcVe/+xf6JgB3AFfJhOrQzKz56aAi+9iKZ6+SVMTHwy+vqRBbC13igHIc53n95SelrR01GNkXuYcxxCqWPM1D1jelu8M/x7xR7bzHfZAPH/r/CNXCy4RgoZb1+Yd0mEtaQETJJxisRtRPLH2gC2masaAvXK0p1qAt5TVqZSd/bXG4iDM3SEBrq8U2tDximLFFBS+ba0P38hcEM91I+U4yfk5ZNXNGVCmJASRL6lMA5tIjCAzkVOgagQC1VH+3RX+trI6rtmyuBDGGovVuc8bZWm9KhPFdPm85vxcTOrYKy527m+9qcoy0ptA3jKcgrys1XG1/43Qo7bh+g35CCEhSF7Wx/W/SEMKHfyFoREioByvFvgfXIBsTcO7in4uLEQj/RjeGCdkke6O3k68f6Wd/DI0KPxTlMNkjvp0YthsDQDxewiuh0eJWxqTCEGyZY1MvLiiFnfQn3VoH1OV1i1shZ9Bv4coYO37GT2F7i5ZXqXQSTaQPjATW8dUhcpUT1K3xqfaghNocB1YljMYaGREsg11Hifj8UR7of7kZTuas+pWnWkRp63R68c4xcEl/Eziz30v0xnZZdYaT/ico8BT7Ca89QYCyQWaNkLoDZz76uNmzsvEGPbDyxhlWmb4ePl3Ht/3Ca4UjOim+LsMVl4UIiyDUsihU1hQj4131r1ct6L9jvfZhiKcs5XL9X+9FpQoEUpxhB2yuT9lIN208YH8Acsgn7EaPhZlx9pqct7vzBgY3rxAJfDbURjezwJpqSE2nr5mruN/6AqF3s6QN0aBhUckFkHPX2Or2VB+knxrfzxfwl7ubzwIDfM8OB9jxEkm6o/IsKs2T3smc4IvNpX2mN9/jxWs3JEa4rb3BF8ErE04vEO21hZaR+mArSyIA99BdGjohsrqE2+Xw2IGKtzgqIC6ozMwHINC7mpCsw5viXbb9lVCLYunhVKNHgsIKXyR3rRX/dS5ztabQrDL3fmJBIKWTkorHje+hUNHNKb31z4zo7Zt3fuSIUdwD16dFwmDDC7r9dGDSZ5U2f9/+ZVNfiVzzy+IF1doY/49K1b+bDMvKu5S3PDoDPNnEsWO5ueJsH542hSoK+0ByjMb4nOL/+oZBkn8pLe9poGlfDP197ZrHaZr57SdV0x114hFGCz7hL7BhUVvV2UgUlUPNQstkvR7Vwc3e86bBWW75r6sahFM1ECHMst/tCRXUUvwE3ohcQi2gKUrXOt2W8tosKsX3DqHpbWTDb1DMBqWE4bIICDPi6m/7p4wJ5lykIB0uRWj77KrLqcXkgE4UybCtnW9sau2f+46aqh426Su9Xt+4K6lv15hYnCrBAGGunzUCTnQcwgY6r1ly8h6LcfAVFjnXpASGBEZIEkWWQ3IwVOAOrQaHrgcBiSZvMVjzvSsrMhgIhSht6i6PgFhSSv3Ix+CrwKyh6VHfOmF6B5Ddagr5y4MDF/7wKsgcvom/ImnKuND5davwu47T9le0QWbVSLnsAE4yDFu7GoyIttaPwfkBrWZgM6MXf371lEHI9EEuz1rIjmO0MEHm26YGomNf1rtuAiGEHEjW3Ju/Pt3jn95IX63SxGbjjeH2Y/hbJJDD26ImwvjN2SZ0iMWMkspwBmfaQUaKhq33u3wYKFpx5AmlKoIITuWWvjpi2gcdNjne+AE16FSst+NC2G0RweBjr09vOKnB615eZnMqncg15GykVwaPmggrgFnlSiD0Vypwp+aQdR68yfOt1weDI7nunzSMiY6T8/gdwv8C8UFxLKuAp8BJHlajoEWOCA1JtLvRz4GTJ1xIsop9XyeVxN70nTwC58WUz+K37EUNyDPANw1WSteqx0mqYhtSe9QhxE5x3KrAFfKFgFIOBzVr1LNrKrYz/68uNBR/hTlHTG6NwqjkpB3t5YWrZxo2V9K0EK5f2tqj5uwEukjJhRDN64XwlYrHdPpuHfNYY/ZMkNxb8npDpm6pf9cvj6Ni69goup8MysIJ6QicfYL2JYJzLgY2l5UgRFA0cJG4J+7wrYfz25xo99kEkW49tuj+ThbEIzzanDy+3Eg5YTArfFhIyUrbSKDSmhLHJE+X+M3hAwUTCtDyfViKzl7EsZ138lyY8HCfqB7NUUurfeLN2o1T9zccKlGHcDTjBR7I8W3xxcxXPtL//3MJnHbAg01Ko7IouSJlurQMbX27n8o6V/07yTZ8wUk3lQzh4jpdOKO48OZpyrshTItaBWLXURDhy6kZJbNBEX1hWWuf60Sh6422Lu7UVvdU9Dm+zkQiw7asdo74jg52Kbm+vVjLO0/UYMh+Ew6n4S9esq/kMhCzn3z3d1sn6D2Zr1ajuBkRT4wgkUoOg7+dHv7ntteYWCK5Xrg6yD5DJt2e/T449yVctfACI0GVn9LlAgbprmoig88N/QUlOrlwaN/CZNqRQ9b5lL899/qtMMSg5LNtukwkVUDUhjmvqZ+ecWFXQUiGonh0pQd9NqYTXCMsRz/F18JUgM4Ea0WhMGvdbFNyieDEqiTZ4jL7vF+uh/L3PvT+f03S2QATzbUTz3Pkv7/7zJMPpsSD7Ihmv8aP6mJK4+vl8Asw85u0LGR5YBxawJ7fQLBtMMyNi0gXVYhSB8I6w9wBF17ku6riclXGi5SQHqUoCjbgQJIjIJxrycpkQxstBJJZQZdaPiRRt85cHCzlCVXX1TqMUTTz9XFHGU3fvlFpEipBmjAcB06FqEJLKBZA4umuNWdPjTwfiGx5r5KkzU1k7WWP9yoMcnm+Mxcs/GLWP3dqvkTJd2D+SQveBMhs6loZ2SV00XQIdIo/PTnuxCWqTBPwSuU68cFrvCakK9joo6K4xqHzypd2hPD86V1b6N2EmTjys8YPbSaNEHpYnhX6bSc8YrLtDAHDgkY+jYBxovnnSlAN6Mx7PictCsK8/inM/ZOSpyXGmNjdyccu/lBk3qjr2tftlbMEGnI75Ll3W7R7ZZnnP0APiqrsdPNB7A3WLCgNqpRiGBiaNI79wI/B33aQAQt9Bky0f/BwruxCWe6cdgChl6Dr5wAvKmfPZJKxrFI6Om8Nowj49fbf2ykSh1gP1skLL/J25tlYQ/eaUF1rf8mKLbO3GveZTWv30WnHSQvI7ZdD0JUgGcRLES0IplTNNg6XTlZVgDOS72iysVoqktGdWa4q88+B9Ybp/8XbjlHWpUAc3F3/4o6HhC8ZEm5JRzjl7HubNkmeZFH0ZZ7iwGy9wpaVYFlt27TAqSflyz3BmoILbW16vUP3C6t/+TstgeTQGKvecXHLwYV11NeY0QoIBjfGi9HoHbSL79VYUpOz6L2Bs1o3SpI6WDDmfE++Nnq4qkoHucUlwQ7nhrv/sriXZ4FlxqtWq1ggYpP/0G6OE81KAilRkLFz5WG1sdnXpJ1YFr4QUjktakB0RvL24/y+xowOm8aaJ2aWsOtbsHx2DF2mtIqdFQ79q0+pOjsHNGsN5byERIpFofatWAecXQkHDXtQngp/FqNiAQb8UAbVVZmxv8/XxdvyioFQZxqEXzuqn9f0Fo1LRLsBEnvucCCVio80Z18Rq/G+a2iuZ1X9Ew0GrjYxcWyr0ozg3g/uwWXFko70ueCGoeHnypf7wgOCzCWgAp9dRW83gad3lt6a88XXRgoCFUGxr1Q3RMzy4A2G0a6sWijRLc85fgDkbbxr1efhmeONzCkOGkSXKEobzuQWL64VbpDcv/IS2juC1KfF4qbrPTo+2HqSp6Q+uHDOnv4y2RWrtNPZTaJAx6/zynrBVXve6NFuft36hPUMicyiSD2oT1O5+UVTvzVehmiMGWwRqa/P5ApwCgbLmGFZC1npbpATHixQEHAwYWWbU+YNv6ojWeiKpYOwL4Z+75FIiI32u9yu9zI0ubLBZKAaA8W+6XnjEZfmN7czVJ/KKyJtlW8KjGQstHfcUoah0LgS1wYt+YeuY4fWN0FJCXxTyCkE/Awn2CgerwpYkrI91vq/HjsTaKaPPTxvUxxbMAGcmd/IG6ax/47R6NpD6nuOjLPilWzQW6Ud9ublYnJOtRjjhuj7AXXDQ/mx6oqmNtsPEpkrx8UeLzVdlH1h7nNUfdEHUHnfS4UypXJvhBIIW1sIE4ZF9aQIEkHFRrcwB+2wbtpQwHlRprYdorV4E5UlfV2tQWubzBNckdqkS8cdXU7iKi5ixIhcsM1/dcm8X7/3Vr3KA6+AVHlfMcsFMcAZP912glbye+LETH9wgjnQpCoHK1iYpSDOxjwxTjWCCkf6Ypc1ys67Axwp6sUtbKa8PhKn1QFe7hkUtQmC6q/LS+ETFShbfSqiDCqCEg78vbNbDkhAy6UTKBz3PiqcoPDRbayYLpzBPoWG4Pv5TB1paBIzl1mN9Pdhxv6zyQ1Rg2DOXAkeQtLOLlUahUtNhMR5nTSLp4KstKFTZ2/IZ5zp7Y1Yr/swbJwLkandEe0MVtdHuZUDlKUJ4aLXZKNy2jPZ670IA7ptJIE4xWH7D8ZWpILR7YT2LkxCU8gFHbLhrm6XA8bwMHbGh/2aqG5oFKsqf8uTywaDm2QO7NO+8ARbulm/o73EEcb/8Nj5nmxR4hmpaptnsbrnJu7Oe7+OekxPXl1OGaknuBXycMXa0N6psYoFNcSAzzH5mxXlZK1YT2Kr+bDrqC/WBj5vin/+/LWEtd59mKKiiRZje/Y9ND2AQ1Pq9MLrFUolKYDLvW6i2dFH3HhV7phTzfM7o9QdUnvB6Xxza2jJC/TdIJa3AlWZ5QKVnG4iyVdwEfrk1K5vNi+B47eoPm22OHTA5jeoN+mZpCGz2XDit4LyPzI4HSsm/UmznVNZ5fhA3JDm+yWsysuCgBJ0F9LN07iRfihD/yHIjS1jcpLaQuXWzad8HBuOgo+0RR2UVRb783pj8VhYHZdTjYsaSNzZMMFKd33Q9iTMh7yMs2W9t7i+y3fr3vrdZEPtMqFqNmbrNTlWWN0uDEeX//920Gc+rxx6KsQNevaWjaysIVbbsKkiPxRA1aYdaqoUcgcG6TfAwsxkEpB3hV+OhxkIPgCAq4NxWUVXxxrlWZSUjrMuZKiLjtICTxt3DwNjGXlfXxE7hKsxa8i1F/Qbdhmi30b6azWjYx5nP4eeaYKGK09iTUyHobiKCJvBhl90mJtvYhJx3qBW86oCYacDl/Uw3+wbkP/hW7FuJBI7TKRKxKowuxBrs3llBXnRAXdZrJlDCQntqOGSGBsYzjK89H8QGzV3R7g2vEebiLsLus1/7iFmPARyzXaeXftEusXgnfzBq1A+V9M8kmpHeRqEAb80XuY5UbNyLuL3XYOfDAs+A+CfVbtrTcQ4BuJprvbBp96vuEwGrJc2NcclGtq7ENg0dux9ZC1bk9wcTsxqdh7a8XFKE0CDr1sYgsq1mTEt9pINnxBZU0URUaOf3GbdOXaFuU42eoLvJbBGzd0Qb3xkCbyzZ8ax7E4+MDmRja0MGWi0ft4l5ps7B91+XH49D1IGi00vH+7kJKmf09SyKeD8dKd2fnhO3jAX7vWpzJ4sUTYP3BSdjN4wq3AizDB92bODYhq0XQNak2Lr53UOWKDeYm03m13MHtWPGhlAOMjjawB+uW547+GkrrGYF0ePFhKX2Oo+Ti786mn57uQvThAbZ2UdfH2SzlN9H2C7HsSDAGBr3GuzL0H2keO1t54DH1arPsM0us13+BvIhWUDR6ynUdi1cvpu8oN8UaUOBVP+Ut4qPX8VZJsSofR6CQjgNU539teUpBxc0xgvzEVtEjX0ag+ysBUHAxy2zpn4AAIEr9euYb2e7MOc2/kAuSE5sgNbwAdSznKqDG88CPL+67oFygoJUNZNDtdKlIQG+MCmjuUKKvZKY/Gf00Azm7Jv+GsBjsa9NeVd0lkbF82AUS9tACke6jbsQg2mLFOvLaynsNeNhJ9utIvsIj/G1OHfheS7TC7m1TmYEcNJemqNhMparyKsaDqTtYa0tQ1FX6h87KCmKjFC8DI4MQqLAthOAM1Rc0qQwQ04uAFct4/dtVdPodHp8tySwVGWBslspT60BHZb6AtQE9J+xak2DQRYjevf02j1CyTyniOjWNdAhGh/QE8GX1SEDoXSUlgWjdmCDfTxcK3Dej9A7EHc2kgzVBhOCbit0/gViQ1efchlq2HDc4qj1cFaxcUUMzZ/ld+nWHfd/f8rbWohp5pLglEtVkRQWD5c27w0FE9iEDShc0si4vk2aTiVENOd3vBxspH3P71sLh3pBpgrjGDbElMydkWWSzwJnQ3ez63tx6XW3ZwobgHovB7yKqJjNqAKaB6fao1Pt3cNiiukXA3g3Bc/XDbJzADeT3n9f8H2XS8zW1vYBd8tkN0wi8/qtG1wC26nFoba6KKOqs3DoM0SCzibSV1xp/EZTSzDpbITsBeeCcTAR8WHiHOt2Yv7DSa27KHTpu55EvcKgS15Aot5QnYnkf3OqdBcYVC+bzBGTQo5RTMcAUQOBNRSI6VRsni+VwWZCWaOAsdb5bb46b5uQE3hGxZ8CXz4hmpe3ilwuGDlc7wLMq7t/7AdRdKgTKRfoUVsWRQZ0D8nvXEH3KpU/D+fr/3bzsfRsG+E7aKDVhAG4gjGyqkivCPGkcQqXiH1SQiZ/pOJIGFbqkBbpOseT+VQQGj62xEuQQQuUmJ4IBSiDRYww+P2M7JHTx+IOmRvSfLaeGq24XqkYYNNNH+qSzJbT9B6uwbrXkQC5qH14H+YwvDTtDg+2kRJ2UYZzyp/YAlE9QZ8NlPi6Ct6IgedVNtFG5/QuefCExS5e4w+oVtNRJYZS0fCFZLY9o72cyTTGM3W1y37SWxsoDiK6kELUxP3jFD1WCab6vD+vRECW3CcUCAmH/9EFEP0pui63ZpYU4rDxaMUItvllscznWGDHmLIphKh0Fup5GvCWCr8tYi9fHHAI1pty8BkeysAxhaqHh5C1cht1O5C+Pyjj3i6tg++gTK8jeMG47KUJqWRU+T01zGukJ1I/EfikQWIxQZNjAqxZFdtapWmSgRavPFwJHfID90d5TRRVwJUjSig178GnJM24jkpow2Nbv2uikrRYoy+CTn85akTr+/oTyr4a0QM1i11A3fmm2D3OjM0cs2d6yGvbssLWw6xJCp0QF6SdAsWmnoPA+BUyree0WYRxIuGBKFSgukAZiGSDhjrjLrj8toW4IF9uP5Z4OdiNBCxz3YTzYS9JhtxvW/UI6PzJ6oxxj4UnGD2VmtIqa7fcQG0nsEqZdTHnbUv/FX4bWt70PhFzteNmDMsjs8scX0N9vjaGIVWzoeSZy/Gtbm/nvjgnBBy4bSdPZigj5/Pgb824u5vMJPxxlEK7T9fCEUJWz9CrwPxNqsFHhSKpqF/LY0LrwZQQF6p3LGT1C+vdqkEDTQ9c5Pdrw4u5h5BeBog8+XlhUSz2KAiSXZRv0CiZAfwsysR49PrjxhO7XjOIFeADhquw8k7pyVwxAmlOUmBBcCcqXAXPWpOKwUWTpGSAA+Lkz1f5lacW0V/FdAMLV9GXc5YiUdSkyQSGTNU6judNJkb2XSAghLyQOtbPPm6FdiEpjhDXCCtmRQcWA5CQkh03j3HwuOnOIy28HoRtjptL2fQCRj8X9yjyGSopG/3++nz/0i9HHfJKUSNt9o6vK0EBM6TURcmr4evbvo2lrZH23mtVVb0h55SSHfihbqjstqB00XCZ8W8rxJQHv27ep6/NT55o9rnSQJdb2HW5QCYX8TDBYkQAU2pnxiP7N1qyENvgnq8t3MUnOffsPMkVN4QuQH/5jZsKTpcJpMfO4Czooo8xc6QGX2weXX20c4LtBBXruk3HK83x6GPXEZ0XfkgmNLaaL2xuBXUQwowSnGBHFd1af8mJI0czOeokL4gnphHDgRszbpwrnx7AZrXOkI2z87c2yPkrMiwd4fjh3ISjED9vxijcfgAG0ZsgIIPchWw3auYVvE8N+34C/M/FENnvvFhubenjIptdKDE9c886q9e1LMFdqNIWKFp+1S826L4r0YrQbfafId/6p1JVRnh91bP70+UXhJiR02rRYWxgLebZYf2nD0dDqplZX78x+53ueiFTtGTh+XAXimD0tQzhoiIqfFXcMsPtgxEpSAlA8xLZ/DLJKm0aBnkkCPf8PUqlxUKYWWXl6Zgzw3LSac530xFeGSSWtUKBcWS8B6fDwgB8eSCuyDZ/UlD0U54pmIs/ZgtNVMJXDYiJzIMOdz075LMul0DgEPinG+Khf848zvjc7tpsqn0R6Ge1nIrgRgAkOjjPut4LHEYDTIrs5/zxlClVzsjKgPMUNn/+yNKM3LoyOPvzcJ1SjmxY4XsfHc9UztA9MabTll9EKtdsT+Fa0lv8BxdyKyOeODMqiLWBhBK81v57ZBR+dTPjCvemlkhZA2LVk0oJJqmPUkXiSc1oZs8OGRIfqYpFlqSZJ3t+9DFNqiDl48bxByeNH34iJW9ubfwg3YWiUmoDlQVqhxrwuoFMNha+dD2KfkEAT/io7rwAlFPcCET6gQcTNVciOty284dBdNqo7y8G0cAVHpKqLmq5WsIhr2thqzV2UcEEoOIDL0HBVAlC0SMqwoP7c4tpZSIr0fRykpvZcstHv1RFn9LWc5eGXW0YV6yIOI5xfoSbUWw5exiu5rY3ThEypu44VvVSYe+sdiYqyP4EXJEI3zefaq32rZaCy/yFORu3FRJ6O8X8vd6z913tqDasIAXqPYRPq/J8w/aMZKxfV96KY7r/J14I1GpIEKsWB8JkCdDgGTOpo9CnmoalO1bnZetr/0Qrj7de5Y8X9cYUYMRheoAXOuJoBcZ/nZS+g592qWe0UIkDNzz4yuGzZhX3YFe5yPs/e3gPKRVIJK2Dsh7ypdmTo22y5N9d83WVXGQ5xbeVroOOZbLKzeHDqamplGD3T3d1au3bbheTIPrd7xu7u/D1bg7IJzE9IzBMQlYXuHpLRi/eLUP6hqaXTghJGwl8zrMzG7t2ELL1aCudtAqr0hImLIthkdJi9NzmUWUBCUrD6wdzd4k38rVF0GlVhPzYg+rHdYtnstNLVEomBLtI5h3p+lBwZ9jAs1HnfaQQbGqsKNHXWSdUqF/GOpxr5TP66NSuUh/kF8DLwxZZCusvDnlM2GzW8Ul9qk4kTmr/F5Tmym1PMGMo4JBjd21q0pnv28gPfOkD3bQYIlx+dlEd0yxf1to6lBxbF2xiXSTWCf/v/D6qz9xH6vXZuaj6HvjmEXz4huPP4ST6tUnyk4Xp+jvjNNk8EvdenB1rjCQRoasIMrD+WgT6URF23+mYCOWU0mPbgKxeA3sPDa4XEvdeSr46/FofTP4CEOvlWoQSNYhGeKtCb3THQ5ZBrV0wi9/CU/UhWYjUakY6TtGSV/PI9Hgac8XoTe9rcQGmDWHj8MyYUVeZ0HoZuUEBijFQ2qk36rrErhQUE0OfvVmfi3SAJfb4+hX3ZXWFuXZ/jLpDH+BVtgB5s0tdOKX0waIrW3lrMliB3f1oHA+XS1CBe7tkIFPnwFOwpGl7HW7PCdy0Do+OLN+ffg2n6nleXoEqi3YUfLy4W6miK+104S61m0hUjphkzJHPSn0Rq5qp5xwGIjR5gkCSRxGeMqHW3ETrNmnFH0p0zkJFrvzjAyJBwf47wlwlBcQ41gjDSgWVqShVaHGc8ikcoD28MIBP12VYpjWV7Ew6258vVPMiS+C7qcEa948nCVUJfs74HDJmMtCEySJHNdrVOulovFgj5V61uMdVQm+tvKEMlVWRetG19fOGmToRFAuY/Np4gv+ihmntK684YbgYbcmtO6YTVsDqoz9/AzUJsouheUuk41CkZYDMTnsIdVr2EmE9dLI84e+gKvxpjeTgBtQdlQyh1KjI2HGH+sVXca4giVMUqP4auWE/fPjKYWH7dISYBSOdD2b4DVoTDVZ42CL2vxaIoRKvcfhU9Y8Sx25fbfkmMiH1P8bY87mnW/sqyr5ijtxZhY8/p/kjmv32SA5A/9/WJ/iBGWvK3QCSMzvetznQFmOrRmxFtY9Obz3M8eEfPVL9aNP56tAeEGGF2hxx4+nzbAgOWBXcf1HqewgH7DwLF1jc6m8oQKtKSOJBiZB4MPHhxInJdZYTaVMa8uJJiMpFfNoi3lH1IcvXOZifdjMfBu1wxUTkm3y5aVocXNrp/8le4Qnk/COF2eY9psie7UBb8Xk86jd6MkxeIYToDDG9SWAjDNKlK6nF41xxMJg8vQ0G6AXtJBkPJx8tRJlb79QQ+FvRlcTWcG1egmpzEro4wQMnwX+T8rWVsXS3Q7kGZiKfyDNgybF3gbSObzzvmnNcbBBoaMJ/uW+AjcFCbowXUHF6fv1VxldYIkC20WOWLjej7SpodXEyG59dgNJ81xTtFMzguR7jnUq0UT/Oi3kjLDokzmUAEHjLAhweVwjQ7ORoF2fvGzrP/4T81JCvfnruH0s0u7jclYv3cXSwyr3ILMVWU/NuAoI5ZK56pLLTV8QGrTYPEjr1LhInctVtJ79/BRxeZ4OOO3fL6j0bDb2gwBpqtCHD9odwObdEb725xzPAAdkb2HndFXYkRUcBy6U/ROX0yGBJHCYBKGcZQmXklJUigwS0PshoRYjjW0JWr0cl0Jm94yMxxKN3CNEtpBtHF4rJVQ7g4dZjGw8GPtwePuU72VXJj1mhoRASYn4fBt/xz7Qwmhrfc8Gpn10gVgGQMQsLQNAcQAoa2Bx3x+r2cgTo6ECYz2SfboNKARm+ZyKFGv83lohFKev91/xId7YoYlyJqer5fOiA7o5pWqMIqmkdR9hrlIRg672TOXFd6mYc0tCYCtGGDXHGQRaT0lYa/ttNsnt29SM4KZe3m7NHKZ3Wv8qZE7u49p5IczUJz+yBOT1xyiOBUNXUBowlYZTC5lFLO2w/mW1HkUiVLCLNxj5k8YLybXivFJMYIU4FYgelwhglU4QhCStkkXCjTYrMlf1V5r5axICH0nkDhCryxjV530wSB+IEm864+JLPEqwy98Mp/229t9Byk9L2hr40s81c2KmB8LcvP/Dvd6aAxafSN1pE54RqVkJSM3TJ1M5LkbDzhtTJ+P8Lnc4vPjUhYyMxZk30jXB/lz0b9oFTpNPR8lrxAwm/eIgFxGOfonk3UOwPMgw48f8qsD1RLR3uilx3LlwdFlNH8EFxIEnneVoYebIdTmgLldYpGmfOoDdRrB10niVkdyTT3R0EJ884L6onHbDU+hvIH6iqR4/3ez/8gH1G+ITPQ4zVPgd/7zClmDGNIcFqCugkkfusoQOuWGTNnOqR5LOdnalbnMMBmKYn4GB50ref4WG8SPRPYHcJHNnaRwoyh+qeH8DmC0X4TXAROB1yuj3Zslzo0h9upowNEey05rVME46+yT7r5M0fCUWwZ/IsP/s+bxA7krD/9WbFwXH6JeMkrkVbYHmJrNRrP39OlSkOrHpjD/v8Z5TJ9evWCn+/SxWPHXtvBKPc75Htr56KSpfc4bjPCa/SNx1k33wHUymdr/r/NKUcDv/dnJGZhwadgg8XRVqddMRChyw2CWRNs2k46Vg5gSOUg8nm7+vaj9/vknUq4z7gEHTTsOwJtsRQybb9ci3doEcGbU/TeDYbvFDcpuGW2w3BEYlHk+rL1UUV9X4krEW7ka9yAMvXRG6ULns4AgbUUwYXNJud5R6fijCcgMW9wUJzGx5vl1OourN2zTIDI6lLwfBWFSKahLpyDi/01g0y+pV8RbRq5/rZ+XsRzz1FYpFLtYTY9p8kGATwmtjRICe47lmThQcYeaV6jYxvNwtDvY9pB5R/8EcStlyKLV6AAZcChnXA7EVX9cxetxdG3YcOJxFH/lQZrd+3u+J43RJIJMjf79CUackOAVbsaZSWCjl2Zdu9eMZNdn+4HLb7o7tOimdoir7O/F4D0Bb6FrDFLpcYxUZqnLMwNpnzEi8OhUidxq9/Ywbyh4VuAA7aLzhqneFr0Hl7DFr1sNJ4Hjoflep8kYNStz8/SXF6Cty5t5m7yHxzkTy8y9D/hXXXcdxYpc/gkuQazO0kQKaLAgbpN1HdiW6kCpAFSti9GH7VgNdVv0fcClsOx937fM9Fcy0DhHmNt5Sb+7qC+By4U5fueiThh50DKYTkmZHHfIOHjiiOR6wtSSHHBs7H98VmhkCsxJONkEmINSR0+MjoaDKWTw7UgPsH58Avh6n9cR9Tvu/MrVDmWaTPNWNjiyOkAszP/BrkjGweH/lS9NgePhuJqL+8xm6KJO1yuYZcFC4x/SDk5VH0NSBsJhgnors3HUQRYrFncGotdKI8SuqyNXoVSCWgycxPcgsrPdY0l7Ro1ciB2fXeWqgCtT3/dj4MIcKBeCy177WgHGx6vjAWB70cXkMOk27qH8fkN5HmbXrERwLrzdtF5CvOltbwP8z159K9TOb9jiOB2RbONYKLH4Ps5wI1SgE+sZcOqEEDJRPQPNvZnaaivmnKWY4eQUIzFfkkpfKCf6zUGLqT0MMo0KHFy8x0lsSRCoWJBR0pvYjnLkJzyCSHz2JmR22+WcLtM1JpF/uUS+Pp1JRGsLQBRDxuyGUWJT7p7Kkfgl3iB/OjSJ7+/R4tmD/LSIMtv+K1Ruauy+iV/h1gyRrMhUq12Zh9zNwAod9jdVZO8aeC/0mgbOFpkNkiwsbfHzCEA81WQkHExzZJYnwmeyj6le4ZP35sy2viUruKqmyQI7BnnQcS3bjhtUZLSKajesIcs5wc5DsigkaZNv0WkheE0kza1fYvANx1rJCJnWjash16ObotyEqowkZSw14Pd15gDOoufgkbLpC4dlgFc+E0YRz+kGI2vjMjkaco0ujngaLRG/O/BiWVu8HvdusY8UBjX2UGdlumsan/QYQAJUex1RQr2APXzjJdceTBC7K/UbuGkYxlPp7wAoPL4YxlZKWplZcgqX6wx/BfMN1IKqnYdjo/XrQExfLKT0RhJGfnpbIgEk+gBycw8yfJEMH42mbeQkZO+u+gdAfAdg+NJzvdmQDQJ6zXxs7Oz37pdYvl9kEBnsUG19luVt66MBkwEMh7r2Gr+hQ/Ny+d2DK21je3oEIG1RXuIKX98NSra48lTRF+ghbTLiEtAwrPk64K5chz6KL2taDfpobd8W2cNzKIJnVkDaHLVSTPLgf1I5caupPj74nqX2lvbWk/OALrVtN9dmdt+wF70PI9jHz4XWV6bxUiYZHtYJ/Ww3vbu2vQX8GGuRB7AmWsUaBN9Vszu409bz0pad0tP9Yk6fdb5fOelV+SrvNo+WEfn8QidTjWst+XPtoV/1STpVZciyjj0oLm8GlqN3UJtUdC9aAlXl1mjyGjGJBfV+zk3GSw34bSvleIpXy1i62BNJXrE2jHOZITbtIizAhEDa1+gmeikCBTgUl6z52LXc95dt106HikUeTWQHC10sJhNy1JUtviAkUK/VQCQ2/xh2rxXE83w7y0NnspDSiFrNWIWlEdfbKlJZyrolJGBApiLOqwzNPOgbYXCwh731E/JKn6XUdhxME7szmqxXCI7D253E51HU3Rxxci5pce3FIH1z5c6NVyCgUNzdomISaBbc8HLIdfn2BTZppek8htqrdg1e1t74ZoXKNHNNekAf2KF6px4pRwzlfNLsbpkvt7CTrK1HajKjaGy6LpTu43qyWLlihgUMmONPsHFght7V50h3W/V5JyQaqt//yJY+DerxPxd4B81q8Vve18kO0CR0s0Gt4FC1I9YULAXmPkrIppjHIzVTph9YV83AgzO9gJWNv16aGaFGx8a0QsLhYdhh6RkY1OUosvCil17WvRLTLPahCigIvQ0QIF2AC8dW2TVjtCewA5j2a4OBwCWt1EyDIqQXNFWj5n6BMdFePt3mmkP8ozvdVJtYcMYU470PPcWyob9cq0A6RSJn0OriQNqxj1AWJ5q5G4UVzI0/redW2w0knlUyRSEFIBoEsbwe6EBuLeLwOZfVgfVXYdWFY2suDjLC5mG2AgFcBZS4Ol/M446+VlV6e3AIyFB/ZZwqgsoKfnbqlKZVTVaRSNZzwmgU/dvac5BHTKj6YHNx8EsN9aY5f3wjYf+E/5/NYcN8Or6E/enkDXypXkyzz0lDfAdPMMctYZb02jKhwuI9KyvBebGXTRFeMIvB/8MsS7hIYOAhGaYzgFX6RCTuc3FO+o4zxXR8iz/90x1UM30KYN7KtLYPVVuHfmDOnjg3wr12YAJHh1txmfY4XLxFCkPof2vc5C9AVwt6+ye4r/a6xV8fuQp0qvnCe57PgECNhX4CND+GdDdwF9qrhGKE8g1oUblccP24GPuhw0qV+bvnwbG7ODWXJHDCFhMrsRBDhXbOkWgI3w6L1RTALwNXwhYQYBFrTS6a2CsucTvMvYXcz4gWQVH4xq5hYm8szRu6ObrgeGN7kV3YyXpu/gh6XL7L1r7NjYxAWXbLtYZ9wp8NdVWXGeGUrvzbDjZVhcrPoRaNGgu5LR9s+Odn+Zu1v/SGHUuOWUBhtb7UKO/5JkIVeOpJc4ll2+NGrO9aY8NWnRz6fDIYIIKQBv/dskXHcJBDF++IoONDc6gtt5DzGqELPbHSgt5yla/w4Ak4enmiGYMaY36I5dyv9VvCrxx71PhnRyWiRhgaTwS7XWbZJbLG1yPHQcrHVOMAp4DdC5HVLeL6KW/7Qo1On7wgVhTFtnClVibTm+jC0RFEgl22jZHlo/tduh81CNUk2ihztf8gDV0TjFHxGquK99itrsUq2NeQK40mWjw0FSdGemsrQPvN/GVDI6KFdiIOnouWzYMvU8nrjRAVvcLMMg2lE+Da0mG7Xlq0JTdjF6LSwv1wfoKwSClg+iaSun05i8jugUUdqECKytq4iGRgNNkp+rlCUPIf0qHInYqPoLzGCQauqgUUDVdkMoB1FweHh5oAOPLBpmfrXo/pTELDRpmn1Jbqur5cFDcK64vJpuK13941mXc7OVi5S9eZc/+0yjzjzwZYx67qGtgALc492qZEGifM7nwaMihig5L3YxjtAX3etLe5/fVOfZLsSnisIoxXHwXE5stVAYC7dge08hdUyYMJaSxlbXxPKRQ7n5FS8lZGb7iWkX7zbfPN9YIM1InB4infoEMH7CNfcnmFu8KeWr58vkgH/ih53RQLnHOzRqN1vrgwxSuRp+c/Udix98q0BnODBoMIMO48P2qeJUwuaWwPpozZECBZWi2VdLqssIScK8AVQ4Ib6LCVcqM8G9M55uQaV+jFu6rvV+DdfD6NeYzXvDATqewjVg44mvlN9CyL+WnIYdWAEComY69+huNztEMNw7GUjqailuYKzge19u98fCeecv16YKqHYjHdvsMUa8DbjIO8sXa8G+RuAM9pIB3AagbgQEtPbWnZed9titZHW200Au4RM=
`pragma protect end_data_block
`pragma protect digest_block
d31dc38e940fd7808fcb3863eb119da401bf5fb2afca1216f496a0e72b04d5dd
`pragma protect end_digest_block
`pragma protect end_protected
