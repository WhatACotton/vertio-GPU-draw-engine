`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "e8b2da194f101c83002d3bc4a5247a45"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 17787)
`pragma protect data_block
jLtR1cZ4bWA12Qz6YmWF4d5eyCyJ3Smu41eU393zCQ11VydyLJUh0kglsG8cJ2kBHUooggOJOMm3uvi35suP1OFhZxwc3/ttahvoaJrZa/jieiOC0+tDShn4twc9CQvo/IUN25wjulzjaPgqFDSt/k8QJoJ9TnmCDTixONHqwLV7vGjE5YauVak4Juy+ND3IIybEeTwhSl/WMgxDmPQ4SA4aB25ynOjkN9Oejf3A7giSwYZNUNsQ/vIg/BVob4FRDMyI6Jdq2q8HY+npcbfNwzdHkumb6uUmjC6eNq+xiRdCrnv9ZrAgIBVsfT/1gHnrnh4ELHARVfETPreZg0syK/HbQTvoWmuAle0VoFKfouNlZxS0jMY5Bu7tenEL4H1JZ5A1LaO2HZsD3TcQqgrQ9cImGyk50Yi9HQmZQDZhvp9qHgCo/71FLsjs4oSVyTkQEDth6hVHqoF0tCAdt8KlZ/zxMB1YztabW2tIkAGFmxcch9g+Gziqao8S+QXRgO8Q6IiNwWNtbw1wxktDMxoj4Y+cACkODnRbVkzTb1CRg6ps6gZS1prHp/qxBDFkFFPLg28+L5nEg4rwJq4ovyqebzYVplFgbNtrAX9T2Guu1pxAAQVHpM6g6xrXdFObe/AU3NcGzEwNUvMWucBGRdFqScaLGmZuYE3PaufyE5X/uLHVGNKemHuqRbMpvOYYuWGqAvuwzMcedV63h9/h++1W2+wsrTde9kjG5uwPfLoghZc0Y7IM+n/nzKn60D7IHlw0bSLOCrNElqSvNurLzzJ2X7KUWq4UUvruJte30A9gc9V7GVoF/rCQcC8H3Fw7e2bOay56yPGZqOyigIqAVClt3l//oPqN/TZ1JK3w0effkL+QKPffEyoeOLYvAXrD8cD3t8RDaovKTEQt1hPVNTrG3JAVXPJGHlxf8sEyQrTxWeH6HqpzsimrJFdle3J9V9XNds2OVDksDo6bWGMN+wzHrsryDxPJN2/uGFAq9nzQVQAToE74T0Ej3WhdzrQusGyQS1aVmea0dM99WOAvNmSgiyF5hQZiyC11UnwjT+t3ZWJcPt6czGcKDnb3u1kBaTR+ve+3vInKIQqCpF1wobIPu82EfPP9kjFP/VuUrR7qzdGIybkH57HIHbOHTiF840lsLY/wUX52bTwUHOZju7yDRMUw58XAo35qSAeibuT5dC3ugKufQzKQTVv6HWXZ7FQNNEe3pkAkUqEQvW91DdoSc10G6EkqNd50IsqmxnRmtoMOvE55C2j1sbKYQcFA0+U2EXJ0Qjtdzvl/C0QCqqCFpDPP03fC/LSTDTpT2nNabJW6EyEoR8DmruiKdKw9WscKpLwlFKtREhfgWnl5vns5yWSuSv8vtr2gbBYlbDg11f6PWXGwANlTJapK+xkOS1Fsh5jO0VtvmaxrREg9xUs3O41TYYuSpzkL9Xg6KL5jUThdlgmhUIHaLFq1+vpsmLfPttTz1gyzLSSfqTG8dkTD35KyNLyMSWluUp0G52nnGQV6GQMbvmEqb1TwE1w6mwOwgPAhnmwOHkFvMF++42pE67CLSQSFULAgZBLm8N5fb11CIBHY9dSyYXgZ5iClEPQan8GPzHoVwc3WfTDmtPXKOgIxE/7fQ/lR10XQDFAG0+n+vcp6uh7BsUWZDnDF3VKefDgXfkKlL6jaX0kBuBPu3e/hiX2srqGawHTCzVXGcHTro438fpBKiNqrUZxVWvS39Li5V28ezT7YpMrC+nLO8ZSY7EQFyZdXJsY5cyZd51cCFCn9xMII1WTmGdidpxNVIG0jipkE6ZaehBJt4Z2sOoINZIPsmCfi5zaVUiBd2Hb/u+bWN4z6K0RdhbhnNf9leplxAjdi5RhFAHTo+zUkXdaWwEPWvAnAkCUNcVhW+41HVWYNRA/2eBpQRiyBWjx2nzeBb9I99TLnd8/Ub8u02YoaCh6I22Nkl1JSsWH2tHjt5TSWdzeRq/eohrPigm2hObgs/E5pNVCdFiRF8TBFPhQo79KkwtCxWEpugQbGaMrbPqL2VGH/ZYpUBd91nsh4hET5GbwKxxy4+Bk/0eOZcl5pJ4tkfd3lT56D8fuRvrLY5PMhQ6EXQZY81sEvvyVNOntWXiTAzZ4cOsXZ7KZtsePpTG6C0YRSbhWELhtTYFTmo8OS1sVKnHHXR25CTmNhTif2j3QnLmOTYePsrzEG8D4+vAgLMDI3+bYkwoBx1Xt8d6z+M2Yz4g1k4SsxU/M5n7KREqNY59hIHpILDwORx+UZA74UtMRFp69uU3nVkmniXi+f9xNjqbzy6qMlm2MGOMpEUygxujXlnGjVYXzZct0h4vPkP7Ba01oHWzyp+alnpxfdppVrSTLh2hNf/FJoaOGtRiItsADQgcsT+3bVOW2AEEiwFQDHjnNUHQHvjTlzdP8mUwzXVKA06jft82KRekjVHC2iq45dc7mTZw91oRJ/D1LTU03FMHo/VSGmXJfDeIb0z1/0z6AiF9mZgDbIGq79ZWYQ/Hc++VcMSx37b/VT6qD6hDdM0HQap8SoAls0ImgyFVv74jAy0muUucjG2nC41UoZaWOl/CDLY3ck6/AFpyY3gQSQa4NI9gVWJSTjIg7fp+MXoyTXnGE9WbDwWDCAZZpn0EOvgEbdI6ckLibymqtmyexsbVFz3+XtyhN5FWp2CSMmtk/qvAwxHGBh5PpCtJtscrnMIjodFfOcKW3h7G1YFSANuueIkiU3Z6swe3el3LkHX1w5hMkTHxPcn4j9PMUPmb9DpJJ6h4vab+lwunbi4u3CaeOQXxFZrtRLBpQ4gC8TWA40Hbh/HSRXvZ7VCykI2yUX/5dCKyJ1lrcsozjblkk3fY/43QmEoxBPjvdHH4UqdMrR5IgeGauoVoI5NFcTui2hRKHdV4NzaFffRDykR7YoTiK53S55er5mkfI9azSG31o6DtrQAe6ztC41o0QVI1GpIcAT0MgxQQHWtuU786nj9vUit/0e+HynTpm3SkQCO17Ui81wkfsR1gMvR6vOjq7qXBG6P11qteNxAQxgvA/XfP76IW8W0BlSBXKzBMEYZRzORHa9pnohp2XInkgD6C79u8DUKXjad8yivgRzop/Y58q3YmwBK+PXS6quxFoBToYk5sLsRtz0AwTlaGEQPwT+y+od2NQ2rCFInESnvUSyidD0xNvA3JMhX5NDl7bLSzQpSD5cz2AsFTYvFRXpcvA/c15ao73I3teiZNhJscxdptvn63h8FeBptxObw1oDzqfv7jd+oVwmtGYaUftydUNBZPpJ3A7w+SfJmDQCDxuQGk4KL9XACkgpdvoTxXOHzNgSlkxSCm99x6zpiofWrXOdbZJZVp/GXdkBblGRiAOCUPPH/tVZ1TSsPlhxuULN8/jGd2XQAt6Xq28hWfM9ExFMnF/F9L1sOBUVwEfSEvIywGmcXVvMOmEWeVzIHF/zPSYGCI3p506MIOtP/OPR5YYUWVSGcJr7MtUSqUUMJ+0/4O99rex18FhyffH0qkH6YE9TDUKfj+927OzV2J9H/n7F4ZcLZZ94pbmuzB2xcSFygNaLToYa06Ne1EMotykA/e2DI4QNhQzpAubcSHUSm0yeuoUEv9wd7SFZJNH8GaYB/fxw8fw61jGx96TTVEdOSlLA43EgyiZlj/1o82zNtAJTngD5xCqzmWy93gwqOZWAsaE50R/Pltt0fKfXyAckJZ1WPN4cIOyD5v7Llf9pD9zNfQsA5T0kZn6os1Mo7NYKBRM6pR/9ztFAevgi3yh/SVZ8fJNXhDqyQQSNv/m1FsID7KCvc0/EURcovwEogylD34J9+k49zUuGXwNJL7tHaoWurhpRJGcz/RtxJWHNgq1XY7eESE46vLNP1zt4ftiv66xC6LRIWKFfRdjTeCOoXquraup8GwF/iAvfUcyFJ5x4sZVUwHnij9Zc+gO0+yi7Qrkqo+3XjcvWJnHaqdwcAnMh57KcqEGSXoPpwxS/4kEqqM31RZ5CxilmVYjKir1N+KFw41FtG0b83+5MTiXRN9x4cd4oJ30pnATmrbiKyP+R53LtUUNIMogMd3nIyeAl8WtWt0AbWXMEtkjtTR4iFNraJMR2N2RfROmc9mOs4uF1QfEJ1M3mPyRiXHWHFBq8n17Sc4Ag2d/R3rs/kZSZPr8+0nRbMHeoLRxTBcleDuqhKdx3z6P/EbzVFJHwEFApd9LTlEvaPyHw7764cAIwyEWJk9TtXNQPW9NRZfVl3+eX66U9pW6ZcgeAza3t0pShKq1o4wkYTmqqHEiDQsT6AkJuDdOETWztOSUz/Ocn78aldoup3DbzvZgMXrctvVGhknqIy/PubsgTBzbxYVjt/Mq2gQX8mssdsoeTXnfa0tSmB9gk5e+ok0O2PKtzB9EJz7ewoIfvu7m6WQH8keHo4bH3MxZ+1OlbakW9svUDwhdcmDKDadoZgNKI6eh4zVkIzAk45w7NWH9P20bDx1v/kS3xtb2qrLbxdVouNx4N2UeS6/akUFSfgZQON7p2xhIVKyaEtWuEHgyRhSooQu2LgtR+eX1TTq48gZicsLzc6KY8joqaUd9ldIkPKXxjn5rCd36fVWId0obZJWWCJ3wdebBmOuCFdOSgmO0xjZustEowdQBfZZOc+rwnmjRIJpWzRx+BO9L992g6q0p8q7zFIDG50UbH0T/2ODgHD6sKZgBz70vIxZxSwqYzHC9uqbDcEClh/s6NU3NFsHDwfHQfDUGOavOlAPnOM3zV6G5kW22vIW7nPYCLlzXvZAj7PBrljz+TETCMCCrPw+pfm9MsLmwC8NlTO7PKooR8ingqCG4sN1e5WFfq4FWpSTpgRgveFGoDH4QUZG+wK5MNDL0dI/EXPWwKwJrM2TnprZk3haYiEmYWMGK9lWf4kFrPFbL/tVh+yW+laiAi+PWVPVo/8WBTxw43q6CeuQLa/ekngxl+GjyHLk/IJcPQpAKNGk3vl8igRu77OI7CKEZKogsUtBPKRvHDW7sUVVKa34ghgcxpGI/ClwM5JV/kv7A5JGPI6ol2aSXVvZaznn+rzJsDFGn/X6mcX9YALtWtFfTyVIGQyWtRGAVsZ8uT/UTIV5RMhgQQAboWzo0K1X+433r4crfs2zGaT4zSY2r2NW3mkUduZgm2Qqaswf/KlWiC1E4oag/NkqeDsb0Pew4nnKMuVELpbEvSbxukE3VNAQ4/3jPgw/CKhW48BRnJoFLz+WJ2DpnhAnbbepQvtWVzvqYVScEn6mavUbBwKjVluQbh/w4YnRFiPtDab+F3NqLA8e03BMmhMXtJO8KhTgV/RM46uSKmI6cexSQtEocKuiBWeh4N52or/dS4iZMNolvuME3vbwvu+fFL0UrDdV8jxV0Ibx7X5yflDXeDyfWDSvea/f+GF3UlxJ8bRrM4e8+OycQ27cBYs/1I6lNvni8qWx8dIWdHCyQ3Pcbssm9ew+s8U/uYVuxuFFo9k9rOI80/vEeO+v1SG270HeJT0jwbvASlZYUZceu8pZiUl4bnX8jMYnz/xgB4i01mXQg3mpF3v8N+MycYPX0oYidrS4BGDIGYbd+YLFC9JvjAQOtXJDaQbTeL+zwLZ9qw1rVbmsc3JbrOEkf4zE59Hb8ObPAJ88u8gEP6MvuZlxpC4cUPYx9woS5eNnBKtEPqoOIKfgh5cLR/CmiBQkf49mCJEWGZFNxOB6QiaZGLJ6djwb5b8RFj3VjVf16GaiAJ3HSb0KQRYdEVESlyEgyyYEERe9d1B0hJERYruWcvVsZ+nkAfZGOhqNXPVjTzLMsF65GTmPDHxZAXxduz/vbx1f9ZackwJvx/2oONB87BMzWIJ5Ck1h2nL/LHlrYhb3z2hWbcin7NYvxAUNjA/p/+CEPSDsVgF1Pbn0B+zdCCbyFf3zFitlxoSHZGgcBPmppc06CAF4azd5lM3clOr8j9qH97UfNNtBpGHCVEPTXNc2Jxc8+1Sn5P/cWvv0E+hT299LdzaH/l87nrEf+Gp6Vk2vjxKnoVB9hXTyvyV1A8TJzHwidaVQc+Ax3zcKU/RRKAhr/9+uFaK4JE3bG/ce3BbYwLX3EmGiID/SGgBgB3Ex3i5iXcboe6F9BHXWvHxb0lfurN9WIvvsnx5mzfqJ2LzDhRcn17SOWgFfOYraweH7uwycjNUtr7wIxKxxeYle9UpguwZ6nu0qypnz4v4FI3x+qsl94NSB21wCX5/B48lZFFDLLD3yxkZSJ2Y6HDy7Di0Dq2kVhCu8tqwR6rwd/vqHOc2tlewQowGf8SNgCaXFfKVfK8dE4a/F2uSuIdB1gQ0CU7aoVVnGr8EROZW6eI3Z3+aU7scogcGnVCm3Pq2PzU08M3qojOhT/q//XhmJMiEkuYRfjo8NbTbli/k2oceDIrSfxE0NoFKTi+dHOSQubzJ+EcnRSRTvGj27Bjhs586dWH/tUpTdfm6wAPcF791VjHAcRvZUKeHRCz/V+ICqEF2nJfxTg43gYLn1dErxg0FeP83dueZ3Cac7V+kG3q5jGXA0MB8p6ijxIdwlL4EHuHH2K+GjZgkyerlAndoOvoJBb2tEYbrP5F+Lb/u6eRWashVON7+jzf9ixi361aNwMnhf78vi2v5FwefRj1Nu6p0BevBStZKvd82FqhHvKcaqqiTMG4ldNdJiodyhxHSG03hdw/KXo+nqh++lZcMOzPC74ZUg568+Muitm0GMsXdlDFym7Xv+/o1D7/F7PbV8uwtvok1/ymTfZNd83zNTRXt+NsAMTICVOqu9v4/nxJdzzxoaPfWP2ooKUdHxvfSYTSbmOqatsyVu+WlJXmCHdlzsIbMkFc7GsRmvdDRk4oKitAYR/iFKPI5+fljY1W6eG8tCH8T3Z0xSAE+cgeBuXmpbCP4NCv0SX/6VZ1EeVutQ6APLXZCpFuF+KyBVi3oEHK0evXndYTwGXCmhSRAmoWr5zFDJrxTkF5R1zvFltRwwiRR+CszaxqzFb2Qb1cjJaqu813nT8Qa0Ac+UIRTeT3SmPLNxJWoqzSdwnxt/EM5uOLna9fUUFqO4ELCNs1wraR9y02oYyx9gLCkn1bC21BiIwYZRJRG4th7A2IjSE944LsRdiBLFJc9yiPPwA4uar8yiKYS+xLCwu9uDSIExYOebcvf1k5adaQzaNaS5n5tjO0rGb6GT47hp0RTHw9Ez53ZnvufBJFOytzMHsWSiqDGZ5pXksnWCxLLpeo1nfFrK5SfxVAecKMinplF/zGsRRrCLa2c4Lf6WSlrdp1LWyCaY5xieekGsKzipN3W/k42rkoEACGFw5K2DrtiJnSpzZq8gYiQZgKERHp+e8hXc1eW2h9HsoWrswOQwqnQu6SAICVOIZK9DIjDt4E5FSV0LSDSKY6yKZsAMruHDhW4nMQWColiXHSutjkW6oQOn9nXpwm04QXZ+V8cNYGmsMfVSXjmblK3I1Ozcs4s8WJ7lspwAC1qG+9p190CtjEnkioJ/AsAEU1rcBSdL+JRqzSNUBkX9etBcn5g78d/xlF04ZDLfqZu+Ox44PWeYAnv1VCXRqU+xo7gk7hE3mgj1pCinBax8vKNUmnXQPN1/b4/b5c0MlbvuXiJ1bmRpycuIamUCd/ZfKHASRS+l4xn2ytR9O4S/Iy99F3jixnPZBHKD7LiLLm9cO0JGzXy6eV1S0hCTyw6iUl+3ZsgNBxub5CVSh/NhDKLbmCG+2k/VtjA/NIsdDgBQrSciICnduclug+JxNftkjXwTUfrQ9NQpHWxFW1kLk4Lvu9qKYm2xV4vibIWf/vQ2380KEsauIID5r/BHmLKeFx+ZO3ZLvxvnrL3+OiG3jhZwvL5P5IQNVeov2ntoABND/o29n8U+rCUkGqXxcsuwxIWrIuF07uRWNuDavNa2z/k8v7EDLqCSRl4RhLsVjyQl9IWIxaxrcLNUgpGKPxsNbymdrIAJIZXrjlSvfKFRHh1ssnJyn6RbhzgFnY5iQT5CiJdavRvvUSkeie06IG6/HJEUSs1Mk2Mo8x7h8m/Y/dPFKwQxwP6HA7O8ULVx2/Fm8AC+6jaO3hkqyUDqVOX6P1aUAklq52C2bKrGfJI9but6feADFPQrLle0MPCz92B+zgNtI38TRidLVS/5C4vpXLU0UDglJJm27Rlx4hyYUDcdscYPWauEFFhEJO8ZJaYrf+JO89pHhZ1IOFrGQBOYOlnC2LzgtxtWkIAGBZc6FuRzTHOyF431dWJgZb/Ej0vHFyfwbWTusBJ9QskC9RAbGbwZT9FTiZiVCa1U/rBriI5ISplbqmsvIdpmSejnMknQYgIJ16PKS9Lv0Cel2nuVK7d9r2jPnjBBH6bB4Rh4BcAP/ey/PgYAddc7j0GGz4papbnpFBExdYch7UaQma9khXErZVQeVhBAqN0HqjUuorGSOfnrDnQ7xp3cWrAYCuPjY9tGPpyQGlbwa7skUZ+4L0LjiotfgqA96gL3/MQCEFNe61FEkG4UzV4YDuw+TMPurJzStGvbq2DMT/PpF71EintKgCEFEr1Zox7SNNBfDVa51bjpqekLnCUmYik0FW99b10u2LZnWMb4qafryeMC+KD4L/0OxYEjVZy5/p0pz5Xz0IY9TmgtHXqvWs2qtqKx4e/uNDuUr6G+mxAtP9fRxoHgL2dyLVxmu+6MxrLIGS2Jtz4uqTCshF7llG1RRTXfNoLq6JN5sJ53i2iF8zfZPxBpM2lHL7DQignQD7Mss+Hw8c/6RG5HwGamgkXZOPW0YJDyLBG+IlkCD3s9yWwFx+hOSelG321OqYNz62I9QplNCMKuFsKyI2AvgRQj0s0GukgYmZUl83jh7RYDgUNS/PmAQgy6F0SV+5aRe4/ss8BQw8s2ujsaNucBMYxUQXI08htGcRpkYICnsnAp17/ZR0g2oWH2qJ8AYFeVow6HDcY3E9f7c8B95FaPWr3UAdMrVFHJT9NSUVp8tBzixe5wmz3xGX2Vfk56Mki+OmTdiPWpeOUpHEwZzT5bHNBA9TQehYOlD3mTaLSWU2bcUhg1sckneo1nThqnru9To9xoylUtPWdCVTpNleRwdgnN2GkG0eC444KrS/H8QwynX1ClH1FaY8Yn+2qDTz38O7QKza/Fty1JZfm6tcgbKCR3GMPLmZkjkZPNNyhXH5hCPoDOhpUUy2gIu18jfNw9vkxpG8dbfU1kQBeoyw0bt/PPOEKNYmPsdm03Hm32mQtrRHizkCV+n0cXYtwVhUPN9MFarls4G9Ao/L+1NUMI/h8AbuY3/yCy6Wn4x0O0CwqTBzeQaSA05HyA6N8k4E+Sxd66T0wTFs8+N8/oDlvM8pjq6B93HNDqZILgl/WiwaiYm2SttY5rw732dZ3IhL2SkmHnRca54QxP1bD4Ri2ET816dpEwyf1oCi9yNJxvIDZh3GH/axKwEAxDPXIe5TWzJdTf8jp6ipvZJ+kRdjQGNxQZcV+n6P7j/jGuN3Svh+ePzaBOpKeLqKZ7iwDuiDW3cclRHH+pSSSrjgs1YouRd86z9Qy/NoWYVrSID+X2plHL/7szjLk+AIH5rNPoozeV0D1jiM1nY7qSoUt4Yqx+QrRMynNyrgGoz9+6j/8YYMgP6ICLC6/ieYBBHjlX71iUtnGHkXnB1k3CJ96GLope8EwfxPFi84hSB+ZMxXctukwFefRWbfCrJ8n442qDTA7tkhhY+j7vI1B6OBv2Tp/X1JsBS/1v5tBIzox5VGeNnMCOxSt7PZYXkiM7rzsTn61Ivyx+JcnZYDyViLGUooOP2F/WwptOyNByJxP12x89M18MHfjQMsoH8m6hj/nPAz3WmxqYE4uZgmRRZoJ1JssTMbc9eTn7UlTLUuRYKHAWp5Szrd4NyHUbTx4WunU4SJOPixLvM8BbRasLTQQ0vhtOQ+hHN82AvnZdu03KNqk6gTyJtSORzFoho6Huc2cRIujz91FWzimkBvYnkEolXFmx6CpfKquJdnMNpXoJTXy5BafqQk0cUsI8UGj0bzoqZinsZPGs7HGUmCmtcU0FSIVJqF++rz0buBR/F5VongfKtbysWawIYlJ4+lPIJP0/FSSqv87g1TGujE5AqWBjXJJbnzs55PTjS0bC+zOUTCsIZDzy8NeliGU/Ay8/RH9LkmfaSqPFJy3K+obzzuIdpKhckmHZxD7WvaQqFg/NYneW3H5TXNM0N2CqgJ6wHbBymlbyDLbhI9FVgGT6kMk6PKUdKSQ81q46h59u3mjuqXMQxcsioS9M48z3V2VROUPzZcsYaJqxvrr6ssGCSwLw9KQj3DujlKbydDUJNDJUcrARZCwPgqpp81NuK/hClYdwbHdAPvJDRu0vOR8hzhQ6cjH4hOIPVDvMPWVW5wGCkfFB3Bi5xLzOBZZvQfPMMECVlpV04/1fGNJFJ6S3wD5Lpy5ug+kUgMuG8vAgV5z7iJdYLFDH6xaYzwI7OqpRxk2Lz+GuiWefPwp3N1m9gCB+XdXQKNBlY5tWprDM7SSdqCix9mS94yY2eZK//Nj1nZc7+NhqVAyI4rN+ZPNPkQ6n39hJUhGy2eYGoiWKbLNKxDe1T9mT2sZN+EbsF65Ebx5CprjIK1E4EbjdtGdRagAsVQp5bQHjGwkcU3yIygUOZu4WNZCFMLhn/fDnKjlOpwSauY9dQXP6R9PkhovGo2i7tFTkMiez7r5nh3ncQ6vtqvAC5Digez7ODakz1dHX0j1fipwoXZab3cJ4RgMh4YgEkWerNEp8KaMYATckDhmQGyMkRxWKUc4wCnqUrsVIhrZFt4tONXiTVXkfeuTi9wGRVbN/8B7xABiqvRTodwweeT/Mu+6YFXPlDndjqgLOaoz7Hv2NfwVB8dt8HQUaRIgUheCa5/iMQxLtuhSbUGSyAC2YIrwBDF/fRieCi4v4xxTKtvlVFxUKY7Osio74Bq90J/8sivcEsC/LBtf7YmkybXsNZw90W1MtCl8esgWfo7STiNYY+wsioMzMwmIuFsq64IQUKkBSjPa70u8mlhkfHRNRIUbEZmz8E24xcTQ8Bllf5hgwJhjGXjBU/it0M8X8DwsWJmEKn4eTmkyHXAFsPnNi0Pjl0bMOU7H9Z+8x0sT9qUch3qMh/YriCJMs+yBXzQfXIta9goPWXmFWV2WgwKOD40KM5kysTO6Hs0tLr8XbhroHrtWn2PrYoOzam0O4R6fYaahbpGbMbJ8PipTjbxsEtNqwCLrpR5o011is4J2Hhb7YmxPNHwIiBUNJUc+64H5HSnU43HevKY0vUp4cZaOd5ATi7gVlnPKTh7f2Z2P6hKqSpcIlmtPmWcGW7ZBQ+FWduXArtxauBWcSMacp/2si5NKkJJ/GQyUhxvPqWBl/8Rn9nrgPJudDwXbD/LvajMh5KtGBPh14ot02B+zx3swKfBWxHuCPhdpnhlewE86gFOPU2KPyv3kbJVaZ5M/YCjapqUZrMzJQtrwWXk6FJbWtubp4trmXKp5MEDSV+9Jrdg0qoCRW8/eFNEHstpEY5+iGQ7Mo03SoPf2SK3KoqqUobqIOn3wt5hTzwHz+HvzomtVx73Lv24PtWFYHxphgN5k6773IbSljSTk5a7F3hHjNIzudQMD/ltBlhobSG7LPbJoPu43FsjnTgpDpYhy5LdjAmlLvfgfvzXJBxbnl4uFYs4Ck8Z65H4BY+oG4svxWuNEeP/3Nyt0jcq7gDrDXAasZDxFAXRXCA0VifmZ9HKTjM7JFGb3oEMfq7nxVLdI5aWQGJFwp+7Mhi1Vu1fjaZs1UUVYDngfAeOYljI5w/ZbxPc762nyFPRGO2lIJhorXEQyJVuPOBPAaXrf1NLZGa+5oblJGZzvshoASrs0ljXoSOaQA+ppjMvYJrkA6p1O8zOlnE1x9ToReVFvWQPDLd/Yn9Y+gOW916CbJOK4w2ufLTVOO6Wa43eAswtqQ9rFs8/o/B9DYz6g4MIL1RpCS3JNDcsEH/RFpTMJR5agaw0RLK1Jclr3ND/SmmjOYPolSOsKzub0pdJA6KpdCdN/pxtYXoMNNU/RdzkUY4vkbn4InKk6uvcLYn65JFjnC5fLRW8/AoyUue0ujLysSQg/IBHXHZZmoTRSA5c2YZyjhHQ016lSyLKM/eiOq4B2xtS0vXrMYyjge+kjsHWdes1tclai4fMM+8UWaOsSmQFrWa+X824bhqr7sZcqZtwFhFg+R3BnI/GAj5A/dCkyRCIjRelBsAadgV7MNG0tAgJT/vo8A1fsQhsZEf6LVd4UwSev5aU12vkyUoPbAvMoiLrK3NY7Bm7dRL+N6D5OAtWGbVeYcg1ENIu3PuK07i9cr26X3prF+JF0a4zUJu5nTLBmAUHUh62QTsOovBU9VTXnmlH681L/nuqz4EuRPW90/xh2wq8K9jXE4+fo0KrKXSn+SsbrX9uz+BEfRwXm5bV+nOEoKj5Yce68Zjfb8YqM2q7cZu6CEL4WOzM9svtmhj7vP4Kmt2bv6edZxg7yQKG3JIqV7pPMGVAeXVTd5BrVCG6IjNObwmLLUisWmnevZDaT6RPFT6M0Capb+eH4nA3Z+48ofYVgM+ROPVTSBeqztEmSqDVgVi0Yn6RzRNQ7a55/qkVqOFBT9UmCXSKoKTaCUMH6RXjX766Q5u967RRYbW4GStk6rQxXO0IFiumc+6PLTkqq569Wc9WNWOQH0OoNb6YxhvCSe2dwuuxVzO8tiyJq156ZYTQMoFvYXb5a27M3RKQg04l8TWJ5Kaa+59e6snTXUNetKPDw1jxGjgsSp8umgak9SzEw0qpDeq/QWLE8yAwR4z0KsUVTjQ+ct3nTu7UPtSTIHQBnuDzl42sfVitsKGgKH8pfdOCIQ8KY62UY8UyLEpyR3PBvTKN6YlJbSbmCUdUwLCS7E3yqZZCrLtZoEPxvkdbzt2jZRljt1+aMVLkjCVJ/SUdS81ETk3h6QfaiNOy8Pey/vsy+2rivAHsjLJ5z/6aUcupd3gmF3mLMGA7tsK8SLHVyVbjW7No+1zSy2BBSK9S0K72bmO5fLjQATuiNSp3pvh+lL/7+vuq/XxdrL3jqJiDQZVR40w+s6EjtM+ahMti6gsgVOEqKzG2/xILBFCY0GhRAJa7BmDO53xO9Pd1u7B+ZgqTITbHKag1WmZoGD5UP/PK0aOdz1RcwmkwK5UuhNTK8kgJAdgf1uLtDh0jlD3M9y7B3WGvnVGI22dlkhnZTxm7WuVwLnhZwk98fRSNyv5efZRZQVpw+pvlBinx1Q8TMyPtudOHJdEd5ebM2gkVjRIZQrRwjSxYdF+aSxqafRwIbPZEckGP7ZImls4cynqyF1gOLRrlUV6U6eOahHMTNJyYinXH4U6fzju36B3OKG3kTQSKN5yQ62YSkCOpJCynwNwrY0EdCXvCHroFXgAEENJj6ODO9WOU0aztW5eVHjvbGvM72NxnvEwg+28Tp3uaEbdyS5/Gdg/6CDnMF0QdQG7yN2SHAbxtYrz9Z47Cwgc8hBdDuwXcydClZp0xPZb3H1M+DULXIJjpIZ7CrwA0eCttfYpaUFtszBEIvHYMsOo833FikFSNvedvFG9++wwzy8qGO3eEC2bQ77wxf5d2AQgt8ijd8mdJ7AjygDDgTA5RSQ6aneLHzrmgRfsM25o9rJEVXwRywcnlASgqkaTwOqAJGPgBtOe851WcR+ST7RT8RYkvfXDILVl9HwC7ZwfIYYVLxb8seCJ9v0+PWEAPMD2Svdl4EoHKfdoWXQNhYF/46/QzuU3f8oFf1Z1zLTP/kNiYUTGCn8nM66EaL6/yZLDA8/z/8FsoASS3mMxWKsf5C87PMxOd1Eg4fJQB/TmxoyhqVwyZSWN4lenald9urwONgW/OsPssPcYSoR2DculBPbFlc4l9SdDchAh1YLi3kKsK2DoVQJBrCFQYunO3vzi83Ud9+J5TO/CkNzm72MQ2PCq34sefKVzDEPO+5sCA0EyvfRPgQPvJC2hfKCWS0G6BiSqIMKKu5pErXWczNBhkcRXiUxhuGKBe7T32QwAlxFsOoLL+glNP0yAxBvczhMv7rpwaJ5OSQmnrbnDjB/PCVCKrLT8IzfpSDM1zaquecaTamnyP4mG1krquM3fndu5F3W7Q2oS7PtHsriKnOlGD9RtQcuWE4rCFN4irPMLNBkJ00PHGYfFXKdPzttZdufqywl1pPN2876oSKleRUC+w5J9GPhPNmznOA3czi+4wa6yZIQFTcj3KVL9X3OM3yoJOWHaxS60z8QMNoiY23KdZqiR13YdwjfG1ARFHqJD0l3kaj8pHGVeHvr3dzY+9n1Dw0glD37Xc/cdOOCNukqImK9cIU7SbsrtuJaYMwafN8bVgPsX6WDynheKxWJnSl8XgXplvq2+R/MPUK9vbweqhtxN4CkklJceKL17xz1sUmbHQWk02aMZJ19NWJo9hlznF3KnCTx9Cs57YFoMYoy78YhFQWEEgAFOYvfP4bEh0fEXAoANd+NjPYbbJYoSipmcimWC6M84ESFh4kT8L7BZFt3NI62jJOeifeJls45U/Epc6O9vh+FT1gczTZjpRIQW9Rn4gWy6CwB1prei2ANCl7O2YCBNjV+AFC1E0PQVCXE3ZYruEbgSSmhYG/c7HM6xsoAjzKDJQEXs2uTbSQag+Ufcf2Cusfx+q+2JNomXWV7dcUS76/qav+CWHA74pQWPKjkJma4TymcQ4yx6lJ6jLhIdXsB9gqm6/Qs+933icIdreNDc6Eb3qJfEW8L2fxxKNIDxgR9w8vj9YFPMiigmhf6Pl9GE6Jy0mxiCF9MlVx7tayhy2oxoW+Cx9IE9cka1mWNNXc3SApJeb7fhuyUqXg2dzDRdebew89amBQHKH6tH2h3/Ga1DleYSNymEzTmeOPouju2XRpo6FuA5exA3xJMK4qPpbqRm8WpUpr5zhJKXhVgN0cFB0UbPfj9nLm3A4MM9jQrU1avt53khA0Ul/Folf6oWxgzU178KwABu7uzBwTuMWPxPObEeXLl6K5FGuSXGhLsAsosP5iegEb+MlaTpDI2cMMx7aY3bntsGhNH7zbJZR5zqJORwIC02SGWf7RZhVGvraVBOnDd5Ib1wqoALUwVI19FsbpfGt/tdHpmQMxIOzGyayn9bo/HzTB+0kv8YzOrydy/MoMB0UIt0930otvBMQgsCs/UzFFwR4ZErglmdOWqiG8FdTdI+LPeR8oA3PcBxSpNwWZ1KRknKDLWwqykcCrX1Ii9aX/s7coih7W7dyTCPXJPsgkr+whVU/cSqTfEoUx+y8mc/QUuwjEWW9hTmXq9+3DDgwmRTx9CgQ8XhllaLuKcTlw7OOPKsNimto8EhH7raHvx6BQqQHISO1gPesdiC+V+3dklsS3ZlrWKwjdt9yBlR47PYQ85wn/no9TiHkQgTDZTAtNJmBqEpcsfjaDyJ73ogE6qr78vrC7z9o0/GqxCIOIXm3wDHc1b/KiNbt0sZKQ9UmST9a23wreMnfxhrqIijRFGXpVS5rIWDCFfL2b07x8Uti8abx7vOwJcD8wHs4ddkg8NwrRZ3mMC0Y/bSo6D4hMSA5uxb6SKIwosvzgRzLyuRe72II/YEvohiB8YpvkDEHXLoOJBGNT9RXaDHB1ozKVxERp4s8Q1YTWKmzel2zWeEODf2/RuT25XzLDqCCngoKKa3Msj9mFhfWxktGqsop7E+MBdVxdK6wBjziZM3yikGsuTHxDCFCYG5I7Vyc5783n9o2Z7dK1fgDy0YCkekdtI1JBXYgdKKe1/+6V3yNNhoQNSZ5RJ/5e6gFswi2FtyuL4jebTJ1cV5x0oJ2b2mJnL4cclDR0ppSuFsDKwvXCWe7EoeCPMUlx9JpWnncjFrN9OInnAIGjjryBEaSmXqg0DorDPlufiKRtofikV6Fx95eDMBl+9Hv2/1Xq9oGuLDiJ3+gfQ00Ie2YOtlyDk+/vy3Q++yEh/jyR5nAshShQ8Tf4hcJmyHpSu8m/umbQsOmzu1Gjue4CwatMDuC51NiciqQfrhVyhB3xT7hbCrU11BHgxhhPNtDVIEsdLkbeudvQpLz/CE1TLEUX/785UKGZhRRBLutRxe/XnbJRfbKqFlszqgOWFbD9M7dKM+1tgsUhPxTWQ/+6Ijcw1c8iQGOFOoyq3X8lHcugRLhj6G52WiyrksWl0doASlqYmAYv27rxf3kA8AtnfKEYBK5WxfHgA3pF5zjtWdYNHOaA/6SxDux9NBZE7F0rfmzxU0P9Qa7a+H6hSyLje3M+WbBNvKnrAvlYJIJ0rlAsZsaB5zSarODsN7zvsLCxkPHcKgKzdYUmG7ZJW8eTIIBVeHiw26LiS5rC+TtuDy44pbljcmOtY18QSVNCkRHx1dOS76BaWO5Gr61LZGeQ9UUlRZ2J7q75c3XlLgbQe1it65mEVjzZ+0+xivCYwtl7RJ4puhS5km3BcO09OI/buiuO1O3/YcP2k/0720WSGtwoJQtKXGc/6ozuqzXx+BxoVkJGV3U2cxeMxshY8fgBt31xju4ZjIdaoMxLynjS2BsYXWepFC0qxCUNjVK69DiqfSUvDmkuWe+n0Q4ErHMN+JgwlR/C3m8oUgzOsUVBXZUx4aFeyzCvwlQaLhfSz3OC8Xq9zr7nv0l8HITBcwQddNZd/hsQaJKRIka32gVYZOsjJj/GWLRIj7Sp17YKXylo09tS0YFPjVRLLUfwUIiofIBNsA6UB7AR8T2xwpMxrNn1LaL+/INGtlNC3fsGtOyZUmelVEH8yeBgYVXq2Q7gHKKPPz3F4rER/WXGBZhTA4D362NNVqI9C0b6aBHIsXFJ5lYg9dx/czykhzW3KZeFqptDJNXcZ6sU5S0zepAf/c1gNEP+EY2RPDax8Djw0EiXnmnFlCKyiokL2J3frskazKwVJNXq3xC969mx2Wad4vA7Waded++UeyssPuZi+hFARKH/nLKUUb/aYfkp/h4sixi5qFKEMvaKJ3HDBJ5+YAYrDiQmj/iDkAVHcffjWdGXVs9HC0GkCXReRV24pTnazHGeDtYHrnp7yBo8YqmlffRAC3pSXc0JuB5pzx7C+bHPTl+hiDYdhhdEOT1KAccMxeoIV6Bz7vE0zYPlyvMH3TnRFL6AK3/CMYOt940xPZFhUCpUGGal5FYnOk6xziR80ck+Amo0jY1fXBbbg2f41IblqnuOlZ9J1E6G+id83zm1bG9PeOeW3dXisZmaCqsvcOXOEM2KrmouU3uG1vTtVESDqxRP6npmu96/VkRyFcG0uAG/AtNbMtyBGnBk1ditLBfrpmwghUzZqkjd5RwwtFZ/0dxJ0qpZodjc4REhZpoaTiNC7B5vFwI5X58XoSCK3HjBagDAygOgTCLkvW5LBGq+R65j7yK3I8uA4xlGKuM6e7CVQwGorPxtV4xq6+GvcnSw0IRxvlgl2MKMjcD5XqfKuznC4meVHH8O7RXIhSrek7LeEl2RuvTbknQBj0jS6jC5o6JgzyDDNlbuCLCikWUyA10JSO0IynDtBgi+6KOaB32W6mmaWhZ4KnwbQ4+VoqMGfGLwMvTvrR/i0arp382UAOGV3M2K+PLSmd6gcwiIW8hgDxWzBlxCOTqnsvhaVLZ+TRNIMd+gavUmbgF6HhbdpatAKf/2OFSaZfzal3s9RPezi2nbOg8Pf1Wx81kqQB0o3YM9ERHP9SbHsaFHTCIN4g3WxXPLGLDYmqLFjxPDtrbfvBEflWyiaYiLf77DOUdaNUDVm4X4bAsVLMnhw/PDP1h1UGsRjXrrBPkpmT6LhMia44bHZVn6r+FFXLphrIwODJ+seGqZXkdfJ8AS3H3ZyFaBiwRpIV+ZQngmTXM9arZz7u+XyMwbqSR5Xu3NnWIZWCklaXxCEc993Tl9dl4wJetk1I7JpyKgg9PBDpfqsR8XlVV30d1oz1hU7SDf8x6DlNqn+3cMGuDere/AjitqwoTJS4FhV+wj4ldoHbW7jgdh++UyAvVMMVS6uqq9UUwTgDEMooC1OzEHFZNfX3RX92tIG2XQ33/Yazzn3SilC7iCovlSyc6obivMgmQnblKeIUi4ldsbpeskW8t0sj9EuxP6SiBKDwb7T0fj32Z+M70DMn9Pzj40u9CjosiOavFCbwiT86g/sYOoKKgvTVVKB5+bdqA12dgPSNJpHEIiXHXCtBzsdSk/K55P2yNsadePFd8/sPdTw6wJLTjwicDQH8xtklwpGgS9SnZUZbwyEClGpGHYDRB+Tl6w5oLnvz1jCMlkjDiwivoWEwqb7Q87AchfjM3Z4TNzgcbYf6T7nimGil7LwGLd+SlbFf0ng+vRE7yf2/ss25BJhYTadDCvVp6YeGoSrK2Y9mQBwqeXJvKPLjzHG7wDSLkxuiqjUUPOP25WmTd//aup5GfJchS17C4xoJNaWEQSXnDTFNyPWQtAWWR3bIW8/fkpSh8AL07UMfV+4xXuehncUYSjUZgWVSNpVYW0pAc5qxhJnUBetBuBQFOJeNSnsIwMq5b/yeMgxmXVHhFyTLILsSocJlid0t+ZVMqxLmuXWG64sJC8L8p47BdpUep1rdAwHcvJrT9DzX8w3SPfAvKNGWo5/V15wFrEjQsBx+QaBvW0ie73uZOAF05vun3e4ng1/nFFA3GoINFkYu1+RgRJw0gGqeY1OFXnQpRDjntF+3b3io3KvFazD3oy6kyc1Cjm7in//suIZjikJ8mWXLxGjcxcVWwkI12M36hL2vUmOokSzRBT891PFZo1xRwmRRqUkH1AER/oy0qy2hy4Kb5TvTUKPalMigmowOfhUo7bkHAGVxwI39Zk8KggQE0COsqMtpi5uyTPGgo1YptBs4YWYEwZD5ZJnFzfp3O1uEgsiyJ0+u930XH0hcugqVK2KyCxpzuUi6jwPNNZ1HXYjjkXQanhtfWG530msTjEgwL3KARz/5Gnq2sThfTprM9PlaxPqrRSDnAgaSzFoph3R98iITEIv5C0CRrMHAh03cHXI+0YPHIRbW/0iqNI1FvHZD94cjyLmRlPk+PPwjsjsdvDlzBaM81WqZffdbEN22WzWOzV1Ii+U4/amha7pta3t9pD+w4qGyd5UxBwKOB3xQYHEXpeciO3LVSRy/ok/6k05hCoXBRFrkIfnyNCKYOjF4xLKFPMEEPOg/a0AlH70eUmeCu95LccOhIcpW2zvAgSLavkR79aLsrK4xD6Ihk0V5os8W71RHUZnvkgZ/vPYJMyyUFm8u3XR48lG5rC7xMRoyvD08w46OrFaUfd8DykGeRMTPbrFIwQlSMjICAAPz76Y1dk/7+fa3s9zLFkbvUa75koZPu6+ZlCNJwbuAqc5LRG9qsIFma36gyS1Pc/SJOfrqO+j4GfHIFKfwnMXKAxn3g20hTLYYzitMtCCXa6ozc6tURip7dC6rjlglVEn3ps/zn6INLQxRm/CrVb2RDyvdqFdQ5j6iicCN5JkVYhbQVPJNI2f2mTyAvtvWscW6yzZhtxbxVQsSsKVtj4KH1SGmwN7/iy6Kq4JQ7cBCgk/AgZwgd/v0sS1UYcOQHd1nuzdYecxD3Ylha/b9toIITcLjR5/CVFgO9oG7078sot/a7JaxpnyaNjnzZWZGu/095vifXUt1ETCSASZaDw3VSYHmcP8wVN9ewyuZKHLZc1VlCSqW2D6K75t9ke1kYji+ys1+CCxo8zs9t7D48doy+9HzMR7Nk9/n3jB4OusfmOYUwlCRo8c6smUNTM9ppyV8eXt9tF4VYKGDC+AAofVMY4WylhVNABXruBpLhxfBvEktXT4ZRZeOfuQkP0KZzex2WPeRHD2ZXnDOrN0yh9ZkTZ4gd9fUJloy2/S3HekyHjyimS2tQmAAb1pWNP2d/7FuFWqMcqGA1QU/PfGvVn9i4QOqhbiGC993y+BZNuRq873V4iMaNJwWgQaORVj4DPOFFsYcmZy2teE6ErZ4y+GltEmShjwmMxdMFeZWTqmix7n07SohdYfFVUF9no8s8i34r7X+XViUMBWdXRL0QH6neKPqJ8TEyIcpZ9JUxNuwTmcs01PvGDfjPe8gkxeQD/mflcjcBb53j+w3rI7371bjPMDqlQVC/zLu7h7XEtT6FQShhG/xai57BqZYj/f7oquuk8KAlsKspGS3idYIE4s7OmbtMIMPb+GKnUpLym93rpQSgyDPOYKNY8JIoOtbHhJJhgj8EMIyqyuMbfGyJp7Es6hvDc4L7c6tKWTtu4FBXJk4wbmz8LQPxu7xhsPxmyBGAFpgyi3grkqs200HwX7qP0VawwU1MmL4yGBp8F65/PILxr5r9bW9OvZdEvC/enJLkL7KxzfYuEN3gE6ep3idfVbK1GJlSCAw6y1J+hnWHB/zL/1i1fEUEDjUaIfjkV8TKv0O5eubJufKummEJfkcSkPMix413I1kA0TA2ZF4QxmEOU6eXGjw44i5WjUDrRjBc3cGBJ9G9d7uNyNxfwV0bVdkyu0O08+ZCKZ1HBILBOOHQrVeI0m21alaZfNKsN+WhaLncDjeVHFf7QPYJoFXunUTwcsnA7MYrYq4NYE7Vr8Y5Nu8qWUXcu1xmSZaly1o2XMSickXzWtwBDZgSRBtccxOxeZKznSFzTEcs5cvz9pdwuSq7wg+WxBg72X0TWrQ7gQKE4UZKxwdZkgpJ9ViIahOqYCE2J2MrSt2r6GPikKaUq5kPqabxIZPDlUfPPVgkCzRo4njrfj+2SlYfO4DcKGzs3Yt0xtzlb4CYb/ylN1ExUUv0ZTrGrKT8cvo7hHYeYKn0lea37BftnoN6jxwNXt9+XJulE504rL1j34rLzNfrJI+feuQaNyGJcMMiYu2zFKDF8JRcW4PxHmm1nhO4uryhdJHTv8OB5MuSxUk3/qexnIHaMk6zUhCp3OTZn+iTHw25PPPWrGw7kl3aCG3hvxljLnCWc0it7453rMIWlKOu+9dL3ah2j0paxnF0D7xrgXttb2nI40nslwqAw8OJUBS4uTX27Vgig4SEmGpvYii4AA/zk5NVjXp32nhy/5pEtPJWqO6VRsuPrSyyEnCieeCeksKRmePYP2IHqJqBMGFcwfsA0rw9j/UCp704byiStjY1Gi70UL+w7Jn5ZdjwwBijUwzavbdeImHAI4/zliK/2cgAd2v1tv3uzmkCdfYBZGI8klQtO1Bp2uss7Pbovr+JpuPMMJRdb2S9Dcf+utQO5vCvpYh0Kd8znCF3FRfQucAtsg/X0loDe4HdHhFHvZLxfrQ3pybaYSiI2JfIAgxf7mh0vRKW3O0mOsL++fcw2wg+G13w0D4zvM3sY9Ky7jE3GfkmspqQ4MHAUGuAPxxBHpxZUXuK0QatIoAeZxJ4SFj0OzvKuE136kXlHWIHOsPzY1qHJ5qIM0adGtmPLQblwtpwUF3+N2hG5nDFMPo+sSAH9Rlhy61lLLWhnIb+H/MAJm2t0Ftx9xEa3qI0YTi/I6a8P1Ya+ogol3bRbO+Zyyd/Yi4rW+uB+h2krlPZ9bhF2iX1iUsUMLfn+EaJzGMciqY9iOIWcdcBiW0p84p43rX0saQtJ8RFH66bFioTNv3hueW9zzvezW0WvN9A3dNHFpBG51UNSSM8N5l2Hd9bluClHezfSg1dTOPedZPVD0YAUhP7MTld89RJUnK90d1uD2+l4JVN+r1mPjZO0W1dPI9m0Q5TDxCjFyjNLnfXF0oyWAfYN9pr1TL+boK7RSCAZgT0REc9tsOhPtw6mjo0mdxruWWrSlEbjQZvx44b99kQeIqiJUtAwl4fDjNZOfBwB63ZcY1wvp8iiP7kmvmylR71BnQgtz1D/eu0XY4sL8tLeNktpgWT2wuNmcihjP8WNry5HcLQ4mQyxUJGLiQIog7lTyOUckaJ704bLwZM5WYf9U2jWeVmM8J8a1R6S6WGFCGo1qy1XH/h2SgZPVVLGrBGYZ++lKAmi3SkfZWn6cBvfBNWYD+ozA18KwR381CP0b/e2uoZusHRupjJ1MkGYJfBljUi+2DrEYOeL4yp0cS4fuzMsFIxQ1XuFamkF77MawmCAAMvBmRB3X7UhGShqnoStgAEheRrNGiOCpMxngIAOavudh2dY25fCLZ3GfgvVeqok47HCV9YS6zgMdts1fgYn1ATLRBq6x4VORn7jh2yLkGJtD3oPAGpwJAKI30wRe9RZjzYQVKkZrAzw4jx6+GyIgm9z8XGBa+EBgaDjsdSuEP4Ao5WJx0Ili/sQae/Y0Xd18jpp5EDLcruin0WoWqDomvlW4dLYjoWB2z4Y+lqSL7oT0G5K6jC884L7YSCPjye9XDgcuG+kzTVeV/yXMwP1QO6WHmhF9N6m2w2sMovyRXwd3H/6fKJNsgLPrzIgmNIHWaNUxEMm8PRuqpo0VpcBUUtdguxTzILMJmoeWW0jcBn/tDMwkPYl5PvdOLay0bFwWIHenX+uItXHD/0+1f00IiHkSy0WmQKKIq7QdHgUGcfypHgCiICTt4XjrQfUhGtkKzg4D1e64tpX1NDlPSTWQgxkaEG//zws4D87lKAsBu1TdpBvChdxoyen/dirwSa8t4dIqSm7w4PX9bRo/c0dHaEDrwySXwF7FtjauYMUgTpUQl9VsWse6RG7C53Cr1wcJRRqX/6x94XsuT8kFcV/FrfO5UsEOmRb2p88qfZCRxWh/Rj6BzVDIkITsEO1zicP5uJyQEhQ2H9saiNsh7JM36716gxFueN7ImQDofXxC9HUEZZ6DNg3PzPG0mWIGhkjwLGwh0dsUZ8YxLu46dnNV8Kpxdz/gVfZLsHHHDxcp01p1+4Ud4tJ+hGB7/1X8bf5PRTbLN9poA/1+wRBLFz4jKqsPBKrSUfzx0s2SdaWOrI6z5rjRkSZZ5jeT+NrW7qreudTmDw29flSYxqsh40z/U751OxqFzPtXtawDccLLyS4j18rVdVVc1/yuicvRoAb/ps6TUX9QcnKgherVv8Mxt5dmPk+v6Xw9OE7IKMj9MuFehXmUCuoewaRMTY3VDRdszIvpa71Z9H5gHkjz+fHH4vhMS+Ceg4l9qtnjxcAOpEL9MD2ek1kpcuqqMYkzW7z7X+EG0BaUSKsmdJtToeXs+gSdawn6n5/j7XZkVMcBVvZ61a8STLvW9yFKVutztGQv7x97mJGtXyCLGCEX/vhBheA8ACK6oAYsW8aczC2PuJqw1uA4NnZ2XeaI5YCerchIqIE1FmV7TX0E3aqQieNRG9zRS8WRTVEMpSlFpwghmp/N34T5p41OVU+BtB2iFq2n9LTOiz6+uwCseaFpeYRujIE3ubvjEp7AylePKRktkG44UqBs6Io7ks0NVcvkqBoaUYBBLdB1FJ1zh5XeqOSRLUXGnItQoWC4mvtBmIT2W1A37Y6haG5Bn1HtEiOxLKsjbh11LC46O/MyxSMOHLz5aPZ93O4/QMunazLsu30O1F6a08CaNLnnohL+NSHU9uzSCrDqBth05wvBmeOylnlsy4mWWnIZ5wi4fkWdjNOcrVQAUsn5G2OzGrmqOVuLcRtjCf2q9UvwyXra1/5HvK1O9xqx6U6JFBiH0gFRANYvNE8nVW08cH+2Sr0Zsz0rUKh0XWzP3k58keCSUpBLiSC+QnqTdXOkyREwbrhnunbbkAyHJlvE7nKC/3wMDOgJXl93Q1rHB5bgP6zt1Yi2zHQcsa7vZAj0Pa8vtJVV+OQpIzOoGA2akMUBWFIcqtML10erwdWHddbSPl9nExGV3uiO1oOiLUXaDbycm4y8ed3sfA/HHzIwLRPsvbl0FOcQPXSAPnbnGc0kUe9orXm1pWmwhmfg7BABO3a+k=
`pragma protect end_data_block
`pragma protect digest_block
d3b4c725c9005bcf5fd3ec2c74467efc47ae836b46807fe6f00512d8db160a6b
`pragma protect end_digest_block
`pragma protect end_protected
