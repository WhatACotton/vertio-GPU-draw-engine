`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 14996)
`pragma protect data_block
SkKbCB1Ar0UG2JDGO/xMIMe6UvoBP9qj7k0ujWKNXckln1IFhElcxpCz3XnNHXWCSif9/m/nkOGCxqAkzV+uH2046RTll1RfuosH8LdOQ/Yj6oYFZWx/vysHFtqM+varXbq13G+v+CClQE8GdtAm3VAV0HjDxBpEr5bg8Va4t6CoNIXdzOe2A6Vi3uiYOD/nEl9NxdFECQS0Tz+UeOFVjkvS+GOX3+CafZ+lbisHkE1t1LqGQ8NVR5hSVNkl918wVZdCtq2wLduVHR6Pli+HqsqDE6Xwhw7M7pULnqKeyPRmOR8ve6v9m66R/cUrNz2kgPLh0Nk3zl/lPPsGBqvzeW4xhSbA9iGg7baT3QRRwYyTzTIYOgxCvnTFhBQ4p+frPyt9T7jyBoiXdmP/9KovQX4eDhmrD0lITquEZXSMoAWZbiutfuehXa4e0w2Cl1APg5F9dQDLyUazstBMbcdg/O1MrPpSNebz29fa87qKV6CD9g1kTrTGvsUTY80Xpa2Kn1MNQBJpk7eed/zvOkuJ7BBi077gHN1IA5rdAs/wOoKpTS3ZkhqHgPXT02dW4oOBbTkYL0RQMECwFxiCDD8JJCFBaNmLorjO9YPfylvVIa80g5GwXqS8Fu5qUeI+fJM3T0WrtQwT2wjnbzVaXzHkHkTfH+5CzzbxHe7AKEJP5CTg+IoGuqFaxSAykFvA3xHvFQ5ADa6L4Snf02gC+hM6j8gulFdGcXDMrY1jZcIXnvMYjj55iWNo9SrRF1bxQ88bofK2nWWTyTN6i/YSQ2q1f9AFHhK8as9456CaSlCzgECXA3sSZvUyHag4fBJmOm/ukHeyRA6ueF7w6q0UZzxzsz+XKX5f+nYv+FAB+kuDYCu18WReZoXjhQJTZ7ZTUppDqNbgafrbjTK7NB+mTSbZDWbvq159/ErirItJ5lOX7myMAKJzssxL3Pmw+WIPbTw0r4/x6OrgYcgSwmWNgGLB8OSBjW6Nny6J597qnZvc/x3Hg46N5aekttTtD3PPBN7rgU1EQBboMmOlHLbYr1eBAianQBgusbtqFyunN+O8gtBdEcjR4+/UDyepfXdUDA5OR5rIL9mpWTE8HONR5wf93N1mwF1PdWHFBb4jtDH1iMEc/b5kvdtSjUE0ixCwEtayGCE5c1lt/PeZ4RuBlvuWtvSeWELKI25ArfPod8UQPKfFM6FYRypQESDyaY78x4h2Ia6BE+jId4tIZm2QBoQ1KadIQ1R3xIR7QmzePUaMLAexm5ZUuDTdNaeiZv28D3crNUHNNiL9jtOR0yWphdZsfZLF1pkzFWTefMA+Q71EgRNR7CDVMjFsvng85+rMwyzJnaWJP1Cx6zqhG/15mNxHhoUdm/+D5oiM6OqxDKziUKPmI4EZh+BYkSavgt7QotK+GZSL7Ek4LEBU8RPVenoqsvS/HGcu+KF828ElLpJu+AapylriYSrjmnKZLzJzxrJ8LRxW4WlWfjGt87FK179seN1s7wENAZxlrUiiVLqV6oMu8S7Eeu6PQqGMlg19zOJPALanke7XhKudOQiHZ47wfVUAKNnlzfc7SpR0HU8+FSPm0BgFJ5757o8XOxuhapEAA8GPs+51iqDavswc0v0Kte23IUuggPlzf3H4Bymkzo/DNIPhbz78brhj/0WPoLFnRIW1952xY2iv3cegkOE+r//kPQH2MpHfIZxOx8a/w6Z7CKCs1rlLMGXlBq+wI5EvBEb1kfY1CeVLsAUNFUuiGANMYETfyCUdM9/zqJ2Vm+puH/bDf6G+kHfdeGbALSV4dyiuB9zzTAPn6uPNcwj871xYCZeAoiGFvyPezFwKFx5wcAv1nGakqZKccKo6Wzu3A50yZrWsV6y+6MSQCIFRdfcobFsc+amxsl4gPTtirNkWdUnj1jvKaibOlkcr8XNdn55Qd76HZfuym3FBzZ4ibRV/0vNERn1af+v2iRbd0F0HWcMbPs5E9BG/Wm/TkgPEeQKynOAcMVeSFrC1QRipZpgH3oplqCmQgATgFNjAbevYMDL/elRZb2Qg0oC6T28nbnDsWB5V1nhYMmNL5hV0+41b2TXbBiilLQB5OeE4U26+m2LhlPHBcfv7Y3Z0hREPvx1EBC3dGzBQceHl2K4aJ8AMMPoaTGLRJU09Wr0o6AlqjjWV33gU0UumumCDTsgchVT9NhYTtf1OgcKDtIZby8/PihDXKibaSOQi6THHmuoEdkky696UpieLkc+fP1d0IEPsFlpTll5coiFgxlgf8W8jeIGX72Ze9pekpqLrvpT4kzbZ/WsMtMYinSMwhGPvCDSu3CB9gj5jji2RCO/T+GmNvEgMQ04mLPWi1O8Zxt05r4tjmB2CCvVrP3as8VyDSPOxfJzbaLu5zQMY75zKKVeA619UqBiO8u4tiGlx/TvZwMkOGunHGcsMUainheK2hy5hG2G495VXVpArQDiHioJDKEfzs2vraEVSMzlk3ELzTvZZjoDpECU23ILlqytEMnLcEJv3oE2soyOLzW2Cgb0PNOwCcn1FVcvCmczYP+CQo0YeBL7jQOV8Bena+WZj8KyHNBqY5iqysCl1kFsqjNPTiX9jJCIE44wE8tb05frabUTsQnkc0hzrFPpLQmCE8PT5P/wa9yWyyroVdonKMBegKMp8MQwhgjxwneo7TzhDYBoc6LsV+6xrN087XBwPDIVC1UlQK3wi5u6gr2Hy8wpD7QMgU1UhRh5E8kI342qtP9fHlIiEZun7rGPAD7cjbofLyLTNn0bdncMcXZCA5LI8MSz0gorI6KhjFgIpstV5WcBgQrP5h5RwhJd1vXCmctTR7IK+ndrGd/YiMMMJ/FP76MdWMROOj+HJ4eF14e8OwlP0sQR1RZN+dxvgIHQcY8eS0xCMFGE5j++cc++VPfLm9zTIF02nIN6As+dQkksNWTT5q+IgGYrhi6sG8STY+7nUiP3bU0tUnuVA1d0cCtkuz3I5xeas34Q0mr7d7YjMBAhvJ+3JMZUxp1G4yqV6IFGrGPs/xvwx0RrPB5gabHsiZiOZqEqtO4wRZrmU92LBM/hkb9AYK+Rhup51TGS1pjYILQ5OhRQVuxsq5JIYz4OoAsAWjeDaLv5i/HUFSkmGm+8WHmnuQvbJXFVEgdS4YP2baCGzOKW3NFyEvAu8WkERHOUxyJEUqlZL+6eN7zClMi/uy5KES2hVwsmgVqXpalV8wQJR4EsEx/ayxeU3LofirgT4sd5oFaUC0V1/ywjXYVKrrTNShTYkne3q4P8TgtZVIU7y+GKnmFmRMyhRrMr1ljj4M9oLNrTnOyZCP5Q6vQhjdLuhM+obRJs7kJqHmV15cqWnVa8pRMuXwKslZDjuqFP/CRF97gZ4ABxrS+mQdcrvYqdASHCx47vEWk2eb12T4e4a17jXWzJaEWKreWVtb9bckMaRIsm0HLxkD+nwNLpMoBdOXh7ss/L25ihH9rlGlVoUMi1k7eTnhMTiBNUPgtgoex6DSF7jzcNrKL8fqlm0gRcI3MjbeLzRUGI1sFhG4Z2/qoqWbTt84Bw58OIBsmaYEDyytq11FA1dKNDlIoYl1wO311/M9aQp2ergIHJ7hJhTwjw++jmA9mOLmtpC/8LMBDhnSX3NV+mOVEVHEoGUkVSvNGyfk9Mph409CEftDzuGFmhmG3bA45u4K5/qd74QbuOfggF6zb6vVe89rVMMus26NiK7lpvipItTZAn2FshzUJ2cHQERHnyHOCVRdrighswdcsm2JFOdxo4xJ3pTL9gp/sS1uIH4kffSTTvhbtd/mquDEo5tNJz5VI/2DTfzOHPtb5Fz66+OapdN/JxgqSnn87cGxP6nWDw5wqvva0j0HwIYdMyUl8BI0et8Gb1Pgo5C+InwF90F4/YUQdX25BWnklcMCURKun9e2mh44q/XOwpnfUNI3UdbyOWzMQvbIICoEgxiG9khYLgRWofW+7ZzzFUCAMSBeXKhCpT2prmRGvbaaQaKFYvK1sEkmtZTRwO9Qrencnts9GwUxzp/CwMZWhRSDDsxArdmM8Rvhsek0e8fOPgWpx17/BCYeTaUDhpf6s/cT/m5Jk2upbdx7x2aGJWRE02K6q47Z3dkiz/wsLZJraHuPnP0erm6yU365Gyp/fLrrhR8RNaSlLN7/GupBlggq+S7Ro35znY92lN6fbI2UiojIGSUTXevc1WZ1/1qurYTWCLvzg1eIM/QKkJi2dNdmjIIZyL8vt/Zfn8eSr3/2j/uPJfO0srOx6Bzdv+kWDEE/cu+yt4aZ2WzZVaCoC/lseMuhYWsnMrDqJgegFs4LsTpJ3zZoQuTPNwJvd6SJRKWqB49X1QvQoeQIZR4olyptweZ/zVxoo7zQu4f1yAhmVHBuzIa/JaqCXrWzDPQVk/bsYTUOXck59YbdtQVnwyjSjgibOHOygGXOv511dFtl6ew321nDqe+cjQCezll2S99iAaZiHBUb6vMPXleLoags9ExO/zeAhXo4PGQocGgFUlCiNAQdfZuXGDS2x50UekxcvhLwZD6a1ugFWg8LsoX22yzbNRzW3HTDn2oEoCoPeMihjRXjPXtRRffSC1g50SEmsv7in1U3VSTrHDWugAtMJN9V3q3+6kixoAadLcXjml0VepgzKucjUzbRj886JA50H4mQYi5e1sAmLm4GnwYE1BIxl6x8V6nr1IpsZkNM+e8JKvz8lgXiaBZLZLKrjCmUAUl8KlkcLhiZo3upMnwKztk6wJGRbyYGez1JTzIkb17x3V/+aX8DbFv9AQ7jN9WY0pgMXXXIJIaMGVt0cTiazQNmflPmCFGvxTxH6Wl39myITYOKsjtoFqqRfbriTjbU1x1gtGlO6f+Xq1aFtvrVKhYyBvcIPq7Jsrq8OnvmNpGnNtDEvidrOIGygwU8dJ9S/CqJbWklHyJdJBsqPTLE+cvSuExSl8WEiel7eZkCuBaSOemuLh5vDI+ovXgFBO1FwTNLmHFN8oykqo6BobzvUJgZGgcR5z5CzMslKqPcZ7zzjHMNfsv68avMKN/RNKa0Kd5Jv38OqO6s/RPhfvEMxdtZDzNiz1G2Q1/xHtAHlriOr5orC/dF0HdvhiFQt9ChVoqA7MZ1o1xwhdZ+v2dTnyei3xqFUeCouh4qvz+GiJUFPdyNhlc94aCUka7HjP/otH1faHM5XpZ9gBeNe/Ae35ba/QPLXkOyUYkp97xm105eyb7O5M+02CJZIY93RfOYTHX46NAyO88Wj6PYQt8N6j9AFKqCWXefuTpVE6EG3isrIlJk2Z3WmgsJlDjucMoRDQaWLkR0u3fFBcRgkKZvG/jgCnYxa075XTAsDl4+vXiPbF88uuRQk6dcUICqCuK/LK5e1AdDLEUfR/EoL8WjQme7xBf8e4cRQ+1tOc5SwJ+WqpjzZiNWc0KLhJD11RD4TYPWr+CuO2ziAlGpphFSKky3R5Ok0jQDe8sDfCVgzdD21dAVYPExpEgM1qVv8B6m1mvHxY6dxZfFbGtZSTdMiPO9EZdyaVWae7xo5sQwu5enwrRjr4p5AIP7JGQhDBqhmhxyPWvwwM1dkN4mqrbJkvd7P21380O19psta5mb2tQ99qHfg9Inb5tILHC0u0MsR6WPhNBU8pqtAw1KGFX8mDEj/PjjJyTuPKildFRbzzqN9/y5FP+bzcpZ0mnNWQGwzXA270tLMi/S5FTfp/MXC4Q8MM5dMxYbsqyDdP6fHGKLtv6NyssNacawjqrK7vlVY5kyMKr/z7r96rhh7iF50i/EaPuv2OIkkRbMU3jpYlV1rFGlKEWtqsIUAzvbzaktRU/tAKBzMiTCVII1QX2k+gaCJuewNTDMuWevfvlnMP46GAUuOOBCArG7/JyiDDBbQiVm+L2l3Mtcydz2hAhw3rML2jlUpOyUYtiB2aRXkzKsgJMSBm2qv16bGkfpyeTPI8B+b28rurtfiuhW9sXxBZCRqFqaRcsmOlknSh6ZNPtez/rG/kbLcQRlL126au1qfx1OXf4/ZL6X6+QJLrpkn85EiZ617k/q+ee7e0MFa457Ni5+fNPI2hxDX2s4/wY15qaneeslR2HbAQqe/V/03M8IMTklUBu6qu4nq4zCTtd7uf/nQUrKsK2oyx6OMmRz6+rz5d/AbkJoqt99r6sGPEwWKlpUtTNizoNs4hrkYD9+HI8VBlCjQBGPgtWDe3IK6ZTsY8H3J/ChfeEeY9it/veQ6qZ16vAKY3w+JV8prWzlsOkBhRqGyhhgxfoJ0pQL/lSOsmQhScLldMZiN59bbd4t1uA3yyEwYb0mF5LeAfY1C6hx1dLE4195oBkeqjBzeI2WAUNzqZvvxT5ENkpKUn7e5U67F3Ll+wMaO20b7zI+Qa9t+ps714c863c4VAv3obQgfrAsXgkaZU8Jgum5WdBjnlDncLRfcYMH0RCKbq+QPZYsuBC00USFbD213qFQ2bB5ATX+UN8xBaArv829vqFRuvo+ImaRbpCskNhvTeWvLptWRAMtt2B1ikdlsJX5ajhMVD1osKVIxaRMXmvh3TTocD8ob26JLYAHE2OCNTqN5nh4ukFQKumAcpmTkCvUqOTQU47lKoELDb0lnLbljyv2DcDWf78R28gnMfO3lrCWJpEZd6Ri7aegpPPFCuGzniyojYvoNr8bKQQakGKR0aTVLvDRcpBZZ7dVdTinVH66M9WqpYr+ZPt4Q3FPEbgJ5kPG48/X6L2x9AcawAJmrVsytyTkMIhK8GgImMymmb1q7mD5BawKfz1W/Ljo5XXjEHoB+SMZlLxfzsE+LMjpzNCB7YO6ZqvAOKD2NB37ky3OStxE1pcBz9stYMZlryvzFxVJNfopoSTxEOj+EE4itqxoh57gke698P4U4r0waeAaVq5Yoxc0FELVBt4uMJSEH+5dPKHzgbAih3EFvthxAI0nQ3gB7iDPD9QYidj8epiBEYdjYiKp9vrVx4jfDIlr0avFoglCxabbhJcch/FIwKgxAuwkY/bj4CCkjU0C1wEWQxJBNfxYQjAUUuRjDI0eMdc5OjT4eeHpPZPQAZtiQBY025s8yUHJJ/217iN9QfZpCAkXgOwrxowmUV/9BIxqhgYdVjG0xdGFOzDurRMYQv95aI90XCRXvDsfZJubvDWI0ojPxOowhpXLOmuRqhYY8ppl845Ci3tEH+Hbn11WzuQyq3CneQMvamP2ny+H3Jzj38mrS18B8l0yLxBm2SVsXBbwITEP8lNJMxQ1fpDukkupcqPTyyidBJrkwHQwVje3Ctnx1t1/B+IsZhUPVuVNcR6XrCLEeD1L0gQ2b6gZoM9d5W7+KN3zs8IGOjiathGq6U3vJLP5J1bBcN9rhyH1CZWOQQkk2sCM+u5dFH1hpFq7kr2YDSwzuC4G4hv8nCEMRqRwN1HXe7WY2fZ6AEJvIabyP24+nebMEfZv0FoNVtGkp1RqFReg/almoNgnX/zusQ0MctfvkZeVmzikAk+iiiy9pHF+bX5S701Lv3YBHPoT3grbBf1uVBIFGSdSwKfF+tHyfd7nyVyPK03964qXioxsmqeQPWtVp6O9D+JcY0kUQin2Os2bgX25bU36dNCKCuI8HY4GeerP6BWn4fzeMxiTonE3sFHacorC4rKiL22RxgNP3jkAwasMNHAU33+43gQoW5PwQKTeTACVykhjUOn277yyc9Gty4adrfXXaGDGvimtH4/BfHmhbDqKBZbSAlyKr0q9Lu5NX77YAOPy1HMdLLatSlepCVWhBJx1ljExy2uescYS/N1EvV+QD+K2bop8PHZHwQqceQ0Pwy/d/UtVyEUd5BB2lUl8xkn/sWObSY9RU3CSWpfUlUdZ/oajO9ynXDz5flbb1YUUITbSizNfzNbrcvbmx2asp9ipURilFtWIj6WkxvXxgrzUExb/GsktrekOhRlkyQ9EkE/OrvKoHBBJH2w3/ea9+BCPC5/4pcAMJhbM+qgHlzvqJaObWUFopzF+49Eb9Oh8vdleQCs5AFJtBGJa3AUP8tcfPbryPVSvJZU7uve3XuFL+9CnHH7Z3iY/IQaiTk+bsBm/mpX7T6jhi/t0lcToLz4ep3glvIE2n9+5RLEbIthitvz5mqnRh+5G0JQpiHWF+udZlP3PRDA/FMDOKcw/guVO5EQDvV8Opmr1dUak2sBznCuo+vYWamnWCKy41060pkitUM8wJ5wOMhvjTAVpGro2ZagWV+aYKkJCjtWHy2iz+4p6Z+k1Iz9zmo83rhKH3zDymR63tDkqE+asckivJoOs3fXtqDc60/i9UcNG51u1JvqLS/+I+uL2XbG+Qrig9hTYp00q376LVQAn26y5R2c7jm+IduHn5D7GZpQGbLOeCtAO7pWCY6zkjLj6iT/KgwIQkvZ97m9ja1b8bOdnERBQngKjTq7bd6jw4Wvt8kmv7HvGyAHFszZLOVtXl1+IJm+Bb5T8JA3tJ9gsh3zJzLCA+kH02LIaxCfa/zxt3MFxo/wVQS4CM/ThBWJHlyK+2XxKgGGiUPzOyIdTl57rHClRA8NwItS9WvtWdTcmlkXa9MS4YMTAQM/0XAlid39QA7GyFdpksxX53JSCwsgriV9K/1tKrdBAFAjHafCNprJzT7RMdUC3pBc02QJFBOe7r+ObJeIltzb9E6ThvZJLcKV6/GrGBu/ABOZRdbEKmMpqgXBKe8Khq3yhi27yWyY+whEiHJiY9o0FNphd90Ql8P/rmb2SSuID70ML6Fy2XUw52Y+c0hpqFcSsN8JrxUNUCSMqpTtaplSvsN+VV+jBR63v//EQdZ7knDPXpKJ+slXPI8ocDIUepQE1CPJ+96gmcY+JDsAeT/heiHUuiJegjps4ITH4NveiPe98jSDZhnqPF2IUmlZC5e+8E+ydHp61d439X7KNoExCyguZOyMW/dnBLTi3exZ1DKyS5JaYaxhdEEhTlP8jlSU6wmkPabIL77duZa6UzDh1YhRkjnINqRpbdvBcZTDfgbGwVAq2zmRu9JzAipvyyehNRpZqR5NImO0nHbKWOsrpdLnrPkiZSRc+JFgfBfkgq8/qvAfltagGa+pXdHOkdX4jErvKXGYyJxBUlwtMuFZF8V4p8kuBEX/M51ky3sodHL0uusi0dPZUgZlRXA2x73jV/OLRgWHR+1XAI9G4/kJ4Zvh+Q1d3Otpwt/R3ybu8qBK1FaaA8UBFAszRsqYWGH1PjJqZPrpYSKVfs44F2gl5vDjRrxmDGdtnfX7AyeMnQMe6ongdiTBkeThFxpbm8DQa1jht4uOZSkoCXtKKrjXcXdjUIiViPmSL1C8hDhYFc6m6LFOF+mlIlw/HtfjKtUYo6fkwtoUQKz8f+zCckv3ASMTcKSD9X90VQnqvzZCGXfq/UgZy7OnzRCCenahzA6QgxSIOBTj7tkacEW0nsmlfBVmmaG61jO0dQwWE57pqF/GwwPL1H2Hyy031yJJE9Gy3UWELYAbfoNBR/BWdAalq7kA22DrTRF/+tQo8QYJSNCYsyuNF1QeK0PnHInXpbV7sDozjCjjNfui2r6VAAxR5SlC+ZEYY1NqK8WJlStKTrBoHUfWmveuxsS4UjPtyAQWTM/m0KKfSllPrIByK1QVLtQkvOBhRCaWVJK/xSDjNzAGqJILczLeL1KPWLWc3rvr8ZY0ulGXgaO/ltPuECpGPar/biLEFE/0S1DMTB5zNnlpNVBe5t1QaoQKzGBYruV8Nfj40Ftclo+KFmrmPFcowClLJz/SuY42DBzi8d7ePx4jS0hSA982h4JClUxhMmcRHS1Smd/LuknTVWrkDeOBvwRECfaE2DbpQNY1pspgtPLQ7i0Mni9hA1IE8aDYDb2yHbLnCRRK87ghYLd6bNJjWyVvI0zOcAfIK2H2msML54gNwpZnc8uBQifZtY1HwsBubDNf9uxg4ARbKIfvwzRA/eADWzB1aIT03FZ+dVe0MlviwgW6MsVPHlMGnqmKXVCHidc40e/ocZ4ae2bcpukeo6XubjbDIE5jEGq2BBezAOoTBvaqjTb0yOwOAcvQrtbBgR2OX8sbSanVy5mq7DXduFLZop5ejhR8jpzLs9+ocSD2IZh8YVE82OST1UxDj9AZU0m6HorLes9GLXZqy8i8rP8h6NFGLUgoViLAqlY4gh8rdxv/ns8qpZldASuMb6lG8OjnF9HJAy7EDmLKcxcO3wOZ4XJ+t8hkMCHQXKglE701RhxrVAk4ev0WvLlA6HlZHMpoLsZR+dX35ItGDLowRx0xiv8lEUQmU2H/6qaEC/xLHGVc/8Rjoz6XrU7dZboAFoOS62TMk+WAmaeH1iyoDaRPT9wWRNLZ9HCRpPVMCwfYgoOLiYP9WpWjzzc0hvLvPHvJjKrwJ2xKSRq5avIKzfFXGzeZwsJIgGgFugWQBLYCLHfeub6LUgIjIXJOemRfBAgrPOVBR2/tShvdGzvsLB22vetDsFr3SRbJ7nA+Y14CX9WRbdfsDwqRJjsm61S5hMdjWTRLoXqwr1NEm+vS4pIB4GXczwhkDRTF5+sN4Lyh6dPh9RJnGdSGSstrZo1u5qtH6ywBTTMoGzNY6vhXOshciXvg/olnMIqmGLKscEyKumRgMpfhf0+3c7JypyxYGh7aIaJq5Z3vZkEqbplzdhZLKO0u+7GfdcrYcI+FiwN+9Z3mOQ81z0jTBQ/5xhzlh+AtUQUjzlQCcM82KSmTW2VyQgsNrxug/fChGJ5ZLuB7UuLI7AEQYQFvWIZOJ1e/vlq65IjKZXUNy1QlwarYiVqjZTZBI275AH6DgNaTeNAhgyEu66q9wHGbZqDj2qdz/TqmDKHPupm/Hg9yMCmCItWfUbAFRufOvppeqEygaiPnFONBwT2VQ1OppApQCWBMkFx3Uqsblb4cZMUpulbghgHEzTtPVYYvfFGnAaPlPH8mUSWzFSl9gwC9zO83O2CHMdz16cyEwoY73yQuC3iGBhV3GjnXfe5MLe/O+9r3rWH0C7T2F8edKQno2r/0kPKlCWOG/bgII/gibW4ckOws7dnKlTYl3UI9oHXrIslo0XtCQ6xRYPs28gt16QsTGOegYkfw6wZg4Vj8cEEKOwhj3X+M7nFCvcmDZch3eKT17TCk3DZvPepoGxbSCRzoNsZV/UTZhpdIbV+JW0bcWRNeZhmnfZl4ediqIO6EDDR3APbjHG0g4nHbG+pNLJ/w4wQV72CHYeTDD1FkMQqxeKIrim2/KALmNVUmWGYoOD4FlVZbTIpm0nwcZYaf0LZzPPnGsDdEu7THpc6k8OMD4DsmqO7TwaMq0bFniYNZQLaCNmiAMemz48pVDx80DtNfQQIfE4+4hpe1TXJludtfaKO+4nMm27Mh5ONyvTnEMuI5No1lE248OvSCmujO2hZkdrw/atoNNJqZETSl4KYJ6aGO15XYksw/PUF82j01X9z/e3envDRKhSi30eup/L97ouCZBF4R5f6NGnVUPcupKKDwoIoyjYJ+x0W7HsNRE5JoorAwlQvb74BJhwgVM0P+kuj41hEszo2OBSijQEwX9gyOuGgd4h+prgYPOQm0O5vFgEad9jr+r9G3CTFw4b+XNr+Uqwdn7o7/nPDGmauOMM5huyStVxlOX1uCrXOJtBbmq4Fu+gYqL0r1fyZAcsgynbNoCnv9mHDUP06o8jJVMZ41jIUb8X8eA1SRIHd9+HQ4Ww7hp7pbGGmz2ca8zeR59G+1Kmjx11TnwMKD2lhgJhiRRCB3kMibuVPQKIsqWCRLtmLrhaNoANLl5tfRAW7H4OjOOU4WApOcEzlKbVX6xBT+kIbh2rOErNWdBU98VHHjyiXpZ38tyhw9X5DwsgJMy6YQEHSYuVEdC30h5gFCW+0uneUhzhObvXrUw0u0AuF0sLfJ766bhjKs3LYtQXme7jBb9wIf3efudvFdByl1xduWCCZiMAKEFp2cq/x050ASgtDkrABYXk5gyLsyWF2nrwVYQ3vb8RAaxgNSWZWNsCqRNVeHWHk2K083TLUXA2bIYWZQI2Ft1yHGQv6BfWnmVlLjNiNvmMH5YmK3I09QUwHhV0itS8Z+7gJr3JiueS5gIO/GdF7/frtGOtMqR1xm6m8DjvKZOSgmcxPEn0GGoZnK9+/LODZMMw1nfFb8dJiKCScmmX4eHT5zr1dYdj29eSiU3JLvq0s5qY4Zk0t1fKWIEWP8eEWuvp1YTbVUhYOMerEoUXrjZ8o6gUTzj+Qwpfxn5dpwAD/wrkrsQT7HRzLkyAKNO0XpM+7gwsTTD2KrEglPWTwF+HDA3/VC0avLnBBQXUTVyNLz0ALCcL0cLI4VAjaN+PfcsRNPWDa2I9jQe2ThB9U6hzBRhD4yq/CA5LK0kDSahszdaEja/9+fgfb8s4ln5FlWvinJRoAXwKUm+V5jcYH+mcPCAWtRmQTXNEsM7xK3GwuMe717zDbpWo45UumsroCXyQkeG+yKBx/BpTmQdLyFOl8PVBTV2gdcATcq7qI3g0tM5Mw5sH2QYnXT/EUt2+ngRk4kB3hJa66zHyBcFoClpo+RZ3pS94aFxp/ai1RmEz3B626TzCeirvo8hlqv2lHpxnpim/GbdHiedd0+9UcXSSE3rTl+GNbWZ6vLJZcgfXskjY6tH61db5OeQ6hf7Gz3ta1Ih1B0xwazShw3nsXkxmC3gJAgTu/PrEkEfXrheTwKDEVY1OdRex5nW+NHa3GJOwyhoA+FcO96qKXpgsTxVEdbIlcu+93NmFTNMLWRnQXZMiUrHH9pW+C2+9LKjp/FdLj8mEpAqe4KJyxYzzRjuwkWlCfeCqKcMbwNTjAMtCje4F0HdbUqYj30kGdSXodCXQnZCmfhxKVy30DnfwwTpy1UMiA6R3O3lEuvR4DSTfOGulaowWE3sQwnn2kCf81D4m/icfzu0bNaaVHIhHmOgnZFKNJPKm3tYi1/CZnK1rWRRIrm1S1WOxvwGJJeMuhCRLooEjob16Ky2K58r/R1ij4WM460yGCVNwG4KnNOGCE+nQkBGxdyZJ07QVrGcW98Z2aBOxN+bVEnZYTn2ZJAqDc8IJmyPakGyXUzQR7AwhR5i1YBQEI68Km+7PqlsvabNzfJwENOOT13aqqrd+dzSH2EzuOL6GBEIsv2PyalutxQzgIe7hABI+6DWe70qd1l7JigEtqzgOEcoB8gbH4WQCghzHgd3x6356wjJ1KS9uFA9GM7WQ3fUpciGJTz4xaQcmmujBGAhRmGi9kycF8U5tzRwHwZTsjU6P7FinPR72fOua9RRlR0a+8xHxjv6vofvl9RgYS3jjLAjMuHgE/QZGjILkgxp/Ta9eybpF15hXvBYYd7w9cfeKXpwn57aAt2I313nThGdUrwyD+R8S2y9dDik82s84IkwxqIKa5uiBoynMPPGIaujMswDGncOO/ajVcqbsb2eDcDOqrX2kjCXY5UqnA5T2tUuz4n1hgrGWBwyxa6wXYnHX+ySc+hOTv9VxeNP0za9WBdFj7wpKA8UIRoWLYSlcLhUixPCDp4tu2z8HgsNWQgV8AfQ3EZZnb8B2E//srsmc8KwRpEqQje61QrNpkYLYPAH0s2PH2MwpfYREaYzR8eQn3SwOvhlfub+71UYcwbsYO+cMyPK8lPLZvmpZy2AT/GWpaebq8RmUsP82NcUigt6Q+sXfAm1ZvjyfNtmSIUSMnzQedr0ag3MBoi5Grd1AUp5hd/3fT6PbjekFcR8+CPp7aMXbpUCx6VjhO0BQV4y0JvsWEFCb2240RZY8NXPpRT4kVvZk9SvTUwSCiGmkMlCMuLaYJ0mr0S1TJir4OYxoAu9EQ2K4PnqkvnYNwM3ntRcoiuNFLFtF2tQZPjoarqTkyhG6hcb0yAVQSMSuaDnK8OclnEKM9GcgKbfzZ1AQ7xiCW7Y3vchd/d9Ig7kvuKyTh0sjIi1SoD9WkzJH2XF0XywmqamjvdVNSasZcm/oFDcoG56fryba4yXB38gRtsLROZe1ChNHmwD6sOYTOdi164K340QtuPAGKYB4ldit08Hm+OleWCLiZmFMFDkrXzdzEkmbxTJbmD0ONxzBtEIRj4Sxp8hGOuLAdZXZnjJxMyEUbKqkiQjwkrHgClAsACmMGq9SrUqPbpnX/zJB4nke32I0Gbms2gKlIqzy2oe9Gzp3FJuicEYJ8cCbg4cqgi8p+BekLiZKdM3+30TYv90RbDDLTGE6cBIfWbqxuGj8B2UCzgCY865ybGQTit63J/r5njyXPabRX70RpQ/h/KhlWbVhlhhrsGbismjhfHYbRWpkefdfRdUXkQheqCXPSw/Q42W+5ahKRvgt6Vdm5YBqhVMNLcjzHddzN2X1nyBIY4KIlKbYf6bscSaJ7kcUARIG+eIn9jt08lHo46EC3JKRxqtYGrNhgtFch+3I2j8sYT1Ohx0vGlmAN54w5F7Zml5a6HvH6TAPu2J8KyvEr2DnYaOD1NXce5Nfz1cz1N/ljuA9rWnewod9S9IEcihSooMhCiUF62BoMcLwrNKK7H6YJNjjWd/rE1NOse+V4qMy1c4kmf9UXg4qwT0bC7jqyIlflL5ljXc4mNrXCh3lzvgDsr/xZOZRgTGmJFKPzAMSeVh2v6truZxfQn/3YVwQixJcco23aWtZ9tqQGyWYphfJYeh1E81M+FUqaBr7NsSvDWITqjqsEnYMmdCo3Y5Hya5Jq6ZU1nkmI4Xk0DqtzISXR3pkJ1czc1wMI5js9bNmPHv79t3oaC9VO1f3BiXablOq56CQ63IvTUIKq8u55eAnOdZhAMlOTrtz/3Q2GZPtTBM3RY6HxDYJn/QGNhe45uFo1G4idWKjtKDbYAigKqNYuXA66Be/9ZroxcUFslCteBMYp7xcRpgYm859DA0yTKZ7tnrtWB0UpvX2k5DxZMEa4OuZrMNTwiM5r9Y3H5FZVVk4sxNyhabZnqr7OENKOkzxUiZOfs7sbrjCPSXFRx+Ib6147OAbtUsgFX8RDbgsKdMLKbVycJ73enVvV+AKa+XfH7dNqzdCqndVG2smCObI+Xymt0HvXt6EUXAyn2bI1btsszieXT2LXgu04wFYJj3dsdqVUKFQu8kbDabFOnCqb+Rj0EP4COiG9y7LNVwTXfzLpVdgE6Ufn5Gb9CQUML8eho0G1vv74MXnn31CNnqkfe2lsKrNqmKIIHfmah1Roe5/zgg/gNgOOvrkPBDnP70g0zO06PKw5Tu9ylhX/mIpXaACsVpMKi7hnBYgmfTZrdLoIS7HPkaqG+WdOakPnCceANv90xi6DUY1OYbAFtvFJOtiB/5vT+rXmfGeIkuKeQq4f11Fjzh8uWSCzRRtfNcKe79g8sRoT4pM8W8UKtPFZcfRm3jAY3dNWU28UOLXpyBrSgZ+Mgwpc3gG8XtSCk5w+3H9AKE9EyeP2Ihx+a/W6cv+taY+Oh0phfRhEGnz4iHuBqmM2IDzP+HykHUJdw/UxMgJ7Ch37ZoX1pJKX+VeVmERmTWSyhD+5veTjcmlWM5wrqVt6KOqz9E9wj3Wb69g2lQOiJkhpPI25Z0drJan/lt8zAszrsMkNxp1rYuesuzHR5CXqCcsOAW1p+xCs59FD9ktaHjKMRCkwfhi645GL3NTE/o+3f9TYHarEcSBSzW819Ewroo7Kqn2uaqnda5aa2cVLMUhJe2ATmS8LypcOjWl2dePEImTdZ6O+sWTPJ1w7w5cVs+2/RBsRIlLOfF1jryGyIM4paHAEY2cveRuih+2/HxjDZ0xyr3tgAszgDkR/ENJ2ay0p+ezvAZpSVQfJjlwfflswXGw6zAk3rd2IYxDsXV2xRPOH2AZM2yMxGTWpEpTkg0f6Ru9FPFiytSm8rDswMUvGYzLeCEJFTpG212qKAz001w9C3by7U1jF8zGjwv6XuEchYlQSousXDCV8+rMesDICc7vo72QlaTvebc09i37Bc6l5CGSViJaRsxQUsl4wWp0dAS4NHC8M6SxD8ss+pjs+XCM7Erc1kOhKuAI5+IG+aITNb1Sbl5M2nGEKeq5XjXnQFPSXIybYEJ03sMVzudlSg0You+UuHK2GkUHENAhXjZHUd04QhPMSM/qWogWV5sa11P9aNl1NPSUt5fypGt+HMultdpFzcu9E1jRq2l5XPhC6Z1RH4eCdz6jc/c91VG83crb7LTyo4pRSr+npa86WMjIB1cB0/vcZ+NvFD+Bh4QYCFfhoTlXJaMquONNI2mDtwXv5ivEa0bLuNJfyXo2B2runmPNiHU7DaD9FUbh2nS287HVeO6dYhQgCvanbRGufgaRPw27ddRMiJSJF31ccxVX2fot5aFN0GN70nFHhDUK/zqOJAC0BCLNCsduDEUn2KiOvViIfmFJe1Ah/HxxlqvEYmn9LxqXN+JjjG8Z5SkfkS05AES/SXbISAKKnC1nJ1hZgZ+8kZj+c+mgc2VU8x7eDgnlKqwSa06bhyQCP0/mB/SxWXJDUxmf16Zzik/4BgNHvVKyMDA1hgKaqRkOWWrMirw+ONhNkbkF97Ajbr1LdTVKKH+ymIZWvOESD83/VlhCe7ziTlxPkO9+uqdMslCREKPr5KKRJkhhEkNjp5Ftrx/4Lk4eFUqQad4x2yuhx3b2OoEgdWuufZxsOlS5ToWdMlJSkuB52shNo/J9Qa7+5DqCQ2jAkJwxnqKJhhSf1z5gpowwqh3TQ0OuUVCc+hF9C15HRzqZGikE7hjSnldXC6j2jU9tLTFZnvGO8AQdTJ8MHr+lH8QpqwoPA4nrb+zrQIz8rF+0InguGvLc7GexBPxtX86jhOLeha3VEaOJThyqdIS46fql9X2DMXvyEZZ4ar8O2hHLKSeXNexfIjE4FcmavBLU7jeBxwLLCAyuqwTOjVU0ASz7F+oEgicMH5mwnyp/JinC6hgukx3cssWhaW7DsQBWHr+tt8ABUQk9qZo7bsmGbT2K9ydGzCGvox0K/yX7CEfAmyOOPoYWks2Ew0zUI6m0mF1BYNwAVCh/5bAwvzKi99TVoNoTV32ZSvV8/raqXt2Zh+Xqrjkb7OXJOumlMYxncmaK7DP+rPv6IZoplaNC/imoMwu/OnriJqrPPtMmMfYysaogCsEmhKREOCpTwgSmlTKOsimRJxjEhT6LhmkErwOWlPtr++8ZNfO+q7KfIlmolFp002lsGTpAnNTbUUzuNy+Nlg4JDfODI6pKwxGpzZMr7kiVyHCHuKMFgZPjflSioYpunQcUb1xM1/yTv9ljyqT++V98KHcYnABGyo2vPPHqrUj+yXMLGXSs7fwYNw8UcmC901sXAGUHtiJbZ7fCgoWSAqq021Loou7PUE97rZDFgCzxEc5kfWOmFfGDBN7+hJRp1BAbXRrYh27wCbr8iWoXCS/jeBIqkSg+iJAZbCJ5i3MU2o+cNoI9TC9MHv5U847n6XPxJUBp2XGfd9cjXXm2MC/U1INUAAyVY34nNa1TeXcZ4SNm1HlWFnpFSvKxO/nkJlrRb4xc4gQo447a6nHdTDeG2fnGHAFK3izy0wgxELk7PS5IY1h7RSt+j3ngLrDHv8CAykxn89PzFV2FtpiyYYSjH8vDs2fhe7rDqOkGer9dOlOO+yf7BQBQ2xv55fafR7szyf5Ung24VyPDLdvb8su+aWX7IZHn7u3UFf2pW0uL+uEH+cOjdkkj6cwkDYkuGAZ1kz0c+X4AtBdrgGrMKDOJuEkZpz7z7Lg1dwz/MHAADd64K6hfP/tVyKj8RtDp+hCbtkcCbaWAD58o3T2XzJIAvnC1G57u3Dtau+JhdKZuVNMpXAWgBONWBE09QZLzIEaNV/XyVDVpb/wm+uSM+TXxpNCo8iKkrWrLGdXlBSPAxb7IuFzlSCkVP9WxTWbjIaVVcc3dpO8vqLzP5zSrzaJnrdN3nuUFLHu7TqeJRJvC/ZYKJCCKk7dNFvlDgFDIs9Dtc5bSWoJ4Yqasgy7CvBUfHMKJYrdyxCOrsv16MxgJtKEdGSWd+KhdyE+E1H6JmhSr47DKLxdw/gsDhZHm4TQn8oa/qkC1O137dM3zh6AhGc2FjoxJ3DhXV6KDPAD2EpSsuH8T8/Z8JXb6rtOBbAmQ7OFp1Zppib7JXHABN7LDjoaBwdjTzJ4C8nl703aZs4TeYKlvZ+xGlkHnqHP1R5xIdWPXDaCk5E/fqEbtk8S6HLyus/oDIgN/o62r71Js2z68SzJLLD9BwURbrTNH7t+EOZCzA6whNgs7SIshmBVDNv+wSja2+ZzBzz+DrJYSRHL5pa824uP6/7IY4N7TOE+upOVxrRmWAoNxFvYM7EVCHo7PZ2mLpRPJVdw/7O9dT8sOX55X+CrhGRehXq4+9QEopf9wKcPAIkad2VV1CBlmqFSX/iNSQgJEAn4QBCUjT+vJxOohNDmWpyrButVz+qpLqL+2Lbt39Gv3jRdyfwJnewlOE1jPPjR/X3icrqVPu3YS62ADdhXDHasRgxDUWYSeC38T2ioJdWUEKTVIX54VdssHkMAcvBKWunX4EniBR1neyu024LW9xrtPFsmK5GrDGnXMxM6Z754LjIwOR9LbQ90AqcKhRBxGQWyYsEtQhe3XMy/eYriRmWfcUoeIsn3pYPR3g67FOUgZbpu3RwFdd38D25+MOu+gSkO/0hYtTltOJbm6eLjFfvQQkEpBLhqt4aBCOqhvBkmvuE0VgXuArLHtWX5bWTIyZl9iTj1FoSuSeFSc+H5Abw/FF8YN07g0KWKLjtL+ftY1c/4NYkwCfaXpVn/Lz6lXIeHg5RTwTHva/1V8XWZVw/8eVnAflMx+cDLnN+z8mEcNvpyfcCF0yF6V5vMeRXbcU/pcN0+E6nRA/Qrfj+BMhfJqGj/rMFJUc9uS5lTgzNkRHkikFWscE0wegRN/jpJdQZ75TchfqPNGgvheceAUnfPca+GXy9EnHJtM9NssalZinjrPvff0Kh/bcRtm1CeuzcL2mtxAkSwtZmE3APdb7Gq5T1AnJyvo6AZ2ZshOu7GyhGIYUvl11Za2bbt3mobIM0VVV+iWI72+EWsyGkvD9Nw/gKHmgz5tXt9WpOGRncoEDwQo0sTqm+cFfUfzkhJaJgwtHg9rk4EX5zZHYMN1iZmI2np4/OuNA6x8bikQV8dJzbQmhpdb+6SmOyLJWJzz/cqRSpGm2k2ve1OR6DbGX8yMsJ/7uXHOfV/8cw5A60GyCHIzRVHgnmm6gZYrD3ohp3obwh7NMlCrGBpshzDg/ATQ9O4cNd30H/A4Ur28S7E6k6cYsiRjjoJ+Fm/KJzBs8GwNFpXpMHQBffUjtwbOkOAtRTmOPe1+pCSXSzCNFqMhQSRxofo+uYLBWDBl7fGUyifB6vuDOl/VjDTsVQYNG1/RLAmdI3moIzHDxXin8uUv5jzf15CDrTHhAdt8n/X3sZXb1uRaZx6k6ETmG0cK9NFeS3BsIq7xftEfeZDdDB4NvDjafOapz4GnY9ijtdiTwWk0UvDvM1MEec1OgArYKXABdCO5KUJ6ot5J7Gc2mnlVLx8oib5/HHHGbm+GEbtY7p1aajlbUmP9tLKPgZu25/vdrH/oDJivU+WSn2oYdmdICElEKpKVU0cRYdxyU2FnPTHm+ldbR27rkp673oGPkulScGUwYgp2s7OkkLbrD0hQaKdqfsZ/KBwE1oxrcZAD9Zd0rQSXR2gvDy8e3n2D7KtQldZVRHds8aofb4ZSQ2KN1opJBJtOLlI7Og0uu4XH2bnSq9DWgHCQdLLynhm6+dUIlld5rSmZYVu2VEsBRjbB0k2EmoOZJzizsJKNgoPXtI28AZKQ/0c6WKQrPeDLl5LYULJ53MCReY2w/ICEOMgGoE+My72kgXMl4DONJfFH4kx3pP0z2nX9iK72NjkmXyJ9lR6+dnSglUzGvA/sADUsnue1aVf9FzoYB6oopJJi4EvjIcNsb/vxnU+plfgc7f27KTR/x7ZI/DH6AoPEomLmU+WYlUXQ5RrbApE6bZr4WN5u00ns3SSHxCGyB1YR71Q82n1h/3CddT+FsUp5l4UTRyLkkm1TuFZm6Ix7RTE6i76AEknm6BexY8oat0EAWgidd6KfnEPV+K6wgwSd6JcLGwwfg=
`pragma protect end_data_block
`pragma protect digest_block
723cc0761026d66b29dcddbe821e1c0248d48de285e1f8152ca8e311e535561f
`pragma protect end_digest_block
`pragma protect end_protected
