`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 8855)
`pragma protect data_block
YdO+cgiw9sxHwBr9zwd2mkDRl/EkeK/vJe9fwr084GgYFOn0meutIAAYR250dODZV64gwXVgKJYKC/yqHPs/Frl0GnwSPmDHgvEnBbzqw3rCNDGsCuF1LJYuUD1AS4MVJv3xHe8PkdS78XXXn66VpkMNsUJ+B29MZwdElp6KCPWDcHcGvqnMZYG0OYmoUvRPTB8lQmrfC/tQjZ1t/gB9mX5Hn0VgQSo8IkvlKvaUKkaTnMXOHFJeJn4BfwoMn2ySFEUAqOr2nUqVPwCtGfurrvVhqvz0PJKM4sVV1bImOoI2pQz2CLsBMg+LgTuosBrp+VAnoBfpDu4tIPqYRRp5N3IhJDXhe5B9s8iLOGwVKqR10rfP+K15ohlwbACWHHn+lDgiXlUzZn4vi/MVp4p34U9AaTDmDRPjRx9WsbNaG7c378kt3+g+v1rJfcY2qbi/kzahLphqhTaP67J+tWAQKVMiQuGwrZp7fGcrAtQga5zZHsoqs9KJJ1WSjPasZE0j4LVQoC9j4Oe5qjsFx74AL6G14/5/6hS4MkT5taEklj54CJUwVBTfaTJlOoJCLsR6G9tZvl+9dXcTE176XYn9XfUjKLXlib1iKjpNHMCgoNvo0kCfOvG5faQUzIgqLcs2pP1G82r+seLZa1hiv3r9OjcWe3I24CnWndEYD2I1PDh8IfVQp5hv+MnAkQduaZuc7w5jOLYg0HeWL8ZqAUx8nf8+qOswFZ4LTosG3v/2prwZ4zfiWl4Y4OIf8W1VmzQWovkRm926g+k6s2rxcsVw1TdWB6rhnZc4It/RV1i2VEorMj4WBPhN9V2pOWsCUkQ1H7P5omUNNYwXP79iPp5xk1NYuf6YjMbjvRfWdJXuGHWbY3nbAibkMyWFzdynUb9dVXtdeSOkopt/2RrkjisyX+kPywRZfCMyIK380PtPe8c8DPgTqDXKKiEFnLplWmZ1IZIbryJ4s5NIVIy9R35wa7PZdifVDK4vuV64qbJigPgUW6y+2ErORmFVzqW/NMPvrHbvcjqAe46yfpwLeIerfBwHt9/CrIlVztu/YDTscvI9W9el/0Zy4w7muu2/9vX1IQZqp1k7hhLajRqhiz3+uhjOwZmCnEc1OKpUJfaI440uyZ9fymYizXhoYg4/Fvmem0ZB6WnUPHOysyL9HZuGy0VwTu+1xHyLglpY4iY6aiw2+v+K8ArTwh8iyQeolTNJIuPvdnry17/I+sP8KDzlQzWOk58RooLmy8MRJkt0Gh4y/PXoGz9nK/gkA3rOB/Cpf0hnY5nfsVBeN/6RGoUprvmTHs0e7HVOuFuWEj4vc/a4Xr7hCQkpma42suRCBUR7STKjdaIEzyY0oNCyYCr6vw7rZjiVLkVLV6PhAMeVzz/wR6154S7sIOn4ltHIJWMqd2ToQLykiUUrVyzaDNpCXyxldNiyJgVmb7SLJPJzTiJhianhlz6vLusRxv3ca5Da9SqAe44TMCq/NcSxzxiRvoVAuriV+EYPAI/o7jmIZdF0CkSzwoCNNOXByCalVYqAZHOBpHXCwSHkV55UJC8kYFYwXunvA0l8dkk3Ht0XLhoii2Aa56aq5mYczzK9YV3mExpDbJ50ZdvAm41QuzGPEMhiAetvSbHQV11Ig8ta2jy6q2EpQNULdLrA+a6T4qTcHLPaBfX6Q2GtHcAo5doB939t0o9zfGEMHvfkMTVyG+CKVqctXI4GYcnN34IJ/JSuM0I5WhjW6wnGmJlQQ7moguzNpu7fmKlqT0DWxYSNFLWNg/ItWE99Yp5MpRXg2v3wUzvhQSuR3eL0I0eoyQ6R5+LBADF+51Wn/+qkLjZp+7CF8wg6FqmTxPdJEfnFogTgS0Xdpu0TS29Gyd8eFvxaSV7AV9uJtXxUqUKqRlWCZ3YupfJ6zNXL4YaluowzEnI6eYv+BgeFdDA/OPLVhwrqootxuA27fT3qs0i5X2ZxiH9jdQ1fSGZMfv3fD8nTpxDuGCCgdPFhsh9Q/w7eXAZLaJmZjnQDUWk6iafm6oVaiXa1FI+dfD6gphcD/sjmNrZS68A5cGlb1vsK60vdCeqN6shYr/Cio9+qNqi9FGxhv4ZwCVtOdBMOo6N2YTL8EARgFmOFBjacVcWhosB3y3JdPXH+V/uGVA+Xa1BUg6J/M17c/OUwWAaQKsXLc49p2RkpQ0Tx0NKvXblbhFfcXZicrnd7dbE0moaZLa2dxBJfm8QjyBEciAfbGcawMBUjplKEGCF3KGyNobCIFwmqFZ4t5kd8IoR0p00Yq7GiVvyeFdOgoEn1hH7judjqef8o1BEpvGG8k5lpq6+S4LORzalFHNebDKhwMwexEptVp9X3q0tcSHdmRNy//cv4jTyZF5x9dyO26gSqCvtMzXwL8qySvHGl8VaUNNOYVyU0MHpMFYg9yROh5PDp+SqsBgZYDqVZ307uljmD389IR77WARt5rOtaXHTUtFLBhyOpXrd0cTJI1kv5z9onD0UecNFshNj0c3a7TqiTJEAMwjmIklYsl++tPotkQ1The2rnFXxHqmxbxiv6LzIC2GMMunhdb61QBnCIWZowVL+CxE/avm6RN5I6fZ57EBkQ/pzP2yaVssAL3eCOLGtn6Mye4A1W8tUJ7cnlmN0i6pdnGbRTdx7qsskcXLWZdkyOfakMLKhUG9BHkYXbcnZHHsHX8Y1EObHUNspvI198wx+vdekBLOdcDie++WkzOTTtUjw/f/R4ot3zH0KJ32b4h0zrqLUGqoUUqq34W7cQMIsn5xGpshWCfoPCOFfnCSzybI3n/7YAsXgTN84qTvUzTokTojSh5zUZAYejgrP+6ciwnRqCQXou42tTHg6GtJ2oFvingdBmv9276CzOEUpIiZwNFon6ykJoAZxWpHSZQUQBZ5hY6QAD8P7kszSo3O7FNXcvRRfkWJjVmBZRXtLyrEuKPB/8TjPMpsghXKXrJVeRP5F6nAPLGu/x9OvmJjGeQZms7hfREyGa2xz1i6weq3ktT3qcfGmRqMWIBSvhA69/fi1K22dSEbtvH0JpZ6WHA7Ky40KqAZqllhy2AEzsrREnKpz0LcbZtZPfmXsbgHRtk3NGDgwIP1L9W+DHxyDixYa8HTfSZ8/W5dhOQv1Vsq5CRa0D2nRP73kUKZk2hqIxSXWXHTtiVWFUo7A4UWm11gs9cJ5gYspl3uyFWjHGyCOHKwwH7c7rIQ76JKXh7OjqV6Mzwgm5n1tOSYBNHMcMKE+jgVJAEoL9oHWyeoR9/czukBDIe2uPK4ysuDTTn3r6kDvUPxCYrHj35GQKlo+0x3YCd2AjtECyhISTcZxMMyFhN+HZMZWqR3WHoC2iddmJFj/7v+bnsSKKoAkbXEpQTzY4LQg+U3vvKnZZiLIZhlA7/lAORCMMmEVgC05tHi8FSRB8i08ugbokvJ/Y3ocqgX67YD07eqoQR8lhYpCcXFuvaLx6YctCAxKdJ4pX0WrzAC8e/bCw0U2Uh4t5oz5HYf+EumpgSiXAdWXI/Vnoo0nrHbtCnCjQWKZI24+PWg/VGwbd3e8WXJAqubPJpjyek/WAIXs/lQBumGYizH4Ad+rDfCC5t+A5dzlfEroQzMLutzFafX2xUCzM0azE8dsUiWsb1snnj7BiCTRZ6mwPf1GLi4ftQ3hndz+4j6wev85TuGa35cazTdxEpUOU4UuvACfM+HlhFv7OJuiXwJmXVutd7sozZl2YR+pxkby9FiEd35K50330fJBkvan6KtyHpHXH3AkzBrLDuBbII1JmEkLPrJcp2YwI2fKwFcGwG2HTrk2k6F9PNWde/3GdEKFul9muMBUdhsK4iVt6L6ZEydQRo0jgenZI8gtDLUtsqmVZLXrm4LDOYpZhGhMvCNn28/pCQguCVcDuZSZW/IweYlPnYBw71xZcsQmMuNR33s9WDNqt4a+O8E5wdMt6Hs4QaTQub0RquE9ZGVwxy8yw2B+e797eiFXMhxUbbB/NnWDsiHcRm+9f+HTfjWiIhtPGpubIgCSHX6X4ugTUB9YtM936Dc+LkNFbGVvK7lkULc/wnmrUF6aHUK76HPxBGBCC1hPMz32sncSQ7CZPP6QUuBGBliJcY8YM1zMA0S+vnFKK1J71sl21caO0UwK+1cpLHlclqtwdAcdXuET8Pq1+jDhnpGSj5/G5PM7b1/S/f5nCu5SngHxqDh/wt76k6c5GmdvTR2vtYLVZxE/KuCxa/G1+qsa1Tc+jtNQ9rmiphX4iO6ksRV5WUQpAKFUOVjyNHTFLVRZMt+d7Y+ECvZYsUv1FzinFNqaZOeiZjGb39rK28qA5TTGxjefAbwcKHKZnkRIcV2seh1FVWeuFkN/2XwN35laqO78yQJXRV7bRUpu9fCjkoYvexmhcCGHRAwGRM3g2yvHBOEqdzWANltYIDw0XBAnrkbs5xo3gTRzcRO/WVz0Q9QKZfM0yar9WQh6x+7Io1kYSbApMkZeemCIc7AEnDcG7fZMcD5LRu2+4/Y5bxkZLI610ueEv5IM9+VBQ3UF+pS/5uGT4pMThOSapo8NekJfX8+gAgSYTINFZfn1RGbFOe5xBlffw/0vNKy1fN+E7ONtzL7hCOof5QuHhfxAhziM+p0Xk/OQKDq/YBhSnLzMI5l2DeoA6EKml3/XM33CrTC3S+cT4/5IWtATvD/erctM9CuEBcZ19IxYLzNGGSxFToBkx9VeUHiQih+xJs0sB3wWJ8o82vKg5xwWnj4qiTI8JLs5qoEQgh6e8YTIVKu51ZhzE/tTmoCpDZQhM2Gj8nwxQqVy+RgwPhKkMzzWC3ybTcgm737mwa7eWNbk9cEp1Vf7DwIxkbX5A1JX1cfehEFcQsUU9baa28h7In/6QpaaDQZ1hSL2+/m6kSGELfULfVqYo5TLz/rEPf04kNcWeRmrfe865nJ+UMEDIAJfKoj8IQmD+SYD+WPp7U17x+10DC2ZCYn8JmF1JViCDGSDEVR6FTAVwGa7KmV9LV7LKZWV2LE+4UV05lMUxJA71BWECA6blj7dz+HjQEHbyh66+NuDw7IEKFvxAHqlE7PzqLtjluPT4uqqusF+v0EjQKK9SlGKi729pZ5Nyxzadx1gKRcgoYH4VJUne7hh25im96CEhuLGN21sHvHrEpHr+gpBPfTTuI7RWbzr5tMR8Y+z23JROPNZlTJAfFnMOfGziIBUtJbTlRtSE/ZuRuItkMe9GScqGHVL4McBBx6OGoV0SSnFbEuy7yp3iKkGYj0Bv0JrSuNiKVjicnc0ytM9hMnlbDGt4GByXuZ62gLPH49/KQ+zgYGp8/2jTbLq1bg6ipymkiewnePYqxARuK0Ii5NrX5kBn6c5tEVHOv+J233qmHcYN6Hp42ZigrH/yG1vMPiqxXFayBwGlaBDOyFdsXOWj93T85YjAdEhi3NGapNa8gX+gW9qmzHrfP/W+YRDmB/NnEathiNkspEWqTnxH9PUcQcm4UUwoiPOWdlQL4KQaH/uMncsz+zeJQi/U3c8BE8JE7+SKHRCn/Go+DKUgvA0nwebP2WTUXSBucvg7uIZMhQqTkOQSCXC+Yh/nX+nitd0vOYTm4hkTJtpKpQek8cuqGS/bWUbsm+Bmg0xTM8qQfqGo7/mNXo9BahuAAHcTT4AwuWupMrQst04fuISgqHCWoN2MnzcVgpU7zozA8glbJPklbDl/tvzULtqqsG8potVuKTv/9P+l/u+pBCXeVG7OAApJPcrmjderzFYnqMqgDjqT0j/+UopDAqqWE1dVFzUkhVIyMJ1LOi0ktiqpcvWvD4AQwhJ1wcpdSdCimjO50kGVb9jC0HIij5KpymcFdTdZmr7mI7AzWZBIMH/EpJfNmMy16vHHpmfBWuQTMKk4tNvrB4S9Z3vJHne1e9ku8gfiFI1pyyjmmSf3Kk1NkodVI6C/aT1TR3GWrg5yV2uQsrBmH3a6Ecn9v5xGHrHL5ZqMXgHEvC3ogAZdKUDwhwc08L+S9dvloRPqbkZjNhtdLFbfYmeDUsEoi7oUUVLXy40/phXLROfSrtTdVjoXf9kKqGMq73QiwC4N5WB2CqicYT7lqH5SCECb4rlULWX395uwC7S+ylbF5ENGczG+SHUg5qiFamu29RJfbfFtJqTWNN8Emjalln8FwrVxbD7Tvtl7gU6sQNYn/dbwtH2vrU0CPojp05Kn5C+89CxD2duNPn+EzLJyYe/m9CGl8v8LuLFmOgV4Qz3M44PDtv08VtCTpxGbxaSH5eeg++jwmsEZ84MG/6YvVrwUpzfdBK1dj7/OXZy9QuUKRgkLmtnmlCwSdrXjBDpopHqV+ar4+Pwx1vZzCoAtg1N80BYZB/ioTHgxD306d7sz5hpAlFABrTndzjBV4uEuguLjmYgqDndetzw8KshfMWgDjosHT63+wCVDWs6VJsM02mQ1qc2tAtoP3URtqXGz3xHroguNEQ9P26BHP1Wz18DAqAOjn9nP0WkerZULaB0ETtj6bDTUo1uoQJ6vB1ZZlYEn38qd0lHYU6ZLKuZNKFGofzY32S64chnFcFYhSfruSoZ8zKSzBOCBqRLiBH3uuHYF1IE4ZXpxfDRrTndNUjg1/0w1UOd/bl8BQJHe5SgwA7eQs2hNVjMtTgOWs9xAfTWzmFiYHWzTnHG5JTp+q0lN1am++IXs1L7HlcqDKYeZongRF1yMnwrBqIu1uz7/wEez4nP596mae5YLf/oQXE2f+FnHz95FqUa9PR7Yr5JAfEkNRQAt3E06leyAZuWXxOLv6x/gTAwq+ESlVS/F4OO19/6fEW07l2pfGKJMklsEQoYeeaBdhqiPD3RZ0/X/qv9zApyp+4ktSH1BJkcnJATvxrNbUMA353Oz/OtWbaF2Xql4F/isbXNk4UhVv7DlbkBL9vdY/Ir+d0XCmlr3mysI+akbXCB5c4oo+Yip5hhbzGObGLGO7aPKgd2Boayl6qgSTFRBTdC7wvRc0F914HQxCy4LTqFmUgDcsjiMWXaRIhfa0ZvbIw22p5F0pHCqhZMZSrWk+xAUO5VO2hoY2svAKmOv3DWFQSuEDNqCk5qfPiRxe8qKvNArBh2g/Wtx9JU2YvTJvn48mbct++yH6M5opqdaeuhRP3MSOpfoTgnDexyDs8aRKlNwZUH43xtscdkUOgDRt4sPltTTutW+EAUu5SjYdQXPjtn7ii7fAXtk/WbihhLXx/e9aZhy4B0biJNBUmohMBYF9+T4BcDkSAT4p7GLDIfimM/3K4KZ9/xW9i2+t1AJYwKfEqBQtuWrTgsbcEPT6XCV0v0oHV5PD8fBLBU4H2lOHNNBVnFygtI+ZRtp85qKN7bzso7jYETt3Q3S6+2B2drP0kP3shYjs35pcnXnXmGCOIBBu0IMIhZ9Uyb6BcBab8r/B2jqXGmVYFFUXxGzwG1qaO7I4ebA3NxHNh/aIXic8PMrHNICT8qXERIkipIZoYPuKEsZUT1+/pEGOkgn/HtJa6dLdLYELqhe7lDE/5AyJiMu8zOLmJlqSoABHy9ikr5CmCE2lqJSVZldGQhpL2J1+Tk47wK7pZFJ3IV5G0NRG8UCTyovSGiGjh6kqXU77S7V5XpHsh9xYOxcvnhaF4KXXslekbxWgX1EfqRFpoIMMHDnbEVb8N5yzRCJCiTYnlewoFV7rgxu9eVc1d2rFFnBFw8R7a4qwmwFidNl5ahbdZgs/KnqDyLXr+suDpMFuhDrS+vwe5/bXJJdAI5wjv/QyyVMgtIXtNiUFiCqeUkBca0iV3MMEkHAwl3Wm4XbXw/4a3Grfl9LqOhm837lzfF4qYZ8zGGZxBNsdimhpsT4icMPGiFtrK41tFDtF98gaJlDQBQsue8IXI+I2HOrLGMABH0aT6E6ymgDLqpnAmkCATSCgwSys7ioHXD0PDX15ITviAK2Sb8KWgG4ukfLD0eJv1gu8pkoqLPpnCMgD9mAyx0uDSZhxoGjCaDIr/mhjX1XKBgcdvAzvXhtYdgYZ1x1N291bMaIXp1Q2+QPHSpncBtIoMBukGuIaLktpLaKDA7RaRDZerife7YY1XNMuA1ogjHFVhdFJ+2+VbAPQGE7HFDMjkpd5zGoaQ1hJR58rq+DPfLmPs2KGb2oVSsIMVZrvyi3w4H5Ava9Hy1KcQwAvdSEM1Cs97xISW1+Q1QqO+ZTb5KN8VietITeFD2VzxF9l9erEYdkmC7zFXr10UVkvz/85gBdDkgiozww8i106AHx+nNEEVB00Myu9pD4RLg3FTS2HF13ZndYKOV3Ij6ZzwGPCGpiZIuWBF1/vM0VWCc3s4jI8bFbw3TxvsnsVfwthaqNXgcB/78WW4QZE2o/5hVza9GBZ8WqElof6We3cKEYXj/afIrstz9VhkWZN1Q+2SGjin26hIwQZgzFGl9BLbPqR1XFkQJz2OceLsXCpyMQYev5/iGJJX/mQjshMosZum7vNlEL1W447Xtk4YHLjjAzZJ+4fz8+0sqTXdVpzp2jAG5Eq35g2GDJtjdc0uWATxymVBEMnarhksR26o184LuaZC1kdJ4gOnCvOnjNVtE8mZKvhfdWxSmuzYp8WZnt+fFDxF8rD4AT2VWZKmDFWGWihovO4lEuvRKgHaKSeZJ2dzcr1GY12N1MKqXjR+2TtoKJaQX4wYO+TXhsZotr5WBCZ0iNfjnwNjLLjOswCDXySgWPUuHGYG7meo7oO8riYDl8qZDIsqYr0bb9p4SnoSaSM+5aiwkaC7NKL/e+z+OIiR62nIBBWRDSHqZnsb96Hbyl0O895M4yorTTmSeQwOenFYI0E5JmkrgBBPqIo6qOMUnk7DhbC4N2S7T0s59QwoHVADsU1xUNrqSkissnv9icyrZzV+vnXEA1CPC1ET0aoCPNLyBC1iYsp9tcsPxOrv2/tTyFfA3wI+LmHSBX+Vi5LinazzNXO5Rz9CtLWQcSnFjW7gHdAsCVLmYkwfWzAWtsHVciHloMjN/vJfex8mCWWgKZG6rQnBtbwER6cQ1oCLjGCkyzy3nu394jXl970zrdOxdl1VQU4BhtTiAYsckaI9zO280pP+JJmUpVeKZPq7ymDbpThcfoqI/AIFYuHLnfoLBot++RhqtW0Rviwm0pCOz3GitV3NyBBdOIcsb9zZL1anR+0n1YUJ3Z2VS/wn5Nwwfb9bQo+x5n0VqAJKBHWo8ufwPC+cNOygLAqehSuTfc+CGfRi9BM4OsNXP7IXc2dIx9hL6qsB8Y1iX+0KH+kdaziskYiUuhhGDJ1lV+9suuHPyAKJ9vWijAdwTdBz8OcvY+Tz+RYAdOiZkTvI4XgqjHA2JiCtDpxkpuJa/+pYqhLuJuRztfTQtCOEN79mWeHFQ/spF+92oWu0uvu45L2Sv62A5FfuxQsLzdfpwQGQnUgsIRI7OuoMtgSjsPs+H3+tSDbRCl9H0fRYUUj1RFaV6Nw+bQwthHnGlCeIhBsi6jGCXSPBbM6SHV+IOBnpMPDOkk5IXVX0Uys5UuQ+/rzkuAg7rbH5xImksDRvrBiUfBZvEZK7/inHdmSFTVgtW2cmAt1sxmgeSOJg7f4PnBx2FnCszlbs4AUfwFR7s/lrvEhqcKqVE/Thd7uDEMnsSNKyczwVcLwx05/d8QPA3j1wbiilk2mhWzGCNEyWisyvacZzA5eFChHOW+hMVqbT9fbqmXhVxW7QtKhbCVTBc7mrefTXQaWXxa3qL4jnIxLYchQZlOcosJHs+aPjv6+HZs4Z4ePNRw1uhiLGOUS9Zib+N9ZVLKkQ7s/5B7d0Jy9Hae9yMPf333NFNjfmY9ERsk8NVmgFHFjKi4oGcMVIQH9Pvu3Xk8vhx19nxSBiIUVjSTIlSb4g4hOsMOb2uu2xMSZeUNjrYOxYgJlO5hOE/E9KbjJIvwQkaUvOCb4vg3Yko39YS1Atx4ZgHeaPtUzPrUeel4CqEuOWy1SOaKTTLZ8iP2VZP2dVoBYlVgLO5Puw6WXEhz3XZclidJMGmn7Td2uFxPP4DRWP8XscP8DUaeo39/t9ffjAMeJffO+DXzWC9WlM62tQfSFviuIHDOnkd4nmUdTCzTqF5nuF1m11ceNrLUeKF0WvSQPO8nd2K97MgwVJLfms++tsw43CfPB36bJdPLKihLpgf56ScooULsJd0KjIJ3po0BlBAfmX1/h5AkAZnnu7iasitK02rNK6KZUzwB/hqhOnoNbILo+49dy1eSXmlGg3fBdOI/XLsKMvQJ20pa8IY/ToR4S0O43CBe+Qx05S7cjA0k3ho8cKJ12zxSCerYRdkrsrLlpOgxWwVGHeUZ8XanSeitp6G+TWOktw6IWJk9X5hCteWYUDazg/lFW7e3ttxo/1ywwdg5UrNzolbTaD8/MypaHtwzUjWQvBSXEYQ/k5dD4m9vHv9JI/XEMN2ITXhMrzS43W5fk2AOvy7lyLZvxzWn/E9hxSyhYLjcU5nUmtsDeAw5Ifvwgp1qK4NP0Fu8OSkhsJBMNcrbHBhXB6Ti1Jab78NBY+6UUpUO9W8k0sJ3jZKBCXS4+JdKm50bUuR5S9NEh3EePDcnYSWq+Uo4l/vXWj8/TDS8F0OgIjIImY1fnaUv+KM4QEH//d9wC83RTvptZSgGjVIbcGR2qWoIhJGn1+a+227QvGpTEAhkLMhk3G73NKZHBMHTwxcLZN4cD+fioyTWhkUWqjUm2prUGtZ3uf15JPshECnI5stGDD2psNeh4baQgfm2y2Y2/5Ptd5s3g9OM6XNR8E+loOjDSgqZPZ2d1itS38Uj1oe6WxB8MwR9x+GJvKzpy2ZAGZIRIyAAnCZ+LqsZKaQlMCtckeUvN2pfWoxG3HqIaOWrzE10pIJOzpbxeVwAz1QCLtzEj56pYdfMfRPpjsBt2mzizCGkoDqsgZB6kiOZu6lhUwrRSoK92A9lNrPqWGtxWBFMSRh95RrxLqQ7Hh1Vhhyy2JHJ+7+eBNIDKK1Rt8QIZ/nrLAeE422ljOv4mG1orCIwOCdp0x4Q/C3HCBWMiiUsT96BPWCzgP3W53FGmus465zz6/7jVbsRusmeQ9dbgUP1XrMSVQJkvnhEgcGBUsQzkm3LIO69m5PD2lj3Aj072DCseVLMYGSRp6hZEcpJ7DKZMzwP++ivORD/s4Jqy+2rGepR7/mbvsqDINEXZKROwPyVjAREtsVqXZJ9oGCRYLnjha8ch9xx0x0JqpwWha5FaA/1EsQe6aFhOBDg4S3r8E30rFbgT9xHdjuSKyzQbhsSF+0znINtq/b2C6IO/ElvDRPaeXYVASrg4ew19G9Ojeeq6EXb0h3wWkg/B4nDUZbFf2D+Juz05aB2Lpn0QwVncXQrBj2Oz+MRRFD/4x1YGOih9hAhjkvhZqceT5zWDze9ea/Yk+E+YNig6y8YEm42hYCcBztN7kcz4EIUP6EQSpufXMZNjBxv7XGlVs8zhmKZeT5dMAi8sVS+PSJqe4fcf/kYvmN9TCZ3bTmdz31aG2nkNH1kIqD/Wc0SeF2eJaxwwYHZqi1hniIKJxTy1stIp+wD+OncyhEtaT7siuLfpd0I8TBNOU/xJ+8C329DOBwwRJwmgegv4EiBFMcKhnhDh7T4ir+dartQChvm4WEqrS4oon4+AMtFsyR9WWsyEjkCTooVq2LIicpfG3GwG+IIREMprY4T8FlKDPYbgxhgk9kFAoOEMLz++pF2C/u7yy8LS004k3wDI6XNbRWBMfOA7y42C8fTop7uLXDllN5cJ3JOUruCuLWEgeZWi4nVsg0a3K3qqA54I90cexqa7zUh6BOqVmcnC98vlonT6etMukVbxnpSwO1lz7UBktz33bG/DwftLDT0EDNXTZ+lNSVefjUywibURMKM/lw=
`pragma protect end_data_block
`pragma protect digest_block
697ff223c85df22423c438d2b960e4d34be55b19988cd23693593180dacce82c
`pragma protect end_digest_block
`pragma protect end_protected
