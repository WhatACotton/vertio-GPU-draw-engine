`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 7471)
`pragma protect data_block
7mfJiylnQTHROHhT1qXBPEkdjtHDpORENwZqmDFTzO4R1bk+9i+KXx1Niggc5W57W/O3aEtlp9Xbw9P1qcGtuUtBb9Z3vXQ5u5cGXxLMWgVoFe8yeQoQLNgRAWzkO/zXj/rdGoj1h5wEMVwX08qQKNVA991ehTrjzrjwRYZ7qoEmq8AJ9/DGPze/Gyanam2bC6ibguRC7qnm3wd2bbXcN6mHKge97CAja5ouVM98Cq0MbURfV7i/pV0JdpOsimbqkgsDYPg/HyiuzTzjZS4n3dgDzfxgVkGQZOiC1LmQKQUS8gii3lrM3HP0WhmFYihau8VtEL/kjsLPlhrQtFX8GGBgmCXnpL41hnlZ3POgLSclt63uGPofRXjTxVYJI+i4LlwZwTR5cP5c2yI49xi+g2PpS4IF8AII9aIAZWzutjOZAC3u8tXzdwOMj+ihfypAo7XLQWw69d0UzqLOf2c6pVbwEGt3h/4xPPC5CMB29q9ypPZ/16AQ95ZqMSdSuNIr2P1pPvdHNkSkz5wQyALNTXBpdVd/0AZKbJIuQ8LWU0xXMvnBGJtV4bjLSpNPCKHyySO5A49SbdVfpxMgzRW7vZmMqy1WrHL+BNiQuJwl641RXZFQk1dBDITCf+T08Y00WIVWjrG/XSco42vCI4yOZloWftVRhLz7hpA2JcIk5hMy1Meei46Kwu5BGKjQKz7m8otAruhAV/9F9csOrIIMtfjPd+wvuLRlOFQAXfwcS2VR66pX2E//d7zQF6WWv+mDIuJXm/laB99QQPHxvHJ0qBK23+VVcQpWVkc2KTLHIqbF30R9rlQP4EWgHd4Xrr8BRxb0UFuaZie+a0/cnRNW0D5zE+Pr6m5bErHQLuZPtvNnJKEu+J3ZWJ1z3C212/FmNi3f2GRadHTbZpxH+JUesxC2EVpECKBvFfVvpKxprzD5zbhbeN3HiDROhXkFCu2whbeUuW41kv7IyqDzmIopsq++OpgfgrQrkxZmkoOxfvskTuyswSObo9jvFg8MOONjwEHobPks+R4xga9xV0JtarglH5rqhS4wtIg8t3CS7fBE+r2XnrMsCIrlCeHOnGX/H/XHaNztJSbmOjByjuA/zlxOoY6+N3CvfoO9TrxQh6nyY4B3/I85NiDWuf5KmFNNlL9TBt+gc55pMHhlGDBGifGGBjao6MGSekXOAkx2WTSHnUJF5C3m84wH0HShfcFcqvIyoR4yphFg6Ll5Td0ehtw5+JePkNzms5LwjXgfYX4rImFgV9WaSc59v6WaJRhOf0AoWgQabB2FABVJsiYNFpRei/lhPyKH/JSBno520SlEbnFNPljnE8IFT3ZY5Ews+B9tqQ3OHakTKhYQSU24SrTVL84eqfETWG+q2LzSV0S4qmdvuD/3hfAANdbLnmBPPBohO+Vwxh4mf2qzk7BgSurXJY1r45q45n7Byb6QZEcca3wDwg7pVl9DZgGIREtH5rSx8FR5MCfPz+H3n7JnZlsAFDNZ8ZrFBmmGr9UadTKRWUJL3gxfhFRrm7ew1Y+nJi41kFo4pooX1gxZop7QswArcgsJBxJwUDr/OZO8Y/2hqM2u4xO/H4jnuPpmygqDWX4JZK1pvlJydCh+1eEoh8/1gX46kUPxsvV6wZUUhNzfW0mBYe8iz346vdfcFsaBYk1IJAUMiNpRNrZQUWCGUMZDyvQwQhKvqJbYXASVHA8zra8kqOpMFd7vZYUgPoFq5vTp2zCZ7RLQj8KFrRWLPYDIquhcDajVdh6tfVJgaG3JAjnVYbk1jqFIWfuwANPM3A6XSFqTRRunDcp9RP0GaZAF/SeH+U41LlZ50KGPvVlP4WGREizvPknG3dGRVAcb7DBgEUk2kFxjThMtYQ33DcymOoqhdSRX8R45bP21imPXpZotgAFG65GnAiFe/zqn/Ehal6TJp1+qbgBIA4mnEqLqai+QEKBIas79sMG2RoyO/D+tBn8fkFiHdBtMJ8v4uDgz3zsZXjmiU4J2o52yMAnK/nu8taP+WrHAT66sZznz4HRh+zXn1GknEHhjprZtjaM6o8GOOvCJiut3ghUbOqROe6S1SY8Nw8IfGonauw+RkiXccGscbvqb+MzDY1c24pggJIgmjq2h8SHQXKNXCAt9DPcqyc5VWxHAsvGNj9D1jSTPucZfy6wby9PQcP48LL4eoym2cQ4jGM9n8HaJ7fuEiay4tT1OJiZRfDc1WPlYyP/+3PssF1VzUpigqWLpY3StMzMy/EboepJ9HBeunAlJ1Oh5d9hLCipFTYa88z6DldW3Plo9yS0l/igjZYkjiay4cpSyTkQFpgDCMRRXP0y2ENKPIPF9K3on2wbMXXeqC4ECJ2z1CnM4BxO4ZmJeK2CmvUyQVLk9bzm3kxfBNFjaR8vItms6SLTSUGI8BTvfpcIV+a/2sLl0zTksJtYZlBhEbaDGQ1+4JWs3tl8MaeCxCOVOpTlGkSctPX0N5nN9qWUeRwm0nEeNswFCB24rgDYXA5vg/Fpqv2P6hvnkx//x1tevbisTUMNJMGcS+H2aFwt3FvSE40O0enXY7NqLpbsxX94wKE12udvz/JfmeNzzQ+2/ye6xCLWgJOfvQe0ItPVdIW7/876ZW9sy2vxlmTT+pZGBil4HKlpv1qQhfs9gvAHyg/Z9tTNnN5oUIGj6e04MYahQFbeiFL52nLs9wYI5cFlXz0HZ6P8CXFZbeRKK6VgyZvbqHdxtGxSWiHL6KV5r0aYJ4TD3sQlktm4yvy5YJIisBDr+M5h/tK5w4wRlIzig8W/aQ2VoBI9jnkzIZb45BYWMLRynOCIKgnwRCGD3K2Xcph1+jqVtT5HHgmh4y6BuonT0ci7VvveoOgEF8U68m1rwMzNnfuKQ3f34/S+JuAxOFOt0z9wqV4dtOqkf0ayETMHfrFohbYI3l016YF9C+0tCRn8llHO2UlJ3b7fgCMftjHDVZbqElSGccLLtT/iXYVk3OcsWBkchEQha0uVyChTM71DUaFvedmSWX0O4ymkuvaNSSK9RUxNutQ71Iy30mmvCAB0RhPbuBOMovjO8HCDWSdrMn8EcqR1z6Y35lTxHHUCSw++1Ucs5qKMl4l5UC4jjPe10Lfnr5gbgYVqmLmekjk847BuicmLS2DgcWhSkqUZwBuzM8TFOvtwKv50pZdzJjSUyFx8e7rffOoKNIk1y+R/XjcOyD3uU6Y4KsCAxxL/ner1tI8Y3nKns6PiUdpzC8igKO7TzHHkuszTtBfrfugRiCiv73/bwx6k2tbsvD0QJTWDd/I3lgit+ruWok6ElCVwCSVY35JOugdhBd968o7EsvfGllkcYv7YcRICq2j2y4BVej0c6+6lYZpjX7AlLTAVfXYOrnDinfekrUdVrm8AzdrJ0KCFhjCNXwxHpnAtEuN5QGa53djTSux1bx+AnkJApdV2YVfXczgOYKB/ilp6bsB78xAZee7Yul+VsD8MhMzTrJbfAeTNkDszSjeTRD+WyO7ufUFFu1ZnqpxFh2kDT+iGcSEFk6sdmtUjZ8voycYgeq9eUa4UZVAW6FNG7uOTDmq7Awr2gFxbRii8hglxFpY8fyoD7EOQCnpvJ20Paz3RA6GMc7GYpigi3ntVa1BUdiHBTtA47GbdwaOU6E2YQhQtumxe5u7izOuzESnVjJzqP+t/aPUrPnOl31mUF7Lt20n8xrB5LiqvlS1yv06sBv/J9MBoY77iXRnNTQR0d+MrBYC1G+AFPCSZhJTcWZGjX8i4BBrjP072T5rw1ol6aSkSJN7c/UYbN6RvJWsWQVPmUVjtLFT+ZEJFChOMXLFeVM5zPjC7vha1UeYMVvzBjk9G4xWzMLaZ3dRYvtk1FJtqeGmpVNQHLFg/w8ZKCf4g9oDo1qpmtls7x4YDS6wLGVcwREYCmwiRQvs+knT9jh33c/LwySaHHKc2jghLJ0+9D/qj+xgnc19dgWHc2UU2EP+BoPW/zTjst1FpZH4CuvYbtetoSWeUW6O5UcFliGOCjrVYJnh6p34qo7XEKgwffrwdDz+IpQYScteCvc9jgnPML+qeYZecVe/S8Ag+OkoXQ1u4rK3xJIJ6vef6Wq422fMmczb94iYMweNJRjs8UywwVfLEeg4hKae3GhRrX/Jq2GOYg1JmN9Cj/eP872d/SwfcNddJHgqjeJbJ0frHGMfK7uR6Rh3Bq+YKuQEwNI3iSE6aEfs3tFWJaqX5vj0m6TlKfitLuudwcB6DFo22w0yd2Adorxa8K7fHGDMahe351lU7D03JOrKuuegsCJbC7xHGbB5rtodCsd/8Yw2gRTGIZ/BFGe2/lfrvBsYz/0sXwbx5/5jpPGiN7YuUF0dj7uc0PwnM5znBdL4G5FsCTgL3nlvgWH4P9Nr5LKkGdzArHIqu0WpHr8pbABwnBECt16HuCb186OXSJlgOZcq/+Gd3h52D+Ut5lbwnEcdgvRlFzVMQwDsGO5l0w5wUvg7xwRjAXxvSe54Ra17jTxXG8zV86VFn6WQ/XWB323SK7eQixPErFyixnOGYRLsEsaYB//0PxboHo8+d4LMkv8QYPQkiViiaqILJcmT3rsBiORF71AZdr/AJl1KdUYqNwZGIYJ6YZ33hEKbc6Cf409JvZuJtx7ji8l5EiuCfrNGmSq1yaAZ8Tb2RQDNkolinMd6yJF6tVxZb9wSBE23AtWBIjsOAenZmGChWtW0ce+Vek/DklJVJLk+hu0i26CBGWmhPZROPE3cozqBJfqcyjnHUUWxKoMTifYEOeDEnihTk/uqrA9eMnbNugAuSH06D/t/QLADRYO6D/Yh2kW7SM0uQv2fI05nSQ4CrFxwmOTGJJmDCJZvOEwj3KLkbGHTax4wx0/yPy3SVUBmFPQrvWG9qzNHdimCG7LXa1GAwDOpgUe0hCrsVdmDYTvjJTYwFzKy6xWlTnmgHVI1HFbXoe4N0WCnIWrCTF1EA5A0iG8awbACKUVgoD4MZIcFpTL4lKpkWLdSEHZmkR4QoJ/JRpNh1aOvw1KWbpGomr01O6CPNfMCIhtnxDhioefvJ4WVHsceVesgAAGje7n+OgSDbkdE895niWYkr6GFFONBslQex8lT+DLHGcTbM+xNKVSYiEA/mHG+FXwYgGUCasxSTGjoUNBvnhaHkf4dLXiNN9WbsG5esWbprUsYgN/2MbCBw7LFOJVtmxRp1NwGbF9zKVUTgY9pIvvzagrt3U4Y2IcGdGOsUn3bm5npsbrHYwpfS5g3K1fBLZc+7KO5W6xSGLrwGP33bYzMh0+OSCEUKmNy6Xunz/Sv59d2OPmN6XH6oK2x/oqnr5/51yZy3dRMz8gI2vjp7OB8SyfL1HJx4xIEB45aWe5K0ORmG7TN7E6zLt1fSiF9kVzssxf+Js8i7GwJEgfP+Db679ZhE8oSCTuDePElpBU3jwROfraKzCKVPdcGiqV2sn7wd7d6BOy4wyrCoAcikL7ffLDJXqFlOehSjxNqunK6XmJ3ly/VvJHVnaBDjunTPeI7ZDhmlDVbNQVab8OBOuXCprypBGO5EXWrhzLaP8RxZb8r20h03wvx2jfvIe0xnXzKKSa83EalT14tZeojMEWvdXDc41+bN02Rnr5xpt1JpPrULhKisSSIwbzjDj80Snu0628GUWO7BscTh1zLmwL81xcNOS5fQtHWn+y0nTOVeuhjnCpg7HzIG+8oW9Ym11NaWkhtHziwTZttEvUrP0cxlDK4pZp7ZXxalkVw08NpCMms3fkdY3INaOAVWcsEmCdPiXdnIF9J4qM+g4xWj9jI2yPcKbaeU4mGxSGb3/GkoY28zphYn3eZfsrGXXPVYU6eKbeN05v42TFc2qY1VdfMJRiVgOIPeGcBCNHeh4FIgE3x6Vg2FD6hB8VN1p7v9VvkdijQoW+3srGqc3TbYOsjK1rLM/CXCQyZosn6xqy10rm+u4MVzrl+2vcbLO6OV3Cu+DSPuyntNB9p+Uc1iD3mhycgqSX6NwwxKs2wFbUir7Pkq8BiUB1FVGnrn6LjMhavMkoOYNKSe5BKRyflSffNdj33DAqEB0z6xTYEbDFkYZiXJ2r9yvDNdxfwnikxgkQsJaTvC9w4vs576LDUFUv2gFlvwNWL95R3qz2nnYIUSXlNCNITnBeaFSwCtpS8F20A2scb5JOksDLpCrGQ5OtA2n69VcW/d4P9fx0eHP8r1anjS+QEEFC+l89BDUTe+UjCvD118AHoFErVZ82DsOMPc5jJKpJrC+ktcDqxPtQ5dx2Rz+ichGAKgOH0RJ+gnl4jjcIeo5qjD1eOP69z7GKH2OSWkxxyBjS77MyHmE9UhELnoTnvZBEEjYxuUO38h/YRNnIQCFk+Pm5//GF2Ij2rDtJdBAzNgzjtqCPM8pW0JvJ5GdU/pCpYAByRbd/MrEBK7F1wrAPG+FOmj5HCIeC+AWaD5h38mLP60xqYvk9bP+T5HXaRTfsUv9zNMnyQHXiZSpTmC4HErv7d8K65379HIGpURbBp1wIge9VUY73TKzj82wp/zPR1SCcyim0TWGpht8mm5J/A96XOP1/z5+GRTiyzLwXeJ/M/uYKuGIbTtQ8ZHG9vtYGO5ZjlzB+NNth6rASXP2fVo4kbekvJ9Y6aWlO9zGE6xSwZg4j93ZXxo/t+PWJ9xvzskK1ozIFEQZbO5frjB4c+biS+mqDTjAfhAWVWkIyUrDKm94S3wP2muCf36kI17AMDbz6CiAii/qZUPJv01s6cp6vmfLzR4CbzrCNu5rZqvLmI9yjcw7mOcFIcLq05PrijkZJYwP24xKHFqJVqwoJhAQNId3WbIYerVW/YB98cxfl5MgOty5QWGgAyAEl5JaRHEp8kuLWxNvJ+zVEupd8HhkV3jFbgxaW87GHWkMHBYkxOwWVywS0sWc9b9pzh8bCpKJUBLoyhfsuQoDN6RNeSNX8J05ZbbK0AAa9Vy3MK+Bm8x6z/OHNf+gdZZZLZRyFaVWu6KjAOFcQy8DRQ3gXvid2S47WV4TuAaIwB4A5kNmN3DTcC7y9y/yZjQ8zy0eP4rkoH6n2R/tq3lVjhGgbMELstf5AAXUEqkQvc6/VXBQxHKvngPEmZrYjfgAFXK/TPVc8jjJn9lJn1sGJjy7nn2TLPTBgeG1zK8oF1ovnrv95wHq2lpDuOZNJCoMZsqTJide7t3yqhEQboukKTqp0xS3fM6WfuqbKn2kDXrXCCErBpVzwi5W2FPrqGL+SDMr4EbFpM08AuO0+BrczNZ3s3vCJR5TQSgC8gkhscNGPcTThKMYRybe0cgYKpKKBWdDkXmUBUkUVnEvtfhmQJaxLsIFl4nFn7Pym3V0mFGMTeVrJ2txBk5spNJ9EtMltt1TJD76LkUo1JN+Etjl5rGfQ+g56s3chdbzxSULTKLttSYXt2klW++sp6G/LRgxAtqaGk0dm0ChK1bxZLSkm8P5Ktdk757KxLU8riL7xXtBzhHs1SsS7YlImq463CvMGBQJra6T2mEmpxYJ9vuTDEmFjSV+LgK704uGb9jWCJSqjgrjVafVnI8+oFIVpMnGq/qLJmEBWa4vEPHS5YQ+EVY7lKT21vlY6vGTToUVZSUnoMh0xMqMyzR10Id/n3CGxfDIaugmGyMABqCm/adT0n1jeOXLUqViORRVXO9ehaYKxDk7iVtzUyFTdw/LSGb8GpNsDUJlduCusTLHqvvMsx97V80j6Gcn9m+sSVB1QmkK9vIiQaK+XNh8Jzja3Dn6ICJCdDeTrBvezkH8LaFywSq9wbgaAgc/IVV70+pJsT4Sf4SJgVBBqdpBc7nvpBx/2awe0Dxc6wuays1Di/1vfN+dgN3eM94lTFuX/tRbTD13/e9Yib0DtXyQwUJHwgu8ILIu8+JBt/rHEFeMcuddfwAPI/oxrtrY91fHicHR4wq+tvv8D/yMnYU3+q0KLX7aFlAMRU0uttdiR1n5e4I0z0z3sqTGRmlWO4zzUGVnSqXtu69fevUOS7JgQEa25SQw4wFwbYGGxE8DlExnvD1w0e18GMmGoIu7FFXs9NLnlaz06W9rubNN5uCx9ofj+eWZgOR/fn7DOsC3gjVJUZXA0H1TXcTmbW7Pk5kAes0zUK3OuSry9YeblF71RTCTK87oQxpiiDxqO4+jVp2uTJVUmwrsZ0+V2pQWjnXC1qhd17wCJSpuxZjdODj8d9wpsuK77UcOwAMpnYjqfuWhb0/okN+m3PQJUt0xsPELpJyX0VKSnrK4INk6sh7Py9lEjMcJyypeOXE5QAqiTj9AeEOzcPNbfAbI5CDfikLCHMbzTAMvwO86z4ssKLfyUyaJEqgk2YepjbFL+of37bvSUMH20wd5B0AUuEcLjY1HlA1iOxbbuAvqJH5Ej5oiH51gMKQMeejhQbYkt0rSHPo4cDlHPHmXw+/ebT8YorBr678bOMOe+Uj9iuH2dnq9g06k/34GLWHYIXo9W/xBAlql4crauzWgCHgrCZq8SOh3NvzpcfdecuF7FFilbL1DMDv0+0Pip4ZUbZwdm4ynf+/tCW53iIwLq6LOOEiKsGb53UEPcUFaE++WFzzI28aMzeauqzIC1SVkPgDtWBiT5UYMk5qrLqIITzUZr8zDXSJqHFyGxW3ZY3bvWG6gwd3IZ22oTAtScktur0I9mLeFVwpAjZ73y78qniJKO8jslx/s7oir6JNq4Nh5vwchQLX0WX4NXiTeGf76V/O9zaXuElGEykc2x8hy4CmJwwP4Y7QxYBYHk73PGKz17leDJCYu0DBoVNmLp+cdHAWSUbd6ZNBgqHskz/PU3uGP4ivGne0iWdGmg8Lr71QwmwUDyxxeLFQ1LQNnpgHv7FhEEr12Dh4KyU5GN9XjoZgVGJx3tAlkxeh1r9C8TcingFCcsXFiaWi32Clt01mucJEsraVd43QHmymNZxkDybYkq4tvQOHUOO/ZyGPFvVlr/bFMgCZ2ZCRwfK8zjuDICO77mFc63uLHdQepKu7UJ+nUoBWwadwI3aZLnYhkjpwERVD+k6+SPZunnFoUM/qPy7p21ZvCDy/ysg7oh1/1YW44EMSx3YX3jSTjkSWzYLgzE0xcnMQKwFNLU1sRttpEL7fWW/8jcUsMqCC2ZsN4b509dWXZLm007pe0hiHqXz28hqxtWzYN6aFmxa8PdjZbmkmwDI7gZrI5C+AoIOdBxA2hM4GZAjJhsHq28IvhW9/aW4NNEkBAx3W75rKZhX6OrMamYo4i10Ys1qMmgzyzDVlioadehgIxURIWlANHCtNwKLt5HLESbSIUKdHe0wdpj3gWI/zEtbrKkVU+3pJu+BCNTyna2scWcfACMc8Dbp8WpGsjHTOgte/5RY5AyQSf6adBoi1ZtmVMHFhZMWkbYxOlfuxn947sxqbSle5F9AVxHPyfOjXIlissnVaE1X/Z/gpLB4N/zbm4SrT37FlTkhwjK0AnptxsuNOmV2FbuRGLUN6VzUzxiRlQO3iA2LQ8sU4T1JCQG+DtxtWbFqCTFuedNpEPzZQxdut+8WdBmny80n0IU3sxaTqXBilF3swcYW2WHmllfw0Z/0aojKFZQufiVOSy2rujE1zHDjYpTVqvsUU3dvqt53wk7O/TnQX4z2lP/d2oWya8179a0KumcArduQcjaHKWrmdApsBjO/zVd/Jmn9ELw+6QOKL/dwevX8QPAmNGgfvjGCMIYr6aBfawo7kdWPnV9MUQ2l1sKswSZGUadYU2NojSqIdXNufpVJH4FaTZd9tr5ZTEqXOenlGBru2d6Flf8Bc68fafu7/1VrSXEudIr0m7LAHgly9fTiSp0nf+1dZ0Wa6zJNuhTomA+l0n6KbLaTzpsjYpgSGoX4QV1POb6gTt+lYqLGmfgEv3i3LtPNctgwDxhhx3OQKs0gDb/9Gk85+k0uyVkZLBAUify/WykzfxnrqqBdjm1fJT3eFn8oGqUfMT6cibTxTKHDUgCH3KcQSuXzYkIbMQBieCb8xQ4karwUg=
`pragma protect end_data_block
`pragma protect digest_block
8915a0c1f869f7c24242bb5ea7f795da9d631151de8cbec566f50a613241dd54
`pragma protect end_digest_block
`pragma protect end_protected
