`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "b8d8feb7f83b43664169bcb13702adad"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11342)
`pragma protect data_block
iogMa4UxTZWLtUA9GFsRWwZVRXJwgBcRr21YFIsDY/VNn3bOj5hzoNb8Y4QZtC97oRiZ9FdbcJrgIrP2Ck1lQ7XctYLxsWoGD3tCW+6kV68SdUSFVmmLcRTd1t2Uy4BTsGXh43DIuSRyJMs0SqNstDMSbGi7FUJvEOzrDdjA+KmmBDRlMF2YSFI2/LC++NozHjnYInlClHID1bvw4EecfjCX9aI50aGZfpzR0iTMTlWLonREfNQQze8zlqOaRmXF0i7pOMWW3YwrBReyZvYq3KWB8NxR6hDayBZUBcjnykYg8boN/FDhzaYtKWq5jnxmRGeQ0g6s8JrsPPcrd6EbHsZhctSrRgUfG7cvK7vGYk73HXwiuX8koXEesrue/GZLiRAeQ+fb/ovQ9HIsKaZOrofjpqa1SL7kzyxE5Oz/zu9Vg7Zq5jhF2F9in7jD1K0Sr3viiSLZFBnAXT1QUtlIYKuKMxdbWhHK8GoDhIzI/Mf+83cfV9Gb3GVLcOrr7Uy8JtKmIUTDkRh7HY5vd6iMhE+1L9YDF8DZCVdGwcEbIl6Fo4txvk4S/R5iM0L0Byt2q5bvILdNzFOfuh8LlkhHN4NtdVE4djfcs1RcFDqwJ9tfcnXD5HyzGLDY5EchfACtMwm9JijDmNrK7woVuCOglu3h5I8MJ02aZouUL6HDf0f1NxePMLPqMn8l979ysAT/RFZ5Hudv6rHsxJvFnyL6f/EKw1PAjrx5mvqhD8HGK2ymroe5/k3k5MYj5h4Whwj9gIZ+qmLbLX3T5P707OH63jfKM5Z4Fbxh1L43MnODFRDkhLuUeK8+jCgpo6UQcaH6CwbxOypYzVogKPe6EmbGlJDGKfNf4UmnpKJ47s/ds5lYtPk78onnOryz95ndobqcGgTRjQUJvWWt7RyVUeH40pPDp4ra+yIqTSIxBmcWPejmilg5C58VbxlPYu9b0ff3QK2yE0Kd6guGBTDtzbAhCWINbskY48AtNny3KEjwU1uJ3LPa3C3CxH6+QbEfv11mmKl4ba9x3OFhivU5mse5cQplGZ0Zx2dsv6dDp0yfMgNVuzcAbuzA2TGEBhKdsR6aKbIito+cARVLCcBRBzkrKS+nxce5L6sFtcZ++PXXuNuITKqOC4tDfEcf1yqTIRotgGZ0j8M+TRV44/fsI0fC1TMBGqMEvGxzxp+f2M6g5xViu3diBYObSJfnH4qEfA1Hm2zgVna3rZsBXnRzKuG2ugT0/faB4KB6SNjvEinfX6UsNOSYjNByR6h/J8RS5WXJBPJvriR9EcAhFUnrd+YFdCRwEvtQiCkjrAJ0Jo7j65TMhClfkCYxPumAF1i/nRZaaHQufMDsS9AlmAH3QcAnhipE5LwlwQ0i94weDGipqyUf/IsPgEBcJTCnXk+MSdyv1lMt2dJa5RdO3bnM15K1d5DD6b3dMUG2de4tUOt+Ejr3ElRlX1XC8CKKgYRMj+EAgwBYtkrh13FZ8iw8AYkkhbMOVSaao3FG31M5nEszjkXZeeS4jmO9CP3evwe4X345vsMfWh9K8omTgPAtp2M3+0a8px9/SxpAPMA54rQ8S/xHnIHke2l41qBwNGRVn9yxvO4MpFio1sYavoNJvLPeIVhILL6oh6BIL/9/RmWo+hUkNe94NCfbBPgsjJco/HYePtQwpqjmNtJqg5kS8GAJ1MZ93wjS5toMCnSxYD7BjreeNGuYPw8UUo7zgpygDyTGDyblrkVrNH/yi42WJmsKZ/0zg9ToknYwYlOPgfFbFYRSvnqXgwxSF25ydwSyLGyozQtdKCH5SNXtNjRyOkQdnjHJ/MsnMe6y505gr9QY50NeW4xDYT4xz7+4d4SULQRHF5YeHTdMdQz3g2X0KxFKxHWfyUJWOE9m2VGUJlRXTTQTRYUT67oLxVRFiDvMPJ8+aVeUO/S9QJLB4dh5W2tMnFE7s1qXcXxrhzG8QIlkzu4ndUH5OUYM7dQINGFqCvqq1Z5F6RKL9RkZh1+0XVqUguK6Eiefh7Cn/fJQGgPIU6JGcZoj5LLk2KHi7E67IuVcQixdPmjTkmxF9+vuIfhNNH9zrT/u7bAyhAMCHC9dwG7LVddK9yLQ+FVDRnuEKzsBL4OYtM6mGBTFNCaXxuFIoNqZ14XECjMHDzWZH9Nrg14hsMgj9tSem4goiZUTUjvv0/04GkP8eoCBvUZnB2YeARj9ZLTGv99mKvXEUY0t5zc6GD8KxnhGjR/okm3Sa4r12qRufJjfPqLjjXyDSfMRkYpjvhuCLut8i2ANp7fxdmqvqYbWcZYxBQR5FiI9JrIDyWjngjhCDvyx+JHX9OyrHT+80844cz/nzXxpAtF8kJtrXCgM7Gby1vpqEuZ911PuP0rGl7bu2npbgpTraTsLmHefl+pFAZLR54KBHkgYEcxD2vNddgacWwmK4wu3Me+Q5gVBjVU4BUt1Vabz7qlEVZyu5EOIP5q6sR302pqbo45gU0k3OkdUOp3lCJPjKue0HtCUXkKjmjrGJoKKs4X8yGPgCWVsuDshGlohPnbo1E8pukMwWi2BDTV8ayB0qv9gzws6pbym/Dw2uhkXnlrfUcZaTm/xOWlz/Mc4kp1F8SJF9yJ84wYf3FCFHCTqttLnaLXmbpcqFR5xCN1rht5TI0p+/ROj50/yhTZyyVbdQoZkRfod3xFfeZAclq8BODx+jifdCST9pVB7vWRBkO8sk7aXNxshvR52jHsf+8Q5++6Dnia/rzFP18r+YXadfw2vbIsUdBhbhM1ZxCyqcYuIPOq9+r1MSOoGwVKZaYrjuov0LgY6dBMFHRlfeIWL/FPP3ATXRiz1nmAuI64hxhZ4ISXdS7P5xM5Ht8mrALnSbYomukx8moL/uBW5Mv1B2dFhP9wht3GNtlCGcFbHhJHerV6AGQ80HQ0C4KD5KerzdGDAcpLO6/IKjiPbwWcBOvbAKaELcNEdxsQ2KGgJ/SNdtNLjhXryjhvGIUkkqxXLURqOOgnhMSYelHh6mookp6T2Fi8LqiSgifR51BRp6FX6C4X80FgT1B71kdDWPRVyDOFfF+w6mTrQE/ubY+L75kkUsrUawR4LMeTC/5hf1wzazv54vBobcO1If551s+Y11uUsrSOKBsZEM+DECB+K3cCiNpj/IEL9TdOpYxo96kvq5j7uuQEzfX1/Jq6OlP+8xus0dRwv1Bgy64W4AUxZ5IIq5hGl80JaBa2o7P7vgiStruOcfv5+gbkVYB2f+6tabXtLDnwVg763ZkOw6eOfzPJseTzSTyGOi5Mnn7zqV04mWKDrQue0akcifBM7zH657Bi6LOBaO6C78J5hltPoazwy3LOwh5DUc1shlJ4oYBgX2OKuR1CXNgMn5AJpMyd9gaXI5/+S9Vrwy0VyXUtnnC7XguzHoe/ALAPFEKHtalCuUbtYy2R3G1UXjk/Gcx0HnQKKF49N4RM4k+0+npHAuVaUO9UCFDAkxD+Jhc9jIBsZpWf9v96BmVX6Puz4wYoD8qVhGFY5c+UWn4+RoVy0+hv7Zi691eynPRumPulfjE8PVlxmJlyhXHCEdozO+mCjED0TN/mnkOsP4BoWyyLTqGOzusZAhR0N2QimYnQoAuKl6IZ+3tRv5zPuZyQuMK+f8euE2zt8UZoce/XYoz4e1IU80sAqPlWg58MDze8rxOn3vfhja4Yjqyje5iGpIHStspeL8SseFmia26STaEPCH5lPQosRqrvXOFvMYb8X6TApaiL3BJzm/6ff2651cau9hnV0/ajHUMX7l8qw/rPbVT9NvSwohmtlk1ArB4MadhZu6xSxvwv7pO5MHoA4ryCaIQ2T2H1Qz30qj4sDFA8ey/nAjxC7+t1pP8vmQ9JDPSFLFxm3mhiWSAGusWcJqcGDcjIufSIOQsVphVeWHg6nhC1gyB5mvHDlLv8EG+LcAkff/b6ROuUz6EFrqrA3L8w5cj5NHA6+6HZhLCZIbwdsQi5texvl72fWAEKII10pM4hgyQ7OpKIc8WfOG4CJOANwUH66kGkJ68Jdy17y5WTG/ds6GnhqzBg9I42SSortnzOl6QPr8Co78uE/e807aVnRpTwG6zlai2oIZM9Y66EyVQwUvC8UNC7Rqi7Hp8Znd6fcRUOV8m8pttav7BN3qv8L4ECkqesRCXxqZ/VvyDlYmPYPDm5c2yqsFicGYjGPuxUeancwQI6CAcBwcZhka9vrtJuxGzcznkvNfwDnGoluQJ2/W5w/emoewPXNg7/J+qGcpHt/nFwDK1WOyFbFIDD3QmP52AnstitAt3JblauTM+rRmaOuENpy7VwqYlcOI5l8uGUGjhB/w3zefgwFvmXj0gflY/S/9DAn+bB+HQMmjE9MtKipCWWSfKa5ToAekcuUJhdGpsL54v0Ls14tzfLgrVmbdTsT/tdzto0+XLXgEgOtgIQq2pqPvT8CtJ+5Lb5PfOCSRZlxyv/uQ1CsdkeOxRPI4CVEXV8DaCyuaecewlj6DOgPg1pf7AjQ6WIoJHmF/BbB04HuwdhL5fa/lhK84XbmrgT7Yk/vh9uz6sXTXhQRrk2w9p2lCGGon1fo4Y22EW1QPDKMor5PxFBGZZ/ASEwAcXAvRTkDcJHG29tKf05GRfH+giRCeSEDZrqm2H78oT/7yKSfSMXDgYVyzHpB9AFysoQEfzH6eryo+E70Plq297h9fTqQBHc/3XYACOtyfKU/RpuLZt9YCYnR7yQEgVBeciPOxz5a7MC7k9LCvKxiKqyu3a70fc4/DfmFFIvtD3d79V5ml8e8sKrHNXJqo6cfdxiIqOOfM3PS3+B6dqEUjIfVrQUCr1YWJowKwDBFzm0OX4gC17A4fdGqdhi/XY03pKk0th69lQRXfAG5AcFjIFDhrySGpWvL53OUCo7HnGPEfeS6XYXlYnYQ9QXE2taZ+FANbuPYJ6A+sLqGJ04m5zKjqx7znHUICpSvT//O/c75v75Az6H0SpGyIr3kidzB4vAGRjzRfXGSQkFd8J4kAHNUlSa45L0sD+t1glCeuq583zuiNOZkTthF0DATFupCbJMfgoVOG1alKJjh4hmcKgkumEoQPRwU1DFcm/QqdLyb3cxRLrsy17uejlmmTEOceRgx/GVmBFeGzieLzjdMubXvSczU5RZVF29UViV2BGUFxGVPrjw91E47Ozeg1rXKxEpTIoBLbGX9PMXNx1zeOA3dOnSJ37mhzMtYlM7/p4hh9fZ2kH4k02Gy4rPkVSyz0muSPbNXW4EnsBjFRkKQE5G0PvvhZgwsrCBZoihNya2PnwXmY7gmiylBv3pyJHe+qBxM7qmGRlzmEDthoY+WaT6Mm6Ujr2kweJaPFwqSz8ha3gngVqJ2yjfMVYQnLBSx5d/pzdfVik9pLiyDT8gkRfJGSffYBHgKWDwjJwF/6Tz9s8R0jzS0gJSu3uddwW/+b22DsDv2v1KvOX8sD8VamtS19iQdhJ/VFZx8nS09sEyzjJs3cYGaNNTnsT8hKV6ZQfpTF8VgtEw+VwboI/LjRZeZcIAcjI9iDbn9Iy8e6ESanfwgipTJfCf6uVYVX46flZqy/72BtV9zz8kk2rjJdFLLkJir6sK56Ane2M4KrPG7yN5Ya40RaOMTl+QeqSRWF/9yiKtwurEknaBRCRUIZpQV/g9X1syGksl3sQ8xd73838VDdbcblr1zDXTuS7lKdx+CZ0kspiqntpqsZUAYJgOSY7g5Rwzt9FisohLEo6rWefaslzQ6KsyEyOPMNO9IxusyS8TOHrj6W2y2WyFoHxNyvPEXwVhHSePpvbNUmrh+IlkIwRqJroNGW24EYWwyIF+mQObFx12ME+dxSoDWhFIZKCAU7xBsjGpd885KftJHtp4jyrflkBUx8CQ9TW9Z/dI8BFcasZ3iwaYRmVU2T8bpbtJ/Rtt9lVZ10tvb0m4uRcAVACNGs4m70SDVAFA3itbJD9MSrn9DtznoEg2sptR6T9INjzpKnoXDrNViC43r/zFQw0rihiLsHuE0DJpAL3znHcIa7XSk4d4y/OAQ2+5aoAuuCJP8ylysLusvpBVeG0LibEoZErCJV/9aMpTV+kWIiK9/EbADT3NAUVFydK9lPOglbqu0HP2ax0MpqjeS6uiapH6+FpTO7G904gRbnF4Dhr+xOmZ7CMLEXPR62MeoaKBAYw9eV4HxSJJ2+ycaafZeYkQQjbRL/BZbd2z5cua/rWOvRVbKSEV8iyl5NFQfi06+fGgn1qEEVCNsY7yb1VqdjNiyh1wkDB5Ck5lwwtmX1jejJ8fYOZVO+NK9CquJWgTWWW6yWmgXgmuss8QNx2q14TlblOxmdno4yBe6uLftx1t++kOoFN+DRV8kxnW5FvpGqBHyj/crl01H5mYTwzx5x1uw0MOj9hLf+eTWUM35W/HBc0NYp0nVN+0acOs5V52D2z1joGcKkQNnW6sKtV7oWfcXaxnahO3HueddDbaLWPSd0p22Scq3Pq4UnISEUKjW5y9z2vFJunvkDgYX7ioQRZtibRen/4ULP594ogs1e2EOeugA/ZCzjDyKu/otjAq9d48/JXnDKWB15Ax2sG7EIFKriQGMX9EfEfxVwWYQseJa46sMuaZvbWPug+/mXk+It+rQJEO699+u0JzJQJz9ri4uLTRIAtRcxVJgcRL7Qy8CqvZQU7buOCTHqIPTCLIPqyWtCLd3YT4FOFl1dXgcZIQY4pjmEqH4zcnB2Z6+tMtSMn926gFLS5b0QpbGg5X1irwHJlVYdwJCnYuKBuDYQCstDO2uG4Ggoix4F8Y16TjxYIdMLWh31rsz7QB7yHEiPCCgs7Yut5FqP4Lh106SxDxcg3Ow84+05QVjqgrZS6klyG8PAcClEHZfyOoBE6UOB5F7vJ1OJuOS3I9XWBf/RI6gkw9B/uS+Nxg7OxijLYRHAnOs6qRzlSoaubU8n0vbuaRFnPn+o7sN+tTCE0TT6GUi/PV8rfk1ncws1QlK3IXPBpXmc6cVTKzCnc+dzATCVMv/o8Ty7FRLMc2qAIyeSh1POMZDYb831mNFIkE1K5jeM4FppTWbmtrvozHUuZLrPa1O6uUb4tW75J6mIe7n1uIMZTjpzWLVENncy2TdH8tlpl9Bad4uvlZuWh7JyJZLxYMzSKdV7QDq3YbYX57TyD3xX6RG8RsqQ/UUog0cchpFdA/z2QjflzrKVsGMOug4+7mOOGc+/nIF3S6qU/2K0shFKv82brXMpH8Fk2gYaT81PhEQhFsC9ASUwEqdbpIZjU0ZTKWnYjLbZbQ/JmysAOIuZWC4urlOeLjpk1lroe3eMWDAfghk9Kevf5WecYeNcGDnXbJBc7UqWOVTXQ95MNk7eUh5iYGNpds+lLxSlUpjKZZe7HvQXHm8cL4Y6iOv+qrlrk8oO7dPLsi1jJR+OlGYGQ+PgKHorlYoJ71/2ypr8Db291FX/V5Ca4ekc2ZA6LZZlXmSnbdxsb3QrnYeLsvHLoFw+VDRw2OOT2yjDzJAxarh26bL8Ng2NgP1vIg75r4srd9SNg3KaeOQD/BZT+UblekiM/xM8EXiM689Og4pNFi9rmDKUHOAMw8bfjRnoUH/xNzSkHw4snrdD3vd5hoegVdu+dp8moFX0KxEBXNTHth4qTId2jRDtjzc5UWlJQL4+A7pFRZQfI+56rhn8xE834Ij771cobJqMFb8BbfeRCOoISxAFbt29wRGGH2G2pyIzAVzZ9peOOTA8QCmCuh0dazzUZXaqBPpMN6TsU8boT7Lmx1nE0p5yck0fBBWJfLFA3MVxjRCggp2ZaE/PqXFzVLOwtgoHOloryGEU0YesN0zh8Q24pyyNREMgRh1BDEj5S7hSFx4n0du7UeR6vRtsX1H2bkDmsW+3vQeIoiHaAahJHiWRamyrrpD34SH5mW4T4LRrGy6OlofQQBtJHwSsleuE/elUp1GX9gMR1pdrA6maWsWSmqqqZ66n+fhQ0Y7qkoQPkb8fOZKkwNWNgturrt2PUr9e9vOJmc7RfTqMwvg1PgYQA3drfM3+u0CXe4Cy/Ypime336mjMjIJP2ewobDXINRiyzB/TGLr/B5xJuCkk9VwXekB6gRfuO+8cZF3E8uP6EhnCwHSRE4x2QCsg7e+Db/HuY270Bkm/t37R9PVSiJ0OCv52B20W/0CTokMRQBKE6rEvWv0KVed19/ew1IzXCnYEbCvpEKt5Q+KFTJ7636qwxZPD3rgC9Q65WFsptcw+xRQ3vC40xGx/OCkuEMBFgtxxXXckV66bqroXK4QaVkWlHCAutN6efjwRLllVx7QYKX1tGzXuuUFYlaFdGsqfCFfnPGpYzRz593OXePBWZyGCdA3BMD/WUB5ebxEy9jJdmcEViEMdKFgnDqHs+IpOkq7EsoZyJ/9iNbPxJA59RkWpuAYgdhptd8KKaBc9nS6uQr83lm+f66AasUdh3/rxZ6re12dUWGFK1+VRU5k/hnsrIxTTPWMsIswCmt9AC5bytJpQCHsvqiPWt8GG/HQRtHopwMx0FmcI3rutnwkeBgnRA82ftwmLa9mww1eGDosutptNRLnuMsFVRAwzgheDfsXfUA+hGqJbiw2UaEB3g+xfUOjY8k9fEIWkZZTXuj96pb8cHgZiEszIcXYHEAb9ekimO+HEEFDgJVemRLCA9/kzKWdt2zXDs/L+LUFDaVWcBA19rZOVR3dCGqDifvubJ8U+m7j0wPB60/IFFJguL2EQvtGVt+4/xSeVuXyRSz+O2zNI0Hedur8Q64TREFBGJoZZzi2lBIRQGrzkm2knu+wXBUxOEF9yaMrcOkTrdMHqyM3nNrH8V3En9QE/AvKuLfAACTc8/22aYVNKURhvrLCuBlvVPUGlbeH23N4lksz/T1vFNs7Vl/7XQ7wdkf7cSXDaFLEnJmB/Bm/FRkpINvBEgWLgZGIvQF6OfLJuGaSDjfv9K8JCvbr4/s3eeZWVVjCQpQ7Tz+qZF5EE1HLl0W/mFgGMK1IOSA6b8w9VNh1DCjE3KFzuBElrK+XNASAecUGwjCNA5e+m7Z8JLnBCK/OnDhaVSh8LS3SnBTWixqaPiQspZyq8DOWGajauu8fhzppsMIufN3R4FXfHIMah1SACwOXK/M/NSgo5/evbBaJXYUXUVn2UWyjE7z3MkXMQi5uWh7XWDp6rFQ+hw++aXB22EdQEqQMM3CZDGUn3pQKqvZ8kj5lIg6oGwzkHBxf25+MdIhMTY8EsfvOR25FdIsi5L3yDoPRimhSapr4DL9h/VnxvxKSy6M7vsGG8dFhgKqPWC/FEHRx3NeHai369Az+OLtlU4+cE55gf01ytI4BARJawBVIlmffiTCEeSl4Z4TJ+ItToC6s4jdxDBx5OmpE2db8nhpqk6z/dbKhrIPYeftbBVVQ21ndHvT4Of3Uc3kNPwGmWoOI6dDaAOw3ARJZD+mJkRa5ljBW8J405hyqabR2TEUs9FoaVVXjZgeRNxRxkQrAhYu8JST8mF35r+TEItN1WQxU/u1FgGmlJ35LV1kfbffk7suWod5IyQAFiKoG+4bElkK0FguPEAc2WwLi1elZRcqCz1Sqjga1hT25m37nxmu1U1Uiw9amg3EQihhMYrsgWepk7sFhyKJXOhSSVM7eMWwZ4tcJzXY6j0GZ+TxT9+rIm55sx6b9UZ5FA1HL/vHLU5XwGq+KaH8v0O/VXG/vR0H87SEEn++/IMoeYJjkgC868kfEF/vN+cgE7IG73uB2Xs5+B0feyhQh30ylHOoCn9c5smS0S4/9msP31zkgjLvJbrjt35iFDz3irM++LLvT3n/4xoSDYbFXndfkoIK2YSSb7/xLg2F4lUPl2uoxXGAsiPbXWSlZugV0s8813Oa5GUa+qTc9PF9OUmUyLQMNrJQM9Z0nuQ+sYuL3HKtef+TFGgaH6oZ3Zqctuyd4rDhx4lkhn47xYF8CojMPfUZtAzFj8Vc3tD4HDGW2L/utQuPeB2nhJ4PpW7CZSEufwmvL7Qq8ZffMvijUmojzNWjUQQiRQgv8q8T51WKTXOszNqitWKrGqKwOrGtuf45BJJ/xoRBMPIHmSoAf2gfTE2tYh+ktil4igk+Arbdiddmm8ZYnXp15vJVafi+3kW1pxTPIfzUjBMsws8F6A6pbztjzR2/zhJNggrh5U26sigLH1rw4lOZMmesTgOTHxzPqjIdTKAnajcEWPrASiyWeMdDguuqlethDzYOCijk6DsOVJFtiB1KI6W3/kcFwwjJjWOWCT7RbacRmuqPNcIg8Z2Ij1CdbK/K8PUeIAhpxWxZRjoZu6j3/ENcck6/eJrNheFLK9COZm9+MvXpTTOGKRD57GOZFXleWpS7+jlpfemz5rr4CLJA/AUSgrMyUef+n1v63aZCM73QHqJhHBEPXOGqKjKbh/DuLThtK4HOQQ2gn8iOm3WYEXyMWwRu19EXx+2t3R6EHWJL3V30jDVgm6qb0GO4+HHag63eHNKH1iZmDqCSsQ1N5jLOfCBjvVw587DwssZNavpHpZWYs25z6Eovk6/gVzDXEFJtUWX6ZM1+tfP9SO4aVjPtwqJ2uIqg83AzYAAu3lh+FqLvxR4L9CNfCTWkEBi2X9CA3V297lUWx6AZEkM85dPLI0VPsabthexopG8Oju9ArrbYvQ4VvsgqKTH4r7IdwKB2xfTceo6ZH5RMQv3pT9vrrSXgTTIs61HPt5DCh36CPnxUwAXrCA44mkoHWvhcLlj6lw+rbRLaaNXOx+1NfjP3IxmvdF4lhNus0i+qa1Hl5ndOKD+Yy5wX2WtdTVlruzE9goln6V+h5El2s9z1763spyksB0TT7NsE+CGYRs3JV5Pm+f8Jn893VFUlqA4j0Yp32mdcHZQi2xjySBvH2YuOaA7xw3HwgCYEtSwAi9X79NqFVrfR7CEu34hJwv9bG2Peevpsua9vc/05LfrMZJNEN41suhrvMX7mU/ufeRZ4nnFWnDRrQ9qKdFuJPz/ADjv8w1JZkGIFAJGaw6VVWJNCqSllJuVnbIhIduoVxXLI3o2zmbFbh91t57D8xFBJxn2yXsSBQ7lRmpjxxO42ueYTwxX1WkCoYcumXOvCUmzychp6iSWhd/kEPslSzSUOO2mUzxU8PCA2hBgbpIdFAY+xEvzjWcs73NUd4RX1l54cm8Lyz6CCfXyktojKc0Es3mmHLceje6WPa3e0bXsJcYKhV8FUYvgLMwkJgC/ezPgoE5IIvCu1vL8reiLfSNk/xJX/XQwRmkFiDwj4hLbVf88pkJul3ZPx3t8j3UjeDnwJaEq3WI7xVl/8cd5m52ekv93ljtiexQJYz8JMhAq6N+WFosdAwFAh/PFB/B/kSbRw8HxD8vUK3jjmXLmeMLnyiHgSvFia0tSWE/6fxeFPcTvUAcZJBRdZcQsUoRb4Z2wL377WimtOuBllOrULwWndM/3DJAjANwJpj7mjFs9+HUWsUKIed/bU+6Sph5aprkSbzYUCAnc9p65BV0l9CTmkRyYOAN39MNhdAgPEFXbEg16qn8CVuMFTYs4UHCL8ZdLF3zRymT3tout3e1GEeVy2/h17rX6zFpZSL8KwxGUcgxPQxoiiu66oynsw4CLf/+uPfC/r7I49qETwmynHulHAZAJLATkFOyC+UnIiACE7yvsfMyXPrcDg4nx/4E6I2FFlIonM3IXh3i+bo5sfvYcnH9ah8n0iqWOCdppjwgNpkDTDR4L7AhXFXrgedHuFDxY1b4t8wvI2Hse6xZio0/FJioBQiRQoJaBv6WdtEWezzY5HUmHog671IjY7nmyxVQ1IPvQ+48gETPD6fRDFQBQJvtmgGxVKOdxbQDAsPLMbhxUrS2+L1e3imhWuyhruTqnT4pU0jPyIMIfUfjIDyrr5+zeSqypVS2WLbic3GCGvmAtLTZuiCqU4tFksa2FkOQhTHOQtuqnc8qcNl68mdqJkiXUGQIeeYRhzr2Y/4ac2LpOh5TDpp8aNxFwlCGL1ovScruMgePRsOiwCh+fCtGNrUxF1cLdvd5kyDeqBjo16hravuiF05eprn6TW4AmZX3Rioro2JVSnIgPpSHXzd8DWyRQmlEGqJlDZB/82i+khwOpdD9Vrqj+pYGP4LIK0F4+ldVy+jwZxnWfr74pvwtAWj3AMAHOM4zilrLvsP2sWowrI7UrnAmJe28yHdCdWl6Gx2yTdzBXkCn08rBuudaqPAq/VGmJ5R98QWmevprEzXioeVVF6HKi1d8HmaG8o8LYk5SNiy6G+qB0I96iYrgeeX0YkgIsFoynkrRl8Y9aH9edRwnjYD3nizPEgFRBXLEQYXmtFQBgBZQ35ewXTs9jki5YFqYCDCVmLt4nP2gg2RfxHcq716dxho9jVBQQR6m5SJ2Hacz9hPHd0SoGj2tr1KV2uWaDr7GDXm5WyIUpg2MCcYLT3X1ndAwpg9hrrjvqstTXJoo4b+BFacStZJERYttx8rFTs3gZeW8QuMsUiAqXSSAv3AiLnxmqcvfkgs8h5BAgoGO5ziUd2jEmS01IF84fH+YK3/LQYt965ghxxCIfnTh3rzxFS/3hNXKFGua0RIKO87HXuUPf0Ni3y0Nz1ftivfg1G+232mZJzOls7ackcaQg1NPop3D+Whu08o0jMS5VACclxcXQqWE2Dc0bN6CSz13isRWTnBrfWurBL1c+s7yL4+hhou3Kby1wAtrTjNgYAhu7j4K99aRgiBpAKlFoGGftVPXyu2L0uDuLFtG1vnxtRgXmMWITFrZ8j42qoCpd4/O41RYl4eSCaeT2KDMoJS7H6GD8LRUiZeenGWJdkEsfm/pPUs+uubRAk6Bt6O8cKCqeetSQKjOQ7A6/XbvKM8gIVtwDdxEx5q7E7V93bDwUJop3XeWLNy94LnmZ8UK81LTn/kz6GlKfmRDu08jGgKRL5DRGTUzvmkTM7fvJZRdEto+GVjPzmdd3Tg4hkNXJAqhP9s6+p4aGMdQf4dOVJnYp46+glin9QzDwBpo1gNOIsjORkViKxsU8qiAEumFuaVBSAh5ALFBs58W3iYiomEWFh3KgVzeMcQMwqSOqDDcwDiPGqqeismoj2Thobaa8aKD1R/nhiOnow9tPPb79IfZ6iaqocDVkTYtkPVyq4sLVOloJ1tfiPbmYY//FMqG2a8oVYHnCY5HbLiJQ3BBmPopi4pMND1yPwn6hxI9F9TuusGdgFWwjTK7YoynrUXI07g6m2YtswKOMLpPVFA9WjwB28ws2h2C4Xxhd0uoPFUiBepGP3DxdmMK+wiixuKtVFxDRW6QN/3qHLnV1/3MjuZ5zu/vb+GJqjLE1KDu5Jj/f7L1CyoDnnwVZ9+rbjnuIrnfb+BSE/9VwhsBwozZeL6r96rFnN2vPCopfnMcgXxMfOdJqHVhjJZnLS40daU5t0BDD2J2KMDzGC/OQhDlyU3PCsJxxv3p/nsmtq0CI+tZLD1XoFlsazjeUn4WIpG+b7JMca+WoFqnScMBHvUucnP7GQVzrjsryo16GIwo2CH++yuu3SR1G/m6NXGm44sYtd3pXEHh5GzGEic3OYYou5Jn3UDcdeaNwDazIIGPHZhaISij5iAOWITvPyq0VkvQi0kLCpmh68LH/6KZpPs9/9hjWbx3OICRu8N0Vpi3h0X3e6FBFyUvJRYlrmsYRK7o7/Nk8esw3s6w3hwB23VmXbX6QH1Jqx9YASbu/LkgtSZJwOgz7UfSkUnvyuWYBm2BY/lIRJ3GbUwFy5J1oRzP/o14INxnpPpFFM6MEcnPnJvSH/ncDIYiVUgrrufqGnjAlj62j+NEs5Hz3CihCj/Kn4jWjjlXM9Yx+kO5FSHJsKiC2D0fnlk1MTCNAu7kGHIMpRHr/DXKEqK64rZmxQiseMbNEBGcedOtkbVzkz3zvdrO4NJLw6bD8L5ueJVeIBfolSUMY85WnAAEePCjHPxlOj+PKedGqY+WSqPlC4mlb0zWQpMHPNMnxU0dp2hflaw9IBQuFwNrs7x5IM7WRsCllazSVMT4yeSKbDJyxjp1Ue7yFPxzJwWchI5PKOdO3jMLAU6iUPnMO05u83b0cGsW0b5srnUB8bRkih6MiMYIoW76F3s/QQJXp3XooRNEtfCZmzmqX2S+ItVDbgQk+2C54yzE+n77/DEJeWvQEPIvITgTBBQOr+JyeermjZYmx8MUSQD+NKYWq7XErHX6aq5gpF1ccYksR2lQXZCCyUllpb+pFWOHvO2E655ADvagtK6Dc/jz4SGwkg13G0dVP8O3lbypG1TpFXX3AoWDkHfAHDr9Vo3pSJlzNg0ZqnQCm5+xT9I7rrRCA1wsR2JqTo4GEBIpdH8RjRWokZAu2j2jaFkCLRX1QzRPDS7MdooGtweeGgnP6TZA8OWvbTF+IVpW6NtGWZdka0goeM9SwCEa/9oUUusVJpA4F+1LeCy1vw75GTq13wjOhoi6P1CxrnlxSDe98gEedK88trDyUWmXFip/rqviIlr6CSgtWL9IocZtsI6Cm4m2eK5X/fOm4NDpnzHnxgS+NqVLssbx0UnCoyXFGAQyzg64jDrw/MbirVoOrvyBnU3SSwVSavdgCCfmEVorbtL5q+hCxNq/CC6hv2LBNUOKsOuRDJo42ubKXfVIK3tzIYl3MfFL8ncoxgB3Jzp+1lfl08TQJITJeRNs6s2Nre6tUFpQQJ0X+sGIyEcTOF5zCOtqvYnYU9E/peRRN9m8UtdgbqwR1Irg4Zr5yJ0iJbe4bNn0wyF1DKkh7uTzxQdXEvAM2EX0kqQ9EdOQNtWlpMwsuFyWNlWwjezPI+IchR+Zv5YWzyv/GhNHUfZ579Pqgzs9nBiRfKrg+SCOhFakL+mgJpFuW97gAFBV8BL3OCVq44TrWTHC0z4xLBKHQCyy2DSuHR7wqHzbSj8hevitxgZSIPZ7LhgDg1SrIy/Z/bCzBB39xFc3MAnjrZvgiKnjbFwFwzDN40lXuSm7L2xIigiS2awpwTmWup4KL1kewQy/nPRb9XSbTouTg0F1mZsDYoxn/9MPUYiurG29Q1g0jfR6LcJyMtCnpPhkqezjfv74Zl+sRahY0pVIf2x56Viv5aoHn0lgPIPqCUE+wDNWGIG8+gHkQ+UrcyKd2Zs/2cLyNXmdD5YDassXs+kZ6DIYjw/+z475nsql4n7ZdBxy8hwtdj2mA==
`pragma protect end_data_block
`pragma protect digest_block
305bd5a4999908c02ef4066d054e179da2c93b79b7c80aded900271834041100
`pragma protect end_digest_block
`pragma protect end_protected
