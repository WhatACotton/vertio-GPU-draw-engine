`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30131)
`pragma protect data_block
u9Rip3PRdaOpurULAv3i5EqH5aWB4pfryBdvF4AUlFfe2YQ8fvc3pIclrtDH/iruw1qvSQ7d3hPXkLO5KX65hjOdu9tXsnE5ME9yTQSUqdaQM8lzy2qN+AaAKsM3BbOct9XDouHCWZsgGioN2SjdVChCxNSOcqhNBLJtklG/tGkh1pYKDSx0gefXfasqbn2NRgrAvOZYUPfVh0cnmH0ZSEAnm1wP6GC2X+vM0fQoL9WwR5WMJD75zbl1pKBYI+GcjSDdYpYpwvIZCco7Y8Ija7cwdKiZsl8rmmOjTBlmgfSNzcUV0QdeCO4tNsoFUJL/Yj0jh16X6V4L1H3FcN7+GueSutYJNobMK7NLEsYN90Q0P5YS+3vLGnMGHUjb4IqsPWK5QFBdQcCOaj0IuNSDiBwOmxuTjw0fmGClwYsOSzXCad/6ySe/sGHRIdxE4pHzdSx0WSxBp1Ni5ixodWe7Hz4x22VLd/iFw4dZC0WF3DdStl5pP3lBplnd/18su+OwA/tjPKe8fYFGSJ89tC+bJQMf2jwQ96yr3ecAVL8CMA7ygwZE34kdiuXjTiiWBG/xnaXoT0B+HC1pOpw+YMvevUQFVI8FAFt83+LBgKHNowEn9vZks9pYIw90Bn21QkkZucMbzfGytIH2QQqaPPKwfUuTdsgiv0oZrBuj6nS8bIMKnnYCerJApTZjo+4cDK7nYBBgpO2xBDfsvvfZXoa7tFfGmvyonMnUhaD7aBx/4NUY5UbR7HLzseHF/N2bnMpwBpFeKosGMod5DJcGYIUH3Zxbr5Gu3BbR89w5CttVNsLct0P/6Vyy1ntV6WGjmCyjp+pl55xTjnpNEsVH0qMQtnlwpOiF/DPl7m5Cv+ZjzF4SFYGKLtBXZUamWz+0f+RIRBKOssnKgHdRcfO95F7CMaJneW6iRvU37QoRWtDYLE3sB+38Z1hpOzis34anJntPHLc5G8gH1ej+Tf6H5BIrUXSepxv3ZflS06Qh4WYDThn1utm2feRlM8NKRLlBmIp7mDmWP+vz5nAFlTwlKgr7OlnDzJsOmMPNbF4W7/S8KBzmJ9PibmOIiMAWxix5/VrfzC9Yzw2414QkhNhqZdjqlrAZntYZqif1JyNNtlR1vTx76k5vNeM1td3NNEzqQijZqq403zYA8jyqz+5eAvtypLg4lCIOopI4+TFitWaTqoCAbjtcaIOe+7TL5q6V/fy0KwJjJcqGtN0JWa4dLE4bE5VGrQL75a+QqElwpk+iLMmONSZnLhVoPXhqvsZ5BevHHExBttnw2nz6ZzTqrhnHPuHPNH6ulfQxPuEmuBPqohIjh0ylOQJwKAPRf6LIKF0v56T82nZyxELya25y//HPW4UUIUqEeVktnBg9cJU/HWEy/etnvkhsrYH1OauFnJyCkBTGosDfXOKdU4u8xLRZc1RFYM+YuOryTR5aegbxeQxW/ZRAP2c4sv0iN3YNm4Gew+gVNRTXas6R+iM5bbIhs3O+3/J3OyuJ4HO2n+vPMvtsmf67DmlXg0gDij1l3jSAMTobotG8Q7RdlJVh5E46vLOobM5yMSicXGhM3xc3zn3wF8dpEdGSydwHDEdHU2/vjVPV1+FxSJL+RJXOD3vvHJqBX1Gd0dGW8eHcwwdtXPyorFTid7/oFJGthepKvtoVKW4zTJE/lcjWBVHZPpCyi19zYiqFgXRYOdIOFhEK8raB5J9jBDXZRVg2LgJQncUoxl+JXgELgNBOrz48/GdI4cAn9JMmtO/oQVqvBaFO8MIl1hZz+QCmSkB0Jw6eGrpQjjrKz7Z4JC0hVPJZeWDVQc3FQBWtI1NRPWKVzisBvjBJQr97qmxMZ9eLfxeiuw6BVfLdjfVwI/LX+mI+eSXgloyTamEdbzdUU3h/LNrUsKa+hQbmC6zQ4ZW4ApMQNC/R00oEWaItqNFsxcWoEuYVeLIaR+XJzQFlSVy9Chf5MvdjONK9F/8URef1I5diX7MOVWZrzUXeIbqk5TkKaxQW2c3ymownhKIovjPnUNW2jfTV1V6jFiLpkwdci+p5ofliAvf6i/8nu1DLOXcAdnt87pZw3GQmkUfEl84Vvk4RVc65NNh+PHZ1fZW9FU3TASpRgF2wG5FUqmPv3ccI9k08D89NpixTWyvz++i47pOu2OgmdzUuE40buG457Z9COLpS+cWwRevaLwyfuko26K4yBCxEiU+nPq3akYmR4yupYu8bwQ05V6PrROkWyBjxTS+ZCkKRXLwCxtQnnHVitW4kD4JU8Ak5L+JN3tS+RMRjULpzgVuqpSKkm1Cr995HU9Y8gYsio4C8ImXmpEY7EErCeYI+HqNFpioDtK0qFrd20MfnMpIY4I4ycXpfyNpdtKeD5V9K03+wU3Cqx2bXNTkpwaaY3FoQ1+5FdPVDub4ZddfEw94x4Q1TMi44w1glGS292auvJS7mz/BodhGw2GkB3K3Tzok/EE3BMd21z7BjrHwuWstcRZlbfyf20ZCcDgdGXuxW4O6VASoxtIeBBsbzGPf6qrShligHxhBlqCSAHbQigNZ8aIyjriWABRKZBiqW5drqFgfaqh1koQXjX6xrUOX6Y4qgF/hdmRFHJy9YGdE1s1weZcRItlfXOr5tQkVWoJnNSVfrEuNhjGkpXbec4Z+KsIP0Vq+V3A9Y4K90flqR96hZ6XB2Y3iOxiy9wmB+vkn64s2wvG9jzSzBjSaEZAHLZykZs5plVvWGF58op4ZO0izoKtURHEVAS30EiDWkqpTS9Uoi9dcTTaJUz5fi17aLIXqfzUSrGHM/i5KhX8Kiqi1VBi52L36S/WQFMZ0JoSEJxuObhF2IMZfDmL7RdTX42st3MOLQizYw9ivScBxNlHnsCKnp9Bn4vci2QPJubtgJWVi0A1C86JXscqbZUFRoTIqkT0lA3Wu9j6tKEXjkL/6dASW1sKCpBJK9Xc9QAmEni93FEF2xnB4kp+Xn7Q01f10fFUz54OXNPLGrn88H4H1tUCqzh3v93I+C5G8IxTQ36EGuRdOjJbTYlFfVj/3RzHmcvsJiej97NiYXXsU0YyEa0tUqnOwqS55mCn95fbmjxD68nw47P/dRo85zOHVxF99I4vrrmOSuAXi56F7CoCYZATbXBrj3lt5X0opGwwU2xz/ZygxHEaRUMR1KT6VezUgsAZQXj7I4JCnBUzv4ibDoRPckfzk5Qjz/EKmwkvqQe/L46dRecQyYvWcp/+6Pm8GJg2+faVc5OwbGY9Aej8LNl7993o07+KV+EvDGTpa5Xdk+ydQ4ZUUk6z+JxtvnZC7nxWRNSgEzua/iazIKg5EmNVYoY1/6y5T3bioakWuu6rFgNt0xPGXrs8FoCUCccvSo+CLe/WszVlObQr6EsGckyFfCI0oA0BL5PxBGP+LlxJi0GiBBhjeiD6W0R0I2BZWj99SRl4z9XzKSGpsr/b+M9ETKLqtTNtPyE2gY0Ig/5ckLiH6+TKy4De9BQxUxIYMVwxgoIFhMHMJ2cMrEMVLT7py8kEoivEAfiT5ChMn0k1BC9gFkSUIvEYLPLpPGncbHyIRz4SmsoEQFld5OFSLWXLbzSvyfJ40niku30XZhIuYMcA0DyYA5jZ2jYE0APKkU8tSqFzxT1/wm0XgDiKLurj1xOBiK3dlnEsiH1J07IxeUgfVVf6nArmHnenuoFt4fXWQlJJMHs5qA+kOj/nRm62oyiahoLlEC0VAt2p4mpfOMnGeOJqQuC5fmQkDjqkTQbcBA9iGaI7DFvYwH7E4jPkJnR/ivABRe4Cmguyi7RrYbBMm2bdA6rCgO5wnoj8XpPYNMH1VWepcTe+vNR7yKF+s+He5026EP1q1UJer/83FkQXWbf8+cK4BT57usNs+1mHK1XDrEjQSBC3iY1h0hOBmOVFqFE4CQ5rwwUFxpmKdJ+ERLxigi8RzH9jJnoavT9053tU5tZC5vX+OgTDnHXusnohf8ldeqNe/F72+G+//eNUCsMhPdESIQEUGEJfcnNMFkPY3CQKY7m1d+v/GMXbGVYv+fQcI6KML4fnkCS8PrLisk74q1sHVkNF9AtIa0p6NQFNf92iciwb8K54rYPYV5CcIXWNIp6IA7k7ovsD75xyOtq5DNGKzoflhj5/7qJLZLn/YlNaMX+sZrae2+eCOGGRc5e2vgfKmW1H/S2hq2XjZt+YPMBf+mqohGE8/91QYvmiP5+8zcwM7MF6rwdvqP5WyUppdqMBylyiOIWhdL+7w9GuX6wgLg4sTRXMObvJiionP6TjH9PDCObDsek5k5JFccXjJCSJDxAdGUNWbzOVLea9fdk0cNjwS0EA7buGhG07uHiCbO7frHrOEdol2i5iqtuYSIm5aYC5dlzDRRxONA/VaZ8zbLpywbd8IzmSXTNBM/7+zI/AGCajOYD6zgbyaksYxTJNzn7YaST3C+OTBRiLMXhRFIM2gtvfWZgeF6P7AbbqxKxjefBzlAm4H59WJ+pqnReojFTH4CU1FHhDQfh/mM/DyXglFABGs7phFp8z0ZiqUzUDPabnNDYBg0KpR1n5Fq8YXSF/2qh8DEPXk92oHj9PisulvEyMY9OYhxW9gMMen3kvNSYT1GWcSravigGksXilKu9zmKfud+eRj2AkKKci1wSAsIDOuVjx5ZalAKrv743OdnTTTmwvx23tVkouKmkSwsYpG4G0tl5ISVQewYAORpqvLmvShUP5XwnigsHF2sqJ0TSKJFngzpQCChhGogLAIKIw17+/onrwW/xbzFLC1Zz7BKxlG2Epv1wxlv9QWju3SCis0Af2eHEkkEymQau8DApBbz9CPs3sogoVe5uMUFj0iZCxuZcdSXqchH2I2PpV8bKK5/TK/ZOJXUKn0KfakWYjbE8ew+CuFZegKcHilUt9xj8LKlvfJ4uJE1xH0C70te+wh0fH9Bhr6DqolPtgpc5Bgn1LcXW/vfAKNU9o212S2hXDLjZwFwryOP4N5W/fMun+YFCgGx0ggstl5okqr/b5HlWgDNkdz1yx5x3fxw1oIJ2MLHIOjkXzhnNp9c2kWH0lgcnc/JrG8QxmkuvWXJrURN1IrgmWDaqZqyr9OhJolUv2T88J837OwS+k0H0lYgy03+KPY7/nJpQQcPgaB3WNaOb6AYUvofjUb+15ybXu0hthWYcaF9z1xZMyBytSfbxy192waKveViy6ne7HM6QHNkxd50Ooyt7nIkW3BwXZffHwSa9GpkLri+F6ciVwLwo1jVmgif/QuSgpzF6vWLNPJ/ErRWo6IuzafV/9YhL9RSjm7MnixEtPpVT8MZy4Nnte7KPdBlZ7mlfm4B5X/mdh6ydl6N8K2rmFaXSsbYq5MZ1sghStd7fD1qGDWcX7F1mDB83sgnCd3rGt8OvgAsftWvH25jR9b27F7kPQCS+8Ay/HsyKT201wjFJtK++wWVRnsZg/Lxr093VJnGC/lNOmDWJ71ZsbdngZaHllfKjE5QGbSjLzGd/S2bMKH0j1KeK2wKyec57jwUJVxCNRRCZgQ5Bmr5RK4Wr+2q87h0+LANT8Ftjht4dOlaXhm6JUcIPb8setMtkZI8Do1NihT97a9fwxUApj1IcnHbO2TakiKqNoChwSS19sFkKba+9F3MIQUayQ4FWWHCMubudPYHjfoqX+zLx1zV578WxNbi6D+9V8yzYsUWRxfSJsG/y39rXFBTrbxomeD4apWMYjrxVjibtt8GACo23B+61w1a3bidppUXEEkQZURV1o+K1OvGPZceKzUpeiOXOh0Vj42O2i5sEEKp4QkD5l3LN9g20ZDKz1X5+DaJKyQX+0zKG0vN+wH5IJj0V5MTJXiMV++0ml9bDTEbkJp+ib0+llhLjyMPY1QSq4yj5Qwkm1DFCmazYO9Yb6GRpT2C7bfK0JNMYymkUzu+hRyiyYwb2dW2IhR2BFdBS+Dy+fMPaCSKpowdhO5Ey6dhAtiXGX1DMLih+rkiXQcsZMH/vp3PpnOkjiiVAVcdeHGaig+ACkv+p/FkmnMfl1mQRuE9pVrxR/64AQ5Xv8psxr5K6wcu/hgENVQt+Q93GHLD7CTLz9JhW3eKQQJFVBTrD0gtqhCTSX98/xzoPm/ejTKykRTYRLO7rmShnXlwvgwuxbCMnXeLw/G/PR2vR99fjQKgoOHEL4tYNSELGQ6s46f+7OVzUc6HC6BZcU0khAy+fd7UQG0N1THfFs/z8bgsPbvhJGEsB1FLSH3P2FsAPO0eb1RAUMocwBnLTpD0u6uoUu9H9Y3zOGT5j7UhiIt8YeSmD5iwJPU4wIcsMrdjF1gcAaCySE4xhvEjOzeLwPO8Nb3AEaZrlXQLwR9FudCpvwWHBlmPS4fovpKSeqNtedteyJlGnAkUTwS1fEKKawtM/ip8zB7StM3ya8AbVykMQUMPCZR0rAaK5YChzoYILGh5ozKD+CXRF1oJvrblIeMUSjtKawwo8p8wt5uvQbkRxx921eIxjdQ8Y4DkQ/8Qv0BXO8K+5CewCfyxK9uLIYqgz5iPQfCbRIdUZ1uMa0jDYSPhJMvD3bzROxQ9BcKC7V5sO7oGB5Wp9a0vlKWrZlDw0YH+uV0GE4CumYsQgs4k2twXnkRiw4URWH52vcCg4enjQH6bwDTGkkSpvm0xEuTEF9ksPEMTbw8SMw5fa4KXBsJ8sS+c5YeuxcvozKNzwFUEl3teKQff+2M16pwd4iwQY96rOxhKhHmrwY86WRs6dDStCUThVAu1WzB9HiCmpCM/TE495TxdJwxSFGPLDWGnDHwP5QILl4sVOyGkR1ik1nF1cC6svG8K3RJscHvmp9HaEMJzGxaO7Kry8Q+AKseiktQBpAaXt5sT7ScoLxie3gQrLGMx0ryQUhNw+v7oL8rpihTi9MUOWtqlJY2w0sRwu8rR3QYjglr7wDY66v3fr9jZJGOpnq1fx/mSlLkR8XjxeIuCTSdw6OWAXleDYKLFxXZfnGkqelYoDscGkpIi19+uQYyCz4yFWmt56FmH/BuEibCYl9WdjQwRV0uA6fAc3morwzsw9L5l/wae7FSVuieXAVJ6p42QuOQybD3jIQpgc0Yy0lowhPfhi+0cIZCPJKS84Xerd3Q8mkl82j3dKpx62d8NRGwJdcGBe/Zz1rkHx7aOqHgChoKKuNZAoYFxJv0L86m4Ou4a3KSrhiMdsawTjbTiS52dv6ipQh5Pkn8xXRVDe+Cw6LrHnMdG2fsfZ7E5xvsqcfR2VuCSC6nJXuVmpIC92Xa8KrjOU/5rp8q5K3PxylbBIlzN+7kGvvaKrcs5SbhfxEPZRZK6KxDanX6wY2erByGQN/puOE697KXVNgrG0l1wbBhO12gdXNvthLy5FyzGLee8yZ0mxBwVlyCsq1cQmbps1O36JJm5GmidP+ZHJhpg2zN9FkrQYMzyvO/GzctgGnN6TUy/XxEZvQqHendNeedzKY5QS9RhqFjIwgLTfug/qyrz6cbqT5yMyTtdTFJMApKamCuK+19txly9ETIRSraMqEHo5NTrqdGp74Lo5fq0DKRODiru/0ydEHIFOKRRHEMDtTyQofRrq3Gu8Wow3iVUvckd//F5t0toIuqH+/zkgx0fEnJ7YZPL2n5F/JK4pJjepQXZeOtNEAkR+pxOma/XcfVZGRJbbV6YHRLa4Jkh7YXis7zo1bzfdBS+na0CllDfkITMmyw6Nd9qgU/f6ZK8GpQzEjjusNEhAjW4kN8vqs43aQ125xzTaUFQUztWeAOEIhGDfP/noHZkJcYUaMnbil/n+W9zoW3ujwxNBbDssUIl7xhmITXp8qn1Zkg/cz7A3c0F26OB66CL2KeqyULSdhAhDg8whHS2f8zwbAr0lzwNXcEXURY+MJR+U0JbF4KqV6fxHNqVnwrvOLTGpqpr8bJLuQ2YIQRUokQeTjMHecf2wQWkoLW+a/DS478sH8/nIUt33msgi5O22tGEufsNptqMAS6cHcoN+iGORPAHeTAiNL3V+yeSATnFSwVUf173kLy9uBYL/jDHWdOPL2DrOHIzgpoFSY2VjBs1rrt9Sga+o8aRNmJiclohXrXH4J/PH3egZbhvrk8Nc0sIi/9GrKarE5lqgKmjBMlr/aYWfhkUsN5ljh4dTeI1iFCAKWRZoYe6N+1lrtb0oyYhY+bqqT+ssoL8/LutPQ1pVzbWNvSeQUIUsrkwGQ26Jmp8D6ZDWDv7Ihvv5MWSkRczRhki097IJsL7Nrg5L3k0RXE0mgDYdKIe6OGZbzrLzzLGUVkV+ruM3s1ZxceD1Ra8q7+/vVELAC3yiVnsuOaQtIFQCQqL5NMYZeHLTfkjOezw0epTxgWSy7hST2KtRAvyORwi1LOkxc56s4+CAsFS4zzFU/iPegcVr4BvN7t9j2SZOKDpKuhajG2h0jWoaGIWJsV81zsx/mpYCmLu7Qdj4wXEUmwOFRuBHCQ92NbaTrX0AuIX5m9K1/b16GJN4Rt57WtSGXwNdvEIMpIMwv0GfJmM8DJus8CheaNUXfj/jfsyNS0L7dFIsDmHuNKde7g4kbgVwQIRL5Iy/JiLAt7u0/vUy70vxNAK3FNfLwXIni3gVEzsn/lgKF+ln35tzJH8aCQ7OHl4PtnNcK0ktpV4dk5lJ7esdVyv2c8ZaB9eW1C1Oc9dMKciT+JBBiVPRz8uz565QYo5syruaYLHmedUTmS9jDfwm3jO8WCmF//gxcEhs+0LLW2WzzI32zntjX4lpI9fFu/rvjmKBzorC+f+u/2ZZWJIBS723PaV+0yTWHXxi0f/Z5S2JyTF+yWnm3SSzc+nWH/ZmQyygqSkXX55y3NRWBhsS7/KfVvn2GaDXH08m12hhV1xCd0+DNdQVerUir2RWrT3850rD7LPX2/7jykPSoLtUXeIbK3xWJUgKOMsiWmv7eB0dTYB5KeaIx0vcnaRknJyEPAM1n7pkSuLMQgfRZ1F8y7qm5hwpr8Lc+eTGDur5lOMh8yF8UNAK3ynmRf6C2i6Avcj12fv4Qbc9GkYpxsk4P0eLIPKuI7CqM/qRW6xTMOlEiqSyOgcLJI6dGsgZ3Kea9d4vrOoukoZnQUON2/JGXLCPBnEuHGTGQLJldQVdsCN+em1coje+8OCQlNuCpfEJtrGIq+RHAOuY1dxvUc7sSB4OIjKzm3+e8FUgof5Ww9pe3SunK/YOZDVvDy8o5qEN09MKBLxORw1QOeJZsJAg8/CeYLM5GCjbtKSgEKbcjLWzahQo8WfBgCIXZttczGIBlEFvNUMaWZwR47CVPVEKufz2PZFVf62avvUKLIIWJsCAfXos1fmaUf0iYOtGSwktKnL3EXduZKz09lf7ciRI9fvMQ3xlN1QP4IsE2pWy0mKa3jZtSrB0yaYOKbZc2feQo9gBJGfSgOylW2Bbvff819uMlXeJ6Zart9Q02exne8NjlSYZPqiHYE03weMUwL1lkmQQBBb1PxAot3jdEhhYoFIOaJLAPdZY57L/lgzKL04W/9Jx84/X05fS8KTFMZJOoNFhJ5X+q6StWUFVjBYtB4GqSj9xGj4YfykdOyNJYuv37Q91txgRO9Oy0VQSKkJT5Zg+Z1x1dNrKwvpkBrMxX5zvjTS50yocFEgE5E++qOWq+rXArPLUvOA2RniTBwZI7YD3wjqmEetTNOTHpTfkQUKMxuihZlQ6yC8z91iU1O3OF4U5t7PNSRC4aGKFbBwQzeQyBo5G1kx/cmAKC2bnx9t6MaipxwrD4Nb77BXXPmAxUYICwd33a7yYVYyg/25MEcsiUWiP01Tq3QCutvQfRguWgF1DMu2Xs+hEMKPjLybMz64txjrCX3oMh0dQiqW5rrHzTYzrzRL/bDpHa8WhLfBREoUUEPDF6x3UBqB9VZ2ljuv5lgcGB/6/34902XqOMNUGGDC+1hrBQsQujcw98gL2NdTKtf3iAuQ1HKkQUA4znsF+ygqYksyskFJOfHClYB3HUzwSxpkaOzCW/3Lx2AggQMMYKQJ+K7/4kI44wqV+B2BCrAflupTF7yq1kfC9hL3CTEQbj2DJ2BaMuX3eeaMd/RaKGlyEe71U4DsHGwuIhdLm69VW19ZdmJDOAo46ydTv7jpk6CSL8xGSN7ydJjNAs25v8BIubrBes7+0VcDXf7IG2uUgbzM2TcoPw6DHdDbqZAQu9HMowF9EpO02MR5RJs5mmHZybcxYNxlFd6UWASUCB3GFQNQqGZI/VsyzvHNpL4zwlORf5o2uHNAByuWpor0joEz750S9UJmL9qa1u3cL65yJgV+JviMSR7iN8kU/vK7arxcxXOBDUAdTFDyTEMSP2JykL1paA1mcKoTRn6HMRq8S0Hup4iCnVFhnHTq4uKXl23Zvbre+kpvD4BmOAt1fmJkI2N6VD4mheaz8ZC9RuXOm3FEeNOmlAEMmHo/FaNc4uUJ/tdB08Nfkindq4uVJ3gF+M3aDBrUMx/iEWBT4qFzvzwmXiUZQxKNew8/IW/l+xyta/Qfy4T4x9gfFaNfJbmMwCBlrITAELNRZqGTNDzBJrVDbzU1MVbHyi6AKtAF3UYQH3J3vK5fYTOP7ccC89DApFC+Z/yFT5w3rVmTKFWeOWbGr1VbuHHxzs+k8lZjKMCkg57ZqS+292StwVYlUW4Vv8F0DzqRGDLyU9yENTyuCNVQkYwLD0Kt2/PdBk1fvrUqNLIF04dczTelZEM/X5RAhrfnvcmeDDbN0e6bxV7cpB1o/LBVFXn1QuRi3WyXfv9DokGkpQkDA7VcsTQnCub9+VU68yGQu1COc3PUl/P77lnMIo9UIScQ0BAtsaafHxlSPFUIRazZ046YgObGbLI4y4lOIdyvOpGDFDubNhRKR/WuQl2beNJC+tcHJlh3OdrMaq7ogGOu4TRIBO6XspI58XN5yZ2Fek9JDElZumA5Y1h3DZZsM8GaerjqZIyh+5tLt4UO1n08vwDZn7hiGSdg8wDIPxqlLzK2oA0drLH/GfEU4vX3PR0oC8sUb4sDiucv7iEBTRj1CPqSzdnnT3VNKPetx3x8iZa/RaCB0mwxSLdt7f8HkRivV71R4Rsmm3xef5P6ZEiAHe0T4uWthNYz+v182utHVRUSH3IRPVZpf8oZwBEpHcHX32e2GL0M+Yvnpmy7e/553DzWdIxwwYAor2YDtgkZd19NJ9/veAFN3UqDyt2EKv1ICoP9FpVlzJNkgTQI7V5I3JnVIxcvxWI7gSFQCTsYbPG/jDg6TPVLHS66U1mrhDTlc9iKM/UWTZQBK09UQfLeZuNSmKs5pKd9OV/21VPgGk60CvD942mImWY3MLd+STRsMqaqJN0lokfhV6yBeIBz13toSnMJ2IzhzwgZNI0gI4RzsyY8s/dAm3c3klNaW/oMJe01Y83E6asFBZf/Fny2fra80l7TIhVlNYMck/Cee+aN7NE8mSUbOFPc3ifwQgc/YnWJk0XmSs0emSsZrdldTnVZoI7MFVf6j07xkVWT51EB+IMsnTAuVQNF8qIyIE31rinq8nxRPFQH/hX8xDZ6/yEPRcWz0FtNHhIuTZM4Om+3MVtZPi4L1+GivEgVBUvXqMt+93IZux+um0FSOVT0RclQt3/z881rhoX00FqH9TGBGzmhHZkwiLi2kndxHuCqVWB30W3IOIrMoA7sf8bUpbPloFeKGB71eDpfDeHIXBqcKAs4OjuSNvuQpwUqJWXComYNVXl3VcIPrl/zhzSgMMSTqwCz2gi0XcMErqykZ1VpOja6YuKuL1et2m89PO3t5/yFNBU4w7Sz0QfnTG6PXR8X9BmFF46844YWsHriTTkB+O10kdTD4Djffdt2rIQtZuRDxG2d5aWqBBwOz+2iD1F8ZixCIy3rkyMpSPttZmGhJpWQ5huMld+TqV8RzoZLhFXYPHGdNfT4zfSAG5X6Drpgm4H+QixNEjM8jUv3HXF8j5LoSc3fIKLyJ8e444xHiz5+wnVjmVCcVXckYjK7kGna0w1vNaRQ7wjFKk9uzJMFL8Mc6glRzH3OBYkBXZaqjIZOwvL8WHvUg+H8l3W7ZnA3ds0ugvNCeptaXlz9lsREo7g/gG+v9PKPP6+fIdM684mEshKF8ufltN7f9HdVnja9gaTGetDUqXokx8W/qRQeloAWCF2JWueRLiybUcGdaVZiGfmGQA40w7gASbOcZa/E13zvH36rvq0Bs3TrWvmGtnqIGzA6FN6ZG5gJvbkM3oxRniH0ze2MrTWn4iaLoyrgTvflydwEl4l4i1TV7CkihnlzBl/MxLHFZmLFsvyzjmOH7TAliveUniOnV9DOlnknhbJn3wXx86QLd928nAHYY1+PtoL+jY8LdxGnZKTVqtLGjlXtK2VWUfIZ2fh3bxDkMbU0DnumD4khoGscFYSfBmsnPZao8ee8dzoRURyp/nGQ+vue+nR9l7m/4IHJTlRe4W+ASF+jT3bq9TRcgfmyo6QwNraDawzRnAHtswmYu3FaB+sYhQd8eVZVvH8CWaIIypgSXyWAqvMMGA6FZQ7QYtbPqgfKseQbfUP4BoZZSrrGnvzOA9ob8csjvNOw88LqcWlyOqyep5cV8aSTxWfoqD8C+1HV1GTd4313fJOG6UykZ3OzTC8M6KUnA8fwcOskJ2MMvUmuD7q1BsjXNfYKUJw91EdPC/eEEVwikawa8uUrI623T8ty/lzZes/KHWphTiSrULUHmkKlQ/6jUK//CKjXs7zvPuhadtkGyF6SMrIlzrOT4NO+Pp6n6nbCeO8I6ISrKMVa15pwGeyq2r8wVVof3FbSX0wDH9PULzJTCQNy4ZL4IB+6pF1fCYTvCcX4G8PlHloOXeuOmxik1YIxlV8wyoK5gQdX6yMT5HAt2xATf3BN6DsfhbRYHjfKLgrKAf4CxxZNW/ptu9g4s17pce/H8vRIy3LNZ0fqM/zvRdvEwpay0HbxzYI2k6xsmzqw0DDeKHI4qq0qiGcfRdU2sxGuRcFDa1KTa/O80ZSVy2tFdM5XH07/0WrEc8nH/LWbsiq76OaDJgTRquTKkOdXHPfs6pQM/jo+1tfWH7MeqWGyrSLPNJsSHj9l7O70eYdk+948Z8zckjnXOTw2J8PjGENXoVHlSo3Lhb7Ki2a3xY5YUI+ogrqq7fh4aiE2cbX8prMyLc3X9fIZhLL2FbjVfB69Q1vnxRU1+7xOfBuWBMIj4but+A//VABJ83yzlu7V/r8EnSyXBo8s6a819gnYDkiI6C+gFad/UO9T2QNLH7ivvkV8iDZc3TwuqIYZ5Zp8naHhDcKhGEfpYZWk8s263adb4ifkvadtDdnRjDN2/KjU73yLLErSdbTA3icJuv8OQP0SbaaYQnBPihPc+kMbYCmzc4Twvwp/CzQ6YCiaIIJQJBBDQjXOsktXQtKKXhUoR2m4BUp4ZArTc8ow3dsFdfOCRuuypB9zlfpkRBeYAwwyfW/olRzzylUW6g2xuk342unJWHvPUjRIHXQG2mtgXbUq01KitHV8nK5L5LwCvP/2Y4KvN0UCs4esK5YmxvLdKhaQQAWGX+1qBadqvTRp3EuIeSe8XvzCZQoGjhU5xNTQ7310PSPJBGn2LO2kGxtWynEsSX65l2JomKgJhO0mLi1dX8NZCWBPJM+HCQ72wNhxVCW6D/j+oVuc2lGMl/2ch7sodjLQvbkfE7ABSir0ikLDlYqpBzfJZ5SwkRPPkqLsZAzdGrDKvuxaTA2PB5OjmC/0MJOKQJuLOy71LWOSCpA+Wb62IdX0Sc1/O8EHv6PpoPzxRQcNXRk77KqpsEjbnmpZL3lck/zLODy1SS1TvpKdPxLgfAmC2a2Lf2eGGeAVee3qeH4Esr4KJ6oc0uGEZtJ2h/JE8bgsmBCgwzzlz1cJg9NGKMk3Qffqv3zKkoYlv5er/ZNVOiktd1c/Rn1SvHndvnq/xyBow/HFPL3g7pSlCfvcgaL5yDgHA8e1o6tOQYUXeyKu/G+pwCz4OTP2J+fBn9EkmtIhBY3EEzvzMkAGzdaby79VUQ2ATgQ9aU3b8lpCK3rjdPica2vdMfT8YxpQSqTc4I43ECdv7QxYN/9lKYh+BG/0Ryr+aBjuyotnQq9EKnIxSP9Py42/+mCUbOsKouwCVoY/cLe25YWiM5mNbik2W2YRjh4Lf8jSZcDkQyGvoGFpkOJAHBJRMYU2L8N9rb8XjCqeQHE5B8AbeGdh/sKV+FRwsvTkL3ccPO6gzxwPX9wbRNPr3sWdxyH+4SAaQTOnC9PJ4TouMWQjt9j8z9MkoOQjZ4KL/Hd4JUokpHkjJQzJNMqO9L6RtVZL/4NAYmu0qzrD6JeibpB1t7WGtPYcJjo1+PEiMtTmmpxcKA81EmMb6MuBj6+Er7gdK6OEVov3uKKz8buELvbQj8p2P583Ri8CNJ/tB/OytvvaNekIiBgGwF4WFtODV9dX7AIP47TH/GM74Oi3+tT4aWXWqVY13VuaVnX9eYRpGQj5evtBYxtmt4FPHkzWubZ91J2GvwXailwUeMD4dCYr6ARZ7vWRSIynhIS+zRPgkp/AUvTCwEyrVt5FC2mEtt4ORVUgjLuUL+htGMkUCmsDHaIHT2JnXPR1yPoiDs0VFXSaWZtohnTSf8iJK1lYFtEAGXmRIIc/gyWOdB5dhB8N7ECyD3lkkKnIEsHgTgSdjlO5D2m/lanFlFeveU6rovqY+fxesdID4iLD6KMcmDp8ELJMJyV180FsNoLQp2Gh9xluQXmeULLYbJV8hXyBYj6lYosOI8BeVhO6bs8/W9Hnifj2pVBAfF4gCf/6/cb6JTHQDgih6w9GW9n+HfSwhhv+Ofq2PoyQD3McYyxC7H44xfWjqD9RkAeibf3SxOIbgI+WZtZR85lHwX5g4WiuOXpPJWLf12B+8kinhxFGR7EZ5V7k2iICij+CUePE7eKsvgc9jDQ7ASlxtr071/OJxxRGfS/JBPL0pziHju6weuH/p8vsi7qn/1Ge0IFAu1WkPRArv4zR9uNN8aOI6PM+f0vx/Fn6t3S5jtB7rzNFAM15aipn5QhPANYZUyR1h/T8F6wSrGfLYv+o3JzBJEA5lGmnTs570hyn9BnY2faK5hvHeAsOsDR/eeUBKpSlOOsCipBYJhTu60ckDinwP7BeTBgv6HmPw0I4BK1LtWQaaGpcSBGQbqNuQ4X2BflbvvDoa/t0tiW0Fcq0w6xJ2rMTevrp6IKmyOn6OwVddu0tyoVh9oO69oy/LqYcaAg3/3r29f+LJzoniRwcmFWhcrOsUWIFXfT3qeIqPwvECSU8gXxZlK5AsRtocsM0wzqHJX6L2ekapkmeI0D7T5LakcOlDVdd75SqJK9jwwyKy8aUQCHAOO4HDCg0DM28GV/JB4quqcrdEMGUz92vyqC3JYHg4fHx2VW3bYytfe3c3MkCjrXZjdMfvOVVZBS4834ijeL/OkwnpL6nS7DdSqt3KL1pog1PhMr8aXQJUR9dexoqSD6FVUY15EwW1xWuhvxxiQBXwbUufK3NpROsd1YCaIT+u8vb9vtTG35LQ4HyFHS1ckfvU/vtSP6G8JjJmtldg8aZ8N2IbphXHmd5peMR3gAi+2oQ1q4JxjNWTdLo5Mv13Hi19cfcYcEcZRa3D3rrSq8+/AlO0ZTddPCyCSnggZ//bdptN6Nt8+yIBo/ASbeI5bC/pDpr1IvJyHn0yc6olJIgdMDj7G9/tUBODvjf0pcJRsg254uleCEze1OrypFgLCbqspbZkbzRmfOYKSp9wMuZ7GtjCydRIHGenjPyqFORuKiubvBVXoQT/fyYMOqLUE3yGDe5iiqcWBG7RE+QI/mPhy+PBvP5me1xUb4igVdnMIxSL71vcnsShHynFRF6egLusGF8zYrJtCVNJmnG25b4IS98/LVh0OlOWNJDU+MeP03SadEFQMq0QTzOxZX/Gi8ptbJSesckifZJ70gwzyLWmrDBy8zKGfn8zGkROyMp8Xl+y4eQskdVdbfAJVY5D79D/ebuxizHdWIk0OFhhv3kP994RgKJecFfdSINCBFdGibY30jBnNAhB6twYuBYUytZT6ubGUD254yNet6hJJLDTyErOpVCuZGmrCHMSWWmUdyV66J4giE6ifenjos56B21Cn2wB0ecvaAyf7jJ1Eh3Gd41lTy4Dv0qanxwBLRUvH0XYuT8PiRJjQ6Rb/Asjt+V8x94e6WCZ+gwwVZ8T7olhRjeC2U8oSxJduqpBq6rEMoyaO32Zd0RsNBeNbY1ZN5kXMViYLXnGg+n4MlmBPYyLDVK2N5C8nx3pe5OmwIz1Vj8wmnJwrKQJ4jfkJckKtlxdGkF5ETfLlU/p0uNKa9rK3IGJxq47s8tWLBnWXx3IwMt/TLhrYWAcYhW2xgOAzjV/AbWLaQaUOW2xH5grLlBIhvaa36Vp/AGZJxXNshuNF6MkLN5AhgGPbdeVLbrSRVV+zhyE1jLXKrxg4Z3q9bGPNVBL+SVkxouBto2LlbfqVNUk4/1vsgX5b7aAAV+FoGVkWytzxDrKl7v2eMPxApkyRpLQ/BRieg9WCXfNoBMcDOi5jHBO570+GesDUc+LvkdfHcSokEQP0DAvcpvSUG18cTaBH7d+HV06MAkuwn8/+qNPz+YR64ynmRQVL9I1+SC3hjk/jOlloUkqCs+UI3PEnjTGoK5LckmILo7yFrBzzfO9V6FtoVkQqWLcKjARqifM1+BpNhJNSDNegHmnqWHbGEECXYDa49vvJ+ns2uuuhxs0JJJa4Uvoo3L9Hw7bnDikvsIlmONUXldWJCt0987CXkCmKE9cUsnU1Cp6jBXSzzbb2sZypz2/tWbbzTFioNTo04D17HEZaH/Tp4mdVs5JnyGg1Y+zbJVAHMmhl2+Merog9Gskbry3hPYok+sQSolAqiPbAcrBiX2kGVOlADUVQtEmFx3P6rk1yi4Nh8VnxjxRo4w26KYCSe0XtkwOBn7p861UBwSHFNXgnLxYiaGv9NZtY+rG7Z/nJXDLNKcrKDslffvk32q1tPuYNR7vjwdwoU0wRe0AHGL5q6J3q9dryRT11CM+MnGIhwTxLZu8Nt71aiVlh1PEYjznmzbhGmJu4UrGybv+iHNzGR48bS7q7XHlfIiRc0WzLLcqv18qnyeD7tS6sbjIr/OF8r5bWvkF49jY5BrNGm9SqHmjnrHu8YYWVDEasfXwLK4wK/3TnkBZvxGT1zWSr4wNI2+dzPi3Ws9qeR8A+IBca3zmO9sl/gwyRc17McRGJWgarOvc5DNpyUAf3rlsO9MfaoZH7PK0LlsPmpsjAivLXafLriYPxAX71j6uK1X0Y7jG+KgVZDiCRJaYTFT+HU28hG/nhRNe3HoR8G0r42I+J7DM/893/SKy9M4l25lgm1Wcxn37C5083FBguV6nQFUxik9b1mj4tqzpgm7OoC7J6m80FlhYiBZQFlmzoZmsGvSWyADdI7p78Z7jgwVCBtINfn9zK7Ed6Kpj5aSWp00PbEBIayyn8XM3aTNC8a+J9tG8D83kCiXYVb3KuMFGBlBp1QP+9je9fdidaNYviadf1Mdy/8PY4KgTtR2YjvDA9T/VBAPfuuur51AJ9KDpb9f6rCH2ane3yo/Y9wzBtGCh2W/ks82sFwBrlNx5NrUqHKr4rL72Dnn98jmz3iMAz2leiVBiSLTHeOg/TyfZeT4TAkXeatlJp340VIpzhoUoC3SBj173L1UTIBmBDWTaxnzvhkPbYMd+zrPmKLzdqrvu0YLTtMXMxF9JnSfSjRgOdeSMVObnRbA1/6/YdN9Spzbszcy7xr4v1v16KPQDV0tUON5Oc1Yij0bZ3WKcjx7jOZ0TylAgzm3OHioXfXpD8iO1ngUuaYrJw41RCizU6zSIh288Pt4hV5KuR6fIsfF5IG1gl/Ce9tSlvYFz5CyhS4PdW19Ue1K4AWD9aUT9EeXgdv0JmiJwHqtVBMn5hF5zijH5XxYOCeYy1cmZ4CJnwj9A0MaD4G2gsUk2JhiyerzjfdyC7A/ShuEV3NIuh3mWMXX/sPPfHEv1/vwttIX1U+D9WbXFpQHfOn4rGo17BwTrHwzXk1dh+fDBylZ4gAVEX2S9gW9BPvJj1JKdy+MSxOz18U7pLbMIdBVnnSRmaI3H5iSu6O9g3mn/vrmrFEgJFAqR6rPnw/OL/ISfkqPhs18bzl+FUIjmbbNU//pPUJJoQQom9+PzNiDDYpSPe7bvUDJuFWEnB58mxwm6bX6ezIrmCsjghpeiM1piPUygdyBXj7cK1zwLgH1kHYHQ4bncKF0DnadUGbjO/4fQEinJRxANPAItKpRbV0uRkHGdYZHmyRo0MZ3mGrrYH1qku8Or+osH9ejeXhn3jrrhr8v2D9y0rGE5fAipVkd4vvWlSySXhvDVl3Nmea0iJ75v6dyU+YTqcdC9ZnizdaM87Ia4s+0im5tRRF5Vp7cJHSqQ9rDpdGMTKSZeODP0tXCzrKygTA13fx2Mml4G3Gd6Mrv15c4mTEA+FwDJ9GdjJ7igUfzUsTHOKwlU45a2AUdHajclBS0J16LcMQ5Ugtt9VWqVcOJlFZ9RtYAgYc23cw/Ac/WWieRPl4nw4sTvoA8Jwnw2XKeSwx45/C8UqeBqFqbg2N+TGR4Qgg7OoiXF6zDRynLJ4P5xlF9fVoiCbFlm07bMQp4EbJ4jT/hbmNHdpZtUPaf3cfll5+HN27YjsmYhGW8aDWkjNhtjj7XpQI0ryqJRQJerwIjfpy8JKb13q1LW4Yo8c5F8tlkEUzhOrjPi94fNKrP0+gQLEbTmUD4DOho7w+BGLNFsRcoidkLIHptBBA2Tp9oPJaQw4m/HyxlMLnehxNMMRKCGJMNLlD90Wck3f1MUXlz3Lfutvc6ayZ6Vj9PsjWk2oZ62PXtDnI3+5/d56z4F85osrv57G+fnsPeoxF3UiKFSSUIXYIAfNDMt4YVQ1RPmhxA+FQcj7NnKpM/K1UE+eGBJ/rIVTtne7yTx9GZRxh14D+bdMgR8lfEqEMEjAe2z8tnTQeRy/UR185/DESuhLmlKguOF5NVncXitiCV6M/GTN2Bmf+nez4vcKGh8aLW+tu6dM6buVL8SO6ujUOY9H0nZkAPE+5nogekO3uD8DRE1gTf1LDJBv+dbHvI3R1GokCwzGN8VodaioJ98ydIW48NLl3QWUjyzQAq+7TskVl3CZEthODZtm8i0myw8TF31RYHDF5nt3VQd2vRnvGQfTPbn4j/47AyPoLq3a7+XZSk5y/xVQlzphoM0/4v9dDb9oLZpYbd1G/awzArFV/1xsDphmK5QkUmtMsnryVDGR/AAeyAWy55gQR8IPYchcHE4G5+y9tQWROZ270/1lTluzMfi77yf9LY6yzMG31VXXKkQuk0uWIIDkLA6ozfoHNdlzFIAYx9f6DYC5iLjIF/VJRbkPVvcFSKWM/NhvqDAjOITicZ4+UMv9CRbvnRD5D41DFYpQd21iwz1AmmjCjZNGhMHvF1kz0KXxGH6Te9D+9EdwVuvOpeueUvuW9JpM185zFl7DdbZu3MBYvLw/AbNcPa+1p+g5ibuUm7NtJ7NPjZBtdGWcM4JhUhAKHF6odMnZxFKBB6wS798nmmcIq55PQXozsaTLb8aSm7MApfYvPAe2DgbbYp0uNXAm/PFBuieJ8AscZGJB0k+TWeKWbU4xwMfYaIlvJluhuIajpt81uk90HlA2wzxzU99cgNiY52139/gkDbP79aj+b3SML5KCet68glvLBsRXdBXMNkJGxDkND2CnqX4Vb/KYUOfIY9qXbSPz9V3/5fo/UCRKfnkl2rzAZz6QEtzOGrxJwwZrzjqa7B489MiQEREscXTsfP2VANlAQ1TxUPFKux58st8cTHcCjPqEGzRsk6g5sCBAOrIem3m9yZFsdwek9VobmvHcVbab+nAFeZznkTsBbm2566M72O8J2dxF/nBn+B18TNsQ43bPotK29Oy8jiL/a4cWNAAxL7SFQnrsd8oToRYhlp/75NxPVo2pHJFU1yLE2K51YJjg92LEvof4t/U/Zuwx1tc9fqgZkgMSFnM8M98LPo9L3y9Mz4YWSbOxVqRM6hhvPVRsEJm4l0HxHIyr8CSGysThvVrfri01iZCqcN1CnAdNaU68JcFWkAqG+zTwR50McQ7d3URIalO1OKcEgplX2/d/X694SQx3czIVbWFuKOmmhbYRQVtsL5XXHoqGHfkOgIBjbb0D6MuWsRcThhMpsdEA5aq39F5ysflKA+qejsrbGlwNEmBy9C/an/LAInd/++LOqCQlPtRbUvwlL5+L1vu35Xayr/bkQMKkjNDZPfscnaYWnz4a7itYu52XMiGBi52YJ2X0RT2fRtx3p5lpQ4D5MW8oxR7QBP3dbhFHjbgB7WR+p2iGo488EIIQbfj7G7YaUpH+qvAOw/6k4MFTeSV/lwbXKPR/y4yAh4z2vDCrkndLmU3PJ5PeKgJpoUuq0PMdKvr+MzqkzDvq62Iy/S+8d0cqzsioGWuydfWHok0l2Bfv0SA7post9ikW1VreEwmMPoHJfZKGfc3nuhxQQDO2JEnmX5xjDTflDsr2dQESCE6UMrnDFCMOXmxSopNPBnt1vhDqjSKgLfz87E7GQS8tmx967wUApM9c7n37186ljAPfOYBROOMK1V4jIFOuKwThhvR900TG+ENr4VBEgWBC5cQObfxjqRWhui9y8fLEvQNmTD+lUv6FbEdiggcp9LbhYi+HHCg1S/cJ/U5S6zptbqgz1UrRDs0wQBWgrOVAAGEyji36Mr5TrNMuc7XTcG6PXuXA2VKSFKowc0S3SCM0s2pQuSmGFrhuHH5NtPiSJ84goNZsRB5oEkqHLaqqImJQKaiMgdhKiGGA+H7Bk5cl8/EewzteoCeEA0COLLf4pv4biTNpFMfZWkPtdidO/ZJdJYX3N9t0WN7Hd5KruvMmjm8p60Hprk9ZXOkzPdorsFbi/cNoCXP4YPJuggY5vSGFvHP/9ajux9qm/j2bbF27fukBuFaAtFJuoG1HuEEQBv+FnjUQvgPBAH/ouplXGGKDS+G0Mef/n/iy26pvm9vgM9+7rIrg73nC40FukMs+9JXPrcpvxJzvVMQPJ+L8lTmtHMXYoNVnS1YdHQ6DHc4IQcgMSdWX8fM4+vS40iPSEeCAFKE1rb4PIOzAKyVrBptUpVbsN2d5teIEiME1lWI7CqAKKdbshkU5xzOEghnHla8Pp4c6MtTB6x2rQcOGW+7+LB8t7bhqE8DKEuImue19+wziKSIIJB4zJ8u6OxqiIKZ7K5I/WkIJbfTQx62lOQtwXrYIz7Ab7KmEIOj3y8DuI+v9qQ50aGaVTqwlMdqUtZUJYdwA1qD+Zxg8TelSooMqsZCBOPFtyiLKNvE+82lIIx7Fs+InIKGp5Un+RiL1zVFa4odnoySFj8pIkLyfPA8FlGMXUGRLKnXoBVl6DKA88B/7RGO+EQKu9HOlZTDhIlIWDnpSnei5+lH0e1e+eeW4J9I3SZNzsfQ+iLJHV9c3x65r8GhtOnquc5pGxDC1dAnbdLqqJjQaHR2AkOnnt4ZhXO8CHQrGXsqjMpdO3h1VVviu/P3zq+/q+LDbs7ib2o8VlluXrxhTLnXSFH6IHS+5WKj+pejJyI2va5z4RPyCS5x8NTcSBH7o9NB2MVSIVpmUb/AXryJIqJQIdGax2EnIA0ZDeopdFte4dK9Q2UUCjr8dujtO1Deo3pCMjCukICWHMyswyDUMPHTs0QyVxo8VPE6iKkeC9Bftze8PwUYHxTeUx/WB+Uo3770vScMaDPLUYAoMeUNldJW7LfN0S5IJDpB52FYjWo5kh9ph4kOO+LvhqTr/FPMUOiW0s+n3nmRCU9akPVpqCt1f34vkRnG6n1UvM5W36y6bhyL7qbUkWT0L+suyaaEpwrLYcVUT6m4Aig3clg3rmJzFTgXB0wg7EQeDLYjqQeNDrhbnx6R50jKgdSXVleuqFBqfhj2DrHJNTJF+ND28I0FZBXdKStbobebfi9FAf5CV8ivXcGExNwzb6Pi8DZ4tViqwJTTq43jzcZFx7Hz8jLx5h6ifEBrKyG0R7ACSIBcThHQMSe+UNrwTYAbXwsZboiG3ysKfhmnjtqKT6v69WXHK8g4mhCC5kmNssbgnDn41eK+W+sYuEA8nFPlRZTXX9FEtTWErq9E+4sDzG8WlEAJYZFlhtMtb0vHZcOgrlXNpAImWZnev/5IT8otMfHH6j1LPjakPwBRZo6+uYCjDWy23167o0QbRsAjuNCwdJPO4taEQ/vc9wzv7Nj7lG1QgANCdsjWhcjA3CjpbzP2DKfk7N9nAtMnwCxjU9TMqY0+Dw44/ChC6L9TKuC1v8gHFzMfay6AVkzBJ9CiD2ui662RgDyTvbgmwNlbW8PiHm2b0Vjl3TifcCLpzT0KKmwlP2XWU+6laj+gaGbqyLzQt3hQk96b51Clax531n6Wj7p/thutZ+KWi/xJDedgc9C850DJrbfRwSkJfX85/guJWvnFfzQXPoCpKSJ/BaFPVsCz2JtQNHPNriG64+vSNjl03hFWWiBdiL1GIRA7pr4cZt6/mao+JvRJs2J1heI/O63mUoeeYOXDreRCT6UuVIxT7NIEzkbGzK7w3qPlBJZHm/g2kpynbne5HmjveqsevxFk4Cjdn9mFtn3zRhBR0W2LjjM8jo9aOTVKzRWWorivZc0ck8lwyIHShtDkoXIJunwHeL51X6eNK1FjqWSmvNF4eR96DjLJxFe7HIrbaNabiXF5Ff1qYElUW7Ah/WQd32mmpGzLtNrPd07rfWMp2n0KCo/q1PB9iJtaLMQXgyXX5WEesT2Wf+XBbPQBGSXOxDKHxYSPCLZJ1tRW74RzBKlcsSXwKmr1zUmJl5/bsU8cWQFNC4ELoxuW2Zl9gnrnCNR4U9cQgLPx9rliDtllYxdaalBCrUAAuWwval8o/H0kWcoUINYEdGUcK8QIoXuWYrP3jHP920zxvxhTDUKBqIQgRFf4TkXgIemhX/Z1iu4OWyzNP3sp3Ppncn0wQA2VHl049tHXYtWtJkoe0F1YNo2sqbF6AYglfznxObh3vR9h6efoMfk/LRATaAH8NR+hZh0ZtgGiR4z6zKzbi+hG2qxp/zYk2IJ97LIlgLyR354YKK272GW7BZECv65MEUlUom0xs/9RGwl0rsfyVXvkX8NPI+eloo0aX15nTVf1asMaMDZkDR1m0knzrp29e1/DYlY7osKlpdghcDZLV2h1FsdQsBliRLD1Q9tephCd6iTgjN/Ghy1YkNil4zQAXV/f6Bz2+Pg+LU5lZgraaauqV0eGtcs216Hlch2EzkJ9E01JEd+rCE2ZskZJKdfnfFox/Aog2DfI6SKudC0bEpztL6wJuLnwNWIXIk0cyTbBUCgYorT6PiXiwUJFI6iKTgakyqmbJqzm9eTr0AmWzflml2tUft1aF34UwizQ8v3h9j/Og8dPwP4duAyBnaszPtChk5R8SgsIgf2QU4tV1zRb1ho8mePn1J+1YnaQy1HiNqvK3oMFIhu4aYSRlECngRD/FzfBXC9f3UMeqs2GcCIV2jJG5NygluPE1a+5YhblnCcVjTpBuSu31aCR3938AOzTLL4n8/KI2XmDFKDv3YJHoiIbkhAPS0wliMCAXFhkolhG0K2r+mm1uWSWIo3/8VSgQv4bQOqCYkKZeqKLd/kiU9dmAEoAXk1vEzKd62/Y1bU3A5d7IpKU0pqCsOFn7FGYRSPRY4hs1uH0IkRHRxOsa7+D05NvGudsewDnTqBKBts6ySPV4BM7KbEGd22mWLTBFoqfLwHUpN6qPyGHv83MfBvqbNrOGjoCJYJ0NEKUxKpGroTsWXFMy4gAFV1FYWED6Kt6oE5sX9DKH34vJyTqphtJ/j3R/p/J2G3OAN7KMYv8f4M74Zh1CFedAK2cZLKOWSRoRQUYjCtfRgSY2R9KIUfcK3WJrHhjj085FaqJzgWu8l7sM1OT791+kjcv/jHl+NR52z87YltViU7ji5dLwQRDm4QDi7FRxhRGTiy1nGKagwyB2FW9azzApNY2IEdu5MUTdgYcLsrMQFX+PCzgP7YAPsm2/Ds26vb+bBTBn6xqubBNZoZU/15P/g6fH4dp2Enp+fbg3781Gf3aL3H6A0E1Bdes2KCccBwZScnVD2ktvzvPha6g6QSDPb7f1uVPROhEAKoX09w8D8nc3NE2qpJeHqqCQbAEHVQ1XD49l2pxwwTYw5VbXczLmm7+xhv0DIHK39efB3x+szrwHNC6zzhbVIj9LafW7nzbQAbKJPbpXrrjuxIuDKATzcZKcos9RkXR1GkVlegeSm81VMxxdyF2GTHVbvbmmxarQ/R/q1gvN625Xd6rPmjsg+c6GS1dcWk5HwL7dly3Fv9pVqixOO/lr5hoTsRn7XIb6RwXTcbzxQoil/x2ibrE9M9Rv2iGEThfiwIB9AI7tsvULWGaLthHaaUXbo2jf3/dSG2CR+xsipBySYmPUlRlGDg1sww2iarhmiFAOqakcJZUGm/isIt8OZ3eOySMB35sceJEWQu/5EgOV/cfj7Ikzwz2KfUXl/06tm7DL32IRfDBhumMtF7zQCeah0WiqvS+gdMYz12777eedTjJP7lLja2HZReMD50XnffVuFYKazbugb/vyQknZEFivcy2b41dSOqIs8ZS3KHr/sljx1Hup3DVkpC64UA84DLczcWVEDc6RSTt2enfIMMSCl1BXREDrF8BIBEpRU4ImaEHOI1AW985KbA+R2ASbua9VNQEBhN2PTTSsUGTyoYMvDokCZ5va5JOtvhnRbsO/C+4IZPnNmA0hk916M3YKjTvl/Dv6Mmt1n7j6ykaR6Nqz/9toSuFbMadu9B1hjsTydlS1HoaAbSTvEEfsz8opU8of1mzuiypdPPJHAhUVrP2+uxhdTScJ8r5vqqCpG14VE04BJVNBKKUEO6leL+dOTdhhnPT4T2HKlEJEno+asm/2gxWGe0gITPiX03l1WQKjSPJE/P2R4Xy1k9JUAEkrWD0DEBKxbaNDUfuTOgos3Tm9ENLf+59xeZjGZdnBx/+3DwSGmQio8UkzCY1stVX3y2NaK4KebeZxvfgmIBomFt2VQkYwykvpkw76NDJQN11fxTJseW/qOimud0698Tc1cJzNGozEXuRoABywEUauAD45vWNaROZINDqHovPGV+qr9zCJE3KKwBEP5/NCMF5fPo24ET40QCwovmEBWoAlO5Pkg48b6gy7B2d6nUIlesgIVH+33WM90uBJGkOZpChKDUAgJfDV2ZM2cAOvlDHKN0EzZ+gL/Sa11osJx7Z5g4Y7svJuh33mN91CnWV9l1SuU2toZ9lQksT+CLB+2roAxHfxVCjQcPYUheHquAge9ajLf17YP8d6O66wDnaT7YNUHwTFSLxhwbcbcCN7tB909GMQAjumy5GmvUuatOmTqjtABYfzE04Pfi9kExrgG+3IcJcIUnNsvQudx96iXIDLUOk8mQOkwugZ8nknDbNqqIZj0LdKB/vFQLrLBvBOIAZ+9RRtqUC3b/JhTtwR+9g290RR1mJfsLNPaNkzsEpnhvi8R7tmoCpmmepaW8/NK2X8c+KHBpkDSMOE4Ebj6owEt0atIDk8DJcXPjhJIX0bibBvL4LfLc57lModjzLYo3+ChvX2HMBaoyoymSUof30YsRybNdiHtv4qK2kwwluWwMP4xyT8bbVzQdybH4vsQnEpoZ9D98PaJkBt8vC2bsGKWfZKOjQCZzWV+7KkKv8YKlDSJBY/qXO6dNr5wNgjYvWJKTbzVhOfDI2S2hxOFQurT/f6uzt8vyCqHyC9y1O010aAQN+U3GpVB38Row/GWcUDks5hkrJ5OlJIgHsc5rTRtsbiK1VS/FJGUPFXtUgP/NrgqeLD/TtrfOPNP0/A4Jjo+XQREysNiiBs9f/hFNWvmiP02SpIlAPCppq6V8HUa43427GQ+c6a16h8qPEtPL9e3q9IpeMUDKWTxDdAtSJFCNAKfdXskZZRYQAP6LEXvcYrq+HLSZXtEaag0/+rM91YYl2BE4GTi2xarcpjCEaaaU63A0VBlOx5mgH+3YczznukeVZQHbvYaNJZdnzau+DxrJWDke4duzils7TB6YyvWN/je+4bw1mt0zHeoatIHnSTD9VhsBMmJSdAp5RLilpZwqMYilbKQjLJi+rswghpX0dfsmjCogzgec1rIBCGeUAoYMp3iiDeK1NAWIGviYrHZaAllG+DJtx1kRKHlLGYnLLmdULmMBA1ry3H8VGbbxoYFHdM2FywtXot2T4a1IvZT/TqXwJz2Y5pr58zkEDOcn5n0YoE/TYp+F2RSxTEAjO+UAjKiNUmvHy82VYTevievH3fPYJhmJJoj7ZHludGqzgJdLZGfdgKB9TaMVnxWv7JjHqjPhpQLvGAIUirlqu3Ue2U3kgKGkDC6ceVorLMhsjeI5cPXEpoU+ifChG9OwXhQnPTkHBrvf6pTdBosb/5/JjTob4/lc74GgVQi4Otpr7Ko8PHnLrEVtb4RoFx3SWUD47xJp2+pRrrovDp57sArUJAFJdFRVQQnk4re4yiJswzIgxJTpyqsXVil2tmUluv6MZsjmkLwCWmE8XhoCCFGsz+CYImKlaX4WNc7Q+d6y4PMVLTDcP1F7Lx7bxSWrXPUrz9pvT0tRsiLRG0Fseb9KRMoMI4ZeTBPINB3wwHtZBPxQCFKbQqgQfPMH+eR9L7MSF5o7ALEQ6GTWVzWyCIlUQUd39Ukvh5sxP1iJxsPuMcqT30vs+1amlNg5gP5nfH1/7alBC8mWJ1APhUl8EVXaNohs9w/K0tw/TjbsuOmLOKG8GagphFw3opH4c9R59rODA3zt1gTm0hWIB1uM+tkkOboH4sbE8TCN2h5Iay8BUzw7s2oXui/9Lx+FYr4ie00FGGnrpyOytcoTpTKwQ6PHtZ0WpB4Q6sBTAlVn6Z34FWfUdCW2LJzIVBJxMkkbrJUe3WxlPVHhelQSZknA4TEqw/BfNyQW30Xypib6yG4EBtvT1ugpXUGZ3sbZaJo1vNY2C1+goapKL58UfeZzF47mbbHVYdryA0nz2VAhw4hFgBpJ1z1El+jSrRDNRtureekPoUotOZQlkqtXcUvPVvW0u7CDP3s/uCBcmQuwKg9csiRb3sJA8iy186Yij0hHeW/f+7xn1XrjCDu5Bf/BLCwrgfl61FNALGFDTHXNnS76OOGukoQVi1Eyv2TbDtqMS/rqPGvD49cL4wPzASN5AmmeAsbViRpaWy2Wz6XHOU3PIDR0XaOucTCfH166dbD+a8ItRunB5oJGd5kRCqPT0tcOSHFlTLvvrf4yFSeQeSLi7rg7ieHC/8d7b7w5u22pNCbwh47ARlTTDfjibTrKvtTvYwNYRTCHH8RoZ4/e+0TGQb9DTsLV/grQPU13mPvGHUKh+0SYLZRekVnPFlkTMV4ch2FM9x9bf7zu2/EKoYib+BHVN/7sBe6ibsdY1GMtWjD5EJ9M9E6dIEWQR1DqbxkMcTCepk9k+OA9rGjvAyzTm8cIPovoi8d9xf97o7kjcqIjOLG1mrL9zwcDtTQL2xbUsDpg19cCOgotPPsys9rI1Hs6V0khCoTPLzQwK5nKFQ70eOL4pVKXyVyDR2v9txvfXIpzKJjKOOenQKTbLHAbhLCOfo0Vs5iGiCwcMoCae6iBrTT3E24dtU3phi9chhivoWnclW72wZAzbYlNu5adANPCm/DziPM+axyc8QmJr2rJPVi4TARLoS94puSm1MI5upVE2T0YsxXXCVCoyc4Eu7qUC/0d9Ze1zS9ExbBfEv6ZO/qf6MBlqWKNJ66ImFJvG6dTZzZOqnm0pf2pOynoXSj/BK3ZE5xqoBeEdRR+s0PZG8ZFU36sE8vilJP3h0x1gAUZWY1YXSRKPTWn8u2FKj1LDEORLXUjYVpzT9YHW0Sg7rePGuXINDJThHAsjAsWGQSz5/hCOh4nAPGfw2IBByX2kw0lHZqLpryGDLBwhYutIV98SYAZ/liJr4anroNWqHYXGPZmNsJ3whiPtd+kLNLzzIcpCdUi8gxABPeFUD1qCeoascbi1KDIKeQXBAaO9YzdDjBNufxAVSBOfPiOL8zvrtT0V6pErS0Yk7I0FHfwkshy7PciXJso1QTpqxSzNvwgHNZjpaCFjaxc8030TAo6QiLO0Lgp++jQ0SOP7tilnqs04ihfbewwzC6yAfLjwDQgNDqCsifCbNqef6+ZaguOa4S1WT3sK2O7Ol2wyCGmnsp53wPsYyXMzuRXan2JzyAjhZZEngOXgwwT18hXBcCww48GbNBqbwKKgevpJWsN23EwVCoqFgBo7GnNZM4td14gLfBpZ3yoROiNwEFfcR99DNeta/rsHs8X/7/bIjpUmQB1NhiFQoz4M4sxxQOk99UxBZpTjlk8ILEDEyN++3nNNXcqYgy+XS2B4gHDBg2hOkwyxvIwLQ1Vb2goTEdfQX7JH7ZZs1LNv9YX2rMl4Fmj4yTc8XPIgISOB9/iJbjDOH+E0wfwaiGwSSEPL3L9TTIVxcayVsXvi6ZI41dzEWCPxZNOya2wuvKQGDe+lRfbRMHw/mZoe5MLzSknZFlffdBROY4QgJcw29bHjLV4ZKVQ0kvj6kHkt4T916c1RmQ4MmoAM0tfqzrmQ/uy6QkMOmwGHj3DnXqs0Qtoi0RVHnSnLTr0g9ApqYKxBa1AR0grqxJhHqpQ6NTrL1c2Fx4gwJk2wnQUDXIVfDEwrWZ+HFD/s9fYvO4RqEIW9wyW0JZiZEuiViETd8Pl6/9xn1IS+PEvMXu0shQmqsYXHexf/d4pzvigUbhvz3GEoA04TIM6LoQqzW1g8rSQqnZ1jrnyarGgIE+stRQgmnE2bGHWlwahE82bvHG6mntzKQc1z/1wayVNupwDeWYl6fR07Myu1VjYQwOnZyxAptQDOhUb9Jv+bCoz1lvKFPhPEvzOQK/P8ZS2MEqGbOwTk70vDr5OEZAGnpKehUQg+jR6c8nXTPnQkV9p94a9Gji0WPNDDwz0SC8HLja0MNhxQNHODAKj+k2zroYCAxkFzlsY4DbIm3hpZoaWHhAX4PUjo4KHzI5c6Pv/vkmpfNq+z7nB8d2MmeaMAAH4KzHLudzOoGBK001PDn8LpgTbjT+deYGDIlzFcXRuwLWrVLFu+8QiZdpLTRToR95VsTOHsunUZNTat8nO/s0VxOFWUy8V9uguWfFA1ztMD/1oiYP2y7xHhP/tYeQw/aBXThz4mXhrq8w9zrVvhHkJgQQj1lcbyxsRNjJrV6ChZkbjKbFYsLMW5WtcUSw8dtwvcjPLH4/IBFiqnIdobUyz6GPZ8sodE4wsOHfFcKv05Q92fn4EtfXpROgwF3gRyqS+01+9ovxfmVVDjez59MtpdQxaxib74xe+y7O2c5ITEb+jXqC9KtOOmdls0TRg+0msPS4yv6LRUfgW0TAJ8mqiN4nKF2yiu5Uik4FfKm9+8y5/T+Ed0MHrnHWt6Tlt2xdFHnnR0lKW2eZzPGqa2+BxSslBBzYWhWC0jqVb8My0LUJa9ZoElqwH/Ta9molDitFKri0Za6uFU+mvD3TiHphWD6aC4/7PC+u4WaHv5LjMVxMU0WU1wMqH1m+w/WdilQpywsFUIOuU9txmLMHRlLYSPPOJdJMG1gb2cyHIfVou69N1gU/ZB8tFmifmKC4kcxDYx2xUX84m7h5Cgenr/QsAxy9RccrKSYYwMtQxoeEQx8Nt4OnPi8VL+5NjklzH+vvZg/Cmfx8higXdsmiRfw7QiH2FnkiNCh2M+rFmry/3YRhTXeYqrznJv9naHQqh1jilrvEhtKOJNRbw7MaT/j9Xc+Othy/YI7fcYKUDk7avfaVripdFsIXYd7olnVLysWE1U6Hbbg1Ea8L9QJCDAsOQbjdEzq5KrytFD/LeKThTMIOAcRc9P7fVMA6waSrEHwi7aHyhSyUKGnigW323Iwwm7p4eHprgynZ/yZuVcgJszw78tyP8M6ZVu0EbnE5UeaKi0ZgGNaf/xkM4di/L9+adPYEfu9ulQ8Klfc738KTl5Mpc+62n9fzlC3sQGzQHXVKqW64uaaRmfmsE3Ue8d4Jx7dyTcb1NFmLFK8L1lfIPYiZixUtUyCY3OcTG6GH7Y23cJeJZFoTtzptxiLHblkOVyWQjISpVLIF+x0xZGJZ8bVgn59klJ9voLgDyQg0i/0pVy8NJdLoqp3PuCE2KB5JCvQYyb+JBA5m0QaYiMEmzW42rOrl8WK1T8H2u/berH20Mulfxl5zbomUJt8Bs7gf0PEAADY0B//bZb/Eho4B5jHnagocedr8ajB6pcjs01rjIhOYJWi+tAMUn34oogUVg9XtuL4aqULfuP+2JuDOhyTKtg2fVx0VWIVVXhm/ViEGrvqFQ2yyyyWZbiWgCzyiTdq1cGoGDu02LVSdHkxdcCNV/v+DL0wdS9bRlLR0+tbwUzmyS5KMG1glH1R505nqVRMspw/xw5N8GgYg+93whUomdqkYb+HhJxB11PArmhPyYUPXgq7lEs1otHqd7jgeHyS0vfTd93NzIfuVDtu3Jg5Ziv4kiStPQga63Btjwyp8oo3jiaYm78cCfnVg0nic6MlMqy59u2ivQ2rMTLpMAXOb2SqoCVJVCSPHlW5zfplT5bc2zmybFNTG1ePsNJkrgZMVpD+46oioVYHFrXqfKsQCcGFPTOkxbjv+ZbyECOJGIX03dpeC6GthUHmT/+pMpEIoIGjJcJx5GT4ZP4Bm54qa5Tj7PDx8vJ9JyHtRn+mXVTbCo+/zbrVUq6JgS9vo6KSX7163wEht54gdNQct+A1vWBRRiN88JKMxN3TpGsVzwWcwtVkBVZRY9LsLCpNvhezVl68Tb+yQT2I0Rpkk+2euCLr5NduDI6m3nWbAyGudIHJWkYUJJXPbGP/Tv8WBreRDxGe6oEga1zkCaQjgaKlI7eC/nDdF3EXghYEXxzmN2Ij3jXRTo3Br1eBslaxtwnHE7/eSorBGEbj34VpMUMdyF1AyQSn/0y0vsze0ogM20og5rx6rLQVLjelIktAcf2yFrzbLSZfRhv7Lnq+QInZITh+PA9bBbwRMMiZqIsYdsK9QF/QeyMc52ZkikRljDUEQYJ55tSSwQ4mpsLol7p8R/0imDx2tQy5w8+6yTKCLETyCjwq5bltpGx3FZCB5aq+5qnA/HpqOrFr5Fq6N2xieNwvcb7dCKy3OwNPSmahUt0MnkhGudVqmB+aw9snUHI/5Q/0dALau5SFP43B62qHQQnxNfNS9pem63v5tf5VLTXAb/1YY+viMHcV4DQfjI4aXhpmlHEJnlbM03Ep+9q3NGCSxZ85rT75nOxeKC75+aDMhNiCM7e2yjVOYlGmE94oqJ3++8A0G01wJGPURDD92dQnteHSSgFV+YQCJIAPjuAwyUq56JH+RWGkG3Q31lZErHtMqTbJ+MZnLMOhJx+4LSIEzlCwZjkL0ZPrQEfI4g4v1t2oDZiUzoeXXx+MYUym3JZaNa42ziEy5FrSupw40dvrEmaMyyfcghp6p/JU5L/jVwCPu/b4OY2PY+QAR2zimOttZacwjQdwfJQTT/O1GH0zVFLp1sCRIeCOLRwobCiT/fvItZZAHTs1M6ZUoP+XuWbUEVnt+ANwGOJjrEIcV9PbRBoCSzWUMVrJg5cdc0dJn7JAe0CT/E7iMNI46YSPRZEm6YNB/atkjyhYu9IjLKD7PjvEfJnck9vCu/hu3YeRy4pqXdSnGsqrhL+seYklSjbTT6xEpJslV3ORs4QgwQURl2OqE15w2mKZ3hc01QnljA/Z60x5qNzPMy8LNKS7aVxmQqOcZdQEOp7KZc6plwLGVB91v7QkV2yhj8/sFYiesdf5FwtEfZDG//PkxkljKXFqNHDprhGQE/sjkdlaTCDMnMox6jPCaDN7KNPrS2vse9nlj3WEWJK2KdRj2lUSU5+uR4KWtfkklMQBVUcfY4CaKWeQ+JoAKaszFVoKVpnpVHEh1VuHOruXRvVImJHUP82VsbYsgLwpevaJCPSu74qoXi+0hnEJVB+c4zGtAqqSpRFF2ic5FKVr1noY0UtX6BTg/dkBQkaA0XYm3+bhWbrL1D83WhGC00Ysx8Gau7t17SrevRolgZkRV7K8mXwc/lcfxx80WyJghXrzoLHcYaDqVIKeQ7QiC+Yfj+pWumlUdTjmcBsf/e4SWvjW/R3ABgY6k1l/CchBnd8wicbihz6SyTAESVlyv8VUq+PBU7d/PnVYd9pT2F8/gODdgfjF2YwjYjA/5AfuZDlUxj5RLKQc3Wk/rB/M0HUeCoGVmjJTziG7UfksNVaKyUnM9sVY4HYSXWcA3419zKQdAIruywV+Xqwnucau1ofEWMuhNhZC41CCs7ZJhCRtBuXSWWbAiRDGCyCm434vtI03PW3FYrWYBJl+ZLXEXN6Vqj+ppycmwAFGpCwrIL2U+3SVfXpkvKmeKsKOZnpwZ7LEpONfx3d6LIlpbmx5H5Ms0tqqe5ytffhQ70wPnZczG6rW7gvuCCB8/dT3wFWlMlbHDC4osIE3NRXLYz6IEwq2HPps1cS/OmmNHOcR07hFkAYQh5/HJNhRA5t66F/S954u6F4w7x+fvVlQONCwVHyoOkQStQgPSeopxwePdldyOSe0yiH7p6c2D6sO6QroD7u4IfQq/kzaj7+bmZSolFyTPZdhGDMi/L2p5tT+hM3syu5HX367hMNq9iSIXZ/Aw2g4GIhLiPYZihdArYhGP0ZtzwwLFG5T5YKTk1zVJb80N8wDlR309MQWK+zU5hNspwmTJ6iRTnIbysOxbs799z3hpsC9ZYhT0EHAaBRvFwK2H8LLQZuGmz1vY1jfJaGEUAaIJSO7qfAUZtCThYPAaEvVdTpKWcLPer4OxOLlKSQdoHow4HtWvDfbqeG7eszVIZM5roC+NxUi16D3+a2IGErlAaXzVptizNim492aRbMPTAkFrPn53dnMWFdv38F+8REzluuuP3bSlPu256F2ucmDG+D8EnRk/Zqp8hgrrVcOup+7P3yu3UOSdUURuQXPuRhyB6vOn4uLDttsv7Q1BstGeANEbbXqCZ375yHe2pwP89R/O95Yh58GQSUAGNljXVsgSgVWMSwAJ2C8zyD2TwG9LG40Ec1wVdM7PpL2LJGEvepD6rWAm6PwymihxlGWe2Rod91xxxbnFK31GC7Pbf6U/RbR4i6MCc4OdjmcOydqQKq9I9E+65TogVIrPWG2r4lYcW31+x2fCrmThaUSbq+UWJhDZ63iqNlaTGa2EvugI7gcEuqzfl+SKvCsflsCoGUrFkUs7k+4+ucBWzi5Cwxb7dJOb8woGoYhN2qb2aVt5/u702CtCPVsJFNPLKg97SV2fiIr0PV4NY7EXaUg2loaKC6JT/K8ruGntVcDYa4/v/Z4rK4seGSf2bNGJ2jYQcfOMohJ02hPC1nqS6Rgpe+rnhaAW7edrt/4h8xbcA3+ay5KfRPoYOR92a7+/LeZNLmfH6ShoIK4lvXIhlNggMoLE5hXJWbSSbM/kjyk3heqKNKMRwGRBPL2IQh+aGGzIeIKDD4PEdLw8Z4L7ItknhK/XXVJSK9JWfNHctJoKHlAo5lZTmBAG94OCVXEplo2/WFz1kNVwCYaGThcd/IK+UOt5Y8Vvh0rQVF4oV2cK0Q1nWozJR8iD/tx0FH14FU1roGpaGZVy2gFDTWUPuS+D1Kqt+dd41j4Cc/oDgcaHIQ1s/7A0yeB/l00iiaxSOB3FP0LPYrBsl/pXrvJx/PSc54dFv4gEZ1SWdLDk5Y82G5Sin28VbxDQcx2z/Mf12/ysShEUb5jX4qZ2oiVJCVFr88scZn7KX+DqB/PqW8ZP6RU9X+JIYvJimwUfUtbT4ckAZrGzKZncA9EzX2jBTRKIvmQ4ntRlrrFSwJpuKjAh9co+wY8gPm1TAtde7JS4pJs+5Lnw8nMbTD24thiefaZasrNiHTw++cNoAB+ipYIUuF/ye/WcPrnyphR3zadXvNtQTI/tw9yErWI1oCEzRJFm7blxZMP5O067QuglDgZLDHhC3w6X8x1bg3zroih6/AwAa4P1RbnDw0Zpd1gAzOjqFe5iG1yadokstJGvHp6euXrGha4IvoMq/Zxy+qnE+1F3Id3EwyG0y8Waapoli8HZOyM1Xgil0+NtyH6kSc03Edy5ksAmVzG92mnoFeUsSzmEJM0cN1U97Y9rf5QrjY8oyshlKwtHrzieyP75pDP0sJCzzLpJ8fw8aMuRbqsM6mCMbbdwBo+FOn3k1NOCkk3UxB4M0yOTpr9bJ5gGzDgNMOeCt5BISPqL9si+R8mrg50OdKkPRPNKeX4VHTUrRQ2JZZ5nulz4OjF8EH8rOL9HUe/SKphFt7g+N7Br0i7oe/9y2T3o6r8NIzUwIcIbO4HGLg8EN2/RhMhXEB//oMIIMKIrG5CrXhGA9io8puWx+IL6H0LjTsEqN0dsM7m5YxqQRSG4tzCGiMcWDsCRYKwxIFieN8eG5UEQ8XlX5J/Ejb4/R4PFF2cOY85fdQYf6L1du0OHrFpNHpf2SSZ+vU+qIymxqjn9ONxDjL+6ltOeKU8xc8OC7Rb70AWfrFROytZDnM+CBUhRVxf6hK+vJTr2UAOVFPQlo7mNSuqttM0ltOlK2xTSJzcld82YrJS1YjFvVDd09fGuGkTmObw5qErqQ2wYGr4BBx4pXWV6abZNYCF4K1Se2BbeahSUjrvozhMBkdgvdrU/FKITne7qDDMSR8A3R5GCKR7FYgEEU9UdquJR3WQa5KTaiL4FSmoOvq7tRhnx6QWXgX5S2edSMuOLPq3+FqwOSYRqluktnfXFVSWOnzmppmo1ACMRGEf68xl4Z3ErrEnsyYAF4ZMZoPNVcKUklhsyLUPVu9wMx8xJU/NutbfNWvwivLzkdmz9R5o5gNjsbTb1jnEYQG85bQfnovSQpT4EZ2hlzLLoZhXQ+wHgFkpcNoxCjexmYc6CZU7D2OmBz/+vafVB/dJ1MuxLCNr/XnJ+KtszhehvA3NcthU7+N2rK1EEtSqrVp1poaRJcftkfbftu2DNpLn0eZDQe1LZYxhG1fk6ODHhov1UQCnnWMEScPUSymXLgAM2FBiL603BcGa7FvjBzGk+60Nq0R14xO0fwNr30O848cLmm4U0XGAZ27HnxSahEguiMg9rC6m3H915T0QkX4SnFhaCYFDAxXSqHUOucV18UxwSmlrTh81frvaF0gfVa55DiS4m2+4DFN+qQSyjex5XdTOoIacal9zpcrl/o4FqlSIjye0H9Y6bBuOyz2/9Gvv77ZT4jy8lx+rf5XMpgoHd7NZsjed1X2dyVzKxUL1Xj7VkmafUhk454r94AdR2Bb1PltvcpZQgpkxotpSxXFF4ZQGI0EfnRy7+wrNm4yVPZi/h+ByEjZCQf5stp+9hqV8lHYFwGea2VvzjceYbo1nNeLvUERiKCSNP0sAsVeuW4cxjZBE2nPRyoxRKSHWFWTJX6H4e33ypQcn7/G09ygGxdSLas0u+mtvWEfgZECBZR2F9/kbRqzHiNaSpgPZqL40hvnKFB7jDfpEg63TW7BC6r7L/FOV2aiqRYgwoFay9Ej1+G8IEp88WRAxdDOnuIMbAOEVJOaukaSszogljM22sNYFXfzrydVgVwQJtpFU7KccAJfZYZKFSYrUDGlxE3pYxOUnJi9NULMuIERzsITiIClo/55Y6UKBF8TXSyRayUiYPvj92R+ApeaWDQ/maYNNjy1ahpdoR7SHBL+jSAQ5ItX0MnyGROdXTayyB5rPQ90mTEveVE3BdciNOACEVWu/lkCzjWflldKKlyiUbmyHZo4Ov8IdFQJYc14G9RE9xbfIzLCfewPdhdxONW64DUCRgmmFghiN6JOTjb9hqO6FXmMbmZBrAeNeK91It3fSwyOv6V/hfZVNcu/7r2sc7roOLNBoMjT8k31jt3BhQhLdZKkfr5nY8x7jCxt5i8/RB1Jh4/oCQfidkRdeR70+HLL7zomeQ61JuaTHqT1mtzq6EcnR1bgvjbRZwUhWSzE9+VPmuqxwm6ZlbezwQeURXnS688VYGZ53tTdTsYzgfrVnFtGeUoKBB0KFETFpd1PF2kBzz3Ynnd7OMVepzN4cqzQOgQguRYZzFvpufG7SBccxiQKAstPgeKEpTZd4yaCQsGEztvT+RBTfnU0P0TAOCaGN28TUgmj0jiMAQdogETDV44KwpmHxGPXuZEE+oF2Wf0Zz7u1mE52vlgteabgJrEhCoCz14T732105vfStZ/hWPhb8yL0RWlRzN+MInYb2vSB6/XxUUX4pj2Ggye80R0cdXGxkkgIEZgTYlOOiQ/JRjhu8XtTvnZTIyQx8Kn0uRnItF9yKXVBrKVNYAvRM1KVCjT9HkauIPyHaN+j22EDum0z3ONx9jhFGuuoETeQL6Z2lztfzrqiohBp6cU645+tKfRaNmC/9RaaM2khUM6yBAB9rKKMurEH3YsGYNWo3nqq+MgneAtohs/l6ZFeofAqoBUSufZq5bTjhiOJU4jDs5148kZKl8XN+9gVu4n7yvQ3NTBl9m9nVg8Q3C+aNH0G1PTyDnourdJc619/xvGqoKBxhXLMK3jSPDPtUEonIcycteyhreH46FWIRqZwOMtw6qCcfU+1+0cKlyBsPeZlu3tedXQPCe/bLP86/0hCKDQ70uAdYRNkbYPCpfSQLuxY+wBJOljhs63GB7K+03jtaiqMJMJtTBdivyol87jWEl32FQ5Zq4VF/hkkGh7QvZwQcGZh81UA4um3Go3IZ0bzmzzul2PUooIKwNsAuetwqAy8wuZvJ4+kWzOt/ajTgrlAZz6MFm7n3wFXkqFiGUWrQ49UuWhslXGY/JCJU1LkhfYlV3rT2HEBbDdKtSnFEdgjBTs/YErP/HA/wSG/b03XOpOC/eqS8GLnRg+lWd7rS2BsAd6Bx7rKLC8d0F1akPYHoAr+OtuG6PFkGtPIjL+RUWQZXHyOmQAER6ek73tdF2reZb69cN6s1nGi2FDIG0vgvpExtJLBDji34K8yxJuVLCqdrmwOrHCqbu2Foy7VjTMVQa5Lybx9XTNLoi3eYn9kcfix7aXevE9B2fJ6NJXiLnD5wRSDGmd3xBzuYER0lM9h3G5yG1pRYCpIY06ex19IlI6X3qMlHInQ9tXJbgG0YjW4Fz7FeE5JvMJKqM5ncZBR+Q8niiXfV80agqp6Ma7ud68Vflqa9ThUv9FVsbbLIcUGilmV3VYQPfdajTdk//sRoW0NW+OtmTM3L/47/h8QtkI13LDhSfcyFzG5DUotPhmx87JDkxSTKCubfQT098MZgQ8NQJum7LUKD+5O/IH0LBzJfPO2b3Z85ECJkY9rutmLrDG+MCyD+DeL+BGm6+ex8aAzTusWIOdnq4j0XBNFufRxyv0kF3NYO5ROr6It0QHb7Zd4dgHrLGQnhawiu4W1m98IJR1aTaqyydLQ3P5u3Kg3dXQAuIHSZjIM22fhmgMQxwn9Lt6OhLYDg+/4GhooIfkl99M0f1bpH+nKrNO1l9W50vA051pGK5FCSFOPbD+e1yKcUNdTSsHizX8T06nHfsM4ys0gGYWbO51zYT28Z6DHJTBcxwHtbSsE10hD3u6TuMMvEXvpfmGKce4fxIv+iurYLTYizEM4Mbo1/qdN5Q/TTNVlkXw3cjS068fZoxLpuFXsRARa9TQOMA27z3exviUZyV8uez7y7SWIk7PXonY0faakLxmyhqNH7+iXEfCWR4tRodYoZCYfIGHE+3a59ELk6bRLF6fxu/nO26TJyfKS0sFyeSfMOfGnQTasQRmOZ+sdHcb0e1NODkQ8D6A+zz898BKcUfcE2Kv8tUo8pm9afwNtCaw2DEllohrwb1azv6MSsYZSTfGC9wKNi1nn8PT6pIgfYBN4fKpm6WssADDIqi+W5L8UEhVpdTdWliGI7tgMbztJVA5IHIx6oge+Y9WBRolpvpML4pvdYBVKVtJ+6wzAzsYAdd0ouofk2Jl4Vwy4MOshc86nk3YZChC6r2hCDETToJ1un9R2Fu3rcU3jLwH2dObD7TJfuh/YFKvrv+DLt9k1ZAIu8o0RqoxOI/PPtJPoEkTyKbfBf9MwWbn3uKNAwH5rMJjVsrzpLpkSqWEy0kEKXUVUdOZlPXY2PPh/X0Cw2lrAcz8T/iquIpx4DrJT1yQ4ltZJqtXKEjZRy6WZ9OegP2KCpkEMhLWugZsD88QNR3ezcZz6wdoWp6r1BeRWhsjPtuQBbadT/rMuIKUMb0TLOH/9CEmx2AFTX75kWjDWAbOyVJzUn60ywjXA8P7WyK3q4cPRzaTFhNsVSIv3B+NiIfqS8Aa8CZ1qJuITa5UTuUvQLp4gz6OroBwNjL5kkCbZlsPfb1lgF+YcKOSA15W7ieYxPx1A6336E1+8zIJW5YUnaMGOHmxuk38KtjH2jqvzYG6ku4zaHk95HOSI/T0EdEjsv7ve5KrTeRcKMQazLDcn3I6QsfUQGKMuYVNsFdPaeHSkUBjC1QumUbNa3dLMcklvsZxZUYZHDf0T41lbaCb/8YBTqW/+aK2ep+qN5229TTTJfUT2zqE4T3FNwl/zGAzJasdQXRiZdKhnSuPR9Ke9Tbxg6pVSpvqWouRNed+UaHXeOfHU8Z7Urd0ihhmij0RSY+qaSpiHVkfSxZ0eifPdGHkceMEE9dD6WTzU1RVp407fby/ufwVQc6SdWES/dFok355MKtSchf8zWDSQO8L7vdgGLMBwu0O+pYIgLI+i02h+NGUxW6lj9LtWLi+faAE10CalLANW8orKVhmNxcB/FQvD+m1LOkzMHLbn55F9Js08kpUEdWzh33Ju2Y7nhLCuFhLALqwHQt3HlmndDFDfsKoTgeODEjysogY9p+39KfgsCQ19pnUM4/M5wPFngIxBxyNnDIeZ16qycjlM8D0xn0QPvK3adblsEg7+CNED4we7EHtzplCS8BhcxBinJDvxzosTmXAFGTIvSpAceKcXCgVvgxZ23fj2HCQJAQi2IC/gOtPv9bU5QNYlN/9S2hj3eSnR1h4w8P0lWc/iF6YammlAIoUzsh6jHzodiza7sJ8ZB084qO9PbELPwOWbVPO4II7PizETmQJbFotBflbXhcm0cPkFmBZNpwyFFa+pOOoEUGSEn8tzhZtccZ3MgwsLWzWeZVdg0GzVwQ8KnQnNolo9CXCWdWZRXKeUCUtreAFhvYLJjDFjRFJwRiD+neGi+FyVWKtVAdVCXWy53gXW5YaPav/OC1rSySFHe605YjP1E92RY8zKYMnTU8juoCqvlWhT+t0ZTIbwqN5hPv9UHIhfsX8DDJhztSiaoTaD9jHCOX1uyjKhmQtG/Zcvz4v9KLFYW0eoT/Dfccypz/+HP8dq9+tuuq9eu+89PI1kOD5o60x+A5h6yXcRcNXaG5LVYZsgjhCJ9gmLArlaEA+5jAQ91y3Rb2VqMgglO5fY81eF3K38amhcqz96r0YuhQNUFMiYOwZOiQVqqhQ8KxCDB9I23FLkUD6GDdWbH2+KCo9w+qGOPhVZnA/Rvs3bc/T2o+qzGTk+TkD4vxOKcR8nwkTo6hHkr7aljJwrNXBwbevHBhjvMsgaDJkf9gxsQW7vzRdwYWEqOyYIFses/kkOqhpNGvs1gB8cicThVDNCpRXrPSFm0nuhHyvvk+9+SKIr2oIuDSLhoQMY+JkCdDFvASxzFSSlHXS7DpDIORvCx3x5YahNmRO3RzuaYqPZjLD9xHBR6NXSUNHpx42T24eHX9fqzHn3Ys8gL4g38Qm9Kh6Q88Rc4/EgRxnLFWn2S1YjOWnCLbM+Bz/TUGWnRFTDH5vbGCA86R2XTSMoXa63FXPGQRxaDpHzKgpcddIHM+1zwn9mveC1XeoPGU/HlQYOKn4gse5FnPAyjVPNZxbGT0HDDvEXs2NDnsGHMZsKQ/aTOhulLbrV4TkQRB2iu3OKMNhwWQOdN7ta5CmTOwznWyZBVO9vuWnZ/v9wTu+dMgqg/zgAipe6eapMNsDlwWQoDxIPsxxNgHDoke87LKgKJLe5CJYYKuwnwmPquptpKImoEF4bDHeGSkO39xYe+7lvIiYGVbCwX5Y8ceCsIn6LyF3PnyOkJJ/qenHyg4awedUDwJXJaOTbfVe9AgGTEnVUn6KHqk0dY/yR+vY2HVRmY88dvqtL0vwllftVMoj4ITiMrPPI4YlGHAsg3k2Sk6XWCK/vQsYdEME92UJZlTvw+UrbUzLSLJJrmoJ
`pragma protect end_data_block
`pragma protect digest_block
7d4a0332ca821d3f3a4f171fc528f8b0c2d55234665a694a39793aebd79c5114
`pragma protect end_digest_block
`pragma protect end_protected
