`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "4ba98359e4692c808939c2bfb8d818da"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11469)
`pragma protect data_block
RMZCpzX+idJeBkw/gMkg1aqTzapSCQdM4y7rQSNcJfTrRqxWP52Wc/kuMUjQcqEOX6pEvHVkOyqbMC4yP/AJu6oEMm3EZYoVambswQ1bML5ylb9L8kJzPRYvLeYRLeYVxMHEzNZFKjkHPmIGUBn3wbkCrmUrypPkGFfDBeGzEK5Yhz8vAKo4KDeS9K2Cfaw1STAgMMgmUqe2iXLWcMVlTBGsRgZWSG+fx7RCE1O0FoNWANE12U5XTK2dDWAF4XZ2ntdxoMoHSbsHvd2KGXlgG+9uXBYTauTvTsFBKlNi8TRbs73qk3IgX3u7BaUPs10JsdwIQLOa99tmcdcl+Wbcr0ZBOufOMVShOf+Udv0VoDdvvaBzoRXRYVBVh12HTZ99edkMoWaZBYK9eiVuLwBoRMSRZ/Eb7qrS2ALbJETZANQL8E5h7d518dmricNvX7LWyyaOAk29hU6x8uSN3/HeSkO0Tut2ip/xYh6x1KBNRsFyByFATl9+Kj/LV/r9UsiNQ/sYKGsf5Y3ChGn5LzZqNLbRh+DQZ3yT0m9H7GN0IIbE8fMiHMd3jX8iZtHiY6nTxvYWOsJByTyNw4oI286gMRgfvX3wDA5VssO8W1AOVTtjDj9FxCJQkN6lXhl4LeCqvUvKPNfOfRVNGvYUnsuLHLWWk7R0xV+QS6DN7vvGerIX6oQsmf6BYUHcDo+w9p009TZHOdAuzDJLqgeYluZzT+KWQK5qmVYi+vgTMQK0BIH2Wut8kz4fSXP/a5jECz4TYMWv2qhSu6SVkwoDa3+xLK4w9/uaeVEGQ6z5xUi136nlvO+liEgg3y9jXcBVEXpv5ZdYEfEfCS4iGuYS9E7k5cBWkev1/TQGIP95+oDHpmjlF1+WMv2JOWEmk5BT9eybZLg2eunvKyqPcwr7FsMx5oXj0V8//WSIdbdqADHjbLjlcuCyQufvAgiM5zwP4OY7iz/2p65KRQVbt5JBb6KepaztSVlWQO6ICiFmIArFK385bmaUPueuA5mNjPu8vSEuYD1L/OmXYBNIId5542f8vW9Q/rdlawy/B/w/NSTlfWR6whxtoWvshqOuYO7zcsmTovLaaN+RP9zk2vhp/2RaYTbPvGAKcuyVZZYjyLGnj0v+9SYmnWItGllIOYJor6RJ9EiO72sOnKthA0SbCpIh5MYE5AbATuMyBmHfRiugsp7LjZhfJfrrPKEdoqyaD1qIjWwQmb2iIbTVzWkwB/QJkhTrGZQxV7LHrHacB0n/QbmzaBgn5UL+CxrdbDXarnoaEnROxmIbF5oMZfnEZbyv1nXiHZEkjAi63VErI3WmgTe4teYuYp9T+b7Y6JIMnsAYn178BsarZkK6+G3bwZABv1/B8N8zbeTrwmRjhlupyhJCG2PnQT7c5DFTrsmmc6JOPUL/SyAlN7RC4OxIplKk4Qg15SspYQu9m//NtRoPOAF8Ij1QmQPaH/wztQ/ivgSpSLnzeIo0+K2R6pO6metNlhSYVhbVIlHTCHOuPqlevRPWoHooQjFSB216tfNhQJR5fNsbPGIfbi3P/FMPmllmvyHj5J35FIc9ryxx3T4iwuW3uvwgsk74IKeLbVdJlj4cjdRYJCOYd5Nx1QlP7HlXH3uZqkFcvVQGxT75D8R0i7BfCkkwmTRCpYy8AfRDcS+hWcJahi/ZYRy0fp6q/24aFzrNVPtVq+UQsntDM9691qXwLdWSYrCgDEWtoijvtnF+Q5or5PxCHbzD+gKIWR8RgLgcH5aTuYb8TMNwucm/F3IjeU/v5LHABI6MS9XszQ6/wKTlsdWL2vUhqnqQaEHDY6s1Ok4+GYn0FulJT5ktFyxZTBIrFHZn6npFDkmFUoS9UrKCk+FAfpsMTo5+7kP/XNJw7RvAJXH0XUadE0jJPbu9N6RP9UP8LBktqQmQX1sHzX6eHKLX3U1J+YQO2OHecxe8dTZGWZmI1z6sBPivF1v2ZsG6fhmFvjPYki+GQbJk7ztALkHyCxkVDbwjMsknvzP7vfNeikBEBHHHdcIG5ulxLQhJt6bWe9gd8wBfq0mTuSyMJllSrkivrOSi8vuHqsy7S1/oCP9pVjaSbn10XOqp/9ZnGQaR5qvNrCg5ThgcXY8LQbw1xZhP+TOpc7U1qe81sxJHbfoN4II3Yr9V9AqTSm5gf7aIeOxx/6+X8L0SUNoLy5Sq3L/Qs+3zKDz7b1bcnkPqiYX4xw6SeZ1wRKMqoqWsJXFc2uDSYlOHJI9DKTgh+XWCSU0XEBAVKyZMNzn6c+VK6vY0xVdo2NK0ydVxJqZ6VdxfRaa+km1qRmHDhyd1CN0nSHUw8IWmrAXcbQe/oMM9Hbc3m7E+mCXbWXBbyJ/HqQrvIKZWukpskr9/AQP7KZXPv7JqhgQ0+Tfy6cXvJ0pI9MoNd0++72dM5qS2nk8jRkchUY/rxeBgqaPl4h/o54mVuWhrPe1ERzZnrYR8oVHfRZtldtjw4kne0zCwcZuIykWKg+gEquyoYr7XNnr9H7I3n1LEVc1zCkJg4yPmlLIdtAzeIve0J8kE7QuJxNKtvKSVczXw02ExWt9+HxzrGs/QVZLdLMtyeqdCGXXx3wvrUA+eT4QgxznX7WlOqithxFsl7Ixxz8iv2bzuy0wSiw5byYPU/6wIIXB5yDH2mauemy0afGeS5TZDSFK9FmWX7oEJhwITnDgUk1srhHzoDXNuiSh/FgdZYXZhcMwk/8rWfd3XLSYeCgfPshJGGWg40fDK+hQTWiPkqhRG4XaBFqvIk/7iL0AtiY9WvU5k3aXYzNn11hLpLvhHbDSUOFkjTDcNAql+c80eyu0ggIo1L7VDuBcvVAFuXpuHM/7AZIyIp6oxmKXcbuzqsWRLPglwl4ZqOkLjp+BJkU4r7NjJY4Ti2J1GMRGf1xlumMJZosOF4bQgfoxvL2OmK7VCYZXhCIarPZHGeeLXDoJnTVWcJcxLSwV409k2r5/t3M4vhC8ymM94tqdqd7B3/YlIn80TN+v7Bmqv1mjDXhylltlwNaFnVpQSekgV/U6ffy6kHdVsaztn9aLL316txwF6STrdlE5wCwkAHlmcSnYOPe+f4YJLHHwZuEQw+QGmd+Q90U/zuBJ70sbx+9y0K/H6W1moeOaPnpRL+2+c/Ln7LJDY2RRbgo5MYbrnno/HfACE0gJo5UKhT7BHwpvd0BUopBplSI5ENkyX8Yioxnuhr5nQ0zxG2CH01rbn1db/Zv2L56DFH32n6YnapnZsWnpe020Dk08boJcyvcy/2PdVXzb5AUBNWTaIhD5O4dVV36j0TmNqrxlTNNW1yJCCIwUZY1t9sSWiUw5Z0G5E7E8KbkOl6FhzO5uYpSTEv555ADM9XS/1uyb0aTmlNPDEThhofxyJLaUzw8hVomcMW4w69NDEDQ53I1nEqIVjolLexgdpsT1yC8kIGQDevzTisapnFVozTXcPS53mqYxAse0X+HCpvYrs8xUcwH1+GqdYmAXp4ZSswcIBVI/eddT8TFr11cmH/NVaYGmDwbzwjRyKOufk/3KvSsAeY2iNtjkh5serJVKgPFZbeala5MdaGMjqbs1vM3c60oxswwenP20kR24bFePrEJJboPEDwCjUDmk/sQMoEkhkG/qINY8QTJa2y07P3oy2elWccDK3UmK50pskpcGsVF0ItHg66WFzhbdr4JX4fcR+eN2kgnVqtSZbUKaH81nTh5tp5TQbYfss8wWaJC3ET4OMGeeY9FDyOTiyp/+3MzZ2RTr0jgh4985HLb2iA5K8niEyIF3cXl7Xw25Gs3TlWqpREm4LTLo9rQt+3pPCueIQZTR2+tm3NQ9ZVvSun9V8PSZedSftDZltyTfL+kl7bPmVHIowd6bgbcpvGlvFX1JsGVVgoKKc6KIMGdTfCqeV1sg9RKkY3j7Wmwh7SyEiLURdSeE5XLIH4UDagISvcrtnIdckwawx/wH7cucFv2TygD998HAsR60wTdD4YWzKv51PIi68KFVI0KUkdm5ksULsGQ+TsjU0fJj7NN7rb5Td/hez79RzEZiTVCvIHQrgopy88+o2jfz5sY/c721/xXwHlyZbWlqdovymKno6Bx312UWuBs7aP2fwWxp2n4HVXuktKAXLJcvxC6IEObjGk71BldtNtRFSoAYnur4abPwBaAGblvMj2236GkaDj2wBkMAOwOSv/9OHzTGxGVgFuB2XA1s9Ta6tw6ztqrv+wPABUz9gFt8ED+QFgtNw597Yn2GrhHyenRuD8tvo607b4yOu5I4TkF9a8kIDPd+Rsn19nCdq6087sPjPoQTqgl4kjM29NzUkboZSbRFnLXJJr7MLySksqFlk3+YG+aCcxs0aNeIsEJ26eoUFuyoNtAj8WNJJ6wQ+S5qin7SegbC2y9zPHREqPf2o9BhUP7P8h1UrY+FNRsjD7oFuPuob1BS3TxNW6fGft5FCXmEqZcmLas5YgmbCFrU2nStCf76xt8zps8OuvEXQBCxYMJ50W7Y7rc8HG7nTCPkNmnvRrMySApYs6N4d8ONZcrWQofbv4uVoNWr97EVRuZsAvNl4G/3ulX8GMbJ9bRGZK5CJ33Q5qxbxvWj7duppePUYqF152ISUca/IoEI42C3CbYdRyV0dgIPDObhT8Haeh9VmE0aR8KH1E+12JwlaG0PUEdtl8b8LsFBfffwvtZ6mhKwW4QOMOnQFtkb+va6ujtCYIFmjd/07Dinp3BdEgBkAJz7ZcMEQ8297kF/mYkdE5Wx38SBjN/S1vOZHRUQtci7vBbaeqK0LNC4g3A8YUxwnKMVxT3l9+dnu8hWXeeHtYFhvgJpLkpQhWmpQNMb6Ms+oUuQFWzuPeUQ6/S/31X9Hyf/6LE8TPkD6sVkoD/UFkQewrk07qbuqOgDbies/B2CT1RnP1dMZlIzCOe2y6QDfO9wzI8RGjGg6gshbcgSwAB+LrG+Yi70Y/gfGODsMRt2T8nu/SXXhLE0SUTT8nRJpw0yo18yktpMFeyYu2eeqc+WqjvaloVwe80n4nYos5PpSo31m16z5niw2x3q0FN4ffzk9dCuTe7QVmWLRMF7JBupb5dn8+q5IBIxlqT9dLuIrrVpjjVRTgtUUXYvRsNbYyO0eA68Z3oBfh2DLlEAKyCNGfdlZiTYOfyaEgN8r1pVv8i8z4L1M8SQjoSKYhKAbJlKBfAo52cnRdbSg9lpDbY+5aKrP7rq3f/6nBIhV5CXFNIp7ZG+tJJztwK83cL10Pfnf6N1TGDUqjiG6LN18hS1bJ1wagtcSENZwq004r426MZSqXfD/kbJJXqIOeBNSx0da21NQCCKBtSl4aT3c9dMqoXOAC8dc9E5Buque/fCaCy5IiJ2U2QfjI8xuaQ4vMDk9Ol1x6VunPmP2blFHyb9vQVsb7SaTRu4yy7DABGEX0+3nF/q7xpEQgMBt8ZNv3xKVAJJqhpai38F6yH1UIi5GJ1y3afsscLPciUUAAfPk2Bzcuza7CwDd5aCbvarGuCJ5eajZazXr1olDgB+L/X57wDaQHAqqKeZgR5hwVVKy5a3ZdufreGidiHHYaHBFJQWughYki+v/cLHaLRr41VKkD6xwaGhX0N1ruf2Fag2ouCsaplLMMeGIzb6F9iYSbn0/T6VQDqdAYAc1flfgVudurDMqMGhROZOl92ZcZ0BUcgukqAA7v4/Qnui7O/9hR3zpWm5wEikvMcHIypL3A87+hQ727rNvZKUCN9KOG7LC8l7sKUBAu2WvfPc7474bYttngeQjEj5B9q/6JKIeRvi1TaKEtNCmzfPG5vVZi0pu+vA6O1b+UnQUotszSJCopVi11M2V2TYDtlYbJge2TxA7Ti6zZWEgJUKMCQkh56Zt1LvokYteKpIJWjk7MJiXDEf3kzstU0gbDIw0rjJG/tPfSMhQ06KKUUKsNMRimSDJAiZWRHF/aCq2vYfh69bPVCrlwr97PVewYDISMX3BPJ6pW55gqvjuBb0oMKcpQPTpB5c5K7Tw92TJxJ/AWMYjSUQ3qqkvsSQyOPiXMVJt2s0wr9fJKT3xDDEP2rbicPccI19/oElH4rtw7rKclfp61SP1OYpp75cMe8ZNj9gDoRCwOYswsDq05I6MWdRPIMCkvj1hcCsVZ6qASv2a05i7inHjUQCQaD0NkGiGHI9w0ynL8pujiwyodB2FvOIAuiKKexfjpYu2K/5DPT1i1Zc3UOqcUi0AEyrPJJSvROgOGiLBeMp2UZ2+8MyRxqDfzQlPhH4eM8vCM56HP0HVtZ91IT7Q8D/Mcu6gCVQts5/hdM3MHyeipS6V0fskLhupdb1Y3w0W4hZ+Xlh72Jazy+3Up2xwD+kI2qrG8oDB51rMU0VcReXxRqSITnpfocg9oJybZS1MOB5/MZ196CfpTreq+efMCgEBIC4aKI655e3J4I8lDPLaQG8UAGNNAC6+dcrsuiAGARUANg28raxiKx/Ciwgh2YXKIsYrtejUPGUZVa1DGPNs/Ii6dfe40UvGZ+3B9PPIh581ihKxLJRdRcxAUTO1k/KjFOxxdLRYrrWCEOAvpH8oXaXY5adGYQF+xaJuDdge0AO91lVBga1uDcvIyhgxQrwUXuTgtkpm/RrQ2hQpfmEeFh0vQpan+Z+ogiwdGDtEKn65IdjFAgV9i91TGo7V4gbmzjdk26+jFtiVcgTQ8UgPkFyrIf5DHgncxCKekfJ+40aS9ADpshpRx59PiGNDb8vRRE7ecqs8nlX30jEZQJsvjf79Y5XN3hKSqcw2a0/K2akZ/tIC8QTS4PhPsDfcB8qnmg1/CJsRgExfuYZVjJHMzIfY8qUiOXuN6fYcmWBEjWrfxdfiJUI3zp7yoEBXn66SV41YGN79SZJcWxe3CpHuiZRtspSH5R8Nwm9SmM8WN9+SrTolxQSpVzbbQPLdbvzeiN8yXEmZRX2+pDbvYyrX0ffdCt8Gx/WRnOgoqs5cQMK/JMQHVzNBRC6VxPoK0TI8eduvp+RlI6pZptjND28TBQfYL5QeZTZzzlrWUqxfKQQGv3paOjfwCTHGkFpO4hFpOTQ8tgL0AFDGF8/TMgNcOiHI72XH9NB0AV2BEx00lyBud97TD/IJAfUrc/UfTQqe7HXK9JvR1EnYxZ2ClpkEiLSI75eQB5633c87dKa/kDVgVe9dO8ANaVTPDzf/LLMSe2aBqRsuMCKfYZzvTLdohSmnZHOcxccJGoLlb/JHxdxfemuNAoHV8Sz16K9rFoVqn3ko/13ewlOLQc3kQHp761D9bSE+EJSYNuXTG5TqqsNhTur3q44SqiB7rqf8Kr9F9xLdWpiyTpOUfmuNEjF3hMV4+catYjkHsChf0gJxk/SLE6RZcmxLBpcjajj5Tt9y/XPC9J93PL0d7dnGtxDeCB3y/bQfik4Y3uag2viTcVO4fhpUurHb3yPUBpm0CNE5yA65Pe5r9TejLLONWyJtX3HAtQAF8rgVzTrxXrjy12NxsKYeH8ryKN1gg0WwjCXbzAthrVpZhDVlCi91qtf5rXPY6S6YSPbscoq3Tmr6qjr1wCMQst3r9QVwRipdG/VURMr992Yk4z3YGoCBQcmyRx8ZTndPIrHB6m6OOjY7+HoAMFTUkHEKfkW4wgrDi2zp+6iifYgrhZugsJdmX7cmJeTzUr4sN1r6jftmaRTHt389zOQUOxmE831NVr7SfjWL4J/hahtU8vN0gc+vcaQmjcn8tneDK8IREZDLFM9KkI9c/nhAYMSuuyOIMaFKiuGmvgH38VcETYcuZIVOWnm6Aopsllbpapv+vCHYVFQ3VeLIm5kvL7lVS1YfRF3uWBDUVjBSzd4Q9qFoYjej0KCVBQ5YNc6cGLKiVqGPsQblJJefFjfGVb+LwS6emIS/xNte36zPEAYvwcToFyeQRH9qK5sp5LOF8bSqfF92Y1ZuSSHVjzKiY9j83aoMnfxDyfhBKaxdhz6Z1tjCfx8d/rQyIFIDJDzffzRx05OqrNoiSpP3B5jgA/7FY7oHq0Lk9VCRoeXIdXQiamNlxuBIUOYXz1yn77hoxPOrGEaaFgvwSwslazoSDU/mnuRoFgEKGyjD8uRxe34uVY4Fok6R4jdY5ZCTATvsquLJRQ7dx2iUOJ36NY187NOtAcAxnjMdRrVNm5dxdJzE8R3EMysIHFYmH4HSuop37GRhBbMF4I+pTJbHShZaQhxXNFBzjecPUp+HLW26qAi4xjjZj9/vpsRRwT6AB7QM1zg8X9gFJvSQh9wQcFKtfxSLHnCPJQ5fq+QIIBAVRt27wU8yDJSTpf9lAiQJ0Y0NrFwoaYaXoUE5O3ajPqD2ZfWjv8Zs8O9P3Y1PiTvTEtGJPJElWV0eEcjteahxQkqo1oanOIu9uRcECEHOGWJtFCFHfISeRw9RHthhYCLIJclmwhx3HHjEDpGH/SFdg9pLmY1Z73LrE6XTQAykN2P/P6g5UwXxWY6qir7t62JdevWnYqZrIMWRbUsXY/vD9KjZm5k0UDlMBecFKp5VrM/bNwZvrABd5mKQ27DO0l9xEQrWO9JTNgMfz4E/EW+/Xr7ZgqCgj+P8iF9FE/0P6Loa/YENFm6ktVDt3KyfsMnjT6OY4OH3jCVVu4PW35hzqdbyYQi34CEJkzNn2V4W9gB9jEcOyYjH2EiCDt0wlNuvYT6P8mbiqNSfchdxjIPOM6lEX8nKlRijhmO0ZdoxAmulOhYaOyM6HP0qnzhmIhImCI9ZtsDHbzVdrFoQ2ejHtrOE68LsC9yCqPUtatzW41QKAetrQnSI+r0b4198nq03ZPE854T82Nw0RdwLmmfB/oi4936O5ljR5QY455uEEHGo8qqmW1m4rPNw1DpLqreDkY7d5Q93P7TJS8JZyfvJttJpvt224GAam+9p/kN1H0xDhDjG11bl4TV4eSLY7zwey0SJv5joSSAiQDGTGN34+6agF/GbzbgM+IvxxW2JvBdECuygm0iqs+G6ltws4rXxU7OLVDZf+fuiNbW0715DNYizd9mJP9ESaS/e9YDDCbTvXJFEAZRUuJBK9S8p3Ikf22ijWpQbVPKqJmPP0iEBC4c+wkhhlxMZYSAY1yGG3zqMvpoOyaQHUrLMJNrBetTF/LiQY1JALojor1YRnXzCsydMlTyK0UHS8FnVk1wh67YGakjauudoa5gOSiMWAUsKOy/j5SJ0Kv6J6vUj8rURW1IjeyB8UwJTaiy6aDMfef6nIqRa8bslxKeIQFHl+6NpinXBRPOx1R7jMB+Ue+OdwMjmNpFLf1XwQc2e1NrjzVlDKtHZpfh2Pfq6SwlilXTTllAoxUFlnyqbk4Qe9rckayHfW5cp8F4HgaqYeeh8x9pKOwjlGzgipYTz5yS5tuv67sqfvJJ3hs2qVZOMF7wZRXeoI4dGR2vWCn3sSwhtW9IeXNZuRQlS449g3SxLywg9TTCg4hbe9GW6THoCvNDPCKsmMVUzDeDoyC5aBfiUXzY7AlMaloOb27yc2tt1ENEq+k0zfe+65x6+/arJG6+DW+MRqGkQ4IlEdbX2gaK+Ifsv33RqAEtYDY7yajuUZ4uHg1aNeTDhGxLR3UvQX3f3v0h+0pdozPTTIKMH2kDDGzCHN+ZV+IWmra5AC0b+X7l0mFzOaaUFlwUfMuBodl7oYFpTcrkQc35XtXCORgvmwTkwkqEvgGmcB465dWm/M3iTOz/M6Lo3s9Tw63c17giYxRM+q+s3IdlzADE9yEr4c7sYhpxwnkCaeGyzym2W8SXj8jRLeZf98FcNERqfMaW/qdAryACahMEQ3shLuAQt+ORa8bg4aipACbkPMSD0s4IZCJLGZiB1QvsS28fOf3UTOpBKYAeb8KnO9v8Tx5LW7U3R7kOCV4GzBsEqqkmtlOS7DAJcYlGfWir9zoe+MZytvM3PXDfyLTeN3Hc+k0xlWybctJl24Gz/p3rB/V2mcfjLTbvOTUIQrKTk/MBFZg2Ucp7wQUP6oO0fy37gU9vw/o3rOj5iVixD5+taXY9GP3bhhcvlenO21Usmm5Mp+Ptiq9xvkj+Z884ollS5TlI0E9uZslhkzqcUXjm0wP90QJ7VriuizxQrS9h0ym4p8bkCtb/kj4sdupi1fyiYMO1FuLl1j4BbsCzBxACPOAkABTkusYPmMBvXZsc7AmdW7RyHA0jWnWo8fTC0WQNifCDgaNSi6XiiHAiP7S/M3OPjRRJ9dzbZJ/4dws6WzF4QQxccs0R2bn7TwZPcJm3gy7fo3IeMo1bmwjCk3fUTWYJ0clyOmKv+v3IiXFyB+eqn21bbbEPVAu69Tl5w6ofZDraStaBgcKDM27vQcNGpmGUMC5r8MwtcGyVmRVLkQVHM7rCmBQw9MqoC7CXLHyTtmoWhpRsINuyGXb6/2w8GyUJf4BqEDTsD4QrUOTvv7NYBTPaGxBxLBCpocCxH7ycu4tHQafBPHxOUQgyPUEAfNLy5OVKAYiQMt7irUyL5YSkVtU3krXU1onizRijK7iNaNS59K5Wu7tIubirDhRxiZpC9Sh//Cv+RFNFCm0vYMje+4rICR1cu06b+zIkNYyXkRf/FHibgRS1GXwsRejQotErR38tJKDhhr8ytTM0dEfs9niW8QbHZ81W8zLLuYns4h5JvYxc7RVYXRTlGzyHL0SFF86AKwiX9zJbaDVNEljxT7YwtijQr6X6f5vk8+l+0JEa1wMm9C1mxBPa80mdQAkUCM2XhyL2vZWPpFA0YH97p3LNgzSMy9mQITEJ/l3hgJ341Db2bTGNVhfynZtZLOFLcvuHxDXniMdoiZnp7uvrG4yMmRAxJysUykQE+nHWu8uLWWmkTrASr+/52JhraYenFcR6aF0nNcm/CDDmcWeUveHPrvMPCk6IS3YDoW8i8/5ll3Qrj5JbfXUnRj7u24QW2zkmltpGIZKOfEddVQsdnRtninSMXpEtUvZxumzqmlWlEz2h0t6jRDF2Er54K1WZcGcWNNJ9pUpeGNNMx6TL45gNW20pNi6n8fyBWgLDI234SP4tlZQlbAJ4RCyH0+Z6aT4KM7z6T6UUZ8eYxjzn5IirpW4ureO0yhshcNcRXYNVkX9cd/h5ViFeFvOz3HUSJf2RJQucE8hbHrRLU3i5cHvjQKMGuuaFLMNxA3eExVkrFIsBdENMyAS6OB3oPGADetnLvBPwV2VGcaAzMLSY5/Yf6Db0OOeE63R78mcS82OOL8FtmNB1WLaJ3lmNwpt+sUecP0lb0SFjBxjambgicwrNvR+NHUv/5ioeKPxeaW++ZuaCXFonFb+i4tq8A6tilWWjTb2zTGPDeFXh704YM5RQSDpILj7RuFOj7S9xIKxKDbU0WT/CM4mzgi7Ouar5JpukWaZN/RvNW4Wl8MK/qWww4x5nzOlrPCbKgPuwX1FU1sKJBSoS3qbKXAhL2rG9yzjRvsFDnCUXNOzF6WAokNkQm1TBgbGijMNKNINi+pQsTBZn/HHy4qglxIgYPQpo7M117GChePwdmTJiw2foaYYOb5oC/hoNBdm5Vt3tjPIt+TfFvk2DThJ6mEWfZ7L9J7Gk/QbP/+Y7SKB6rxQXdRFO/+wgE39AFlljSbYNVZ55RzQzC4vgwG8M+r90ikKzcB3Iu8f5mswysE+B90GqMGvCGIhv3mb03Pg2wm1UViDBMihYOMajlJ4vTxn4EWNYrDSirBx+zgyn+DjYItyeqa78HBlu8m32fvbq4djrvkOuZKKT4UyUvenOj9wMQRbX7P6ZBcGlzb35LMFy4njR3MdAC4rCj8IVwNMbOGU2P2lH7Ru8PYSHHZ7SXcHnEAV+xpVQN3yVZU5Rw/K36ALwPhmyAj+GKaPs8pyFF6khjaofdHNhehKUtikLC9HBjqQyfUOae90E3NOcfcPrNWFUpPQ9DxznbyyaBppwYKeRQIMxCrVAbGadtqBF8+BYefXYKGNqIBaup4DyQ4Oo73tNnhVHxLCFfrm7nxwIcA8oVSn9jTw8SXCV5SFQMERVUWcC+xXSal6iY2J3lRHUx4DA9TjP1w0pxqf12A8th8AFT3C+YL//Y7E6bCf4syD9qAVTey+H/SMRuw14kesyidppLs9mF1Wr7SM77IDMkbbdxU+G/BV8q0JBwxIKjzmDj9W9mUZZV1fHWkxhf28huCVUqvCLzp2nAYp8/1I1bcXFrXGDBhuKwTaMvIuosavUyEJrWNL6es0KYqD721hKU75p9qIEUT39fvyapL7t5NtrPTwihqpC818Y5vO8HThZoPwj2P3WiJcvkENzPO1TZ3VtTLrWSMiWo1uHvk1Epv8TotYGlo/TAnCFnS9wQ46I+NgV652bqdIO5J34P96c7/b2GZiiymHXPqYs8zQNyz8v085vpdSDHSiIed2mfz7cMigRFmG1bxqER1JQrV9uzDxZf01p7UweeltKkOx7howZZXiaugIXCj9Wm1NUNfLY7DN1l3xGw54zBzg39LWZgHVoiRKGyBn2Stj4KOLCk/PRZrF9GPiTBK6SbHkC26S1DfNOQrLN2lBKTMZjVI5aXdrz0DYJVT4xg1ISn63YW0gjmg6FX4Kiwbdtaby0ebqA0JXocXQqAf85eA1Q4SKsnMEucEY+Qocv7s6hyndRUckmcvSpSiOuP0072qt4mY3rfXi9XBK6SC0by6+Zr/R/e+2pkT1ziD7oXNL3YIwqbK0re+9RXY4Zthl7OcpHPk985ZnicLmNE2dQulkDWwWTyHtbF7yFCghwX7wFZluZ4k6rU2rNxJRsl3jOrVY9KqqYTh4ATe2K4+ck4ot3Ml3rDtKfFatbREATrVUdcs/2AhoiRXK4C6UELDF+AdssQlNuF3977JmQheEtXSAiQOYUzbt8SoHm8V7TXwMPzFkqggd7+dPQQfALAcICiji8b5TyRIxIBLKHgp9SCwTs0WjJzS54r/g165FMu2JiDurAnfsLhhYV0KeVryGBqisjoFMZSQXrbk91JKY0k5ScGdBqEsUULf5Fgj5pZlXNend0/vOIocaKgJlf5bR9+0zqA2/SqcKe3nvmBOPJSS19iah27H3kIoLl8sbjTaR+l46WZZjlZT7AB1x8iQ/4ZzxRh+rTlJcbc7RCf0UmT4RoocWOOrqm5z+8eIK6Nl0rwBRklTVLy7JdMQs8ZlAhI+gj/0OKHfQq8FrsHhKjSp4GkTm731UHWw6DqDvEGttzCs2wKWPL1Y3otc02J4jWsVInYfz8ZH75uAoa7qsRXjndEEQYU9B1kGTLbsVK9W3tFevr4zeOe74GhTnzZB6zkSLWSCCM0LrTiHtuuT0TvgJ9/Mw7gF9Ire+RirBWRvqizZkYRa0oJp5Wh90rX7GydYoYf5R83jnDN94AS0POwJbQthTfjgf3cHuTnjB4oGIsx/806dnifT9YPCT7AOAphv9UVBrfD+M30sFHOnCVbCV3PcEFLxYvFeFidC8l82ksxjyvHStSLFRXihFWwHYsk2v/Uchs52BCQn5Xhv2Npujwbnl2EFtX/6Qc+bLSpP+HcmcacbB7zKqOa++Ir5GfbHwUz70sVX/BU3bK/SKkXTkPmiSNOF7zm72CE2xUV/dpPp9YBmBObAlnOEceNX/S4zLZpFyYQmUk9+5gStfWcTJUMAq3unihBdtH9C7PctJS/00k7kRVOQofXZKY1R0t6Jk/nBwOnioujXgIFKV1do/j40AQJB/SO+unKhNHxmwBDif9s36sg1OXHoKHEM5M0H9pNrO3nUGVYih1ttBUod9rptyxGlyAs/K0Mgv4Bi1KBM7jGMA64H+Go/qwH85uVmZXMZamjxouEXaZflLQEjGg0DEanGX0hvLhAZVTVt11wa83MDFmWJFaRNQDcrjj4jCbivAvL3//F0eH9877bPweQQEeOeXH2Z+w6Vs1jpxRthrHLJMj1pk47pOer3JKhvPaoZ7Uc/y//WpzLiTcT3jUpyTOOI/toSAjslJ2AroBv5TNEnEpDFvJGvVgl9Z+16qMosVnvEvEM66HwsXIIhgAbSQ7ydOmljefbIfIVgvyhgCxPkmKFJT321z2ngmnav9hBPHJpOVG6Ql6Sox6NjagHIM+1fEL7GbJ3OJFoFjLEaNg2hG4bGk6t7bdzaH2Aq9qIN89OZtekGT+4M4DGOpuHDf93a3Q7DvQj39tgtrabXUd07k4vTK6nl/RgOHH2kc/WozlH/CwZfyeRPmpVx9Bm4GaxvpsmP9hXcEVpCP2aVBI2XQfZsm4FVzgt4rZr+QpWyfijOY/i6H4fF5CU8rpPrpxeekLax7T7sVZ9HW1conU3DzSBiDGEnzpI+x9MLkyozHO+JwnD56tuoyBzpMSlF9Tbd+6fbVUPEqBKTfngGZ8KkteA6cnXdns/E8xIa5U94y3bx2xvEMXoiSQFHs3N0MZ63ou3AeXazLkMht/WvrsUzhKWYqIS9AYPLFkKlnssTV06G2oiM5r1E9AOVGsXEPeZAAOLVoLHOam8YlfZ6UOUqzqt9SH9NcUfqLQrtsZyNbyKC9jPNeZUqowjUx+hWU5Pg7e5JkkF6UZu7VQbrpkfGzgWuva0NfG3230f2E63l+GWuEZ+azEaxLPWAgFSeGZPv59NrBU8jPu4aAiYSPk+rbW7A2/u08cWoDvzXDYPXC0LonSbWBT8xzUOtezEqm9tCpSBilwm66uzJZckKHQjxRal/kZRsQ/29Zn7KHF6nH8dIOW5dqIC20+quQW6YmY+3GcdMwN+MIPgf/z5A/tNxny/JwZK9cqnWiFIWjxkravPvgIMmiHT7uze9YTFZQw2McnBpFVKj657Uy9jZcXPDl8LdffZSUTwWCOycjlI2TUJf6xgNjm/6GzQnLLAgrylxrU71UCSEBf+IUQGaPC0cvMQ6pAPYmPg+XJiseUTh8/c5j65Fqh3juGfUZtw9KB2zf9HMM6o195Ph+W/NQmBK7JQMf9IWop3oNPB6lGHq/2ItQXRkD2uh6BnICIjZmr96uEHCO495xAkUf3eQ3SDxLe7JqPJvQseru91+gyAk9UAAOH3m9uQCAiE8EFZtfRfp2k9Nq1bZmG4WmN/5PqF7nKxQ+b9I/Z2RJDT1yU7oFAq/gzWMp1YRJcFFUrzgQnho7r3tl8oAiGIbwMETdXppmg8IpAAOc7ZJptUdQsHwVGbkVXXnm7sxrvYbTMA1LEHDGGLD/xVbdODS14GqdgZvUaw8W2j7gNQvd/Vc0ap52OExn2xWnhoaV0IfNXYHdqm7g+/A3f77gkYAj4B6ASRzxGpEV8jgRAeofKe6u9e9NoPyCsCp9RBWfm2Y7SntWnDrWQvJBMLj3hCFBYs7Y+b6wSP9O8L7CGYVi7LFNezwBEHYOxDzesuiaWsyrWU
`pragma protect end_data_block
`pragma protect digest_block
4e6ca3d2bfa243849a5b3e1d3bdefdae76f3d159e399c5c9d90e340b852830bf
`pragma protect end_digest_block
`pragma protect end_protected
