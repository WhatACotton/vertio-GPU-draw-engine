`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "3419227e9e67a0445698376d0bc55b67"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 10637)
`pragma protect data_block
wvoAlgnxQDCVD7SojnIr9TcuVV/rpGBSd39N5sSsjSeMmgASKenI7eXK06oQzF8TmswP2WwEwIDqF9sQ5nvZuQ/V1rWWf+Ypzy0T4QyBMTSVXMo7JQrWc1xwUlbRKbMZa6Noueb5LiNKZdcP6Pb6ZnVJqAD7NQb/Y/J1AhbYbZbcSei7uKfGKBR6YPyZ6XHiZ7XaXqh1LsptBUxmCHPzLbKThTHXwiWS7EZ7V7zQOWzvWQlPgLsSawCLJQoM8fvI/ro9yeok4jW/cGDvB+nu329mdgGOb5t9x0MCA7FFvDkJrr9B/z8kkAqZPR9xxdIj4HTrwx3DxcH6f/9MMeW768i8rlcDF29bWii3sEL7lfGeJFDkAgcGUGS3jRiLuMn0KlUbYwvOof5Rh77Fi0PCvun4j2bkqQPFZHBVm6QpXtFuc6vTvqhvDw5wnj1c+raV8aWMPRrETHXCC+1fkzs6NzQSaMQZKSNYjGVA5drbVi0kV7Vdhj4btojN1QYLnDcFW43xjF+/VTEh+qo6q23PsfRUTqSv5gJFJL7VUhYvDDl7Cc39sjix2EMvebKUfWN5rzAhy+Y77X40nDqZ6WTQiTP4TJNrJrmfOKq6ZKIhKXFXEwVH6cSxnmGiM5V5hEg1tuBmW0g21gdUdc9oLdePpbo0D6ESbiNUn+LE6FT7p1y024+Uf6vYg81vvFufrVrnRtQoaS3lN0zIsUO6Sgkx04AdjggXCgL1Gtty5n8z2OHocGwvk74Lo85meqncaSFGolGFTvn6VAWo7lt/hYTvopSgAxn6VbUaf65K2GSDpY9f3pvzGSlY3+pc8tsjGL7b7YJvJuYaF9WrMAnIf0aiq0ocnPVzcVLaSAQ4QHPMOnbsJSUXj0t4U/C3aaLwrj0OAOPgJQ1vjykWD71SbOkn/7/80GSuthcUdQ/8e5OyjWcucHXdy8WVNAXSX0//JQWw88wYYz/Gk8EL6cMT1jwUlJH/nAm35uvm9JNVlEGFxPpACbJtB99OxN+babcGNDpAc8IRQTTaDNHaE8UYS/uTfLLxmjVLKCM3Tkyw3+5+7/pp7/djBQFBwUjHk9T1S6tGwMye/48MJy0NguZxLTsTw7SYedh3VRlbWrAV4JLRAIAS63XldMDxH+6Z6QLPzouuvOBvYKiPYK+mcGQ46bEs/u8euFrLH1se7VTXFhhjnIRMOAr+TCLJkMI2MSwqssKQqoPDObrentWuknc4C3mmHIB1bQ+CJ5DZxNilKZFMxy2RwYip+45eM9OpTrkTzNSBxMEzW+4XY8OF2kBm9awkzH9r5WPEG+PKyuLMsV30KIN/UEz2ckmLGiiWTW6MVyLTbSTnzdOsMQUa8X7yPaVpqfdGC+3hGvW8/eBchsdaN02blMPIPQxGBYR0CtY3sYhuBxuTeEnS8yki2IXVsMxnnyKImZPe9bPluDa/Et9VLOWFUMKiJNBucArrVMLLLpWGvH7EMXa/MiaXB+qPLvQhjs7+XdMePJYPuy4Kp70VMk5iBDLjQUOAAyqZxAsbgFCUivRwtB5MlTnGdNJDMppwqYgp3MIQNAd/GHDIqBVlL/4DXysyMg+/F7mZpR2zQ53lzmPlk7cEqcnqSZ2Qswm2cyQ2Fox/TSrZN6XY1D8sJ0jZBXQP8e9I/NmpVrAHiz2SBmVEAKZ6Kpjw3hqVj9OEPFp2DX1Exef4lGr0E0gE+QrHCWkiLCf8DM61n84MA+hndlVVU/YMm8stXpalTqkLYVv0eaLDLcYmNX4Mrp2WXPTX9Kh60IwdlarFsQGtv2D+Aefa1e3r3FVrS1esOwMsIc1ctGtWyKkC7MsunirRcfFYKK1hYMWJlKOfBnbBzmE56A5QVD9GuJHZN+GZbbFUbpmQSJvA3ckGgdQQtlvcx5LicrjAaM2q4vw7jF68t16UR6NiZCCnHfVMLHyMm8U4ykN1c/0SNHDq7ZkX0RtZTZo3rL2xceGbkd49MZVVcHnk8GdEVyorxtKZQRsgi4V1AZJqGBHJGXP2ql3P9tZ2gPTp3fIFGqhB7Z67zXR4pR1pSMzixEYvlMItg1MHWtatJveIZ1BwlAKMQJcr92LHaHiai692f3APbvXCx0pI/gkmFR5paMcP+ePDGuwKIn2BdGhY1G41upWHSHtAfmQx6RssWJbF1mVLLNrC8qhVerYt7CIQhBpisWflh5ZE7DDFTJsMxjnRCKx4RU3bvltkNII7SOT/qp0zGo082Gvze7dXul1R9onMXSlTluEXqvsMZsKsaJxQ7XU8k7V9Z86YQu11YVSjhdT+Dlxv9Pq44yxxw0QRUpofvdv3NNGN6k2wCOGgSPYre5+2iDS/1WF88gllw0wCQBcGC7CSBqN9mrpjGdZNlDDExWyRstZUGRdq/SVY2CyoKoCvmRo8C94j1NqwjR/hwIXRQQGSY4oCDF251QvED16yXPrOH5/RAmR5IKxfpCqjAq+DQc0EKj5R/hjdcGIgmB3J+7QLypPUNtlIwTb5ODrGXUQVjz7Ss/VP64khHSgRMKhhK11gVyeStPUwMatzTM6yiUPQmkmlbFrXMVqAGVqrhCf5gw5WagKFu7vwYeAmwOBIx2zoED0vwf+cgT06fqMemud1it5wx0ELi56m2t+tmjTPE7fEp7R8YqcEGWdMCtsVXsEbEmYvzNfimLAqbCfDZgM0NfBVjdOf4HWPNH4UrFO6QFeruBHT3zenXstHGvUA6gWM5Hb4rMlOSXLl9X8PLWQkOccFFTCprG6vCuktx4kc+myLsLtuzluiYzFYOMvD3g2nodbTvCjOnY8mszY3lZc+pluirZ972wZN/PBtwlQuLIMoL1mDTDqChmc4SZvc1xzm+yzelmIkuMoQF6Fd3OyZJc1i0IYz2ogrDIO/L6lbtLyq+awiajKJN+smV0ChMpAwFuUSjeInit58T8yZXJmwptdotKOiS9qjZVKJeHCPFTs8iHX4nbx8njktuS4rHKYfXjB8e5sgL0R4zPwWTG2HOdnVT2GNN7bhjoKp9tOcWDsm/T7aDiE5ML6DPVePgTmVrdR1Av6X7oymHod6aqduB/dNNYPY1Ax0vkfXsPcZVfHn8DqbX6U9wz+xrH+Wf++tRS9ZYdaoU1z0c9utp71yaUuGBj/RQ3E9aMNNFoM3CNS2PQ1BBI7fPin7pApVqosLzpwEuqz3KtXvoxx4JC9J6FK+bd7cbgmb589a0S1MZtU4OiaH5dMHWTvGeQ28ZoJoQ2X1fDQkXZmDOQR/os2NqZRa1NtxqIFyI4l0xp+E+WypPjOUqGfxVtB/LABdHifKtZeuatwTj+mc1u/mk8Cyj+Am/QMh6QZotRCTFBN660j6DWc0NuQMYSBpVodNl4gpnza9Y/U8gEE0B7UPYWWv3TildO4Xo0Mfi7M2sgtzXuWZ2MmUzCP8Pwu/nqupY7Gt49J5xGlFsHCYfxy+X+G1ZqYApp8kSXyu9rVwWuLH4gLM8wIFaO0+f1I9SueG4OYQ+pYmCpC3tic6F/FHPpPqv13GYYjHYXU43NKevU+mRJV24USzDROkpVKNfY+Foo35WAoMsJTsr7D8y7SFub0vKAZb9gmQOfLpg1Bm8yYhBZXu3aJBB3DUKjjLkl7YL4OLJ0ki0yY6hHh6ADzyUOa7dsSpJ/yYXxZIgs5aeYyXGz6e5gQOqBtFuqGOuyOcJBPiP7HqqZt0e2T1mlYVzcO9My7blHAtwsJoIhrDtrPikZYVw+Q0IEpZJwkJjRHCQ3jxyf6BZLFbe5O63nAqgrJftwnaqZOnU6mNY00464ZYRV60+EKLcTxSkWeWiK+UtH75cmIsmLB9T3mzcV3WzjPlA6Rx8Qmc4P2zEJdwl6xsytYC0U+X9Dn0x25998TXZUJhExoXbEMHGQn/e97V93fyhkY7PDr19mYOEiANw6/IQSIgF2kmZM0fMaKkcRdYV9GV2D6k+egk8DQ87WFQApffoHZgP96stzYt0HytBK1yeulY3QXWKYqGjv38NeIFjMcnTUhPdE97CcInQZ/s5o+2iUGpFpv8H4UpZiEkBtiRiKZZAVvfNmqoMqYMHxh0KdyOiqDpiOxHA/ys8VN4kEqeAJ5TPyF6ltLH/naNH2nEPHCuSb24nORmkKXhVEkqLuVVFb/vKHZdMdY5tYzUu8MEsQiF6sAAipXA/zjTrtVQvQaB7kRBuDCWrXG4HYz2RbLMIMIi3e2kx9tid0EAwm9uv4SXuWmbm24P+CCmMSIEiMgotjV2Lt/OPdYadJi7EU+zhtU9w69mSZRIpXbe3LXCQQONdX+GsmJdyYicbH1KLJi3KZD7ssbdeae16fcTob1efK7yMmPaSMsl6PGZUevDYhPAf926lb9db3vXRkxn7B1sJS8TUkK4sZlfS/2HgVpy5BVjgQkjQvDM9aFZIlpTWwNQBUXDxkxKCABzSHVMxvOJDLAEjvHGufQV0dLSoldYsGmRsozHHrh8kN7Z0Vj3tYwL/YWmA5hWX7UxlCE57pHHuINEkZPCkkTNxRZfKNu7BwF8W4carYkF1x0qm9icPzT7Fd7OKUT+VPESVmGTrRzwlHbLCgVC1HKZB+z68Vw5lwOzJ0tVecyqsudDHGtOwVzcjmjq1URhc4de61eoUXxBUloE9j/omrF3bvb7MEYM+n0FJUO4K3/c6ln7JVJs5xNMsDA2xvo/IjqVPHI92RzKaRehtCuvYZnIB1viiIfRzEsrg+p0BbN85uMik5rvF/LXcmccwoYAb+Uyp8vxgeiFoHO+H1I6WoH443hJ/Z1Re6tNoppI4oXtn6i5RoAlp7LT4a1Wzmz/zvyqMryUkwHQJy4yL7fTtako4DoWBVZlXWqhGiimnaO/rIhKflq8eu24ViK0SLbXX+M4guY0sJSQg2ACv66uV+vUkqCzm2O9qOEjkg9TzDtUIn+F8UMvXlAZAuQj4wkef3DciBArvg7A5X2bhHpU/hq4m0HQ/VxLRJUgSJ+QWofz+5oQ+0Nzepe4SH6abaDq7OPMBIGVbqgki7HIeBwEfVJUmDzAOSXzxohOadADai1lurf+i60s7+9mYeom+PqFg5ZKwsSCsZqw/NLBmDuA4gQiDG4yOLwFfhb6l3gEam3Boc1v9167FE674DX+hOReHf9bCMbZNUIgvc6RzOapc4iiAABcENzjEPj7PUfodEF1KXb+Mazuwi3XmcksVvUFzS3x0z8PexEZkzKtUgiwRmB/Os43IbrzlOJ1clIyA7yFGo8VXSKFwRRpWx8xte5VTBYVGPu/Hcge2lzKjBCd3hUgDN9LCPkLCZ6ss7Yv/XXciOwa+MvvXRGYp9OWCu/Y5dUOdm8xb+aZ+vqAHPQoJWzxORqQnXqyx4DfSH2+sfuMir4NZHCSvBoK9wWub1eFU2n2BXuS5sFeQ3y5UKxa4jPLaXVEOO04zB3no8kB8fcAMfNwSiJXbujGtpk9BiCPZZj3y86etIlAXNSbTGMKggbR9PKbL51uCRsESv2cdaAIAFECOJplhLrT16l9aAopLK6Rlg1NfQBzHHe+RRGQUE6QKIflTqGt7GEkGhVOd45ImhrN7JxKtYSgaB+uqSy6yPaXrVMnnyO9m9cL/z8Vh6XCvcgobaCNZjmqSHethe2t2n4l1AQ+5lv8JQefPlNKMOaAlC0IHCD+lxvpYaSoD+Y6qSMcTNhRs0IjcUahHJOSK6OZMrHdUImsqCFMokTh5TPO/6QwbMiak2aNkGM//raIfGJs34ziSHxAQv31pGScQeT4IFoYZpYpUyx9ssz/7AnZ9D2NP09kq9e9UUr4Mv0y1PBvOwiYr65WQYqFAzT5wWNUjL0WZY5wmGQbno9DXxHvTg7tmjl7MV706+3k+5xMz6XHlZn+vcrpR3Eo6JSxYsPX5e+upJQRACW6pAB7ElV+OpnaS3zd2UpIJ2ZRdcvFhpzsyYEiPgCGk/suuW8MvfEYnp7pPblKmfo++ZQ0SbND94VbsNtHOvwC1vaUTAoAzE0URf/5fJra5edfzOHJz0khvV/VNwdkTUF7yDF3bThjLRdW6lyVykGpUOtT/IEhYVVviGDfRdxsLRqNWK8X6J4FCNcGMckbtOK3MbgK7xGrMA5yvigqbdH39nrsDE1Qf1tGofdy1fPCHjq72jhXSEn34k1yAW4mi86Edj6vRTbkB1pF4bZTxlFjjEtKevhPX52JkzroWPqMqWAw2trXEE6lmxSzHnynuU3/bVgCWJCqB/Ie/+T9SEL9fw5ATfjoArlDfmPNlWPFpsDCHdfOLqHh+d+FfbLmb/CcWTVH0QkYKktJTJehS83yzB3zguKAmpLCmFfkECI7usyk/MyaRBET20a+2x195EGXmczesTSsDSATSxJnj0lBFnfeqCFyZaLAJoHATN2Vo4b4gf4pwk8CQFjs8GavTLmOijFdM7xVFFCpUTsBujn7xXsKTfDm+wW0eFTXSTp8eYDEogRbV1iq8bSIgToI0KwdhfvkhDkHuUUiauXPO6ISRfWhA2MUfDslpbnQDuas9G8O77fzg75QaKM8JDdLc+PeLrbsAW5nyAB5eFfcKkIecEQGkuRL0yUj1yJJk/FYa7wcnGtDRaVqEbEyOumAc0VExwspWDNEBIBslfxFoLbNJU7y19CBQmm/Qmx3oFAgkUetL5aWIjxixTeyJ1EYmFWGZ2IPbgVPTsf7bZDISaMuTk5CZC4YkEYYYJ/3OkgKtPdd3yYkGnvR5ek8Mx1SDvFM9zWBKFRGfdufLvuE9DYAeYQqSPEjt4vJqg+X7AqFpolY8UpHh3xVvM2V122hfpapGcUUrbxDqizfQPz/5gqv+WnPNrUmofz+Q3eJPUJBQ8R08u3sBPue6I2ucqdLAQbMcctcBzocqesY8GQbgtrCq6UoHpW8FY4PDzet1fuZxy0AUsycu50otxoh9hhS66wAWeWz98AfEeU/VF6TF/M3nl21aE4wGDcCjykbl0l0F2xZUVxzOzsgBNvz1Srn1oW6HO3c4bJXNJHW5NdzW6VFBDDcbiHsFyRL2Z5lDUd7VhJ2HtKuocN9zqF1sv2Bu7sMwDnUw6ukkH4CKKUKNbG4hVc0iBV5ehEnPsDoDeJsdxaY2GLFeB70wp4iKAhwGvGOgXb/LFVvOikf8Ki6DsTShYdvNYua95cRQ8RLWe3O9vZAkmeJHGSaJynHi3zs64n/vi1sSpM+mepVV+9emxBa3HQvCCy+DpY+Zbto8ALKJ3HmWqxIwHBy/vtqFMl0qV6QA0hqZDoVfD+NExuICyuz97aEKznRQpgLIs5WyNNdXY4I3IfWcUtsow0AieBD7MFnWa2gLR55tKs+zHBzDeKKdoRR1skT7bTj/lpV0aYsWrADuC3186lmjIYl8J/qi9wrQQNenIzK0sZ+Vz+QWrAAmYRIeln+QvciqVu0C2jdw25sOJT5Ht4e/JLgW7erHpr8O9eB7xuZmM3iqb/zBRuXPoJ2hs6IBY9pJLU6TkKVaruOtm11wW/NzDebN431ra4sH/7HZ5x3l0l/KLF2zc58foXaaXuGfIwHHjaofEyfTiVi0lRvAkrftxIyVa622rKgTYYx7iCQfsLJMPZetfvwXqhzuxFt5oE9fcylC1MjNsLPbhYfNp+soroUW3hCLqP97yEtK0FM+NKC1W/QFw5sNpbx4FNmifvn3jlPiqA4OH7dAZtmoBL1CEViwl7kYI6E72Ke4dFhWDY36wnL2tSr95NSanymO7b7puf0EIn8bXDRloKDY+uXEMYeudLyqEtLJHQqNmxkmWlxZnuIn5zKmIUKJThlK/Wxq9Iy0bhjaqMJSsn9NZolBdCGGIhUTNoC7AmJJJm7BO6K2h3S4SXapQogjdlJ/9gCcZYM/B4piVvWNGPnKiHJX6MoqkGyxLmWeff+urSW2VnsTGQ8igObiBAoVLSZNNXkruf6zGuQ2v2rAwVNH3MXD4Quxyt+T229ASxSsfR6l0ZspzfBt6SL3ZOuZ7xg/kqd4ZKX8lCGj4qj6/OQwKPwKZJgd2GFLnLOsOcIO2DzMESAb6z0kqrMD2hnOKqAXP/Fn9Th+L/dOfj1KOcCcpGVZTb4hqhysR5FtbTDvRqN/S5ren2EiN/JGrgXv2xHOcWJimTYtyHfLzHfdhLAt1O6U+8GINy1VkLp8bPPCiElEXjCFqkBIQMqQlZoZx0vgbKc2JhoH5daZfWgoL9uwnx6F0a//UdBlGJrOH1iS/eziQ/xGpNjJShkSKWdidv4leKSObfxB9CC/4zySWT/F/9uwvEpEJOKPzWzCsdhWd4ja06jHiyi1imh0VC8AGlMW2SemPQb5r51HYJnHn4zXdMTXfz+2MG2LaTB2YhGTx6lyIQlgjxxDfimdOqfBSaNHo1dhbmZy+GKPbxiPxIhdzXfNcXht6+YmgKVOXaD2cv1tXh6YX2xaqR5xEHKxVugHX84/nIdN+xqqxKmg/KstGkTiB2HH7JlAyAUGV5sT43ifKvRr2iJN/N5vO+iFb7t3YETWP2R7nSQOGIyAhILUZOgRZ+zSZfCHlMWtsuPO8xuS/haISUR3otZdr98ISY4d1Ja82hlkFbmCcES3XxUoyTdwPdayiM9vrhGMKqoooBviuD5tSzi/Y/dYbeZ+cA1f7ib0XFBLSgNVnLA8RkTuRx3w96NzWzBSE3yDgUNhQHwLCh1z9ihJ1iOiM/+OYlUHXZU2zfVFie+JGs1uIgxwrDmv91N4mGt3/7Oyi/k6drXhfQLO1s2d3Ftbe87FPIgFKtoPaWuGvZ5mC4xu63M+y/VEweIJP90FDOLrqEfatOSUg8XTymUyvbaYSd20TJko9K1aAARk/xKdw+EToOgrSnsp7RmoWkWmN1OaGaJYsPdc7so5JzkTl1ozxQqKdQ/s54UaGDhzSJUt+z/yCFu6/zpTwbvKEVo9tPzfHJTPz8HXggYCURCfU5mIdrLrfmfaXfymWCnuvtJAsFQaJg8TvQYZPvDPZtMqI3qm7KlonFhb//rWXBAC+TAqCKq/G4lRmfxPx4x3Hh4//FO69fxsUOxexguV2xIcou9VeaQJDSdRMZy72P9Wi8rPk60uefSdwFfC4lIo97/fvKSf+vgmVj1Xp+5tEteCWFktb1FyRpRlaQQpvv/9ZU3yWpWO7lr5V07Ndb3SvXH4TvfKopEEToaxmEptTxGf4pH0f7wIKLEW0brMudWhd1Ey/egaEkIFEHYavIWMQdzCXScZwPRFqwWJAOGHI59LdzSCL5GtddlMNeo0dTHARpZetkCyHwmnwFoUg9xyz73nRt4TzISx+DGhb3PjmJ06ZKk+yAI2Dc+1hB5blJbZPZGKkvkGzR8wvOIdCrInq9LNSEVX5quizTjW0Wx5a8cAnV/bJDSu5vufSkIJaaTBSS3zkUpCHqlMXbQGpnWOoM1DOmKCtFn3z2Au7aoLVtLLotjygj6vF01VLt0Am9H6ApnwH/b4V5HsxckQtCrX5ZLuikst0MVOBNJmzFjj29oCYERDNJHE5escCLxq/98zeXDGbVixiXeEceZyZaBsXNpHaPgJxEep0DMYUngcdjE2+kHcQ44aw53dtYBbhCahgYjGcu0xegEt/hrsmFEGTxzMMbG7zxCg/3bSxu5JiUQRnhIZ6vavJoq26rBeXRTXZJ+/ay7AuKbUzbg/VmrOM/2iEdoSCUWCT63SlE4vsRFRAvQEWgSNCy4SimHQNiCPEVNzur4StLFQApt+HB3ABhBBYJQrrT8pdXtZVv77e/lBqX0WzckRNGcWyaQ20OP5xhd9nvYAhEjHU46KJDcZEwTsx0CONe+pj8n1YM9jVxnqvDQQQLU40ANdovmlLTZtq9FWu6Pc3GaChjO5blJ8ta0WJkJ3NgGDHRxHSa/Mwl96AmW0WGBNHsJOmQZYyCmK4rf1vBF6f8qjwMsNaWELWN06nFTLVB7slUxwDbcibxuG+xLYAhpUmFdjuBIZ1TozkuMLx4MBQNVdlhLDBbwJqZvFbTimkH6LbuXwdFNItHWAyFFYQ7Kiyb7T4ec3RkzkRvGHvdtIFfCz/zr6mam7/XfZA6Ij4C4jjyhGbuGHXxm6KhA/Tcd9yFTmwCfXQs1rG3exMW3gstCT+kqih8n29fN2XdB9fffNohM68hKEUbZwNnpae7dAs4Efj6kbaAyx5vkj0qRBovSPNwZAteMMm1WLp6agwa+OIaejhe0zWdd7/5T3tBvtSvQ+RVVafhsSUoTD5BLWKE9DzoQ3Oej4zSKlbR/cWaPfFCFd+evCzwxBP0MF0lA2kPdr+28yDZJoBzlwFtan3lP+9uZG68u7T2ikDeEBoXhzkS8toYXAW9cDA+V/RW3chqAPVcxkDq2x+JIeTt6p7Sfn4f73BIMAXQ46GvoWUUjbA/byJfSRlIALP6u+VGn0y3quLZ4FA59Rj7qO1GAU88Ub8nAj0Q1Ii7cxWozsj+uvArtjAFK6Z7TvZa104r+DJjzs5DVKeaInwBStZHtDMH0IQxEtToe8btnOoVvdOxOS3OrREilFwieUt0+bspu466WlqIDdt3T7/Uv0vRymEmuu1ucZtU1RXRCbUPF9xqfKcbXrs6/O1t+qSBEKopWjOUwkR5h3PP7M0FlmDeTK80a52H5YRAkkfR/1GaXdVw96CwpYJkB4n5SHLQ/kfzmaSnNwP+O/rhAxiac1UydYPS+A2Vvcp3rGoFO8efBnLAUafXy4t1h7J6iZ/CkRnbLEZVu6h9F9raLNvlrM6M9Fo6+ope4GOXtZyGrwS/DTReimbEcjiRscSGPEeHXj/IRADuwCSZ8pq66OWJkEwJaH8uf2wzIo2bBspT2PfxBFVFfka6VuavSiFHk4eR/3k1TBugEADYxjXiPIJqwqW6wmnT5SlgRlOwuvg7sYoPbym0LPwGkpzUyrxMhAL5lvmtHlMLpEdpfvUpfoo50bk/Tlwp4wUuruyBfXGbJmEpNVXcVNa2+mQaBdoupAdsiFj7EAK7KhlaB+3sJJls0/vjGt1XVD3JSUpWtbsAOYiqp8D/b/I5I6kgXLH+hTk/SFCMNKWRat0Pz8pi9LMac0cCaizDeyZzqYMp9u0TPmUDPaEF5L0jfNhf2bo6Tc0UrAi3zOMRzuvM1/gSwKPVoObjIQDzWRALd7D9NzW238JoUmV/n17MhD5QYJ7YanonlNvS8waz67oh2m9eNzItPr2C89NF8NCh+egXtSEMME9F5KkyZNONve5YtdM45Q/J2gYlrPFkP6HglCFj5KCPdbN5t8zhyHPP4V4kd7nj0FEpI9Nxg+f4/BdMHzC2NJWmdrkcmarG9qir8kyNXFxaD1eIvNPEoJVr1p69pN0Xh0RnWNzP7PQ4K/8U4hltWmwH5xF8MJinzTvnQwqTNYPuE+RHNdVwlcqmZG2jJG6F8+ExaffNj55T/DyZuYqUr+dQbuV5fEy/viy1an5vArY6kVjVZgCDLlGE8gwTcPdKvsygKivV7uaTDu3UigEA1jYWDkBOH+bC/ht5NpOr2I8FP4ABu00DhdkVO0z3xXu+EQEhgCuN4qR3gZIKRwqEmVemRYVu21R4S4LzTXSAGwI3lmcd1YzVALLKEjFcvM0YhAQWJWIL+U6T+ibkk80/mPraPjlkOMQJpxFvxI+otdcRvbJh6ieDDMYWeAHvQkqoqTwSOzjA3sdIOGC/Etu1CbiqSAlNOkycVvph8s6eq8NjQqnVnFEdgkzc244iwmI/A6Y5rsGowVFM89hx0ugTGBQgAnlNOzhfg0jmep/irn0OFdrvjttzchhT1RhG+xDnAoZS63CuzDXNXFSuGg0OyRNA2K2aRKiV9Xy46HPaCAcCvMzOqfhVLwad6OcYaXonR95R8DmDL/8ZxFQmJvgWnQxUIpaBTrCQtNzPDa3bPmZryyr7tlU2gpbHh6l2c6SkEKxjSmev9S9NFDotFb5Ui3M9c0DmAy/9s+YkfpWbQ/wXJPHm//I5EGNIiXuXJXC1LkUEAg6j3aOYPpqdlh5wwmAbBVBycO+3taPA4ScW6DnSHBFbIjLCkBRZjbT01NyrMWxVRgohBIlwk0UOmNH0QNKXOwTLvKD2YRqEWD638YldeWKP/jrt4NrHP9EUQRioVCRwDhrymOSs1Cv2QjRYg6jjns3kQoigFwHWNMwR2QQdF1C3GHQ2Q7YV21/ImgujUSaifOx1cRlrDuHUoZfSYQIga+/Et1CxZdzdE96TmYP5DFnpRQEiHjqOHPqCWaOqTpKkQXqBlr+yiP32gnDkNUXHNfdzOUxAm5kp2faTujM3hn45MNlDjP52MCkwxRVTLQdzuGSPoQK2Lbgy1b4VPyctM0kNmUZASuT1cQvqeFcOp6VEHth0LBKGs8NUI1chF63dXXlNiY+Mr9Ib0xZu9AybFlCEbBxmFEDAUA7LmbW4YUL/eF0uH33pxGhXjL+fRkcEzgw2HlgXHjeTGQWCGgjIljWcPfTJT2rn3uT/GL9ozqf1OskRXlNrllKk+vGEznULhQG1r0OmR9EZyOvyjNsXIrnscyMbLHaaowiPOhJhr7FtBEDGV4wGVUQjcQnXgyO3KFQMMvKlifbm0GOJFRJNBavQ5QLPDZwgY+QlG1/z6qLV9oYJ+7xzzRSkq0WEBKa10thBPp4xrSGmNLZxoO2Lb3c5TYNXhky82/pywGokpEsuxWkClS0aznmUxVCH8JvcEINes4crA6bDX/EJVaurn3rAnbFVPaSle0iEf/1Z0oTqiOHlTdI+vMM2nshHy+mzGFKe2fwq3Iuamj4Z3htW5W+F83MGsdVCD3IA74wLGFaARcU6XterchNug/zmR25U3bKEfrXHXnYz+rIOva7HA+HEu79utMGTxl1RFr3ogTPq5awom2wfP3Yp4AmJCdxT29+mmjUVxP9bkE30XYNoOzdOZWeeQRKP928LBJiG3K+rgk2cmReV+mb8L2w3MvY2YGCseSp5S47FIbyL9V4V30o4JHuXs6nClvDPR5VlsHzrNjAX8DqcWx7DV3AZUE/B7WhXgCU4oyDvxr80y6jF0e1YMF43sc6YxrBe2yIJAO/p/660nGK6NhAGZ422qRyn1+V+C+zQ3azWVcNgzYELMexPiQrgk8bGVXctSUYPfEfUZpz2o4dCQucnhaoYXYSiQvVAw/Wu0bqbpatlBbqEB6kazEqU0K0W+w23fzbQVEk1BWbh0gDnEsoP5HKVPOU80y2oFcPfftPkOMo45P3fC44NkjoE65R9uHwzFCECgI98gXyfwMOszoCV2ka/07cD8ClkSBOn/oGfGRGAMPScHk4xR1iHHx4jHVMNvtfoSa+iL1oNj4KZsTVPzzxD1omc2FCiZd0DHDqs93/oAlRaUMrr6YVvGxBB61Hr8wRVIWesGkzNKfWCBIZl4Y/GGLrd3NHbQ9m7xmCx/0C8HqygnCuL0jsl1O/5Qj+JsV7ae5tg3L6HtnCtQ8R47Gnf+fyPKXPuOgXnFElP9gJkqh0yxrLLFBQJgYaleB4W1ESBPXXyQZIdxsxXMuZpAvW2fdbeK8ctIoLmkqAel2sNgt0zTNg8v6kHS/DgZfvQVDEsSzbAEgTpY/72pr+axYodn/qbH4KK2jr51guv89NKB8Isc2m10DJCDBVrTNIy2wtq0kdhNmt/lkhFJT3fnzB9V4RsKqEAUB4tirHtJXSU6LJMVG/eFD9XZ9Bsu/AriIEE5y3TEkux9v5l2RsRcjCQMC/N5VUHp5KjrW2unu1jjRlwXkoxqvYAJrDGPGag5ClyFp4ESbp8WzkApZpPcyFjhEebyRsv6Pq+V2L6C9pjLBNO7j6PGx4Xpp0lbzP/i0JhR7N1yomWYFX3p2DFAwsDmc3kG75ULYP/9GcuZdqhrrQ6AWIuM16B5+xNgjE12a9P/oCiqG0dniViruA8dgXHiQBEyN/IqqfPSJFNYAOq5a4xEcKmh255YpO7DTsCbIrPx5rlF7F1BRcsKaSC+24NTCmwrGY1RiEcT2OUA5vQTDV2afYGEjikDMpHvxDYSkdahDUuiilUSzLPUtIf/uv6o94t7bgO47A3JG+Ij5MSHRDnY+nnfHHJm7IxT2euq8wwF7KUtkefLD4EqccZ01QqTIEo4r65cIVGqltf6XctzJyp1Jl0TSYsnJaZxR4CYlh4MXam6ALsMODnr4hTOkXkackX7IYwZVZXZYdFMaV7yy9s1Q7iIAtpx6o/6Dw3w8TbzQrFS5mLGOghmgVeRndFUXHI=
`pragma protect end_data_block
`pragma protect digest_block
dd879eab8d654ee212596ba46d9a7caeab09571a432dcdae12c3d13f7b258f5e
`pragma protect end_digest_block
`pragma protect end_protected
