`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 9629)
`pragma protect data_block
kqP2rZ11n4/mAFL8j2IDlMec3bCqaw8+8jPaIvl/LrxrQsJg2hbsjva3xmSMfBhf7X4XriHbz+ldGnuMfcQXwR+nnoifNICl4cR4zoE2pK+XUPATGjPvAtEmFmzgFikZ98M37umZr0upbTFbgeJ12BOWzF6glGiPk03wIP6qFTsXwBoKuXhqlsFRbYV8O1+RuS9de2hZdf0KlpnajjU5VRFkdBout0QjkZ0306/mq/8sQ6NhW7P46eXTyip7P2ip7QsL9uGQ1uMKMS+0TUbosPh3R84BjuzI4X6sEODzLY/VyFECPYeRFTFB9qYwrMKpQYhgiIQrwZAI7+10T0jS3p/G3slUfkJMvBWy9pSKmjQqQGKMEnUWr3XHpZazjeV0MvZKyScu4wXoWUaAODUs/zHLqsJh5DXtz0ikc0HoCpygKamWAesaljm+fnd35qPJUPAXosove/S6GyVQS4VATSOQEiR9qwDwORrNqjQ+S3R7eHfd0G2UEv9t5yMqqIgjcAvECj/hhin8FY0HF8nL+miCswIEZPOcSrcJPaGiNXALHj5BT3cE3QMoz+4Czz1YSZjz1Haq+AjT7XiwVJeYeTDg3gUMqmJGylVX/R4rGqEm5N2Q1kYdLDUUhnV2mWZX3wr7kDow2JyQ+Ha+Z1JGdgVRJxPrnHJmzAug7SnU1IvG8sF8kR9m72PhkuNhc34b6Elk9u16B3+3ZA+6Eh5obUY0paFocD7CjwANne3NSgdsRCs1NEh/JfhM0nmpQnmMU0wp1kNjWcD7OgujZJ97r5aprFvCveThE/oOVyNHrUpz6OkNGBUdC5P4/sc1X2HVBZD1gt3YIrQXCRWSMrmwnEn7OCZMyIO2btYrIa8wpNQKG7uwchd39irdftOAeR8ucnjKqXFL3h7M1NyYpTN7Ck299zViRlcjZANGutsPyWg/AdmmCBLZQv5Ux/TLTyWbljD+aJsHypcRq9mvNQlCHj7LNr/vPsLBgN5OH8h8qBiE5hqBH+sL+jajmuu+ht58y+UOQb2k/bN7Cg8DzEY7Ck5rmF4Ih8MehwlQwBP+Xki5X1JfdhTiK45IYYwwf2C6TcBgRBQ2/8048erohrnYlmxOFPhcOIr0h1mypAsK6ZLBpSm2DfHHczlwRrmfpWBYhBK4btEyR8agcWmVCqI9en9TyWKAC6NoyKYxyzrt0YJ6QRgjklr6J5nDVVkIMQ0/orbENATp/mNvvX/p/ykTkCTktMQ+/Mm2wrBoXXRFzqPY8oCgH/eTLJMTh4lPFTzVIFFoZTTO3qYpbVyW+WawaCFfRQQa0SfGjPmKeYK9sIh029rF2nWKgzXG+TN5Oj/q4uFMgYNP4txnQEF6YLD7PZs1KuOwCoIzbpXXIsjc5fGnpbFDNKn9BI0ZiMg8RAv45ySdVCikbAkp8Od2bOCqBBetaGBygPjWYwQyFSLPjn3Zea6dmkHj8GmMmIbODAxiI+SG9Cz3IDS/bZ6NizUnwMc2pN5l9jxRj8BQZ5LkvARufy/NiKZCsWHjeI3KyEwt0GkREWkUZ4G67wM2iY+6XSymJuOJDdLH/hsdwgQ4PCtzO1i0897a9Yx1UH2gzKPLvVAfSG2Nsx3AnfU1VGfhC5yjAO+VnUqqLOGwSXx+eS9RcPx4553T/4S/qbIn1ZpePWpLPXAwoN5rwMNG5u3OEH5oOfgT99WkVY+RmLgMEzEYPx0ZBvGWRtGJRWPmUWsIXb+ZnkLbEEGF3DVS2VzLFCyRcn96vHEbJvubKSTVkdmic49zUqIFp6uGCx8uA3yWBoRq8umrKN4ViU66SBLGhOjCEIBGmwgxilrup3z+LeCyg2TFZyVYMh4o2pBXpwWFrit4gOQ4KEFVc1mHOSymIi0fE25PKdZin3yawdO7d+tAt4KeLmuKDZBD6hdiSlH0XXPSch5r/2w8mfiAeBQoWRO5m7BuR6A618N/zbMSy5vzP7zHsmRAibCXQ2F2GLqZLaEkNUyePpxgF29QFF58OWNa/LqXvNMpWwLzMK1+AQwQixc2TJFKnzzrYi1+SRVqj6EX5hEAsT7wV9UsY+19sYnTHmNk19iPecZHd2qrTaAC/iBC/xTSLwggGaDhHSip1ZAdPvYUmLrDc6qKjFJQmSwPc45pCDI9INn7mpFqGRfJvhCRnyhzzokFKIi710+YJny3WfhhhkIeD+m8WYalLn0Y/ijVzFTmqxey0o0Z8SnJl2td3gdnd+gicnwar7wYHl+so/CmowPpMbvsjMJ95Ax5EQRDxjgVqVknvKNErW1YEAzq96aO54/PxNLTmju1ghMI1GX8Jd9GIqgUrGTAWVqQwwELn/GXcSvCHjjeqVQrvS+njmD8caFgt62rCZG5vcTi+qFKF2+4fBJZvuxxnkjfm9wlana9czadMLW1hsjmPrbLcucQEantQm+MuQ5oz6QdlJg8GvEr0xawRHnbi/DoFwmYPMnjTG2LeQSs+aanx+0b1gulZz6RGpG2X1nynlZA0PB5P2mIBWUuREtoLCy5LZKMdm8vGs4xY5DvmwD3ZTpIkaycAjg7yWH73aKFy3EIHkcqilUM4ArxkxMEAn2sZTLEcvi+oeCloXrV35gjqNLbByCFpi32Pgwcfo1ksuG838a5dMd6q6eIqEZVO6sR/0LvG/fQ8KW0vWG/4Pl83hMeUaRR226kbuSQhesc7GX+KCgQ1DfDfWbNBqCrDNKK8Za0jpqdzyX4lKqF58s7891xWXTmbsKlRt3BxewS8Z4Z/f2jviPD3jCYJk46wwNy2nxdQTAb1Tz5SmghWlCrvrQQfbnB5rBhAYontGnB/586q2CbIgRMX6KInLiW1bOu6FmXi8DoovNww+x1JPQ5lJsX9VJ0/GnVHXl6UH6dLXWeMTdGMVmTLwVDjKyIiGfRZbP2eC63ACvHnG8VPsuH1plO3fKdQ1cdFnoF8/vt2+9EDx9fDAkanyxPdHvwF7s1LRy6HnYP9RO0mPkxT+7k8VqpimpIfXMc/UMkAA95x+NCYs+MV0F/0fvFPms8HXnPXrbeiTTB8fvgvRhr00tAITIQ42yArFXpy23Ctz/1Rl/RieDo+Q0AOpF6h8iNeQmkVDH95Sbr03PWyT8OxpxYnu2kbUuqBLPg/REE3iHqyjHJ4IUrytZodKcqhEAh64Cgo5Mv7sj6XNCelmnNyydj1gq2TqhzDeU+UlBkuzfSLDeWEy2eMQvK1I5Su4cFZ+rcsQnoOvWc5Ne3mF7WrIG7gWR2kltcoamMPBi8+QTGNVpyxALN6sh1fwXwtQ3Y23JJcOw7YD/duCG3ic4FeJP06wLn+dyPV0a+QWE17tSTNaUUSrZ4ZUNNNJainexX7ZNxSJbC66+3Gm1jNmgTWEQU7CamqbRjyy7pLrPQFWKUD75Jlxsiv+HtH7WH8k5hVPZBTj57/BB3MYTPiyP6EcRgLsLeIIfg7XF1hk2CCsAeLWjgfdtwOF3ddR2F56btbNIpKaUfrxUOAcsB5vZMafxog8Nm91/kAvwndxLzFxhFfxLpCRpUOMAeK4FVzjpjUP7xNjPPHRfmylcsTAWyJ8ZzKKB81W1IY+D7+9nSOCn6cSrCxIVb9/5Ft9BzCgKDrqhEXiHUzqpHRUKv5qxq1fNlusUG32jtb899iOppltDPC35F58fvPtyo3+D9JVjC4RrEZh2EfWN3oNv6rkD9L8nZp2hD9yIFt508NVF4WWflYnamyjsK3Ad31PosGEij0nhkA/XZTh4eNJkgyAd9KUvCh417QovGaOA4CggbhbKmasu6kP6mH328Ye/vfxDYfciPN4oJa9TtH074u44c2Cb37EPrWM1Wv9rx2cwaboZsgCihnrq9jz7y18kSH25V/kjaLSLX//l/777BreNKlrVmo82RYmVgPrlke86Bu0L92KW+3bndrKQqJQt82mJJs9ZkaHPZAt5Tph7Ewsy7DQNTsLUpDOFr6TBWG5JKl1zbqMIzhdIU40wsXEiuqnaINBYuAYLeOfFrzqJzwaUzIrmeKcEUfk9+dpjl05z6KUCaj96JAWo6KTuprF0ZZk0268zAF3Ds9CZtUe7DY61jVeq3HSAd52Q/uwgKbGCrT81jnqyMF93ROEvVLxW4a5OCzwXibWtV5TJBGJGg7/Yycbf7ghSXsyON+PUHwbX/kI3IjQKPBKOx3wbODqnrUWrzHbja9pYSXKhlC3gWdalUH+uaMQDd+BEuMWt+DODK5xdZDDdDnwdy/1Icpl+DNHApUVquZlFlAHnYSMNfae4XzduxHKs501+a+NQb2Ai4U/n7PdmmzoYvd1cq5l/6An0z+GUvc/ByxFG54OwS6Ptai/RyEKuqFHLjvLxld6tVpJIuDn7krTvMQk3bYr0WEgLrvzDb6ieJxi8cUz22+WDPeiTQ2Db1B6z84LsjEiCocEnBeAJmuU5fCxEixEvFNQyacbZGhv+aVHlHHhBo6k7V97qY7zY9DkaFnnAVnxj744qUZxK4eKp6C6Zcr41nfSOuBm8VpJUtw7ZsDXh+htbqgb8Vlol/AVuDhveMvx0HmZhpkj03yShiPp2J9x0g3iwatY0+97zD6zkRn2TvTfgVYgNI0TpaoiFtZg9vAMCBLj/jhq49LeV3p05GtE/Ou5hETzMeBrQc4dNe4eUYhZnwSJVd8aW3/8DJl2TR8Aw4IYlBvQfoTESNfJFudXnFbbLhQgPTslIte8NGEvciRfIHjWlRYB42ZWbYHEpdiKW+j5bYFTdX3Lqgz9qAFfATV6DTpuPLLFcAT8d+nC+0QmLuhOGD5BMuqFPVim7hcVBRuD/OyUspIQjT+T8lrFxa+tSMzFZWxY8FeF/H4bl4y4xoRL0UUmLU5sfrf9ScLLYBqlIQ+fCx76W5yhJOP5S1NO+l/2Pt8Lv8BQjEgnsuK5Wq5z6t4e2y/T8KkO95SNrh5dAVeUmpAwq/mjVv8g3hVsYq8mbaqK2JGWdA86QwzVpvW33lCpBU2/zHjkob38zpqGJNwH+L6kjCKDaH7O1854X6cTrdV6q7Axn+m/aX+L+pKlJamSv4txYvLXMIYYiwt1Y1xweX4kfuijS3rFaGvz5Dc4p3G1vpc1ZcoG9B5xikvzNVw3Vr5G4uCTN/NwCUIAsC8Df6MLM/K5MrH9vvdhhO0RX7MlmBu1Umo+5jNtcijwSEh1I/cI3PUYK/cwvjpbi4zzz1yxJzzwNF0VHVFt/DIiJC9PplSYnzoVY9EpIYeRTdnezIl5nlxiwZLZjmbzk8j38oimARmJYRhDvC/2n9zAn1LDgTp0v0aQABIY/c7GhmxqSjM4cMLtqmnUofp+6yN16HtIWnbIbzaLiuC4qBZ1YCj16FVFA/OOYtOo1hM2IhSAb/zdyM+fRdidiEVhLxi5QtwthPfjSdPO8Vtt+FiVdn78V+ird4VVps8VUM0augVcLMTzlXg/T0G9alOIvn7Gk4rauJhSEBI9sEZC0JXCTm2ZCNCnBRmXbwteF3D7117IE6HrP7JeB8y/Oiksjh+OJ15sgRFjLRuPl2AxUI2yCWrEE5eFkMcrPlM1DdweZO0At/SdpqK64gDciSpgERg471qJDTw4YRAgrhSabBVrurAjBUDpv2+5sB2+VkpDwIBlbUnLe4rB3y7406iXzdudxlOEybHRTWLXnnGME/zq9f7bgNk/LbaIwI/90D9StA3tlp2bCzEhOrQPaqynuqOk1ku7Dhev//5Uerxyzt7+uSUOXeETh3eZq+LbObrlJgog4pPAfp+utvLFm5HbaO6GR1gSMAL08kkOG9m1ceGz/c4O/5rAWTwtQ9dyhWkdLztv+fR3LO8TAZ+KRYkBKT93cvlGK7BHalCzIvZ4FHm9GzMm3yjaP9SBUNr3TaU7RB6gIOBJwX/yErFzRny2g/GOQkIVpTSPyoWFAGa5u2z7MhRVi4trx0soVBwW6qWRvLIC7K7Aks1h7XYeJ37uRHpQ3zVJpbQBLaktFuM9GudGYGbpscEYNH6VSuWNes2Exi0wci9dSbYAHPmjixoynEUSDJGWcoBydEmoQHxVjEqSesmmh4xlwb2sPmK34/1lrYnNhP5FUx8T8KrCz3MSSeCaHXjQ2Cj4gDbEpmvZp9+uqDQSwOwseQjci/5hGKbNAexqq4N0SG9NP1kOPPsC1qr27rT53kankIY7RfognHZEcft5JAffIdG0gFb/Vl63xGaKpGjx/1TBVZ6Pd6e+COg8vMeQUyv0iSjfgpJ0e8BDQbVUZOH506ipZzsGs7K/Vaffi5LTTPIg49MdhQgdLFkYLM+Tg0BgpyORhN/Y8pyfzJyRmxGUIKLy/JgfLanY3UpK1zSRKNPlYBtdirU/2pjxuXwX37qST2pVo41TT/Ft2dR0dvVLW8k4alf1GsOb5dpRWr4hNeV1ynVuud8et7y7DCYPqhW35uMOWrfIA69H7bGoGsA3SBk7r8i68QcNCKDGuuM5eD6KsciEOAYfqe8EAbwVXoZdSspc6PHb6HFwKc3NTBIcy/YTOswX0bXhjZrRL6Be5rDoKpXXKoJwkkeImdGUHgkTyeIxYsts004ksHejRP2iC/it8f75nml/liLMQuh3w5XFcrJYdLZ6o7OeAKgwiiEYi+JZYANUg5DOcwRH6VPVAs/SkawDdjnnl7eCHy3vhiuM6MxYQDFt63dBZAEXE1QJQGwptG3WPBc0IPFhoaWXtCFnX3iF9nekGfj2iKaHgnHEyapLylc0xpGp6S56HOZB6htuBgYpJFo0tvWoYe/upVaXw6d64zNXvWNQtkSjIZVhQKJCBEQRBqGMEUowKcZTf6jXno7D4O6hAJ+ue2UwCnaHhtBv61KWiNjbSKc+MCyQ3UIUxnZjYkQF/IQSeT/Cl3PczOpl8Dhlvv6DFhwZDfPIOvsUOIoQ+M+4nTc+SV5ypzpM4cBUt/rYWin5pz4pH4VSkqWIBdf1KDFWUs3w0XJILeTiL7iUjx5ElnuZnoVGWGRIYtVXGLU2dabdynzok55dZKoCeFIYNn29bCNv1DCqZyqvBzgzU1qUZhgFjXNhW10AbuHkUCPMlJSFNk2SehotmcAip4xbxGshfwlBQiyOvtjzFKaEVPz0vc3DNa2yNRpULrv3MQ5EdVAxUlTxYSnreQjjZsIXmln5whwIq0UCrKAJqv8LhWLSonhAjIskfJPmxuwxzXFnlkt12B/8+IfnMTDaDcMnsMYHnQzLymUrho40zYd0MmiAbl7YF7rnRnLTm4ivZEgwA0jWVasXHeaqDbPN9vtAdH9R7O7eH7EL/PCXjheZB76x4oI8Yve3sdHRHJCe2bm3wWxavYKhX9Cewh4vjJNE6vLUPgC0hbcZQPrQOnA+XbpmgwAtzo+uZYiNrKin+dhHi9HlayDo6eiVnuyloRgKt3YpzF47rr5GjLx4QvJjfM4U/GgVUR3s7mm3LsJ2dQ9Q5wq/74VqY8UWuu+zxWVO0DxLxsVTkz/o+OO5QHwGkALHZwEOeQqiOk9IZ4vVsoNleBDlFy43f/5mlRnNtIEx49u3E/7d1b2+PN1H2VW/FUALjarRM+sssrC8UesZowz5OAZLXxDvmTq8cDW7lt+d9+l2/BTtTlVzTinbFoy10bH868wJTWBle8zz8dxlTETuYI83adhIm4Sb3Q/VivCze0q3pVj7o798f34EeSyyWhY8bQ43wc/i4SwC/94jYvfedfRgOh8I03Uco7ZFGkpBKOHQ03QgnKBwf6nIhsqMhzcIN990FGojsegNaiEo+C20xTT9mae/lVeheGj2MV304nwQUwr7xgOKVcG9B5G9HPj75i+vDctz6GUdYZJKAMD4OjrR9eXLFjZix5Ssa5/yB2FicUYW8dhXKwSgN/M7zyS1alAJcnHjKD+g3WngnLGNzJ+5WTpN6qvo9bqHNKfTwg0a11fUfWLUu2MaMqpRB5bf4loaSemK7ls+v5mKMzN4YJDdn1LX6OTudEfKBhtPH8I9lz4yktRz1UyY/jmCltlKcDK4+vXkoGkh22mmfViBbkBdcnwdmheMdApnurC8sh+KQ4cEVlkczfelgdhmBC7uxeqyldTNN6xl4y0AjtxeB6x1nwAmbZtcHbz2Nt0kHKlpHbi29KXtknUIKN5+HLhhGd162mwafg1VDcs8OZB8leYlI0kMf7frpJg30zLkNklR6MK0JH2omSRXgEjaDxeeuTafHNG6HvE2dmRc7vDvZsbl+F6/02VgoeFMnzir7ipV+9MLhg0qP94HztEdN0DeYNfywnt5zQBa44bOlJSfIxSgg9ECv3Y+wfDsGMJKqEL52nwmBqDlRb3XEBm02APb+e4B/mh/FpbfFXYlxN3WMDK6QsWhDLaTUh4AWDTC7Z9sNSnpX25w/fdq8EgnaE98FLwj8R/zORU76wc4rjArITL8IonPHw+LWIR0ovQAaLcdA7u+72HQTcvJU54nUNNuarBbOWYObQ2kpE8DUxy9C6/d2w/DxDNSSZm2BRE07CvLhDqcBisjjApQsYDxKWdDnTVAyulowePO3iTcbifsrgGTxI48TxVZuel1s3YJ6ntu3oryVyPUy+o1lhKeK9X1Q3ZDQIPyJwmLIWNYCgdE+v0Pqq+PMjkbTeOuzf+Tx9pKIWCk9A8r3dHn4PZcYB4N/SfVp8iiFNdJhdwTZLTGvBRsRdYE1z1hq50+c2aCUIxLWb5zyQR5hZ1dX6WNnayL5zc1H4dmd4ZTlQnLB0axiexluuUpzUmgzabTNmHXmxF/94LP2Se+GXg8Vzmz5jW78EVoaLwUzXPIq8Oxl9mnAsoeg3M1hKfANMCcIM4urgnKAt+72aW6s1ardThpIH1xPHROCKCgZRhopKJX0dgxJxT7tZsV+mzFabFE6Esb64xFdmU3A8VayHZYnGyUmo0+ezO749Tb0yYytGOXhhx35VXFAD7hetNr8Q93tDARDS/CxLVVJMqdEMJZXOp9Ne+4hW0pW6D1N3S0E/yMvcREPplJJPt05WsFm/Ul8QpAMkZtc6y3u6QhEmbZiU6wulPptHpHaWndDrXNV4BNm49ZUaLbOIFUQFAVDBDZcR6ZWHcziajAtY9QBie3h2J3CHsUHgMrZm8OnbgCfWYgtqHJ5fUOMgtVrsfpqOgolCXHOH/LAB6g2onsdli+18gkYcDEVGzqrIe2qrmS1z+NwZCBwxlMBoXe9zZt17kmnDcnKgsQisWUfMcTerPjQg3KPx0wunmFJfXimny9D9tsNWJqDEIzUeRhCES7TsxWGF2bY16oOp6/yefJn/jL3ka8a5yK4lMukryjUnFxnIaTCB995wIIOsLE119IyfhBigh+ASZuSRP4cQ9sovVcqzfonVfoD37Ssq1l+iAzcOt9chAcfIl+RAXJtFywvra5sQmARTNofnKW+BK5iyjVxelI+JSH2efAL3W+x5BOFdJa6wW2v1tGkAu6xeg8/47EWqa/nZSV5LXdzb692N3HRtmBkdqXdP7xz0v4oAtZKMi/e7QKmvr4R4TtHsDOhaM5V3G3undO1MJMfUje8pBX+UGpwA9iAF8c23JEFpjBBgRD4WTlyXhBVJIHpBPY1aWezAyV8ooNthaUn4i8LDAS/rZtjDRgbvPH5E4+QN/jlil6JHd6onxMTayM1E/HRygZVJ3IO+N9952mUmSn6pQ60WrliRDtcy/yb0fGgb+zu8TA/UmCE8m6aiXbyqRsp+9G2j5VBhJ4cZME2s8sEixCu9Hvxtst4logN5UYoLu+A7JYcDc6RE3oKxE5q4lF47u3RDazsX0IHnaR7vo2DhYCfYpQcJzuuq811l/Wr269jevhnpCardlJuGsrOInsFocJC2qK2jqO/AcbOJqqGhVwS+E4fYwV8avfRP2KMnVpp8xQODjOqnzNIdlqUGMfror8ld17fgTSJNj3092o5LLrnZ3BMrh7PsGplDwQUkkQd1fW5iuJ8ubxjFVAi+6TXsZY+ahAtxi1fbXZ2ff0Lw3KiYPb6bQx4vytIFKUfiG6FhIMjkmGYMXnIpKwNoMa2sWMPvEg2DmIwA3UCd1fWRMQ6Y6AeB3ToW5bslWBSP5nb9Qq6giyK9qRR/fDU5ji2T+C1FSLjQedUEVi7UZvrOR0Bwyj88xXjk/SHAu/bOSbCCXDkKlSNLH85MaWBwZsW/lG2jyV2JbekGEDRVhVxIWBYHI/1RSjEr+GX4s7BtsB8IA2FmEj+8LT1An7iH9lpzBMkzz7shZsOCmB8cdLMtUY08GpvJ2Jm1+mp4eDt4w9KbuIysX0y0RwbDYd37k6j9836HxyxoLKWtUl8jjnrDl849R8OvCP4LiJ3y/yNIhgD/uYJJ2+n+Da4zNkQ2JCrtZ6e3uT3DO8mraOQS0W24AbMSZPMCEI3LqZeu/1lNs0B7Wwu7I/UM8R3H9sPDchDkBTcT4i7WOzapIKkXLNDeoTU8mRCcvX/jhWSvkJ0MdOswHymq11ymK6cgibczzl8neDLSWzPH8NgiKs1PuE6VkHfF4JZpNDs76k4wUG2EFkmbMhktrep5vq57T322hJcGv8sC1id9EG/K4pOfAjBOoBj2RBWaYTyc1JEoUhIdWRaKvjzz+eqPZsKD9OjFmm5kpncIu7DSF/CnZHzZwcnZMK4gT04TEXRtSooGQHKNs3VxF493z/ftMu+Nf+f0JhqmeXBlwOz3Uuw4tfT6Gg8wVVgOgS7v2zfq3iiyuojjzQDxkBcX0Pgr+6zSt8r4PS3qco7uKfN1ccDdwoDlQ05i7P1TPKPH2DZcXmtv6IODTKNZcuInyoWd53Zaf9KZD9LpTfTDvMxyuIXMgPM2WpbNd3texDVwtAivVXmdk63fdi6bzuC5LuCvwkBlqixQAv9QTWSkckD4D+q20QVyxKW4aem497K+s0ZlYhJxB/xvCs20pbm2W6Tr20e2hh/fpqv5zhMuXW1HM/q5HbwA11NhxFf81C3+yI/C2fXsObOPBS9cjauTw/TEluGkDYSZhqoSl854WLj+o+5jVmWJNLxROq2QKne7Dlp1TeTnEC4DcuyNX71XyS3D36zua+AH10bkaiJKQmSIn2hsFzfRvR+4W7AYdwOkuQ18o5ChQwCBMt24UHMKlS60FXYjxs8Jv1mnrRjBCbhvoQp9uCg2s7+3GmsQzf5Is6MwwMqSE9vUqvqCqv/Mbd60dDHXzQT2GhB2E91ygOiiguyN5RQPBxL2zsHWrWKvDPpyZWSZ0DWmtUHTBedHSPrTZhSo+9kfenqnZYJe7Wj2Vj9k/+3l6R3G0KrD63RoTQwsT9u41iB6qbFPjxXPdUUxvd8yB/B7121Ukhgyu65iEgxz4rBawlYxbEaOaV+FR01dO5PkfHE/X77+FS4qcOysTqJ9geIAQ9qgPgCHIb/kuclBVNfSmiS6RerXEZTlLiQdBN0OgeF41BRXHNkjUP6FMm6DKabkswUPc8Vc2x80KTqjz3A6I8UabOPrjDtAjGXivxxFZbQBIXzpIYPlTUSKrp+B9EYJ9DHMCfNzfFUxL0AxgOJXkJi80fONSzhbn8RkMEQXFaeGr1MANdVF3l+vNop+DX5Zf5V5mmMV7xIcK/WPXLVJzbWGgOPRoIWBmMcKEIrhWEh2z2aTgnHR7K5pXw/JdkMN0gFI933kBi5UBo094GqdINPyEEBs+Uuuo8y0vOaUe9VAWBXso+pkJCwg6LaGEh6UeRXvRIXnCe9lPUbRkpCBY6GxcJqcQEHrANa40D3JmmNckHP/QIWZX4zObffl0WCjxTlu++itFn/ubJ6PTLnsdEGC2ozMhjBrxIfGxFVYwECRVBm2VZ1P6iDds2n8poN6pAjAmvfGd/1FJVHqRWVMbL5GA3BW52DeLR9eQHm/LkVzAQ8mCAmAwS0OaS3mL6sK/ej2kRYzZz3dCsE6ZcMj1q6n3f+CKVUg05KsY8l6Nf223ywn4+YZ2rbUBqHSbMN9wPDrbfQx3edhZk4L01a3ujXMegfpQP9xsP5mKdQxZkm/4VXQxzxEDlGe/Y3J+qJazJZ57sp5MnE/SBoJvebHnVhuQM8uew1YTge3qzWtIDC+Ey9OUzmPd5eLzvyaTzKr1oqT21aqzI69yZl1NPG+7mQ4xoovmXSZc29/FlF2FCvSEqWcNYVgSPUebJrR56vKGvS/l2nFa/51HtHwgMi9U9JPsdAC58W02xcJuG2q66tnZ8OpqvnwK9FfGf1U2q1q3OJXWcriQqzCP17ByC4pb8tDbHSECmyacO5f7rCN1b7/+79W6vIF2zfsC29TytBLkvDTTb93uOnJCh52KLacu1y/JABK/5LH6WnCZf4nBfWkmgJa/Ytzw+OUU6QeuuK6FycVAm+9ZbwS9fczPUoAZNfhyP0AUYFJiv8Rz5zXYNZEDzc8QHtYbdcR59HiPMd+ZGiDFiw0iTdXpJzWbWhR+Yf5TQlQoXZwYE8fTQdPUZCa9StwqpejwzPJx85UNupA/VSeOmG2yOdl81WLPovJ6pKJMtnCbz5xol3MZnQepl3xJPGlZiK3ZV9fm4+DH5uEKilrcYPdBIS1i5vBsjnfN1MLh/wKn2WJZXhhYns36ws4s6nu080gzozAX/cKUWqcoju9ABvL+faFx2krSjn/o94rSRYNLPxRnTfPTkbitb5w040Qhc6ZFVmooJvEuai8jXyCTrcoH2Eet5kdE54ZRIe53k/9VRirW0axEGySLDkIzs5YtYCaRLjqCanfYlSxk3wNXAXDle+NnMeKxF8otwv16kZpVFEQxO1lHa7v/rqOeMcsySG8/EF8f0AEa+cmXehovcq/SEEAYIFl3FQct0csMdz25EiewBmYnRUf4db5ydNYQfhdkpXfcSKag5MqCPmEYGMLOALU10H1/RQ5tyCs5UGQUcU=
`pragma protect end_data_block
`pragma protect digest_block
b11a511dd7574d195e7d504614c4196e9e73ab6fdf24fc4e9370b312665a40c7
`pragma protect end_digest_block
`pragma protect end_protected
