`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "18438de6b00f24f5a2c68075a02f6ae4"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 11780)
`pragma protect data_block
emuDIhoU7Fdh9nbs6IVL04/cIEtl4hZ7OZny7C5G8IplyAqLQ/bwgLIOBmyM0m4180WlVcB9IvJ3W9ZhdytyEkJXV99R7/bANjplzx/DhrImBnwz8+16BbbMvKjmfeuEPMrQ9BnjyfQXf1TTvp8DiRC/miiFAFPFP7zrXKG5h10vY6wdcXxK+y+JrASuPA5mHnp/E61w5N+T2I8M889DysYnF/6EintcZWxsahCUlVjckcrUv1Pq1J053LoHnDD5QLTmkMJtXvtYI4oVYGqDiM/+l35CzBh8jquHoyCp+CSGJNzXbNmh0/um7aFGC8Eu5dzOcqyzmPwE09r+oy5pXjUUoAzQRHaNhkMDsS562WkN3NYFBS/Lr5VBabMBKXACVgCav+d/2HgiFqZ9w7OZXUWTi5Bj0y5OvxAFpGmPvc1WcIrZqXO0tAZR5d3FxjGnjsYEqdhJvr/az+EYjUTQvx+AVWnztHdZPzZnxWX/cjDh9/5PCNfxWzm85GPcfw90xnQzf0GDvtB0uKtch6f5yvkwZshbuSCutENzSPQY3z4k3ghBoAOQJ3dGnm+BlLxAaz5uFY7YFwQvnZgss8SV+U6tpMTKvRNM4T9x+zfDEVo1LCu588z3o3GRaTKeqf/0wkMoVm/U7fiEqZw6J1fR1u0ylHpnJaTFz4WhA9H/0rzjL4nU9Lh+MKoPE7BN0ygAx/A9nFWt0/uKu8C0eYFc1BSKctfgEIUITpvL5xArGR823KIt47tIaxwUHn81CwSYMvr9dmgZYSHvJjYL+rQV0P3z8dwV5nJ4cPuFj8dTzAetUyrBovBeS8BeFnKHq1c1wVKWvtsCYU5AYFyywZ+ekUIU6bOxy94J6VObDPzI6PVQb6xOaWUf+bwxF8wA3XYjJbViPVe4XBW3VZeiwmleo/hHU313XN8l60v4z7lZKahQHh5X04k4VZ2VCMPdSnxBzKRP89hL52v9w28L65O7ivq5Sftb9j1ZA6iXkVdTxykj2FFE4VefEEbzu5+lZux9FsO8mvF5msdWffsffFcMdB5bajnNB+qty0RNdJrIFzWqzIyg1JWWvi4vzn5vaN+o7Hgo31c+KlkXJMtBgGEr0NZaDvM6YSjw5lcZDK1af/HZtCPXpqKzIC19NQjT0QDXf1XwmxFZ6evQ4JTz3ahttKGuA9sV/PjeWv1C2j7vlC4hu/LdVID6m4GlRW7L240Oal4JDjlw++mvMuxk/g+pb8gsZWTn2y5V7b6dqTTs3WXvtWRBMT5aF73i3mOXEnvt/sn/oQNPkGRYxJO0clY++Ua7BCRewo4TGOZpbvaZK21GeBidu5ytTjeRkLGL5FWuc61R262SkDuQ5bpH5PLJJlwa/UuCsk3617VGI5+kWVf70RYCo8wHuz69U/sYewLLtrIeE0TOKMidLJSgaSJc1KW1UoDllQHanfR79bn8Q7j7gs8w3JCL2dj13YaddIM/f9AR6G99hXyhNjm+PZ2Hs/acLl1mEx743XxhsSvHKeLzHpdQXXWKkuKuEbVIkUi7aelqLdOM4SV31FqjEL4kMknAAwb/8PgkwDvivjEC4v+FB5/PxhqsYlnv6OZHTtHFXsGJd9CU7gjYFwtgRt4+fbztypiYtwl67sT5OjPcisSz/wS+nNGzxObae5nQmr6CZtJYlmkvcWx8mn/R9veYGC9myjmcvKYpaMu5a/w4XMIKf+aKMC48rcFNxcy/vn8yWcSJpIZjjpkQFrDYb6Y3nDvJBOc9g4oJGfJZLxgwcM9k3qy4xfe4LPdkpuBEVVgBjBBXlpNUQkhxccS+/W0WXl6Lw3e0bVBAZ72zMfV2rgsPBMMQXyv8nXsjDY4MaE+51uVvdKOsgjP5dVn0ctrDCmzOcHmRnp0VjNC73iwZYS2jgL2yVJYxFA0CC9RlCRZYJyII5G4VXodshpPfUN/r+QsZkDmxFalko5h4EYVV5hg5UopL3vf+0NN9JWsrW3zIYTqvLK5j/RR3CV1kBsZXdMIcJya0p7pIUNu/KHp0JYsyrhsJpagj4xfz8zh2UTvkjFMG4r1cIiFhskxTqCTI92T+2rX/qPzNIQIxP3jPC3Ee5NMYPJ++8Ugtlof4bVvlT1pT993HSWheX7kWwg9Q6zFZI/SlcbrgQancsmnV3O2ftRUd//WKn+yPaxxtEGIGsHorXA+q89EmaGoPrQAJA2yySuh1mkONpDX4wI2CUvQXuCcrmk0LQohCXKkIfJzk1Tg09o3QfzdEbST0vTJEZg4DeKzh3qBkNbvVwKWfr9WOeRU1jZSWZE9nMA1qyQXXLyH6HT2q1srglEwRw734mbYywb8lzTBw9QAabfXjVR5tEUi9239nABk73OFVye4Twq/sXKTW49ma2V6ofgP3bQtOtZg4B2c/sdTMMcWEHk1JS19qFIsTqRYmOS7XNXJ2dAwPoJCv624+wC2+OOtu95GVdjZTSqSWCZ6B9l1ltBWCM3939g3cBA4U7sxw9YcnjtIm5ATYNNK6ARANVLR5Ah6xWG4teRbNntZBbfxm0UJx/ht6QnujwL+XicWGjJYw0bvF3hpXEbTQnr1ezQfJbcvKj+faS4TtT1aKLi93ui9ZD2vqdXAXd1KYRqKeF7eiuuFQhWn2Kn/JHce25FXYnESMdSqVbR5+fFpHqi8QJb7Pc9ZqbL/rskzW0rv6i03hfR/N3KjHfx66q3Dsun+Ps7ob0uCQFySJk6spjJn8vQAYywerIzIon3XWto+cD8PS6vOO1vsoLe86Cw8QoZNmLfvRaQZHFfw8grSg9rBYzwssYR3GGrfqx8hWVODgtMH5+DXKGF6fFrPboeR06ZAcDzBrYQf6yqnzfVBmBRYSGErt/cuj3CZ7El6Vm7REa12fuT2OCOqfMHaIJYsXbTDBgypjtFZWzcCiaUY9Pv9Fxa75M1kn5OrR8arCk198w3CwaqefRGItC1E0si0pUScMzeYYsdzwJV2rbWh/8qXw6G3r282lZ7cTwF91rCg+rOviqO5RNz6O02EtRUAZ2C2ePfvnrhkILKb23KacuNG3P6Lg1sb6qAAV+5TyaA07SiXKPDkdDGvrg3+0oAi7thtP0XXzE0r1RddVNLVQAgvaDD1/Cer2zV8aKre2WrsNJ17ZdYvZU6SsEyoZMhkG8ZaCpcMGfkSJ7OV+P9wry8K8kUwQ3vxlfIQc0AK+qgZTzcKSwwYrt3mIaFE8f4IFML7NvfUZQcjaTU7R5xmaJNMKrGwX1wyx4OuGPQzcfwaY/xjCaFYEXHdZDYEhQJuwIFIo7m/5mQBES5I7HcOCFEbw+fT5HazJ5QcpqC1MA0U1uPkUt0P57P9XiyrCAhV522NgZMDh6/XcTLuAgSC7T5mBIGTlAi+ZyxmmMYOBm13YIoJDR3Oj0jtfXTvHzo8O3sAHAYljQWBbBFRqSF+SZ/h0IM9Ml5ApeNR1E7FsM8xjjxW/0/i1NAQ8ryhogn+4kyv2qCsefXOV4MxxiW6zDtRf45sEbbh+wQi969gtybxbDsNQ10xvP9zBbYf1X3lDwA1duToySQtz4G+wDvHU17l8QGji4iHNfVOD/0tWbGAdlJEs8MwNvGcvbLXHSUjPwso1Kq6uVHRcnK7kjYvvY67I5yUs1QLlJqVxUDCCiL5YunGWaWFqznze9Lh4qPKBqqL6ZTzHRo7+wNKkTYEFw7ryCY9Bgv618tIqW86OofZf7F8FnK60jAVl1kwZNokUCsHoN1UKuzfHWGgSL9JBMg6MHygMK8StH1S4CGoPCJqTBnGvXVo772uF/iddNeH0nXPQ1UpMCYH7tASteKVIgR57xPBip8jbPkIgD/k57viljpYvXgvUmhCwJZMtAgAV0GBpQUeMIlisav+3jwf7NT5V57WjT2ndpKNlGoKSxiYRrCMceVNcIhmI39UffTEkKjajIiisWk+s75yVxi5RQVTSLDhm05LLbl8/oOmXuPE5QraLXFuC7orJg+PDMgKSwUZB9WeSGRvhCWVlF2cWbYo6Rzybc5KdY7bLbMOH/Q+1decVZRrDnDqGPxaEa8HmpLPf7/i3SotmKPoAo9qixQIhvXRsqVcef39f6dGmRedgOgc8rkVjqIcL7dadaSEdkqbovVtvzm4KgmV5cnC3/W6tnSxQt1uheA3CGQuWmf6oWZINbqEe1bTnGy1h0JginnsBkngv8/cwhMPY3ohe5sn9tlqKL/xL4hwhbyrR7THfZy4JT049iFxL1cVHUobDI6MvWtU7SPRcEZjhjjtxwoyGk0aZjfuhOE/pTkFbRUSLTAkRHo2p9imTF1RNpJBfZg6Yo3H6wkGfQMqFMIHhNpNcjJK9ubynDoMAEvck2udjFHS/uvfDvZQIQV9F0zaiwgA3DtB66QS1xv24W7KeN7zlUK1GasNEP4Vfz9g/u7eLnBJ2n6asvocbp+pya5xOwmutQbR2DD12qzs+NUPLH3iaiBfhAN/dwBYU6pXXvwcoCXX6VG1cLewo37w5nXe79T9brcLEms3KcPwVFf2Glaa/tguQnERdF7tmfdnCb82nX9Hl4jkkXjYAbXgCaVNBwexDJcJO21hQ2lWF69kHLMXdGBH7KrmMbTmLUWZvLPln/fP2zsoJVs0AndzeYJCb8pubxj8X9EBiv09654f5ScRmK0/ms1hH43/gnV2qlpl63za72PqnwBJdAT0nNDlvQ3j6p+0uVY+vRRaAjXNPWDAnbhD2sm90n1FQXznMylLH9v+BAn9xyBE7d4HDdBmN4hLyWVkqn1ekF3SUDQAIiupoUg41CvA50ifydaldGpfZTrPpGuuqzRHgXkWIphp/yaALrIsovqI+PcNLofiGmLOOesf+txIEPiXhlV/3SWBe2K4tLXSPNEtObDcbtiZw91fBkNWyslM3u5iaCe0bS1UGxHtta/fCud2/fyuL8to3Blinb27hIn4CpAifnmCea2N49/OYU1MFpwpO7wM6i/MO/bmzvDdFUocKGX9b4LDlZ1QnpMrVqeDKMbLxLJo3Uj8VO7sY33V5SyiMCPoFysbgc10Kuvsvqxn83r89g2IvF+xr9Sm51pBATi8V6EfFtatR+VGgDdFG5y/M0BoqI1xFYlQs8KAvcMytbJK7E2QEF2zN+jOzZ+fqrXqRIHfmKJePCJ2rVeSRy/cC8ASDgmKzGUla+VHlVDFXKuf6BMOqX/1/Thvgf+fY7LAV6/t6P5X2+S79EE0UQr9U89vkUI+FDfnb7lnaEXd6OD+xXPeRsC2HzHjyiXamlyeDx3RwJwihbuCAV7jM+t/enTm4LXaGfPE0MCOw+x2edY1V0gEw/HfPmqDYuaYoIVAQNtDNk0myf5rYu5ixX4hFSj6bcQ+lgeF7/aseaWgWvakzIhPidVpyeH7NgsIup7PjA8GrXkT8EW9p9TIEN/SW711D1XAJzB+1HRnCi6eCZRphm3fEgFfbhzhz7cRKQb4R26HrgRAL+lR0KM+HtsLp1P5AdwiQoo7ve2HDetw+75hNCb2msZ9RuJhRNeL9pEWweZBgjuEcnTT0CVKiRGdDoZpX8XLwZfU+LdeshVzZLl65Xs2Y5UuQ0e6jvRTx7ybAFL3KL9wHSad+lW6LiS1UC1i3i9o8sc78rBhaMyHE7Dtx94ezhFNNxbmqeQpaIs5U3tczqimWjSf+MErvNiY9vgtsbuC5xF8lN/EvG7siEur4Kr2cSjP+TbADiYbrCsScJvPQofb3hlZq1u0f7grImjb4qsWpkoqFMs3TREm7Bm0x1n1IEdAAqMn3lwg6028FqX9VxmaJnweZu1OG29I36ffe6D0gIDGaIShw5iD5VCOqQ6L1/LPQ/8BhXXhTdE//zgdf7mZOtt++nhe60aHympEOzOSjIlRLqyrHrux/jt6sGxO6tqup+gQUsY+WikUkqY5RAkWrW77m27j5Z0vJolXw4HV1KE5q+bdL27FG/9WxJk9lMuWrqfTr+9ACkPIPRIsj3aEUHY5Hkifbt+yQH+m3muDsGnQFJQVMTI+/cjSSuAyrvsXa0fXEp/e/xidroCl7d35MOW35yyUmpUE/2d20f8TzYSptQ+TKds/ZYRR9G6zMifD0v2zWxnfhk3o8HLSXLmfY2PWttpMdZpWf43zohFnWA09JOvKN4d1jFEF7wB2wKiBAQ5ApT3g4BtRdm38s+DwtxHfZ5OoM0aSoMfhxhiY01NamABWZ0Uprw1u1h6ZGDRCOErn6oRsQkhHRebqe8OXHgr4yL0oemihVFcOoxYhi/e8ZA+r44edrIz9OX6j+9UgkbLUEfGjn7CQIznmdo8Gl/sZ3H+wS71IzzUE10lc4kQYbl0QF0h08RhH4ctP/sLHWdNriwTHUYBurojtLGODqxkXIjLP0lt6LcVkF6qW5HXtNVVXzLCvoUty93YqmvzG3w9UD0X+u/5ZWIdrlhzTlLjRQKWT10mNaIhIrmgltcwqpYnvL9zKlWsp0YJ9UvSeb5MMaaSKwiNATe6i13CEPtBjerphpFxoMZrPwlHJ+djxz5M66Rl/XcI6ELh9kI0bNLtEja5lmV0NTFkguGVyC6XAeZbZGwyPLCwb9HpC2bFXD/m3AwARNF4vG+uLtduuZMor9ojhkAesOHGWNmGLeGpYUYA/6xpWG9/fnBWbd8nmGi6i5BTwhNTYamcDfTG3swX8/D7W/fzMpBf+4oEbO1PRQAA0QhvYXRghZu4T1aw0shyPRiVmxqEoQCfn2VDq2YqAj/MAlPcyNXEF/iw+qvjlWg9aWs3JTRRfjAC4vzrdFrMVrh8fikS/cX0Uklm9ugFUHAu898rFS9QvQFtmVhqwD13hgMjoSj2K9oNnGim72eBsTqQgXYLiswhVQiHbOyG1egno7YzONKn4j4tit/c/s8lMK2FKrSUrNT8o8acfZL3CBjPfvATu99KMWW5hne500xIgIca6tL25wmx1WQZRnk7SQx0VlcaFhRh3GZSCcvjrS1rsZhDZ+1uOQHl0XBo8wBf1a2poYOqRIxzoWkdvMRV5I29ZmWYtmKO8h/UEXa4/4LeckQNpBg/ssvUgcBrIFU13yw9TwR/DJNeT1xP8coKMv5MCfqGOtpUDP7hrjLkl6jQtAQYXDmVJrydblm4kNYtxhUJfvHwPoaVdhpoU6glJyYxW+0CZfy958EIdsLKc05hTHHEi2OjsyswcpnXpOmzP7G14qVxjfKwsJ9KICJj9ycJHpMvKv/bkBnqOAB2dkrCT3aZf7VisrbeKND+YZ2hgxieWSU8SOAHoYyIG7sqhLLHBu80S9uFjeRWTx1i45k8c10zUlxX+RGkv5wIYQ2xMRkUbqQRZuv1vBPlJoQQ1S567IjW+mI3X99OqWnAIEkySBjThG8KoKVyCsRGti91l7Xn6uoSQuCYKfMR8p1xvb8Jo6tskB6CZq/2/pJ2rxbE+jGgOfGLr4VXb5x5mP5rKyAcq3Z2OWqOOk6GgbZNrRDIuQDE1q9wuGkAiT3D5jlQ1H4tUla1eXljzGzMjGxrnigZeqU82zBYhwklnCJME1NWc1oVwe+2kGcVOYAzLVcNqYEYyDIacd9OvMvK/t9/djKqHmdF+qESPfzpg5SOSasG5JVVoiyNgI7kM440moDet6H0kGXxZmezcitiqOmTViquRb8Md0FVXQmlp1CenjP/B1pSILcssFANqZeqZHoUQNI8+agYUuERJExKrwtEmLiG+Dpe8hTzLxjauGulGt9qK65aT6/erfAYEpfrHaHbq4ZZhQxLAsFoMJbh7asdGbgZlCup90UrkP4BOrOqfmeL1af8R0WduvCE0w7xC5fzknLEk3NgKy/6kf1PuaJax4zE25I/wnhqzIpvu+ZpuUdy4K0XX8VQtbRlwdlg4avWh8KJoPgepy2f+HeNsSOkRZVU/xauM6c7nkZiRcDhxikwbtLf7RB0wFBWAnUI7gCFh/9F76L3dEy5HBCE2Q05lU6Ll16N5XhQN3qEAay4HW4E7a69TUMHVpWh7dTcp/3v7gOdIWqRqF+nf+rJvUNamis4Ah3J4ZlZcDgh9kjaoR1Qdc43ApzJ9T60PaWU85rJpLfWbLa7WvkhIryHScE5Cz4VFaBiK8k6AYr35O6T4FL9qSu5jpBP0bJSh/BA50H30y15ujRly4eQleEFiOO6OaqdmLu5vWtCn9pQ9DuGmFjxWLHXyDkUg8Q2gfHL/uIPu6YzHbPl2TKRIK2DSQYTnCH93ybCMcezBguRPgXlY3UWGm6k4dzwifdDfZ2H5uDvF4WYoX4AHcul2wqDMO6HbjJoxZnNBUpxbzjBB2yXyYp7/cTsrHXBn3uiTvGhEGnKHVtYuuNsokJZ0w/9qFa1qLza6EGFtciHimGWwsKBVyoQ1QbZLASuYPs6ile4hFuSZ5a97U3UuEv/zO5o4CkMD429hpD9cZfRCQwoUjFHeKWSWyTVLhXhx815mwRgCk3/PSQtyiu3t/TbCSNbeYDQZ6VZua0IP8CFxcRMyxq3G17CQnD5Nl47HsAxFgswTgWQHIrjKZJ2fSx3r6HZxzFhi9b6bjt1Ttp2PzxUUNycBu6rKG6H2ch6OMAWiymNV08Y+9DG5pltwirMcfJ8okfFc14VNqvWPV2LqRsx91JhcHJEgdfqcHgaFraWbVKOLF/VU5jt2hFu1QxMF83a2RAanj4upL1eCLmZZ2TUz8/zWtzX6jWeb+YVzeDzk/QTvgJRGkZ5pgQC51zZ42GBTFEJAvk93k0eMXw+5ea9DMBJa2uZYV6VWY5xM5VehY+fMSzJYAvbmKPbQwRPq6Pm0vwOsa01J5+kleu70rtRj9JFmosel95B1Es+WB/wJvvC3INihoCtGYYJKh2+gEb2taQECf/TCR4NNYjA7EJzp5NcJKQ4zvxa5No7jm7TgsGG4ivIzkYrJSvWKI2+6+kF4P3ymAUBHXI9ybLxNQU2s76C4MqzwaVZOXLhYkkHkgai2vDywOUDys0fCgxIKJ2XRcSlEQmfj7c9kDZO+Y7jXLQoJ2hssCuEGMmI6VELgOy0gFyG4wKIWbe5IzgUufgo+J8M0OmjEOj8N58jHAEe15yGfRmfrrlUVigl/ofYquPx0uyaxfcmdSfntMQr+cA9638SLGqaQRj/637bwWn3lDv9iHbmFp/2fqDp1h6jHTKoLjjccz7b5c7zhFhb6MB+2cZNI0UZy9WdOEYl8aChghmQY3Dc/tYecUYfT1OSdzMdLsQwbYY6wmzRYRgutADynuG3h8qO5CVSA77CWvmvDBa951FVLE1AiWD85ViDsAZHoixfrdOVJba9t9//KSuxiZcKwgRIb3DF1SkeGY7XIpqLSCILYKNM5nxa8/1GTUGDUtVtJB1IY3qs30xcY/w21/HY0N/vF0ZbQDmTkFrQN6CzTaBIigZtrboYPLa64SbR8NTg7jvHknAfHEG6GF4/+pwmyUeVu0VHZn2OBBhb18O0/VH/ZjfRF8ulyEmr16qdtmSOqsVdof/Cx8fVu9JWQ8XzUQg9P0fUBGIOSdUrHl22bu1K+Yn4p7BaWyvVrABjLGOEp1YRRJOve08sXat4Yy/yXZY8zKUDlxdIyKYVDN5eZYBeRgB/pchQlALQTASVpykq6lAYqN+7JqmySGH1JTt4NSFuE3SKFRbtWzEgtp//1p2xIIpMZxO5HQRF+Y2ygFQvEgx/XagUCDAbPOtWd/qxIk034fyMQigChlp9L+LU+pUYvza1EPRWEOqjFOKiSnjQLK3YdJG0N8aUYuRJ6roIQDGv1i7AsEr9JWtPod7MsMiZcqBEZyqWv5wJArwzhz4LdhHs4FpcBo1ZKF5gZqLEKXoyvESdxuSDR97Zk3Yc5u7sxgupY19fElCrpV9P/Rxem3ALH1lybqJPDTv3cy519tVcDqYOMTt0dC6D0nlHzeF7QitEbyJg2IVlX0OmxYHeVYDYpSYPsdP6lJOsXuPOJg8sJczy1MsX005PtnCEy3GRjt5QOel2wlCrn1JwAiKG+2m6aA+6qjWQP41R2pudPr1GphqQA+WbGP1+MC9KtdZci6AoUj1aoYnNVl17yLXPOVyGGJVu1GFoDL/GV1YzcOgQLzDgql8z33SsI4nXjQ9Qg8Vqh36M012tZG5nQwERIso6Lz1rReGNpwSfo52u7xRZ89iI0aez25V2ZDwFb7+yoE03nhMnQJVFGuXOeUzXf9AbawBI4GVvt8sX/0tZApdul66TrafV+vHs5BfegOnmN/yVUzPrjg+lLuytC0eWOL5F1ZYq3EaozYXCr1gBPWl81picz6YLYohfu9fH6NvgdD1bZPtHkM7jVhbWava2i9v0RLTxNM68NhtpXiDQhcgGn7w+Z53wEjFAmHjDZvYuQ3AIlnH/nRYu2EbuY7dOdrQM/88dT3OweTp4MMaakTKb4ochO5D+uQN5Hyy3NmluofJ6LPaZJU6WdLGqQLIEtGurDtt7U7EdP8XVSVmJHnRxQLlBfiupMfEBK73g7pBtfXp82X6vUUiqSfifgRo2I91wY+qtnxCVbj627qnsJBs9zAsAUi5tJ/m4hUM1lC46u7WwlahdHa3B6bn6BibD26++y50nT1MOZNicjAAiy2W9Sm7u3QDmxCdG/VQ1Mt9kWSqubLxdjaOaLofmOj5vQzfkfMbt9zMDZNu+qhEVI5wCzF1TH9ff1g/FbJOJvRNYYXkFL67/AYn2+6ZKucuHnmORItO+h/JdSiZCuJOlnOtPG1BM/rnzGYuInPqIvx36iiBw0rz+TJG51R0PNsbxtthqCA5GzcO4CBtvaNiHvdMhh4i9zrNJbpFljjgmWKwBZxh4bWQQG/b8MAuxqR4UDOgwa3CezPb9U3E94TNDAFk0tbEIguC4bA9gilAYHxuXoWniyrkdg1qle0mk9bWPLmvflCs2Z97UFG7w3KXPdDcWQJh3A7sJ/uqJGRkteXAPOys2mlJ6hoam+wf2MEdkSQnsm3iO8o/Dl+miPKZ887HsBcmudkMhzVevjgTNFbo070ndkn+VJrOnYczWHfcGNY43atP10em5SWvKUIrtsOORss+YDrXyHoBZDmSbqerYbOOrHqocPkrgY9RXq2Hnj8z6Xl6MiZwvWEKJRUkpF820kEN6gWwLc/hKKv413nclzcnuNquEYKD9YZbmW5IxVKVMzKkEOdM3ax7pUw2Yfo/pD6U90Nvv+7yN6AM3MxBq9SL2HglHPvGv/vmvt2VtyPXv+kO6qjdrbDYAhIFKs6ZBFn3JNGjWylrBGQZZWoEYnRcqQDFCudYpJWxdBF1RV//HHOqCX6OpsCxYgOlQ2oEu4z/oqznQOrTt2WdXkjKsxZwqHNJHISAdGyejXOt+O/UZ2EvEd/s8W2me/GaWWNBGmqqRDamNJvlcHI4ggFfRYT8S539P2M/wVlRiXe1yw9WEurTizdlvlc2KhWbS3bbBgE5bcdBMwQ/ievnf8wn3I/XIrgNeQH2OFZk1lGkojC2j71zKdw6rcvcrv+eAXNeZ+sX2KVOdllj9JOCGDiKE29btyWRSK8Q58qOqjXa8RM9e1+yHfdFvEW1IhZfXgDrNpSkiHvjhua4h+Jqu/6jBwGpgvZ4Sxm0PVMTDlYlilB35QNKz3B7/VitEPzyavBs7yaLoJCv61uhkSfYcspMJbaP8O/cXGzTAGy/+csTSs63WfVm54eiY4ceGZCCZhd+7SqRET4Oe0qhjd9DwjwLd7OzxJZacqK2PKGJmQjknnRtQzCZ0niGxh4B7T+hC9Ur53tBat2WRlXTIxcTVuIF2qTe2oc35PHQVBrEheazcZbIKKycs1c+KvqvOj5zxsB4i6FGYZc6cRSc3G4MdoG5Ul/qebw5jjEi+SKHY9ZW4C3eYwwdvMuGwpopUCBp2wWXElA+On7vZ77YeSSZODD5HLU9PDCie3mjOnSp+S25OLqq0Xw8DMvkLJ4dsBR+Nwkpof3GWlbIi9Q8jjQeOnhmlWml24Ktcw23trSm8ApfBWhsBp+lKh2eTac6XE9lhpygp7W5WnfeNJA+Oo13vuuWLvHKR7gvwAoqulw1+797UB5n02xeGeuhnShaEg4CFntID+E0nVoApR2U3nzcPR+VmCpbp2jTEuGrZrf7+FTOrscPxeFGgQMMCLtOUj7wF0t22222/nLJIfD6Jh6M/EiyKGS3nX74cMcABEJhPWNOAThf5iXr54Ns3DwqYrHt13D2eOuJHxeFo0W76oZuTL5MRAaIahzwlkICIFXCcgmBeA9sFZFpcYyuqgC2hF8i0d9gVjauGy7yzXoqjkIWjvopfdIzuAMkfSM1GKjRWn36H2vNSinOd50ecrh8ffyBsXfDTjz+c5rIm3hl5+lXLtTD8RhhFP731IO9FEcILnA/c4uhe74O3fkCVj0d99IgKKdoZQ8kZ/nTUhzRpVJJCeQ+s05YUuQcZd0sNkEjdyX5dgr/cw1FjYsUIiyTTW1l+ApLg3JW6VrPqKhVJhelr3vYiX3Q/CBvIHKSUSpdMlX9hf2PzhrIexAzAxV22LcmZjs6r8BwO/+EVPdSD6PaP65kPOvjgCaGCzTkdj3xJj3ge0WHPOHgrdWKd0x1knlOPdJDRr69itsas8CXZAu0IS+Z4GfGmpIHLSCzH8GVLhCEH3TEKtVqDPCk2cXRDKvpJFRlz0R5v7Hrj1TTbUTKxZ9BqEHLPptynald8mw6WzXDkz1EDhPdUGzXKJZ77JPvkdyicOs85J/8NgtdIrQ7PBguHV7kJeGwVb+CC66kg4O3LZS8bRX52RWF+AwShuP7Wxsn4JK0IErqyuDtRQr76WSTs6XwrCgx72sDQKD5vDZW1mUtNlwc/ThX7+KONA2pnEnpgxLdYEMgh5cTKsqTpo3hTMO5OElcMda3BYvR0eUyqsfa9JMybDiutrwsYbxEIobTHG5Y9Uf8ymlogbJYAC2u6Vz+B6D0Q6yhPZMDbNKjD21MVRYkdPQfbQqTNS/d7J9SAT4FUdZ1H58N4j74EknbZgOORLaPhX2pKFKMc3+PBoEoRclv7Xk1rILcGD9tWZwGXHzkh/Hf6jZnt6WL5Aj6z/eR1s/yeYvLtPOCIMQdP0IAFBRpULcoCzUmRc18XpJHMUR1yJ0yougMsS/NmTl1zl7aw8wJ5mXDRXNW/JATOajgIF9JFJore1vZjgzLiRQMVQS+tuISzD3h8q8uV76uuK3X/TpzVuzVOGgOUJS3wjr5A98r+Ft4bmcaMOK2PJ0PQp9sODSpqIqoQ9CSrCuM3pkAZf7VwuX9WBmX8YmuGfY25+Q4I4+4oLGSCyiMdBlOn/q3blV6zAUbB6GjXkacwwY0uaCo8XXsqHF7TzEJ7gUqrYgMnEidgwXNXxMd/n2UXEcQFr5dHYo/nZlx9kvZmZ2U50bxft/JVnR9yKjbsLU83AYX0ouPEuyl4owpuqWEKuSYOijEmrbk/zA3THgyoRX3QVw1X5Tq2/TG2sEEMZeVeQ94QfzeqEjpMjHaWnjT9vP0gm7IBoq3Uh+wsSFvqddvMmfC0G8OgMTOGMy6Kd6JKWFtCUwuqm6wuVuqiFMUceF8lLL+VEo2pQYybtl/N6f8eHk7r6SRuWQ4RuGYXGAckERqAz7pvrSHAFqgVBs9afNDK0L5OLKGVSTCw41ZDlpK1uRTtW7HsKa3yVUSRTaGo8kSuzaRWGAlXhUQ3gEOwr6V16rTOmrHK/k8u9Y9OsYaGf4rpoplRWog5IZtCgPGPK9yAwSsoVKKyBmjrRF3B38+BDY+CDMT2YOsRZRajP4yvvorD1Kgm27ofkS5dLq2M3nl67iTss2wmN3xjQgd0D1SQar3RU6J+Mwulz6MfBPUg9CScM6h+obd/i/LmGmIF/AnhZ2tHMRjzDRZLVQ3JnZfjLbSUk3Tl+HdxTrI1zHy7GToutnA5rDFfSRjqz3xYvPGaAmT+cBHP+cJOSi8CEI+UoezSgSIhzkz/wBQR14+G7OiGr9+K069J1AZt1uaV69QgvvmsMJ88PveeQf9U8QzB4POkPxfCiy8FpDZxyPq8dmR3QstUoBrFiULEw1f0zReStd1SzeCYio91Re9inq502tuKdBwE9cvhMr+omBQV0ctDTq8Oqdxr8y9JY1YSJkofjAILaF5tNWNnGXqcaTsIjfBP+cUnQX1UB43XRuSpgOMbDgAhB26b/zJvmGEZi0E5w4gwfd5iMP6Ee8wgjQwmzRcgBNrGOTY6g4zpJFxQDRGk5e4mAwXedtKlYoCyp27Ll0iehoTXzort4NMfTECIaMn9blPoeUJOFicbWScJnjpTWvn4JVlNUnpEEyXIUZ3CwCTawYDnggwadwrnxoKX6jQXxGFlXrIkqpTJBpGLKGc5Op9ZuFos22DllzrGUvRw25szKJAk2w1jVUijlXHYA5TBFBuZlsLHEeYtnIJA/t69USpqpOiVoP7fdaJFeHyqp+CRfNCTeeHME+AaU9HSE0pOUvpyu0KX1e7GVzdAdhFOBxR5KX8y6gaUF/RSxn+9j3AOmMtlDA5OjKd/lKO7QvkwZkXyoUzoL3HwwG1UVmgM+L8i/WQ04q8mGFjQr5xYG2HMveqPcj/cip6T39Q8S3Q8/7CSyazijUgCt4IeHNDCXLEe+DhCI7qt5xTzvbzsVoF/rh+SS12cYoKyiaBe1U03i+AtKu2tiok9pWKW+sozHrPXHewWQj11uhvvWr8mdvD4r1NUpi8BB/IGRP1XrTBae+Sbc6C7goUR0DDq0J69dre2X0fV3RBlmIuhYDAivgtA5TjDh05/tHnYkpsHZEBWhMa7DZ7KRbDyUws7yQ2MdiE00wkGrVFVoRdi60Mn+4C6AgtqHhq8U06KMhXQd1jQoaWYPS5GzpjoVyvh8EoVqzGKvhdhhDJvvQtTljFeelosDga03mxk4cbXK04Lf09n/BrEMCgVJVRiuGTSpJmXnKeHBE1JJv5xRsx5A7kyQKO20gFlY8iMwTFbTm7NTVOXSFW738WRfqG02ioFfBAoEQ74byxs+/w8SfJQP3FXCB6TUo6U658co4myLc+z1HAN/To8ovk4CVgqcyMfaqlmXyX8hIM6oSB75zKvXRm9NQZ5XHJqnvC/jitb56+3lL7vHLpqqIA2RqoCUm1Iro+VSH//rj/5m/QlGiRNitGv1ZJArmxFtvE86nwX+VjamXGUdjZOz+vgD0tKnk552g34MM23f9savd8iPJfap+0HxlAknu1oh8qw49O2Cb4oJ7UdMFTfCm+HXiC9WgHWJAQBflOAhKTIM/NIlRzlCYQvDFicBa1nOh2lPKbkO2b902F6f2EIo8Ev+hpQvC4uxd3/0ByR/bejlMadUzPmmOEzrnz51JcAYDPsjGG0HkxjRSOFZ4nqIHWTyQEFHfv3nU4h0kMcD4YBoYx5pMqcuAhKYYgq0JoS7tFo4HUQOUPMcTflM9ggYFFjoTm/AuSBfEMHZYNJdeMSzOiYq/vrSMyuk7TeROG96Fi4YrXJhnlzm1loDRgfVkSx096mUxDiC3w2xkU99wieBoyGq4MBiVIm19ovIJPDxH1EDNRBHNeA9mXLRVx1zV7x6/tW3Vo8kUXkxZbhbRbSEhq8BqGft2Ku7fWs0qI/qlPXkeAaXNPH9Rwxyzz4Ybe7EsUGWzfm7ZgVejEKJ2gdaLnKxGv2WOPjbgU+QFxv9HqcME5n72Wv/mvbDul7wH2MV7EODu55PYJiKpwvq7ix1ciiVgihaJEOZru09nx3I1BhAwbcTFT32tFUQ8vucrJmsVaDT4XEEMsNdLNXs=
`pragma protect end_data_block
`pragma protect digest_block
0b70b1c97461f1836f5416edf70b137a9560cbd9243b6b31630e9c8cc774dcc3
`pragma protect end_digest_block
`pragma protect end_protected
