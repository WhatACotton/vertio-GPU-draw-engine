`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "draw_engine_product"
`pragma protect encrypt_agent_info = "AES-256-CBC"
`pragma protect key_keyowner = "draw_engine"
`pragma protect key_method = "aes256-cbc"
`pragma protect iv_value = "0a45606de1f4be41384ba9e3fdb4938d"
`pragma protect data_method = "aes-256-cbc"
`pragma protect encoding = (enctype = "BASE64", bytes = 30501)
`pragma protect data_block
gdZcIDoqegoaDBLeF1ZEfzaZJeGFFW64BXQc/DCgQSIuDlDgNfNKNhV7bks/hE3WemtbHJagVYORdmL6L8w2cVJnoaciabHwUXksOK8lvllF+5Sezzq31AvNdF9S/oIDjv92rkhw5+s1rcVLw+HmjS14BjnbDToQnpkscO7gA7duZzcykGnodd8jm73r2U6q25pL/YZoTHthPHSeGQyUGGm/d4/yGfQm8EPtDI3cEHnOra0x4uZIXvLbXlrErBrb2f9RiwVpX2OO8tvq8HzDGzxB3jsUldg1Mrbw/NSrRDlZTM1lfa57X8Ae3ypNeJWlQf78NXX2HShmT8SMoKifsIOlsThKH8+yzb/xaOYwpyYDJvyJPAXR66ostW/xtW5zQ+0+vBLM6znrDkIecWO5juCgCDb3O8FoE/vPggIatyVDFuEPN8cZCR9DWS1HWLJ+ZDQqk274HgWDEJVDG4fyolfrRkcb7kKFracEWMpQhF92Yg8Zt6Huz1BD9yBHWGl0f9bNQe3zAyM3Vu7PA7X3yl+TcE6wVOZ186NC06MSdpCbMEU3kBuqyCcAucJWDkx2Yvn45cghz1JTS2ILH9Dy7cFHZdYFOLkJ75KVZWL3AF7z0l/HqTDXUTThQEQcYPP+kJdFjTiUbKL4cLhuRo7E6t4lmGNm85QI2Erfo9bV5d0hlv0zeVgmzy/mYMzbHumxpJQGtDXIgYaM81KIfGJY/pxnxJCyxSH69d8OOm1kKCw6dPXYXrv6uitXse7q1NtCgNOEgBPmFuUHM2meM1GZgoqjg8tHuzdsYhgZ3xMmbdI5yFcuHqgtqgBtIs0UZLxd1s5CI/f8afNdC/ujpLG6owQubPTEUygrI7K8hEcHN9wsgRX75uIqnx09Yw+wXGwTONU3cNxsvh/KtAlKRpWeb4ifB9819PKx0hTe1jsZN3gVczf6BELGzyWd+M7gqxKjnaY3SzPULgwcTQykx4j+j9yguUR/3J42dA1Enxw6Ze66R7Uqi8J2Dkdy46grwiXVLv2hshX/1YaMlQQM3sltnZTZjThJ187XHj+zgMDXJCM7Kgxmy1iXqaaOJMFjCL4og3C+anASt3MamWgSbAZ8XXUMaWAyYzm7RZRBQRIux5sUgJJ0ldYT+xL7EC9wzkHrtkjTxPjrNRYGrvHdFe5Q+nk+CJ9gQN2SEqjrNpInWWdOgtHikdNN8cE8dDDScbexNCmPdMfATL2I6an9ZW7lU6mjEgK+9aBBJSRoow3DZnyQ7t45djH/7HsoGxXy9SfszUzxTbsbFo1g/cRTG7au3bZ9Hso9kNNKWi591SNH9zWqy8aritKYmbGaaaha7k3gG6f/wiEv+e/nFzqULa0aSfrQ9l8BMlKv06opCrkxGkfGdYSztsf6RkS/58BUr/nq/kNpoOsQ2xnBD7hoIXufFrGQbWIFHFqp+KI/JBIyTNr0xSX2V1dE4295ioO6xOnbR91spCdC/vZViUJWJPAfa3xhmNfynHiL6nZhpfY0zUmIJy9u3t+Ow66aBJeJ2LTeonAStmotHGzBh5RnGdF/1UACMpuC8YHvF60IATJbgwSpAHJ3Youtl9BqFDcwDMrxdosaR/UUTRd7igdX1TGWjlI+EWESRMHeAFlzPx0ofUCbfERHJJnyJSev0uf3dwA+QznV+wn32rqhqf3B1RKLnY88UPJxo0s4kTIgPsVMrQFqCKhvvbo0X1A7d6VOM2/AnzyaS1E9kYhjOr4RaeogGuVPrT7STxbeBlWExeLUuOUXJ6CpffXlm/RQ9zjDwQEy8PR/BacM4OHf2FNQ13WAvkrWHDXoSzIGrUomvkvLPpQhA7hYiCF1/ymsD7BpHdjGtl3EdhcBve+nTpWlWdpupRZ7b3c/4QjvOoGPmkRQECJ86orXLz3PKujVvJty8oJT9EezHWrdCqvRUjO4tT0QNqGTCBgmRphmXwki1q1NhcBI5SzdLIeCNewpOilZ8gRBYpO2dev/ffq7Z6tuNHLGeLi5i+8xBvFaop9AYPLIZij2bzxZsL6OKQKQRo38rgxMnwQeGGi8SjrCONfiom3UFpE7swY2NNh/sOU28MVVSwX9XSemDPt0aSGDSJrQVTBjATSTFBs1uai6EOk2WQciDRzmpbBLthGxU4AmD2XWyWtwh/l7JA9GoYBgv7Hw8Ukc4z+z+tUvTcGZDRmcaToAhYDqnm2Pxtnq4q70GwEYyxczTy9dp5gb9MwRvuP4A9LrqMLveBwKChasEyTgvBNPeKNgalAnQ3R4q4DGrTHTS6miv8uom4ks1sL9IggAxSRsz1Jqght3lJ72zQO6NHviWLmIjRp0IJcn03KrKQdGRQTwFfIsjUuWhOvHCr8/GBXz/CMPykYrb8pMFG7IsRK6FDmfX/mCBOogMnfGWRgv/shR15QUDujajNvia7AH3jAi6fmEKkrxUdp+UmKQYerFWPAYEHkutu5WYjp7gQxNphcSLjLGv8AjhJVf4qTmSXSEwiAVor5P3U1R3KbP38lsU4hGBTO+S2bJFLS9AYujxjpWKnkBg0c3pZNkM4Tt0G+OV39p6P6Jm/8q13dNyUS5Kwfo2zL0qjSeojzwyjK+96VdO/w85fVFDE68+ktaCETJEUPBsMWk8S3+DdyGTQE00zsluWLzeWJ6ILSUORA2bN4LQw8an78mRjrNGbkVroVQ8ZgiVkYrN9OLQMwaWHldMqyEqTVR9/C/LMtnAejatiIigqWUufnJmCPY6fhTPm6jv7cWSXFefuvWieLVAz8d1Z/67UZDc3cYtu5qSDOt26Px5+hNK2JsvLIZMUfHX0Zghg543xZ1rwX50Ge0ERB+gVNJrxHAZ515vuOEf1Am+bzxfTL9GJd/SaYpbYCzaOrTGOTxrC1HP9AwnUaOnI5WDYdMjmrJ3KpBXoRocs9IxluFgX+BexszlIRV5iJiHYqdold0cU+VU31b2RTE91yd6OuU2rOGYwrhilgdqJRYzOgUNau8AZMo5Ka5mBBl6yvg9JK0jicdMLj3cLsGrAPiFO2QgvIFwKu4Nw2cwv/DFLRL98IL3HU6bVBXUwEZjJolIz/QnfHem8g/N3VowG2Qaq2+oA8kIiebjTE0t4NxFw7CnYtVU/rVG1PUfY6WSV3KL2Z5D0B/n+lhLFEdBbx+X0SFTLEMmh+jo/PR8g7qFuK6ok+01LA1tVXih2R+oUKVw/ffYSPz51vz427vRT1YJSi0f1upxGr/JxqSt+jwkfjGviPIleEwQ+iFx6dp6vAqKHzevZsvEyVAqMsPKIJ57YPGGQIx4gQ4BZprFbZjhZkWWI30NuZsded2KazJb9tAGrZ7O+2gtOW6zOHOHAoIn/e75NWGqYih0KEXYmvKUE+y9tMJi9SST5m6xAXDFiWYv9SyaoiojbaUChWLPM2v4504+RNIW28glLlzTtshQ8OGRWeINpex4RvaxmhDUQdnzkNSD/qT8rJDAtssZv33u2mGHJTtzx20+OD3GUwLSAKXKBLVeL4GDOJgfX+iZuTp+4pMO9Yb7mFc/xqudehS3XPkhUBZz4+pKUIGC64MruUJk+DZU3IXbUpqWI9Pjfn3wOyIkCtzPJOGAebqh55bhVUKmSxtvwtRPq3X/92e+1/58d74qz1SS0YaLGXBQMik7asr2FQ8IItNxhk49tchLkuMkgk5JpLVQjA7vCF3LqO8mfBmomVvkYkH2iEnWSrSN24wnVyPR1+gzGZqDPvVSg6VxcIWthC0nHEfT7WgOcNVBAO92to4RcMyXjtAqtnw8KY3XE5jd5sMOiVN+W0k4rDbvjkDSiO0Tj5UdOJH9HLV8uT1KdlAXI+J7QYxUq+DKFZldRBd//VyCA3okTxIg6OqE6xMUNY7Il6pAKguL/EXHR3DAMMaKC/cH4qyIhhUirc4/P5IcfHETwd3J7et/FCv0pwyNtd3MZMN5elxMM3rV0nh8erXsJeTcvSYQO7qsAFGn3L6dHXfNwkhlcYEmkpjN81rAjxLYSBY2jxJsvnWJD3QYlFtrMsSNOC9yEL8vt9aFlTSA1BfjsIWemmE+4EzNqdxW8bltHS4d0kyWCWH404vm1Ee5nj6Eccz8Av9zzNZWa8ihFor7MLWdX7tFo28r/Hv9tlNVjmM4439oFqX0bS0f+xYXga+HzNSrypM5Jw7qatLtrU5bIxm5DQHfMjfbIHuI9RTSgz2E34bnyVM1aLSIcJGNOqs5q4dkoJUSrO9HUri5qDWgl7Q0R+PWngm4J+tKb4WfCj6U/wxIdazWhZmf+IXV6UXqWRRBP56HMxfswaRwPXgsLD5det2WBGHceAceplRS6jP+XAYLqL++R+QXOncZRtDDEZiE1SWw150rUIcYHEJ0EGUHqnwO4seV99pqdaa4eNAAsitWHGaSR2zScWG1+LjByBvxowyfh1UOrkMNQPyKKTNiCqKspi6GgpomJOHLjrG+4SbC8PB0XHO4atzyX2jJ1Zrae3Q35T7rdepGyfT/rA8dHFMYWjTNWcRB1ohPdgxFmiiZdGvZ56nbMrYpoBzXt3JVI7VQcGeh368a7EjVSVH68XnAw1xFqzmGwDGfmsXKPhWeZpvLbXq8/nZOVl8NkGAMHVzLixWhFrnHQoII4/idUcODFH8Hl3MuLQyx7TAAPVzL7WUP4unwphnYt4jxYARxM96Eug2ko8Md+irBtlfABAp/d0BAOBPwTnfyF87tPXrYgS2q0nAOVuIxIsyvWJDx0nWBuORwEatzeM3c8bzH9AiRP5gpwZyeL803FYMfZlHGgkyjcf5qOJol96eGQXbbhpWpgiODnpI0TqzAcz2QEw6NAqhnTDzeEniDo6FO0fPX5F6qSTo5dQaYAX82Q8tXE6HckNwg8lij6ysoPbOeijMUnTpP2qG56dQEuTgsTIYQYP8FhV+Gv/067g68OW8ILRqqbPnKDfXNglqF84A5+pKVMZnTirRUbMehspiOI0+8s4QB0sZks0/coyA5c3hYE0HnPvmvEk++zXLd8pPRY4O5dsZbGFw6Y2RE6t7pZpdDoGRz9QBPqUXhy5WMi1nUp3cYOgQA589aKjIU9bbFG2SRO80mN7tVzbsE201/cwWHNu8taP17dO8p4JCMrrQ1he8bSFIBgVvmOkCyGJAiIwahwu/ZN6jyiXQU+NJ3vKF8KaLHNabV4WuCvTEcwwhIWHSY0SUZI3mIGGJepWMrOtsc5pau3ry85lZ2NUghnRSjjSLpx+f06kOSUWEM18CsS5TJnwKuLEWFb9jHP1xj+PAhPisMZyP9F6d6zUUkfQ7VWZ52sgVRJFtt6IdpD0PgGWm6eKWZO0Bdru1UBaUjX0Iwb6RJE2CE8UCIYm5js/ZkEKY5BUCwR7gD1vVy7ds3bxJjNVkBcMBdbUVs0ZRmt8/ImKzg/NN7x0q/3Ts4e9JQ+8qJHuB0YGmMsTM+WL9g7L2SjpcBzBBZ8m5U5rmOr2/WU+DispMJghZHQO9mrplYeN0fNhHCAJZ/KjPeHPLRhr7xbDRSgbI7keHFEVDw9ETO9d/9PqopHtLi6eJfz9LgQyBEDB7O1udX+Fqj6BLwj5mWTWCV07568hsxAEk7ZPsFYCZkDzMtArlmdugWBspM/0zotqtTSs3av07voM7rO1AICz1ySksAS+It5WbQyXJxZ57UiOCfFWJvtESeAg6C+0Q1E+9pk27oGNBaVPeg3xCU/xfvwR0y/E9mrDDMWvgi69LPx9JQCAKGJZWlRlGvy1ef9HECTsrg5+Ej/qIWkXQN7PwwUkdJ/YBAq/Qkpoz6DubxBax29mhKgG6S95743RLm4DJWMyIfEQ5e6awkVlh1MxsJbKZgSEc+ZMe1+QKWwvtAy6mMDKoy8zitucIdod7OwuYEKPWeIrGn7ywlZaiSsCLZHOb+lT3oDoTPnM38fIR5YHeNEn2Q3wda3d8jI03NyV2VW+C7giBDPPcqYedF0VzL7qp6I4ZpIMmej1WyXpv/nMBvRIrsIKciHWSNseYnDWDDzJdAvNrk/a5j7EFFmO9J+WpB9gPooSasn6sVtoOaGlG63RRRcxiZSPq0x3mT2huMXca7UajyTNj90GOD1DNFOGtB78YUJNdjZTWbzqnNjeE3MkkFEbGQc6NX5RGbekr3qEvkCdXEMGyzWeVtbK5mYzCdbrOdwl+NYtkWTEu2ME825FUHnW+rrXYVB0VaE/iUNvTPv6+LbOYjq15jgaxveeVBJYb6eXFmvyiyzLmuyjp9YxtgwLN2B0AzGmnwl+4c5U5fpwawUzC+u128dyQagQMvyD6CVD7REjbxyWymj2SW8r0lJO2ef4hLO24dIvtA3/ckGtXtY03HARiZdRAkRFS6c+o6uOOQHumdCQLzAZt6sHMU0WQ4wZTxfW7+VRB5cU9HX2fjQ6p8j/u6iT/6WstzHha6lZGaMLBQMEpCI+BtV1dN2SuCtaCnInohGQ9GmmpuMg6892ygixR79UVC/HLIgd3NuIZajgr5Iu6RQAenc0gupgH6IQeGMLO/7SB+E/smq7VZcznPuD2aNhKT++dkaybHgBX+pyoQE4P1lCIG6abKTj3HIs74K69f+0oEIlrk3vi1fdmysfl4DF2X+3zTSzhohsOnJinuok/wuvAVzxnGWBuXiCcD80G4T7u0ZKfSLQMM4h378UtuOJL96QaCGAPr725L8CkiYHPaJV7RchrxyVdUYuAxcyxEB5KTcchZxcC77oo/Zt+vQRUOq/ALWzGd2kn8O9GtrdyscfboYbBKeWhb/kSdKp7QCFqV9oVSySRsrNGKQ94m4JJVDXX7pCHJZN5H/jnS/6YaAdtGdwTofEHSWYkcOWAcfMdBr4HgJz31qlsH/8GIN8n5khVggtpUHXBWjVzuKuQvrCJjB4PSGAvuRbVTENRJg3fQq46jaqrDwyjaqeNcg/sX6Wm24m8jzVXLw9LEdhHDMEI7tHSfmbqT8O3fauli6XusoF+X9RZWjuQYHCMb3IlWofDRQUanxPqGhbpusPKKy7DcoHH78qY5xQaAk4x55dA2Mrh8qCl5v5TOsbwGJGowoFlykq6oVQXtgqL2lhwCM/3KL4le++0+2EWwz6cgYU79NaZAsFCQc9NjYLMJvZluLZYaQE+lZrWXLgeNt0THXwW3rucxMF2RqsFI1gAj3Z+3C6lCaeZ8N+aIeT3ic7wwOuDxOqppGIyPanTolOVYPe2FmPYo58WVcIjeRuPn9HCXcJOpeDSKcyEJQy8ARnDyUCpsMoWSqrmRWzrbx41WYa94hnnDg9ZTTG6mxwCNMweJX/oayjWqbzfaLnPpHMQxC5qUodGrBZEOF8fC2yGBUqHuxLZTX6Lq9G+0NrkWwxEv73X/uJSY+D/v+jbeb0WxrgOTCVNkznSoEH9K41sVkkdrM4GffDWZ1aWYhFOuRbSJsMeXAkSWvSikTemMzK6lI2WoLtzSvLuADiB4joJz5n8wxMWTTApvTScFfMVUoga66Qh5wa5/JacosLxdqZzbgIVAoG8o2SNDE9HpgBPcaPRurrAjJE/XelcFZvMNZ/ee+KQ/bg7DAESDV+tlmh18EcLJRbT6MjEUUQGHayBZbuJ1KYUZErHiZMxDx5U3Va3gbS3ZZxaoEnX8PBEE7kXOGlNWfVNFr0ILMmRPJjboNGn052ze/VgRFLfflEH9u95wTRYqK7eAVVgkGIbk3sZkkCMq3xTTPXAiYdNPJz75sWePzf412qwsZOjirwJhxwhXK9ozpL8ZynePVv/uyN6/SAY4amUYHEJyM+sD9+CDvL/uvPwCVhitmKnlQhGrmfzDMetc2A37V78cYmh/vEF87lliZ4a45g1zbl/2SyudK1z/KziHKP3Pi6kPqUo9HDnoL/eBlx57dg6OZp0lTg1VkJHhk24azgW5ueSvvcHCquFF1/1xW6fO7BQdxl/D1drfrIvfZDbANAwJZvhaOCsJ8282h18thwCl9E0uZ5g3HNhZX7lrBUFivgEgkTakJV2nPh0z8wxA3tImydjS8J9zkBYRuxN/DIszBSxPJLQE+ZHSUhw0RRzfgzCy8zfbWdjHrkM+tTTnMDA9OQAE5Ec+3w/2GJm1nnr+bRkfHLaGgqwY3zU/5Ea0R8LgMagZK9eGxfyrilYT1c6Hk5ADJuWS/913eLNkFcETORKOGho5492LD2nlob+58IMBuAUcCxTAC6iuEWmlYkrJlTB+xh73V33ZMljDWf/80g1a/kHXcxFwCLbjtfYm8+ForQaCU59w1xcCkaeNLQ9KM+bpUtU+oNSL5L42rbqqQU1ozf3qzfdBcre2pxvBXcsvht+GmFuAG53z5EEv4hW8JGdO96OFb2MSF4593uh71V61XlhgxWL2lI0IyiYdu3zNjRxOqyVxsK1G0L4e7WrNHW0d5EBdqxs73t0OUxVkfFfek8ToegVFH1ZN7HKX1FF2PKbHoS98kqz+KQ//72bKQlyEUI78DYvDWSPgYpZz1EopaElInpnugKXWHJTf+B5LRGbQw92EImguckfIpEs25db3rb2pEWR1e9rSKaKAso8dn5R/L7n+a0hfVkZlnEN8LNajVHe1zvnLyvA9T/m1RkrdFbzdhQLjfM3chFwHRu4+DwWq2G5nLPci8UBj4V+KcasATLNuDQkv03FCHh9TBJ0nHrike0b4387K614g3+q9fpvsyL/H9QRhslm3S5kzz9rAwvA7VWE8p9rfoH43S+YBVascGoPqkXg9gkK3mhYRD/t30cObm7BhBJVMwqmt8XhgPcQQV6AfL2lN4OdszDyxq0T5AaaEkryPgsmX4skIqR8H80Am7AEaqPznD99oja5E8z43NkCOnYiU6yB8m/Vka6jQ6bbZ+Ikke8BhG4X2kaYsnH9A/yUWbANE+JwCSQe9yvfHoid9YoxZNx3o1mp8pazcYuvgw1gYKdTaj7TdjMCvCu1VAaUH/DaN7HbMlOUZHVkriqjoB2vNWH8OBrAP2e37yQzeRy19GjSgZBrNpe2cv3z4Qow99mCGnvbdo+W852u43rHc4vl0aCP8xUnq4n7SAwf+zu/lRG9joX/qK2nhVcTb0EdJoWVMOwC42Yy8OAaR4HirRBf2Mr4yz9e8Ch/UPLBqgBvzJc3dgmQMQQ3hRODdQ3X7aocKJOpFZXCUQRy+sqqtnEBdZOTmW3s6PFasLlr5UOt/U4Zm7SiEH/CHGXvrpdGlLOHpFPf6TOUjciGoHntUtYLLXoAqAitqAQqOh1TuCScrAHu+09huThx8jq+hXgZxoxfKda0QIF+ks0wVVH8TUmGOSJW25ceNTIr4yJFQ6uS6XfaOzyPYKNqtHeXuksXzGtgUUkbk0kF5bbvu72g2NJjLzEOVT/qTLg922tHYRtl0w7ePd+3AF4ybqz93CDaSftmpu2SL/bw9eUo6GRwYegF/ao/JvT0/NK6Uj/IIfKrhD7N1QtUfkQEJrJhuwKiYMxFmmuCvfOsObq3HiI/OhbSg0Q92tZiIKfgSu1dGIb/Auj5ao7Xwg+YvGZwH9ArZmcnyTgWIxlw4ox7cfRG8m8527rDow3LQGJ0K4peLkxBFmBCf8Rj1IVjzotgA+AsTdze0gRzMvPW/qISZd1fc8YeCBJItXbLs9azWngKOR+kwCb8PIfnHchOsMsLyMu/XQA9EnpTvdebifqBCk623kt43fCqYUfIGmyXOPQDhCAotHYb0gzA5S/vyEIpMmScJwIlGHx15LWJ9CfqzoLpMpg7+03CK+IiieOo/Np5RL2kbeYuwZP42ZbOBY3TDBbhzpxnPPdmPTT1jSZb4w7Cj0p85KkL6vrufdkzHjSznaTk61/Fe+WukIxU5Tpqnhj9RbB5srZGYQQNmC1jrrTpZyubwMQdG/SQCsmsYKRaeIMhI6TS6z5aS/xZaDCHeY+diQrspO6m9Eq1NItp0mzvmYh2ZWit1C6edI0IH1lab3l06ASWh1wXm6BSBaAqkP3PBeh5Ig+yoffW+s1J9LCBsBiaZwdMX8/PBFqtJnLR13IZWNBeyjRE+Mn6wHf8jrcW6lNwv804wo2hzLddgATcTtEnK1djC6c+py9wiT5pRFqf46Qg7VgkZByuLn5U4CHDmbv0ywl5RuAAdH/O2l+3Lt+5TWj+jJkA4nSirdQM+XyDbpMvGsEifTUC02aHhEbKx/HbQUwLlnuLyciIa8e382tObXjMRNeeJYnGpAHNNGkg3Eratra8/yCCFfyrij25RJ7bheRDj2w6oLSlf4LKndoRt+fVoYbMRcsmolhioVxyy+i70lEPvIJK1jB3zk8BJbWQJSYfWYrSbepUbbxApBKg7MSz27hZ1eBr5+1YNs8UwPWvchrMkhmZ41UujbXPQuldp3eFJMRd9PceLIXjEb+El9BC2qvltZ2QEpJ6elnottS0hgdln97BcZwUTDDURkRC0HYJDx3JpS0ritOu33z3vddMKChmhXt78gaGP1efbqqxl1anp32zX6U3a9Ndulusqrs7pR0z3Z3ipkLqCin/koK1Ga6FWjag4DPEVMbOLYBWUGIdmsPSlTeLIM/CVhtf4iFJOcJA/+LzNLPHgCHNCY9/L5u8I+D3q1V4Xvoj0ImwpbE6DIpUzQ9gHYotiTM1lFhQJ3HSprmTjf/ekbfktHjg91tHP87bGz847Ie8PcaUl9T9H4QUtdo16MU8oNOZpF6hCHoGYODj2GmIdL7iXoNSXzEKqSCoICGqpDqp5xHiSju4u4nTAJqAUrxkQyQ7jBypM3CeWB6HwGWIGVnUxm6jEKNcyfA/o23HpgaFdX6f2ZsKRP6kIbhLJPr1UD5NiW/u0qZAQTKbGpEwA9dzNNNDLCwEInjfvJxm63ba4rZWCy78XVQAs1UD86SJRfComiZBVTl2AGjUC/GMYuo+3NAY5dm9u/OmkWNKgDmakVipr7S7SPvgnvDGpIlocG1W1AIyycOIUmkYfmp8LfJYQ8NnSM8hlycqYWM6PEuTa3a973HV5clSPw1KUSbX7qO0cCqAfTSgFgJ75K3M1VNUL38XQt1V3erwKtNT4wmlX6uYAZDpTtWHFDU9ZQ+U2n1XJKXWsr8Oc1Xrxi5mtbeVy59vVox3NMxb7ZpCEHbTWaz22m2/t/BgsbRG5ysBXYX700PM9oHg5wef03XocaehKHMZw03qFkNatbrIdrlPhDvLdSE7RgS3+L9V0bmtW8zs7SPsWTtz1pi/5qc80LE4btWuxrZgjs3JJ5HfAOGT+lPJ9r+azE7X8w+12BOyDFQaEn14IMGUPXJtUWVjQf1+vn6muzvBi0jOzoIXdxYiBed3et52lDbmInD7niAjgCnGMx7KfwAoJK8qXvJC58HgvsQE7BN9dDSucK4Ev3dkhdUjp6Goh11MEbG0tRgZ7jGFqeyRE7g1PVjNeo2A/vEKglBlO1gPUBffQXVZD6DLKn/enN7vY28L+CpoNzIOmwn2/sfDDtH2Tjf3szido9MC9pFpRlr6exJoDGLV/2zpFElYy2f/LQ9WsYB76Rc18cMmc9A8fGN78zHzhATrWeFVwL9co+p8AsqWXJShm+WZ1zGA9LCNVKebSc2sFCahASQQyGjoqDlEIft2oWw3pwVtErNfiA9UiHaQpIx5zmtrJZE/xrvkhulRBc93xPXGU4CGc+8goO3SbOrU5UjbS6PGeMiU+aY9Nas60BRXyEvwhvuPnbB9+7S1OPPOHCaV5f3HiZaC+YTb7eQB1cIKtUGvWFdQxlEzups0lq8kg/QWf68ptt0IgVjwhtbITN95C0wC30Cc5NrYTOqkZEVkt/znxM4O5dJZ+jSFr8JGvlFLYbGjrjwYWFwNzjLVnweTa5+OkPY9SxlzBHcROyY/khaN3bZ8T6YBp88iec79dWdAocdkpDeN0JxtAJkq33vB0X8A2QEq5JGMNK8f+4EM5v3iOgQTkDwGRMTOqs6ylRE5u5xOWHF17sb1p9EwtlgOFwqnQfAh1Bao6QY5JqFqWPBv12VeSBco7NslEkBwHdomU5cGQTjGH3CFmVsuE8zj0zWIzqVLe5mozLdTIYphrTIhuJJE7Mgt60IhlGuh3f6H08mQ7WZc9t3SxUXL+kK0tKImX/SMq3kAp6UmE3B66pwoXc/v68xmaBKAn6pT1+mttRsr/B3k3dT/eYyW7y75ZE3A/BEalBAc5b9t99z/6eiS/b9DVrhyW8A0SedIhclxB2XOuuBMaMEy2v5da4L8iL16TpQFxEDqpAyN+HHhKyby6nCqQWPAc7eX0TXqLjY1OALBT7wA3V3EjK9eikdNeVnWr9b0urvv5LBOXxG/63VWOKZ6F0qdmRx+UG7ubliQUKQOZiDwkm028k0Au2b3kDaTp1xvQnaVTUueUSNmS6BT4eD8CAjGVxFy71nZhnzKubGBEPC6nl2oy3MpnZsZF1lGnX/q2BNbarkNeTAn2izuOFm3TiuprD+BQ/g38oMA7oNYxBAwXo3Pw4rjzxn0NRkDmFUxltoC4+zJk6z56bVKVV8ra0zV3LUcKXQYVy7ZAo5L+ltmFwBczX7RTQZIaYnidWwhkLhGP3IY/3XzwZQ8/lhFz60oCEnYObbnTitjCgd4vSJVOfBwTAx3pusjD4nk75197XNmKbIEsT1aj2XjBVzDdtItD6hU9FFIN4Ky7aQT9f3DCLBQ+Zn6ehGCEiryDWBk9FxIUdXfYSZGQjbywNafsOTgtUfT6HCrJq+x+UBOnU9MKxFHu1XJML1MmJoSlX9+toOjrBMqGhDy43iHa5qGJ7I8ieGXFh6UR31+gUOS+KucO0s2q5m+z5MTpNldmCFrd4fog7uQyg2SLvqXwq8vZHBx9qLLXBJtzFawB/pwcyVuWKeWJ8lhC6/imvuX4FjKo4SjTObDbhM0EP0UprLJZ2y/NSaa+d5xwiAKI0SEIQftzvMHBEFyzLg7zLW0P9FfmZoIbRBPuih+2nRdNPcwY3tobrcC8e0lF9oOiW37hSpx4TO/pXYkL7aGxXWHqJaE3/yLh5N+20YdAgm+uIrtW4ENX88so1NkSLXMmoq++Tujp7YaX8XxhK2rwj3uXXpKlV4RkxN8ErevtMV8hEW6Yvbp0umyt9uLuI+wQOuFWgwR9ESDKR0TXT57pjKkeujuOaQoHCR6pO7QGYrmYZWHKYHJGT+ygQPk8gaCuInNWOHHqMby4WAb6tSx23IhOMt5diugrpZb7SFGWwLjH0x5TQ0XntspgoYKdFeg4wAXdL4B6hX7nxoY/bVoRqfdsFdT7aWlQBfT8vhHzbWDEokoGwYLYIghVAVXKgmTm+c67kj7bv4/gk+zN/mL24C42Vr60O2Hsq5kokt2jaxApBaDwTn0YCg0JONLzgsFeiongSgtG+oCPbhmz9mF13A08I3GOEcFQPyBTlyDzuT9F+aY8tQEjl2KkvTE4YcvjLuXjfcfkCF1nkhAf1W6QXBOyAh8K+DS0OxJoaD8l4PdCz88ZMCxtZe+sgWCDWZCaUmBsjl3fkan3Uh/+KEbfEJ+Jcc5EAefFrBymjLOSq892FQ/+Cjw73OieDfS8CN5j4r0ihKwDT4gii9xwRM3r0PtRLWsKeJYGAlT72Och4cVn9P3x1C8m43H+7UcrC90TqODGnJ+wvwifPH4fjbZAtjZ7PyZun1RODcdByFFRh8uTlGESibLzK2RQudsELMux5l8Gw/ilXFrUlXeFjcRkPAXPLRA4XRxsKHgYGJKU11f8mtk8PkfgGPqJNw5hfTm9Bo5ZyR/qW1Z+ArNK24VVY5deW7+ra1SjZn5ibJ/D3S1PUZ8tNA2bLKsabWgoZC5IzVsCALYS4MQDxP9i5T1wBj8GtUWRNWwNYs/mNL+bjZi4rieh4u73e34mtuGmrp1MhSwNDlW1I2jEW+3THbzWBAqpAiW/HGap8UvtK6YsfHcbS9KxFtwhvSF95ggnKU03eiOqUvPIQl+Hsr4ELcnfN1YtYYxnwIZFkQDoS6uTm+G7rgNEBKXNAYes06McgJ4XxUA6wUNOcoYdAtm3GKVKXdBDOHPhf4YKc/30dwvd6LJhuajlhqXUceqn6qQeahe0dCYdh39SxehvS5RPjrKT8fKhgXJ98gYSDWnFajLHeF6CeOsbu0FNs8JkfxQHBtvQ499SCyOqRsMzQLY6ncZ3KY29D4sl3gmLEIjrfMn/XdCd+Yhyn3HVCSvVw8L8xvd8+QVwP7CZIp+bkgfEJPUNO5dDsEFqP8x6RGgFUqFpDLyeXm1mMFqb14kTMkXWjSsf0PtSS8jHMSCo8wJb/Di+AvRn3W+g4G7rgIqBI/Q0nckL1cd4VwTMzMBu6s1EiAOz1akYycKusF+5MSfo3psLoZRIECZ7yaBWAZjFfmWkF0NP2gasEcRnkAM9lPsfcw4KfGyNgkxO/A4cmJ3Gbv8de9H9qDY2QCP11I53MXs+sW65s2UVr2rbna1DeJfzvZ3wAPMecm/+mjL/22NjUhCDmHPuIqjU6BPX7UNwV0BPIk5rIo+zQnQFKaP55nUTPympVuYEO3ZEavxUCJJJQZtUNw0j71Kv61ySzzgkSfWD2TLR7cm3AbHdywIe0t/sAuiP0IQMyVb06xFtHO6d1th1vLqTuk5t8K/Y3C4tipm1Ge+g+E5JvE7BByqOKYNTJvtq2jsd5ZN2NpdCdgHHWycS1LoZDdLUgd6YMBcWMb997ay+GKlPzhPkL0PqQ7lk+jTOPided5MaNnIzzKGLMBLPx7yQ+lZEd7ipWbXSgqMmgm58TSoOS0KuiSpMMkGTGsusICLQhiV1CHY2dte7JeTAZlFabj0rDGUWzQd7qSn8tG1DHNihHt3Fj8f5QquO7qnkA+XPJHOGWVRnJkj4QZZttmEiqx0EQQPbw0Qk2nvOZDrzm6djjIpdegz9WHwVRu7/fRdSNzVsM82X0mICTP2WaaPEgew6ocWjFSs4quqoN+uwhJA5qXx+00N8w2qv/cFL/2g3ixyhyiVasWR6uYXD93rkv6R4320JOJ40WRyLAmXgDfozLuvRG9S9QGgTfg5bwu/HuRYL3t5FEE/PmeLgn0aTaGPE3+V118M37oiNjh2pfo1CWbH20V7DqTtIkJXnCbhl7oeVqMVOtSjsd4EaFecxgvAGsQ2CtWIIA1ApJbP+a5NQftQrBsFrFTRMXy6JXXFhdkvg2Cm2bjE7ixfyygf8OvDpxxOHS81K3d+PnR+5keKgLGY1DpdktRQIu68Qb7q1KmwhtFLAbhtwJsZdsWrTgc5uepFOAgpLHLs2XBAXYs+4iQ/5CB4+YQw0KSTGaQANChjZkkxRUHnwUl5q2n3Il3STXdLCa3GNh2hhSUt3vy4jHpfOW7UVFemOyXiCatKp7/56zpBxy9wrRntcrn1pzdntde6FMq/gzCG+Y5v/iANNzkkF+uB6AI9oNTPGmU6qrLD2237qKCmh3MD+TmKUrbTKXzRDKy5e1zF30012nhm7J8mdSsAus0P348wYEtegsHZ5G6/ENtv7X2UDNDWBh5T0Y3QTti4KCasb0hVJdeLgelEA2iMaUSzdhaNKl5EtJ3m9Tj9/YZFNaV9W5RR9tCfPqLwGyhbt/ClqJRq4UcsWo2zay0qy6NZCkogBj3Gx5r1XJQsz9R+oHec0g7PLS5W3Yvi/5Hq200gygAPhXDpr9x/ADzhs98Mmgrni15NUT3I3Z+S66HExiwCsIGGZ5jTTGDzh0tUZZiChNCfJVUfndZFdkpj1/GYJ5Elr0t1/W+iymPNiERWbYPBl7YgC+9Ptb3tmGzZ+q4/1ARw3Hxy6Em6S1sHWpym16iie/PgUkkF3tR1xbyVvMq+n2xsEKNYNvBC+UCkg/LozJyoW4SHqhEclrLvEFoImq8vxW1ibkpH9sRc2SPYOW+WS3bH6bUYQD2Xck2Fz7Da9F+8XLlcTp01JhoQ/WULDQoK+T3wJ8nkr1pPtidXBMXeh2CZ6Cui0hGVUMEFLtE0GCRKJUBlsg455bGhyETzgK17ZKUh9sCfb1E7lN9s6nAt2osoW2ONY7XeLcHRgWHueaqigm/A+vrCge3wcIFrxyMTEptvu9XaIOwcz9MGg7xnBx2LrhYjWhjY2Ma728huowOmiu3lTugZXTNWMhJiL6j/DW6TngV6qC4yWW+vYMUEUWIbV+uyrlpAiUXfBEs1ix831D3dhktlq6QyTuq0Ov9g1NvmcHldNwgBgNw3nxAZg5BbdRs/bOdFJ2FUckHgqCzpnyFgzS7b+3vpwohcyqQcnW7xvIGQA2t2yGcHA4ihieyyxtUt2106kkAfAsclHyiTBe22nwuywmfpiG/sjNxI9acnTgcrP8LFVBuqoDluNACbrMG2LKFrfsZZt8fLWtxuDD3mhP798T/9KOqGvRftfqJGIPeAEHBOfF+YCGcoTr0p6JhpVFJeFBqIGu7ACXMkP6fILZxEfYG9oWSzxYlgtkjp/4tQFkwhyRWFuB6/Zlea6HcDQ2JB4ZCzNLveibYT46hU9K+pPU+g2CNDW9W7TtnTh5xrIbIJwecdDKpJqibxPp8H71bR6q5uPeWszlTzAknEhk5Cg+rsunVnuw119Mj0CCC0JOR8wfePrd5wgimyQ4rbKpmOehdwN8e5A/xwE6BzTxrBIBkM0UNkN7CZhovVY8mbBgj0S6bXWpHItMAjYRMiQsZ7tSwAaxe5W+xF/Uj+auZ8IRpVPinrgS/diWuRXsVx4/LEnBFyqMbhOsNxJGYtKBMz15kSi5ojArnSj+MY6ss65PBHaGzozpPlUVmOXfPPdSGbRU8O+0JGptI4l021JoJpDtVUYiESlI15ZDNTCTGVB36j+BYU2TY5sOemk4uc/32R4zU803A02QMY93W3j23oIGwDpSxWOYsYKD3yuuRxoINU1v/5/nuYENTOr6DnjZWQOCqCCmM67QHF7t46do/md/Ms4TgnIYSOtvNi9pY7atyyzb6i5qWQtZ75dQhuJ37zYHGkIvfGZVzzYCj3gKkOAUUjvBZ8B7pguEZlx+4GO3smn8QgHazROvmSX03dDWN0FBO6p5EOa/BFrfbWVEL5I2xvZKASu6HK0KVAQ+aBhRbgrH9cVwj3omr2JGmBTqw5PxKfIzuhI5+AzWOKLlB94IdRQZjtjLRYREMIVuRUiCiwJnmv2n5KK5oAatT4n3YLYU79cjIXkhS6BUagpDhuO1eK7czs8stqChBbqikWtrb8/3AN6d7Bk7DBHtzCdEnR9CmJUkMJy3JPnuyx81sfbtc5PGknH8OYmjg9SmEv3RTDMBJMuNVUUNWFAfmQFmA9k1Fu7sfIPLm+oV9vsloWL+yZ+5RVtbwPVt5I2L0qvYuiN48hR5c4kP+wTlQRSTFqXXuEAWWKuXV9kOdBplV1v5mg8w7XfPqZ4865i4ZYIhrUgSEieptaDgGAH4wlUteccBk1RosZ1mn1/3JQptMsd61jiESpTsCm9A8UHOIBjZsJKKqAYMET0kk2vektADgd0Tvo5M5AZW2WB+G5/Z7+4gVncFXA2xyGQ3gAigFHogucFcUMj6PnNU67RvYWH3r5c0wzE9J6QwiZS1Sh7yMGuxxhyofzsNF1rZ2NJRU73x/dWzwSaj6u250jfWwibXeq7D5fXe30iJmdIC3n5y70ORBCIWJki4+vmfkhJko0FXyHmqZnM9C/cT7jrMoUVqRIQiS+8nSgAAR0WqtG7uOEm1sbkWpooSShE7ivapj0G9umYnLnjtvYYNKuYf7Sw4BAXrGBjKAW+hGCjq8kieHM/h0IIyrlBjGavZ4u20H/KIiJBiEBtkMSvnUX8ivlPEbyw7boOLsVK+igd4+6P5kPQP/SBPkHsEJytuqQL6esZCvY3RsMVTvlFvjZ4SN1Vvl+gOqRdUbGahR4n5VbAaty8W2XxWB/1mOmGk5aCcg+gP935KfLT9DrQOC1rUl9nfO1UF82muj41y8+rw6A04rVej1hBMCdUPFzVbLM2A35/l58ee5ytbU4Qp+UpiqBRPTdymAjg3JwITCaJm7MNlkQQrlQHujsZHrcyg6tYVm5jeXuEGSJLCgCR21LuK5LQl84asmJiyI9bKeNC2yx4M+yIPn2bYdTSePNRlcp4+XASgS9KO3ZEEAveqUZlkMABEpuDbwOrkbNOkFuiEHIOKXv31hxnSP7I/eFl69NpEHoA/PZRD+DuuPg+feKzXQzrm7QvaFtR5ApV2Wje7p8+uRvV5ZQvg3orT2wXVSech4DOKSB2xETS6sqpF2B2BidP3vs80090kLS9yYIB+2MSewHuCyUy++XXSK0JFUzA5OjBcyw2TVtMrgenC6uunicKbWKneP8GNjk6xRm26kzLtGbkmkd7S7nm99INqUODOBox8hBoY6TEAGByJR/yuPNWfzdbz8lIf0ZCeXGU5JPsV7EXf3CfW2Grh8p4DbHSiqA6zWTVtW/yYUFLren8eMka0Xy8MMEzLzDoboi2Mh5mzUd8299wFDDGyJNGELbdKOChcxZuelmCYvF6/CsDwft0MyDBpqWBAjeE0tOw3ZgQzl/fBF+US+VBPM1U1SNOOH8jvDdnEU1cuvqbypiFLjLZHGqlKYPZzUTntQAqT6vlinFIONjan7Xq7myrMj0hZC5wQOZIq3ta4Yw/ItjhFNYTWNGYwP0qx7Hcr068OzG04lRD6hkWgtwMxH43UzNqrF4/o4H6ayx/uJNpgJBd9PKZl1dBcfiEMkmO/CJ9nMHBswhdeLBaCLr74m90D9l15LvR6JSdrh3BxvxWylPlwAsAcWzCyt4RJwm/M5vTrXTWlIZtVoL0y++fZQQevggQKeDycLYUCNH9rUiFiJF5nTZRk+Tzn5orsBYcS+S5/bCntyDrypG9AezKuo1BDFjnPQJwYMwVyE3TJ2VShzM/oMarP0Wn+gaomBQ4AAZ1n3PKk1xyJ5yns/8pJJpINUUyE3qeURurG5ISe39ex/I0ZBb+EKg6CgemGPKyH/IXfXUlwof2UvayVoSicYRscF6MbAUqdRzs6qY2zQhT/HyMz7tvc2cCUcrua5vCrHe1lVAvhuPgQWkTp1LEwPPhvdTpaP9PyU3ybgzxCXWXkH+HTN0il2Oyvo8sI/UNJb8wKx6y9i1NBby2ZYovFZN8XGF2KQZiCK4tBivMW7054SrkkxBf3M8VXUlNRrJWt60SqS7ssOsfGmJEtI1WKDwauGySnhlvZI7IKT0mBzNOjGzoh8S7l3jfP5eQPrdTflDL3s17HuWp1nOxe1mzmg09Wud+8G1+HEz2BPIIACeGy9dB+ZbOgllatgGIQMRoDnY60JCaW931hEjnrGCGZPXzAcoXWH9TKiL/Q8TNsd0yhRDgbRb4mKltjSX5wTmnc4rgD/TcvQ9hXnyDZfQp9kP4zzzOBHfDYTnLYcv3yOAHLK+BxFg7F4QxxsTyYWyTXNia0JbgPvaDOoILSheltzsAFaEBqQlnPn88/4YoGlDMYceV/Yv+lgIT+dG0aqlXpBPCt/Ox2XDpFLQ5K0gfF2PE5YVCmJchyOgMwnp3aaSzPIzPMS3/0aUzEUG1HPP0HHlTj7aXyajRlYT8Wf/a/5smWVG9RROBEDbRavFzRYSyxx2cKjuJK/mGedSc5z62Kqdb6cvvjEOI26n3kzHA8DyTrJN4ge2txOc3ORbBT5Sfp6X94MrqA7lZmSmqTbasxNqTmnV/1VLNPXGbn20kbGgpSUjQO+GEmIaKvjGT5WqSeAOoLZLlnT+YjnZkGpYdzWtD59d4nOdsNYj3/jRmSTqoH9za8rIiydFBPKTgCXRm/x/cObPrzt9hiRCGPoEJPz8tZPnsEUpnB3RGA/DmrZ94FWFYzpNlPuRVKTyPdYh8VTDBcQ5XApoZYveh+C6357857wN92ertE4Bzi4hVJ3W3PTfyfwPy/yID+lffwr38aG5l+TmCmi1xWAqJvJuHVa75DlyyyO+hDCw8X80XcazZjfKk+yFX1uElTklBJEmjU7rBaphG3sftYY7cWDXC/93v7HFLAzf4tFf2nwYn8AEgZDcipranWjPOQkl9XLcCOczi4c/rn4WgiOhB+KLBZM+vhQQ6ymV/Rv5VP2r51Z7zVU1Mru30IQjszsWgI6HfKBitsObbyR/+az4U5zQmm073OL0JslYg3yYhATJnij9YqjGMApYg/eZWGp5NGXcL4iuECQ0q1kiaeqvYlqg5L1oBJfsmydSOjrUR4RkzMbfbALzXjH7UBir4wjmVkz3aPUzpkZeDt2Dtfkk/TL5pJ/Kk/LM0ruDcubQpQDiXPr/D52PP7yXDxqSXBgaCYxCu23mPy65YUyPTNCbX5HfJziWpq1qyYS3Ttqu70+Eqc2i72jynmPQ0rukYV+2w2djVcjfwCs9MeD1YNseU/O1dTu6RrQLlXxnDoFZmC1/Oo3ERzDfcPdQJoTQCoQlS09dv4S8zcCuspWZCtfq9yli4ps49bJm5Ix+PcP2jT0sjoC3jjyQgbhW2m+7q/z+64MHue4l/dqBDTqN9XYSyadp7SaF3skXOSpk0NW5CBjlJDY3yq9LcY1LNMUs48NXQ2ozd+JKxCT8hmrnKvf3pR594azmp38hicrppd3vuyCL/0X6Sk2psTV0t+puJH2l4/POPyTbGrSKn1cHueKsuCmfPe3VvVRAxQE+uBxaqRABo6GhczT7pv1EclPjltf5Ah5LRGjwFOCDYeYBoSb8dxPq+33BkvH4MB33GQd2lHXF2uKetgHQvjBhWmMB7DFv5em+eYFLPhZHWeJJ4pvGbMo9OVmLh7j7sZ7H6opQVrfaYDAhIAmWJKPVt28wXPnmqkJXyP3LA/I5RvzZWOB+YdnMVWSY+rowuGBA+OZ6htFHWxj9Og7mNi1gyzly3mv6lth/gAC1FMEBpcq8BKSCewYljYwZYcXyC80px1JsScLtVK2ly6BzCqg2wFtWzH+aHuohor2wTU9qyJQb2Q1kq5W6m8sMP87tJNLgjQBrH5Qf8FXNlZve0oHHAZ38AywJqWmHzSOrEF3YFnQkGQpk2mhrQ380pz8qtJOT8fptWg+12pdHD0jXsZQX956x6+g6yrrWRNWwa0aZzhaK5pXBDvZhFmi+H7YXqj2jinc39GcaSVf6K/Q1Xts5y+xvWTK7EWGt6hTHGcrwUWcu8AzvdRlt/uziXz1JIsIIu745YassL6iv6fOD92i8kfZVJ44YGK2ZbZE5PrrSjkUgFZ9JevhL3PYNORFMQ/M14E2wmNLiEcaHZ9f+FtNXg8lB47r+LAXf6dp++RTQ1oLO/RCsShr+OJ/L41eZb9XhizDTRDmE7F5R+vDFWWMsCJg6XEkS+3iZVIF05tNGeGF+UyqWB/vN8kp5llrxwY6FuQLN/ok9P+dqDuHce7XkvB70Z/qyKShymo+lyC0EEQdy3nX4jl+PaL8wJqFvv7JQSdldXudCL1E7dHXFH+z2zKZ2Ibh0HEb3Vga6vB327hhV/0omzZFswoAkrAc3lFnyAe8f1C/mP8Q+DVHYFgAX+TdqJm8wrpXx3gbDJOOTM/Wk927HWc8jN+k1F9gmMq+pamj8sOWVYgmGyv+phLwEmmTJ9tesKmtFsEQHidH4zfnD59SXp7tesnWYt3/HAF/CH4AhKB/QM0ECgYETQywYuP74W1iIksdtt86pMDOHq267rCvUnZvAWYbaKASCFWaeajhpmbfNag9aSHe8nnegOVZzJHEb7iPiwbMpLBtQqRK/ThIhfcTFTQn4dHtCuYbFPMEge0H28XOPBB12hzReKBRTXChTnorr7q+DA9sRPNUHmLZsAj+I+bWkipdxO07SEGIxum2Aegn+mWNmp/r/oZ9thOM8Tozm33XJ34MVcqMniaj9afbdDpDKq/zg8FUb+vMcRC9nzogBY5AhHKjL1D6L9xmoN/U++lhQkFD0G+Ezv3ClHVLjpouBzq7bHBDKc1o1N6OWHaKhlCK2ovAFro/FZAmtqQ6m7srE3tUXonVbZ5mhkl8lA/gAAhjMR5mZlwGcV/NMc4yckVk4RGUMypEr6RgBMth+CiSBDVjICBbLqRuuc6j07feOEY2H+JF/EudHNUuoB4+gi4Czi4f0E8y9eCBimKM2YWubu5XYFHFAUpDihU3JgDROvdCljJq8fJvBzxyL8gay6PqgpYSCjL5oHmem277voK31QXMCxuuZa/Sd0/Cif4aJtSR08DFl7o8DYoeF4qOlF+/6Yi7iNlD7YY+Ol6K82/l0udO2/q6+gmtADchwB4JIUO2JtdTmyvc+E9iqb5AJeqLilD46XhzrcYsvj+FitCwY+jvE5x8ahXsGOYLppeqY+9Rs+CA6u7rBcoGv3sMkhJs83KlKF6DBk6BFFXAqeZ2soAMdizWfyRDsgUhNDArRzeBGkWPTLN2K1uhoy3WJVCHcrR1OJkb8V8UckzAdvWcyyIfYlvF6mxuZMO7gegHe7X98uZGN4/R4HK6uzwTxNjwgnZtq+xxGVMd4yIiiI4Ckr6N2yXXYN6CY7l1dr91lXgFXy03pDNhy/5vX01jM7lMbP/N0IEZT3Y6uT4+ep51vSxIEf5w3xWpQ9guK6iTSxjcIkODzayYYVfhUyCJB9J3qLEGzlDTwkeG0sRpFcdCFD/tNbZMBVOwHvZyM4V8f94AKRHuQYOEFHkVOpGVDvnMVLjXlaFaJstySP5inoxpnZw0yXHafTNmkM4KcmneTOLkjHRhKCIS2HtXdADSxt8ZFHrbw1A5rgoRg9UWrwfipt/zpFhtG7IcYYCq1db/Z0/rkNAybvmMX3IfxL66DCWj5a/0W9TnkqczgAHxjP4A7cLRwwEjah97/ht7HValRpQXkLUs9KhVnbzvVKOeFJ/OGWs3tzcpyG0ab26XQQCk2mrOWcKRSJOBnAuXc3J7nBEpyZzKGcOelc8N/cWzWHIWehiI0a7tqNkEwguLZ+KvWmf43ND7TsqZwFmulNqR8ytSF7CqOy6mlkkSDABMh6GHHHA4rXRkiu3uyMKK3Oqhsp2iTTUnmiw2v6NOGwf6dcLMixgznBwBhNd5n9bmlohkDz3/K6TP5E+bT0tSmPrC5rsQAY91ncFuXdGfTmPQOnonwhcdiYBEJAtxhT3BIXes34VhevfFXaqwWSpX9M+1k5OuhclWZZciGyDVCdyTryiOxhibJrc8GlK2MaN7BSV6hSf1/Kih1W4JNLKOyZiS5gMKkZcaoUuR8fKCSf4dyjonH9L6aadotzRASOZ580l6IMk8gV5v6cW24E7MuPtVT0dmjdURBeaOjKxvZVFaegE2kjP7+jRSnI9HB2Flo3UVAcJcqekoTnJnwjssBygq/EXa/ucyjbSDjPlGelhP9CMAlM9E6F8HsZyM46HXJw/acNwjXdIcUW+MwpkmX3eeDcoGvF+JnaBR6DejiZsGu5wqMQs4HOJ4qZN47af5kVpupFz/mr5dLJ4vA6XvAyyRVDgPNbd2bdc2SweAZ9sFQa8P/3tG1IqllPe5Dwz/L+94gt149VX6CjpwvGWyAenHu4oqWalYxpQL+P3XnWxb4Q501zoX6dpttuJIZzp57EAZ/4oNTvOhgOeAjmX9cJghRtHV8ZkZswdNcTzuR3/RpeMuj95d62dtKpHf0/95yoRTs2mfP9uS3SZhZzn2xULdZrFik0aw1ExRisHVWdb75Zm6LpP9CL7GUSlGtwId1a6XLtvVux1Hww/wRSdh5WcnfjofcPy2hJ/WxUXrNighkxr7RKCUI/9eHkMOX0X7uQyEzauvGAUh1bNSWgFpffYqgypZQ46nz7Tg/szSESNQ96jxlghntLG4ARUWUOB7z3NBYY1KS7SFDwTB82aizggh7Hv3d5gI6ekEsQY6gtzdgriiLs86rZCiFo+N+7WZIk073HYhlRomfguv5QFwnIraf4hQMXEds0Pnf0bMmRI4ZGIEGv7OxWX6RWbHblMn0U/DiJunASCmwAJS7zLECwdj1z+ONbv6QuYcNIa/zmhyAbhGiyL/fimi/5FZiBWzRmI6s/LWG/Ug1GQc1hAGEGGgdXtHhv1U4XXF0wA45itOnXDFRMv1UTn5BdXwE81WZibNmGAj8LjiIFOeqo460xkemVotptDTMP++/tAFFBqA3QQXgsG7aaBr1FJSIZARrQPebPYmq0MgStPThxeGDlO2IzCzZxZ60JkJcY9xmzS7/wGwP/9DANvgFUVaPcrfdn4Gze1/5VNAS4N3jJ7ZpIn/q4q/KXzc+rglgL+HkUSGl6TTY3Svfbdn/6+UGNZal8Fzw35MU5eGHZwll5Hb82pyXFTmhK+8syijOY3QlX+mEZV5oRzTeBScZIy2dPF6iNrjsb/0bAfd1uoj1S6TNbrq+LkOM1gjjcnzgFzDUn3Qf4zQVJXKawxguUjJjGPYAwnvVRluIs+9Sn2jgKBgMPP65ek99Le4ImKhgfLqj90zh0mjjS9+8mjpXmnz5TA2e3JttOH8enFO4EU7VXtj73kGzlKv9Zc2KlPF0aZAgIVJAyrjHwyOuy/AFvevkzpZMgtqjJKoMuprKfmc2mdNP8l6Vn6KpXw5luXTcQ5m+bqCnCNC4ZUEM32SiFxLQLIBGxLSVCU2j0ky7WOXUiuZ7riB+KBjlhgkoIL3hWT/0lZ+Orchs3a/NmrSh9I66adgUvupSs0CLm46i+fNpX61I8wk4N2IQ6Ltw+Ujga8ke2VVwf8gNn8C/DPbOEXXHw0jdUcfUYVtqpDQcHCr/tKEYHWM6LRVYGa2gL4M+DnSdlKhqKLEcAwQpc2neWKfRWKyVoKHns6CXIWGZYTnMk8teLD5vbEgEpZXUwwt76DODoy9vX6jl1s22qVWdY+RwcTeIrvDD+3XmiYuxQE02WxPs4E80JMsqfYT5dYYphlOrIRSljvbaqKoplhBxU+DVXlbjoz7PR8pxej/kKAlLohZnj6USZ8bHJTWrXVdipZy73Ce3w2hXPKlEDXEHDO5droPmtkL32iXhe45LqgSh0saxSGW0NV1qgzVXH2NvyHbylkVnHOyWlmGRLJ8tDX/1TkqDhN134XoRAFp5CZxQY1x6J6/69C6p/o7wS0hviPMLejPMEqwaaAzpmAI8k0CXfyFwjk5MhlfzN2lxyUVCyBb+lVz2td8wjoX/FTKW70Oyb5TkCg2lxI5yJ3E8yzXI2SpRDmjClcmNeNkM4CQd0Ng/zhxq8M50QWIcO/19gnryT2QwTjsGQd+z+gkq2hjZfE2hCkdz34jdlZ3GuoaaJS1gk1tagwvuzmQTYj7fFJ8GPgI9A5pUTv17zYW9CAwRxvWAUKNnQ33H8Rv7b00ss9bd6SBRu8EsEEghurY8U6ZTmiykrBstd4JoVJ9kwklkUolSw2zY/G7qV2EUAOxiA+mpxSqNM/kwMHzGsxXnlkoKEs3o7Cbdbncc0sbpWPCpqRHiMqdi1jLguXptBxwGURHEu7IX9/aEMhgC1RajqGl9CBzaEnGeH0BB7jW/lAp3ueauXGjcXiit92z0m8hWZ4lB4D8O++SVI2yGTq47a8Xt3UFCONDLJmm2+21UV9A3KGRUHHMnqN1i1XtDfkoQ7Y4AhcFJg6Tkd3Hzszf36EbUpp2EJ9JoZHvQ9j8jsgnr+QeRou7dPvXerpVYoiSgfducr2nplbgMPTzTu9cs+dhGsVLpO56SSaXK8FJ+VGkOVYk/SPDC2/nvDghkq06MokgsYCNpfm9MoqhgHh6g5enR9Iif+Ia6JS1yFWd334qZR8mkovyZ8/yXYj79mpKS35I7YxTsEFap9Y6OLge4EYkJXLbHpuReGB3Dgy1YsK6jvijRKGVH2xsbif/repmvh1+9ucITSW2HW9ZGLvLQajTOS+WwTA+nN8fA0agDy6fSqEDROkEC0YZn4llGNo7buFYZ6GwdXTQATsLwmK+gQ9QElJiaKiieXS2ART71fSA6N4fMn5swCmhIBEbor5A8kpaZZ2gM3YXDcWqKmdKIO5EtFJ3QPDnBTgJTG+YIaneU9rdl17Bcpa3jOIpzbxXlBk+2Zvn3KRZY+HZ+2Cue7Ci/i3Iw22Q2FKUUcuEHPbAGbxP1A5k1VDbu24G/VHcvo4bUhCK+84dixmwinayc9wFeiqWE6KoA9Fr6qHQrOR3F38VNkTzh+zKs8kozFr+mZ9YzHbjrF/53Rl0/y3cLSe3lktxSF1jrKnmmzTS3BTYFCQXsr0KcUCLIq0oM5y6LbCQ8zOuF7Aor3laQ/gzi1hIxv89yHCOpzdA1104sZ3rK+8dfdcI5XbShBzrAb+bKodXfipqgaMv6nO94zBDrB2a79SX/zNy63CHlsXBo3q7MCwU9y8tWbVMW+JEd9Bab3W6kpyfY1D2KG3aCyC7VPjqlpkStvSzU1Is3tfAZr0InWqtOZM0nmE3mwkF+zIbjpzU/B6exLj9Jy/w2C5Dqp/Df4G8jkZj+5/UWduln2k+CltUPNemUKGzLQBqC7MrWGStHU4mP1bKVGXKwoU83x2PQvjy2luvyKQvfijdP4tKUeilz2/VfDTLKrEf+IoJtgj7BtEz7xnTCv6igRq8REbH0jXK/n4YTIlpJ3/5kBaG07nQYZ+OQ1m8iCrlabXme8y2hO4l2UhWnCgAH2JCZfWNxk3IFd/F44PyCjn84gYJXOr/IQGKimJidQ08uqf690I18VSZmVGBXkoyF1/l2QYPchPsW0jO2aQlcLcl3v9H1j+X+iH2gZyA9BiEvVEuLdiWm6dNdvuzMUy9c2jj5xh6XZ0Zp34HpgD6N1RB53RMhQjfK3vX94siyf05DBme1HE8gghPiXgRNoOHrMxn4KwCq5hhcW1lfWCuvlCgym8+YQbRaJ56TbUigCHZGgOs4HixkAyLkl05C80vytl+jJsehSyrhC44uz7oqoiPgbUdwUErEEW8rBJqfYsvSKM1w9zgWVzmeM43Y81vy8y/sUHgahndmorzab7dsQFz5pkGC2TwX3yhEfp7/XjD2ZynvHOVCNmp4WM+SKS1Xu1NEIl1Qn4BnqTOjjkv1AVBSZh1ZK+TvGdZS1/lahKxFv7E37khQYr/UT7IKJq9VuIOUoftd44kzp4Q2pT2FVz6JCTrFuqPedpFUfqdTaSUgJcoKBPqAxIXqeAF7WQOaP/vGZyfXltZjuZ3YU5krDceeWTvxk7gkbBKFFIprzGPIiuIqMNYAjX2icuVFPiipClqN0MVfMP/QDaVPHlREwelTNASZdDj2kJue1D2MxqTkejfxmoQE8LnARZStjzWC8wJEitZY2UnY4OejM0Te/lc9AnEjHsYzcRGP1rcyRxqnl3c9UFIogpQ+e4y8KB+DvaG70jr/KIgFB4FL3HBe8L8HgaOQQHdehotj3NTWff6dGq2ywjJm2sGSrxPYa0TwSoE353OfcNUtOHG+ulOxuE3yRC+Po/5s3YTzlx5AcyVYV+58Z/oduRVO+trGUCAYL2nhmhiT3Cm12D2kQOGCkbD62uRIPcimgMT4H7VP3B6r2qAQSsleJeU660m/Acqvu4AXWkHFOPErO7IwVZf7nn6ROM2byV42MebONu0SwekqvXQ5DRRDDBbBMrNiaeL1YxrbUzTh6VX6VkDWzt84AeHmeBHMNY6LQpaONru9DlYBMwmtwLH5yf/ORpIwq6taXKjrqI9O/QcQBDEwI8iV32z1Ceid/Gfn94IZVJ+Vpu3Ap/0k2Fh0TpEtIZUcY5rq0qVUHIx23ewxQOtSZlcj6J1WN4vOSCH4exXZKqhYWrN3v3Bk25EcVU6p8rPBoS91RLDR04wPzXI73NNz7XtoFSMz3pU8CmuyVtldiXMF3fwsi6x8MPVYJGYJH6hdf1v9++Jl2MsOeiiSe0jNhWAz4yW5WX/WcZsfPoqxIOlYJhxiawuKKCZYE+/xe2vgIyeeWZ/TxZcG21iX6amWuXKYGfHlaszqbTSOTz5R8t8FfMVy3AVYWyJ3f4P8ExE83IGyt21SWO2D9yRq/5jsYs9lQK4KVl0lrS19gKe70JdWSqsUh/LOWQuBWg/SUTvP5UteJmd+ATNo+7z6ZLHPX8I5yQ5e86Jah53TBZlWdlJJaVeXJxLA+0UXtuKOWd7Nu2DAhexBI43h45S9RFYTNFepoIad9rmGIN9RTO0bBs3fiy9ylvTaw2XJVBmkkb+GSXwL3MZQjj526Vgrjl/FSZAsYvOHkpIMAI7nS6eGeEcvNqyADwCq5YLpznuB5hnPHQObD39n4415tjBuHk2LV93VFh2mSek9f93DRWwtdIhSnH1N8WYVdaR3bOB6JW8bvTc4Idm97k97Iw++caqz8YPljLBz9BzS+gxjvTIOOhLCCLdtSIBDSzY4thzJ60nA5JEgCZEwqZ4oUVUrZHxdqzA4OcoaTMG7w4DY221yp/oSI3bf7KCN7YaFfeAZN0wR4YGjK9dUU/IPy8tqDnidu7yheKUcxRn9NQ09nfFSSWU3LnO1Z4JaUWRn8jjZjsVBFnm9COSsojMIRO8HZYlQWFYkx32QxfNv74bVgdTRXT7xTeZe26Z7qshQ2tlFtSCWZ+nRqatJ3I9zMjzXV0jvaaO7ToL+ZegVcAtyGkx7mM158csJK51mAkSXGlbBLcW1A7VWYlMTuwNpt9GyF26+HI9ukEaiVXDPpj4x3CfhDJgo1rfiBMH99PQ7e66wR8WFs1nu/Wdh3tWLxd++3IgucQ7rR2gXkFDW8nAe6bAla2BX8jPsHOJeHh9WJJ5V0WI9QsgjsZNvxu4YWMOLG0FvqHQzgI6SZ92TwA20xfA/RX265S8ZZ6LRcwom0lCz3mo85iqtNCxNsIJ2d+fueEjVWiAmJt7jQ/uuFoaR+YpqTt7bvI3eFzv8xqO/nlECwzKXEpWubkGHyvlpsu3CXo8BUpsFrCekl59jaz0n+2Q0kdm6BAdfVOt4575mxUTv6opsp/kK2p6p15MQmnWYB2ztOdqYJKf5BQwVfehy9/kyz7+3aExuAkAxLm17EiZ9bBhSPe7cpvYtUFfN6qZ/S6QNK+qiITSvBO2Z7/CHDe+kCiAsiCUmlxNDb0R5XkAdkn0cE/HS39J5aJHXslEGUY1plimfg9RG0zHFZB7jt9HIdolT0VP+Kjqe2dxQg+7NtnV5sU0hlKH/ZvEiCTNkwGdDT7ejU8t+/ivAJuqtCvlR9F5h9zcfjO1TiUsAPoyQ9g0HKo2wMHpl3+ZVbDFK38ixR5xFqg/glMGd/auQTP24fGQN/fgSaU9WvBhLDjMC4AH//yM/kac7Gb9BD8SMOgN/9YHSj+Vc17zSpaX3b1QPupIZeuNb60ngehfSDurqnt9G7tUGvR8D/v5b/+iTt+yz9VLZ2zDep+6zFkw6OO4ZPVNXCPjueiyFoXVAPD8hB84VyUj7t2O+lM46E/n96jT4Ezo220xE2vyIC1MUvI4hTofQdeeCjxFJn5m94osHDCRE4fN2/9h4vOJRwuCApb+YBi5Gpg8jPC91vLNwMny+P3TlLssWi/kDj04teXwPpKackKMXBg99A1oYhevl2DxDe5o9VCX+U4tM8esba9IBxH/R60gS8CS9/ZtR5/toRjYxFjhSu5kTSbz6KLHGNtvGFN/UDKLsSpUa1rEfgILVgIvDDS06rjtHorkMoyKyi7KGNIIzQZkiJ1TQW+u9g8orzkfuVVS6UxRiYDbcvW2JmnSF0KWzgsT3BRspVnROTBu13KzmruINx67Rqh3XeNAPaYXFhUh4NJ9Rv15Sud0YZY3vejGODAk7iWf0Xbq1TwFnLtob1u2EuZobSImTZHqTa74LAiaGwhRUGfSFzoqUUY94itbwoms9Fu8iKe3lx3j5Ex7r5ybBwIdglc8nRkJW+qBKeEuB3tyNLMe7QqUv+pFKJPHBXDL5FrGT4DZgeWgnCzraaIIKI0JG+EEvJLMBhJIHJbXBMDY3BUn60+0CshaF7Qipg8W8wJc2qzRLn3Bl3EnawWOKWZGMIbvhcCHwSNV9w34pij4H7GAF+D6XFG6Y0cMkPvW8kOWSzLPofPmfZq7Zr7MfpORVXGP9z1O0Of78GKe8GIE49aUh42BI+gq0vuebPUEdRijrXgsFWXaeFqp3cUnQin8uV5Gq8lR6hwX9dV9hv/J7kXRf8bQ/22KUUgw2SNxG7OvvSfOrAaB8qQXvDLfcMerc8dL5iFR44CRMxuk0keJtL4BzcszNDIuFnDVBHlvMHmB2Oa12zq+0YxcC5W4cN4vbCcXjgu+H7X3CfPlZhuZ+cqjLqAJAZVjgrnAUBUwSQjQfOEZMX5/4Elkdjgbsnm7arO35UFM1QeMZobzOix2Hg9KUu6DhFnF/BJXYvPAjO3a8zDy6/jRSX9A5MplUqXLDH/nG3RC363qRbu9yrhvTjnhNC/FpWHtBFTNvI4LFp1t9CX1DIw6tdElZPQtFjLEQiI7/kZslxHjvxinOuIFLte6RTKojJLBp6fkycCUqgMUmHib/FteEIsBmGd5XWZt0SLj7I9PdLJ15Lq7Y71R60FEsMGqnLbOe5iG7PTxBpZfq4a2dsdvpZJbKSpVLRpDzAwBLwTYxyCbHKX939W/MJl7fHuguSRbQOe6EtMSkbTaYcNWc7PKMklCeDoDerqkhi+HetOppQXEYH/h4yFSymunER0a8tTF2WKcC3VUz/EsjTQYuzKwAx7LVheFadwLm0waqqh5LtjdON9hI9nQBiGGgj9u/LfZ/oNSpZJhRs8J5mEAGqlVnzItv+skRkMw5y+Lx2x3ppPuxclfHy16gibyH4R1Th+HW0G5eaiyJxz4jLSakCxm1aimZEuvTuxEMnBzsKg+6HyCI8rOtlTCP7mN7OP2zhpKgKbJdVrtUXpULnDxi1ozyiUcF39TDFl+YesvtARRBbaFuASO88cE1+ON7pnLsauoL+Cz/E6ZWxoNVWFc6VmM8U2D8uFAeK/GU37YsGxTiRO79hZyYew0/DTeELjVwLtzpjuR6ugIm/oyp0DZHH4U6uUIyxdgUPbWS4bLRD9Xm1GmDTvq6YSVDvRXBMKZlVWPeOkxSxBZXXYAqKN5jzVO+CcQAsShkw0WtqHW2KrG0aSzrO+Ddk2lf7CqGK8Vum+hm5G9+r5NM1Q0Vs6qAlRvECpA/3e6eOJxPBhMuQ9CZxq1g1TCvKNi5I9qWG408xWf4xt3vWZ9nZO5Zub3BAHpSOdCVSAegLTGXeZVMANo+Exa+4mAc2EYLIOrrYy5paKUSz/WMn32pgJwEmVvU3au7qX65IbPq3lRLIocsGK2/IkkcVx7+OmKdDLrDFbUflzZjq6LpoDIuuKd8wmM7YC2eT3Qe0Acib01XorNu7Prbf0b5LY3x2+QJ0eyw3H8BMGRTz4nuIZ0T5nXhk8/lY5FyngxKIvx9XgxIr16HcdbdqJZJX6hLZzEGrXUNCXdNfmKnBkJBIR6L6GsIa2tVqZzxYeE5kkQ1TS5AD3w3H+CjhwUmScM57xLTh2VrTAxk/c9KnOxpRDXLlEXk1tG+A33NApfiGEPaBytlx7gw0so5hGI84BHY2GYkjSgLJ0XsDKbb6Jp4ybj3wFRw/fY0n2mogC6XXgGjJrne0PTZNMXgRasZcGLtq9URxVGvsNzx6EtiM69TsO8eNx6WkOC3hiMY9VjRChqWLXsycHYrsTaMuLcrjK9f8EM+gydVDnU+z7fysxDzNKYo0oUNfZwUH7W+F8+inOBBMD4hYmMx8ZC9V2Rj80zcAhqt3Jw20jDf8Id02m4C/C4laVVGtUcJygQrr9U9T2BIpBjdTsDbUPRuUOtnVRdFTalBYS+qzFsUzyMXoO/jLgrtCYSdcjC5TApoiPgzLntA75QWE05Xx6XNR8WD6ewN+btQkKjQTJXXCqjwZBNdkRN5zssEBIsrkOUomfAPoDr0Ja/YjR2eNvdqkwd2HiGUvtV/KBbYgSsDxspV1RDoMWhFi/d0NL270Rl79s9p33H+7rViIBv+OhyvJxaONHgTqz2mpkRknW4ykosBySwRyPUrlTtU4xcjtjKL3erCpmoCzVf+LL+aaE/ps6QxA/dx/XYHXsPT9TV68YZwSn+t+J5Fg0o12PVgX0BqfUQyQIFBP/Qwc2pQmm4cWFZD6jZ8SzHJVXJ4fV+XIktwVdL4Zm10Nm4P0QcAjzWL8GUnKI9GSPMW+97fag2546Zxo1cIN4jL8v4EprNikQ3mCEEIC4VPWw5leKgw5oPys7UcPuNJXJJOAvh3JXm+nBp9aZgC/Erk5Z0y4euxJBVPq+XOJmVsdTxfljTjZUzYFeuLCPSQWIF64ra9YDHgLLLMeGdCWphaSPvQ37pBQEqV0oKowSBY7fVqTchWe++BI9NGNepRQ9sR8tR/2nV71eNJxAJsuewc9xRBpbnlzaN+ecAAeTIKxvEiUH8hGtxlPvDvpuXS+5jNGaVFMumRg+5zGr3NRAq6puXO9I3J4AnMxw/BPeItyNAL6QbV9eY+Iia3BPRzkF88MsmZj7vs0MiyN2GodYf4H60Z02Q44rODR9VoZ/AMb1bY466QQHb0c70HvequF7A+5smipk20YmpMu0H6TgA8dbsuQ73JEgxY/S1ywBlXkxI7ZyJ3i+1CaZvdj3Xl9ZRP9IfnZIn52ANkWwynP04LGNDUc5m7Smp3MLFKJ1SPmseY+6PP6zml+XP9247882as5zLgmo3lnn6gn0H65V6p7sOO2HNFv6/d71/1aVjccR1nLH18wibhV/Vj+wUUEK8n4smX6M1hS9aHc2rVO/UFPLU+cnV/h/R8eJiwLsXAaCd9fZMNR48PlE36lE5MHp9iCCdFNTTQRONa+x9wNqmuNqmp2+YB+9FuC3fNOQ2BAagqo4RHa5bASxT7+rK2wWloK4dfUJTSB7CKF3XfMMeZQ/wFbHQT5ct9mRSw61a4GnEI+yI78oyN37IywULxbFOlpoxPyyykI7iETMWJkuvAZqz4uM3oW03IooiYZSyS23AysgwuKdTq0Ww0pMVMOvFejbseJYmbfHGUNzKczIrN7XlgElortqR+hKYQwIHkevZTngjf9XMBUny6OuniY6v9EZpQu1TpqTm4LOeoag3BFF4B6AHrKmaeHzzCYVQwStqtaeBR3se5P+sAb5cOR2oMoN9EZRzcRpwSzOVfIGGlIkyTLWuvoBVG34EAAsCxHCBz2GB6ayQiPwUl2b5RuVhuoxsMSpo7Sg1AnuK3tlBum3hXBTJKE1Vewo1khCAUo71aBbcagoPJl0eJnf1vq1LHcp8dqx7aD9xVoIugEW7hqaKWCQz1fMYXZ8U2tUj6Gtn4n7cp8tmDGhsmyrtzBqnL+yHWLkvkz18zwGGe+6Kagr4zHLLQDodDgrgkMzppwiFYea1TIhzWelLtP2uYK8IdycvpLTq90ZQbIllkQvJI2jL44lRM2wLKZc/kK5XPjsZ0KQldEvRAFltVZmmZLZ4red335Z95Hhp3tvHs1M+hfpGsxejPknqz/X0/7AuhbULHS0Bivq5/zwiQmqnMkd4AMUi5mLgZ+YX2c52qLhNd+M/1u55P57n9Gf4GGbRGvU/dMGmAOIFVOdw2idfezUhSz6lnvRXtW09pUlQKCVHyzgcUj8f6nz+reyruBwOAR4eILSUo5XDlIohb9fprkyqAOgwDKC1gyYgxFGNCB7v8KhdbyT5eP9u+qOxQrdPQCL0N0/VoL41Z/3R86LmC6KFOL/UNyU6DIglADsW0apQtZt9TjXViWeLcl0VfuYZp2UNXOSzZlxLF0Mq5BlGN8aDJf4xwoOHvBXUui23K9pDEg6EyxISO1FNNXr8vl0K5dCo0CH0gSK/n5JvNvidJs5pEk53MM6UqVYnvf4lpLqUGIhjy0FJk9LCUM8Fn3tveM5htTBcxiUtEWIWo48H4Mn4koGJjR2mQk4IYfFRgQHEE+5aPu8nNr93YuY+zv9UYjI3CST0BbKFuf8TFXxIvoHTZDqz+EQhM1MohoTvmVpClrJaDdziyIWvO3SuD6ozco6A1QeO/HXgE+yybc5GjSnK0mtlc5bCMS664ZoSvtdwY/ixFZpRYZqqXLKXqX1n+D1s3m0Qpjt8P5L8P8aJmDKhCundLvkv+8PwtmqgBn/ZJjaA8lTpjd0uXiHLm29tHycNxKZfMz8mKID30UW8eaEe3omar85VKMKdFEkN/zr3ncegvL+QAYudaA6LGGtTFiKyYvVHERthKOZobUfEcSf1arQFk+qu4ICaDESwg6ROFl31xtcWrDuSRMVJeA5jynZKBSo+o6cdUpw4iWTjPsG6WL7/Y7qDT2xT4y4r+Czl+SR+yOj85hd8a+4ZPmNWmSN+gAju6xTP9A5lFaVCRQ8EP3QMGjfjDX6FMYPrEeIyXkEZofjWVK80Hy8jos59El9TGZQtZNRwmI3mIRtQBJebltpIldaKTqnktRqaE08bVOtrH3fB23BBDcKu2zjYq3ZKO7xBh1+N0q7zKXUcpVmCx4DjSJaRoetLPJreVqZLT3jYzYxccAgr1z6++SQIfDSjl06oL1QtvqVYBizZ+HlGkehqMg+pfOA3I7r05UGqhZSpqEfEz8IkuZdvdZDXX8VP5j0NgYm5wbN7/73Iitw9oz7dSldotdtnIb2TWBrt47LYf9CU/3KcRwtfjsp17yrL4V4CcI2Um2jSl/S6KkSeaoJcD9uz+GWm3Q1igQYy5sC7ihjYCUnp+cPepkFpQzbfb8+U/82G38P0z2l/LWGYMI4GKvfNK/S6tweqxiFxn6LpQuUijbp7/KIJBsQVZggYk/09rDexG9oRNG2T8w6Gr/soNUp0JzCXcPeaooJa4sE1S2ksW6UWN8LPCpJ86FTNU6ur9AbVdOuvMGvFSgG4UgweG2dK+cbCRgotO5H1cg1amUF1KP0a76r0yn15jTbI3dTDMGWfFFNhw2esNRlnuDEIi/iTlABiKBQQIDkZuHMO0f560GNilqFMl5oVN6Qgl0p5QeACfSdBHctG1SFOUnlWkj1o+bxEVwwum8FDQcypEoCx+Gz5wxhXw81ACOTCBxpmRrFUmdghYCw4XsCkOovvBFKzdeAkfpJtK3fcnx/zw9Ar2WpuGzbkW5SKVjtDHNbJKud0h1U7KnXwYw599IPiIbn9V+dsh1qrKm66NLEwIhwLWDUJ3xgVC1G38enXW8nREup1xDrKSCOYKx9H4c+LXeneZN+x6XkM8Nw98U5Y4YOatAZV7wePEYunRVFseZimrEPzZY3AEUD/Gqw5jE2lBjG8ZjMgHjwSnV+NoL18qNFrRPNJDoCvam9NEied3uxxFqyEf+0SWbDa4m3CCAnksGuVBy36MDauPnTwNTGFVTad0i4vqz5QsN2ubAYBR8BAc8svDKSdSUd9oJvf5+OEM75hgMgegjzwfDIZ1GsYOKGN9ZSRUMpDur8hhGLWwuu4IDhXkcbyLanYgr7DqTKWPgHSL1O7/pn8tfiJSVTP+YRcqbqBSC8yzGjhV67/K3tPjNXBKtnwvOSL0uvHQ3luwqwW4y5iAhbClLxV3lriu/Oy7v4WPxT6Bv23ukGXX7/njO3aEFFpv9m1KwFgY9hMm8u8Nf8ZynhgNXJ2rziqbc5YOMP+0oxzFiwB/+AViSZt29wVb3E6srjnZGoD10NBYf9tMV8ik9oDImudRG11d5nhwMMK6WEsTAnEPljfKDlv8nVSeg8+dNbLbxkIcg1bnJYnuWGMxOZXOCWcN8gMwJ5KtXwg1eC94sOaa7okG25XnRqtwN7UvM6hm4Tx4kM3nhRqiwgSdAjP8R+q9CQRStt65KkF9iAnc899NNKuqcQe4L2Shek4XZ9EQwvUvF0jZzpaG5O3iYlga4XGqI2PrlMhSX1MPl9/g5XzQJezf+PIxKL+wytbPn8rMMA/P9qrmrWUlTmteSBaoztGKUXGZ7pnOApgdsI328vAnGx0FlwYUGKJ217w8vmpkJEpHV6vXhAl4FlKLBaRU6C/k4RJXp0VP/SOufTrOjcAnxzhZkhH3xi/yqBSrwf6C5JwOmys/UyJPj9Mc7p5Cfv7kKJX/+yaTNoLr0bsHLN2PfGaJJWARTwdHEgFeBu6IKyAUxSb4fMUVBVpUz08k16XI4zALI+GpQz/AKp8Xlc3D98vHsbiIIfn69HJxWJ9OuQDnTToBW3NJ4KPHGZc5LpQju7RFsITPL6wjF1PusrObSVci+KGVQCD8FlhcPc9mejnVZR/gdVWkh8zb9qmV6cGL19uuMU8+NM+oO12mKpXkcwf5Krt3vs2ViI3opZ8VlDEv2+NOZ8RNVtUPVTNxR2qPLtKYDzFfcnGkwY12fsL4dXQFXw5N9BquXfDFokLyzpK7u7UVhcbPi6ko8Rgbxa+gpuITaduF+mYDGwsBiRYR51YD5CDw0TRQD4x/OKLaSGQBteobQLNxIKzqHpFpT8rQTGie9sgKVzTfh7wnAvz/vonNYFtYruvIEPitwaPjcBc/9Fkg6ISn/xIhsRq7hEp/LR33CUif+qjm/b8QcLcSgb2OpV8+mSjSXk20K8ZnkrGZborN/3AA9DMRMv6dV3tpTUtR5IVZEr3i2zxxipYKcJwAsFKCHITMaC3yyaR2x9w+cPZix6C0MSCG7Glwiq0Qh06d5xnMkKzZJa+ahZc2ngNxrykoxDLPicjZZKcQ4MmN9kcd7DBo11fP2G1xkVOgjXiBtZNkB3vSMo1/04j8+rOzucWwC+oz8FgYVBb16K0wGjaF2cayOEpErgzx0Cuhn0bR0g+Uyb6Ce1HbX4jJbKfJDHAJrGlm6BTxI1/gkCYZTgmpo1brKiJeJj/QpixuAnomQITGqLcAKq8Fm+1hc6gjUkTPuMp/pJCpF9MSydKLhs6/kHqgty2KO6aeSa+xe/Ru3KZfUhaMC/c/aZzW3XeEN9ZQK8kaWQIpsThya8wwxpS/weQ/enicOgsDgN3JyDKfJxPf6kIjtjuCcG3DuynkEoVeSXyaa1uWIiJVXVn87hXFQYazPRlz8hN/trs1n5AIu7Akl3/lYvLlVE/KJc7Zx3OAgrq/gMrJwCCCYW39LF8bq6sikhNZqyji/z5VyT0DzNc4CA4gUe62IEdIVaP0dxvW6h0k4mZfF8nM9z0qVKvv4tcFPKFDthFJ/4xSNUpwbfQfhRH+j8D/wh1s7A6iPW2+Jv0nHP4OElI9SA/dOrll81BAE9GFtNlcAKmRQpG5wu8cLmFIuG19ehTT1BJ7ajpCtr776Hr2iHwfCDfnfZrjWTUkgIW5NBfF51kwLJ3+YvXV68SKSQYLs0mLhbX0FHiEJMYFE3pQkNNfpinAAJSvssAnJPzmuSooWF63F8jHPpcMZ8AVtiMi0NWatLpVcciO0TsslzTqqiQJvHU3ct2wAvSPNjXHPwU0yCrxQTLETv4poBr6uuC8HSswGVbVoMaaeIp6v7GosAzsPLxIv68PJC5zE7RK6XYZeUrM2nXyxxAC7FPyn/J1a+9OVb6q9msnwCI81deTCS5PWFQRsH3uzmepFlDymvjdg5JrJlOwsidHFLZ2yuvbOsqeJO9n4XaVZpgT++GURfHIgzl6XaQYyDUB30qd3fT0TqVY51Wrkwp5OK1Bfsx+qde0hxbbpl4j7Sz3I/Lkv3mEpFSMW3fbmaDwytheRIIVE3heH9RMsR9Ka0L5q1BZwBpKlDdC7w7OBKq8BTNatYxmJx0FTpAAxnAKG4SEI+Cw354WLMEDo+GQ2dT0NlWjNouXsg+88l2FETzOaq7a/m+hb1dpaq6OP+MZQvTu+JyWjORmp9OpRDPaBti2/KVV9abZB4e2m1sx2JSQJPTzx92NT9dy93j04lngN5y4zMeI0ju6gBJE0y0XKeCV29AAwJ0m47Y4vNlRKLkeLr306MjzJB+ukS0+0J7h9ry7Ze+cXIlUZeY0vUSr/IMeYBexvrus+h76VJcbvdfUuJBzSvYBCRR/HZbOGrZepfPMD6/WOEFcGQ6EnWnT+NqHWIxixmeaa4258R8yZLtU2XY+SCK44vwJuLkq5fdt/3+bG5mW/hBvtwmLrgFOzVv69XWC/xSoSHTYZXghVRYdhx56MUeAxOn3z+o5VjFKjUuXk3toPlvhUceH1imRMN0s0RJGPCFpmKQhH4TdZp64QhqIJ+H2PqOE24IH//Va0ZLUpT2BXv/dkpXS3VUzl/PRaR+f+keYxl+uJL9mRFi9IPJglD0UIkp+IqB5PMhVcwHkB0icjpH3h24BFcqM6lpoG1cqnlMST6VBgwK6zfBpnd5xrHcmAwjAm5rxc5W+c1IFSoW93ts+ux5khi8DcFD7zF4IFTMVAAtrjb51JRvM+Q261RGfB6DUD2uYuGxal5ahcKktvkaFQphIf20Z7JG6SdwQuFyhqXr+eQp1PJhVuii1sYDZ+CXdNgyLDcvkGUgTiM+qZym5Q1vcbhr8EbOl9JuGWoVgRI7RxIqtkkxwLaSZCjHyszbGtVI8iQFLSethjVxH1s/eEpbL3bzsdsXMvRRe01Nse9HYlZ3YouxPz0770SX1c8obiCSY0N3/F4g7V1qGiL42Hk6wpzvABYPmHA50zqdq9OsUa59zrIUNGsV7+bBjrhZjOAP3rXU86/fKL8E1zZPUhAPyBcKbOColl5aGQWLFjcQu6Qjxw+cM2FC1OAwkWtiHEJctzIIsgYHIG+7FgOoK2SPAW712qF8EExr3bZOUQ8qHlr5s0kEmFvm4eIloprs3B+bDXjvuuvJk+YInjXnXq3iuveE1LxpDHz8+bCKZBEriLdk61e5A33JWF9Ihchoe3TuKU9THfmdIHac0drP8nnjei92MqB6/eLTEX1T1OfN87AMQyVPQjOH7x/NTaXOjXGT8J5V0f6b7lAC/2HEvTqpfvStilXj2nn5MaT1/lhGOZFkHAH9ap/Sljykw6UZ7WUadXQuCbDyO6K4JzhXHtFIom2n9EN1vb/26OlUdu5PWxMVAL/FW6Gu9H/zWfn9cmOVfmTdFJI6kRKod6u+XI0EDN9mMfeTlihFvMiseU6/fQwLQ3sbqb2FRTgitrRY9N/vIsljlpfqcCgmhtsbYCPIqRPLIROcLNurb6svfWmud+/akmkb3hgeoV0JmJfBCIQja3xDkSddVepeQH5QYiVHyMlgupsq/4OjRbgtMrf7Fx19g10dt0xhBlrS0JmSNspg65JNzuAjKa+4nS5d30y4r+488M2HSGdV9R2NJdx6+maQHld2WNumouTU70sBgUB0XiM/fNifMSitzDRvx53cybxMPB2t6hvCorZxNgZ592Ojhs22vCP7y/kZLRGeAlJ60nKDfDgzLYQanxOB1M+dOZ0htwXISpaB5E8H4xjb2VP/bvZ5UZ5sxvHceStzWF45/1Tx/Q7kj6Lbx5k9uNhbz+GdDcDRBtqFuQuhAYoKeGBNkrfbZh50IULrAV5xByWCjC73t7v7cKsi+/ONSziUj3RsifhT4D1E66EWCAFPuyCkBFi6i5sdoGnaoemTqcqOAZM2AcYcUPYmbYqph1TAhgjw4bAEiTlWSbOCFvSVjflBuONLzLzY0h3TTCeRNqsmP/i3h7M8cIuX0TIKvQ4IZ7ETRK8qOW7Eys5OJaz3RdJODfDIm9WvKDq+iPeWAKPCijvkCnafadppIx9tXM+265on7HQqQhkqCyej5GN8muQJgNPGHubKyPkja+raxKHLJPlx2kZ2tPCm9aXSxtc7I0WInlblhQrktKsAKwNOH2IHSORmF+Xm7eiZL2YK2DhvpSuRa5LhevQpFgJNpwL+iqHmNLv0NVcjIlFv9l5xsDHa940in3BpG75uh2HB6y3kBObYLHjFfCE646OwMsPcWem2useCO2xX0GPEFjUFa9jhtquBxzcZuW55Tnm2KM41Se/gve881dLqj4eypYLvA238DwYfYHNiCfuJcVKUFmp9u4e0MMhnB0Mk1FSHx4dqCOI1IdaRZn60EqGn5To/tVTDxyd81tQbFHxHNmI5NRRNM6M20/nJIKcqS0QVkXGYLYivum6LducNGmU9/Swof5w99Sj8fgJZQQxdPOz2ILNYrS2iYPjty/zoZgWCMmqO4o5WidE5M7PKhBklKAyFO2PmgNXqkLopVMhcBUpy93yVKB9/sIJC9FujQl/20SOWcqoUKsH+DcrN/QRaopF26GVD3+RGecoHey1/xoALdro2D/zzJbHC5+SdQJuCT0jz1GGkOMW28eI8b6M9ySwXlK6/uvNhfki5nGcFcyLcqHXoTammjtMvutoq2cvXcpFDJkeom0zJXLDmKfEGztTMzhDT7uR2tU1PW9NoBt3xMF8T4XL5dxX15x4h9TbhyJDdozxpE3kLzYN8gaCu1J/iRdBRYBC6N+tPwHe7eOlAb6nafJYYZlmSBLEQNcIsw/Fqf6FSmWh8BQtSGkHXB3LKbIQITTtuhPHlbvLkUsaFi5Dct/kGFfbKeM9+n55IBS7I8tqDLN2HpY1/lEIkBaNiKVT1QObyYSt1Y4Fcx3zS91y8kQ8Qm8jLLf82UkcQt33owQpCUG9Ab4INNtdFFzIL8lg4uR0/Ym7mDiM7lQnzmBhifptqH7JNrMjvwZ9uLJOIxuwHgCFYg3/EG+9GBUZTWeP4GW8Sn/qbP0xdJp+WQ3QIm2xOmNAmRgjbLz8PnK2mHat9Tz1WZQ0jz0K651qVfPwEa5E4V0qn4XbreIEsENjzVtG8X7/6URgu2WSJAcFX3t4KI2dtJ94mf0g6ZZstng/gSZ6U2if/GMpPj214W/+Dm68XTcr3c1qMZbRtED9KnVszO/BpS8JtkUxyZ/VW9iMhEmlJ4XIVbgT7wo/3NLPEhNDizbg5NAWe8IZ5vP2hP8ss991c=
`pragma protect end_data_block
`pragma protect digest_block
6759f066ea717a8711c0656c6ba6ad4f5ed6431b451575cb492dd13f5ff5c99f
`pragma protect end_digest_block
`pragma protect end_protected
